VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 11.475 203.925 11.645 204.115 ;
        RECT 13.315 203.970 13.475 204.080 ;
        RECT 16.995 203.925 17.165 204.115 ;
        RECT 22.515 203.925 22.685 204.115 ;
        RECT 24.355 203.925 24.525 204.115 ;
        RECT 29.875 203.925 30.045 204.115 ;
        RECT 35.395 203.925 35.565 204.115 ;
        RECT 37.235 203.925 37.405 204.115 ;
        RECT 42.755 203.925 42.925 204.115 ;
        RECT 48.275 203.925 48.445 204.115 ;
        RECT 50.115 203.925 50.285 204.115 ;
        RECT 55.635 203.925 55.805 204.115 ;
        RECT 61.155 203.925 61.325 204.115 ;
        RECT 62.995 203.925 63.165 204.115 ;
        RECT 68.515 203.925 68.685 204.115 ;
        RECT 74.035 203.925 74.205 204.115 ;
        RECT 75.875 203.925 76.045 204.115 ;
        RECT 81.395 203.925 81.565 204.115 ;
        RECT 86.915 203.925 87.085 204.115 ;
        RECT 88.755 203.925 88.925 204.115 ;
        RECT 94.275 203.925 94.445 204.115 ;
        RECT 99.795 203.925 99.965 204.115 ;
        RECT 100.770 203.975 100.890 204.085 ;
        RECT 106.235 203.925 106.405 204.115 ;
        RECT 111.755 203.925 111.925 204.115 ;
        RECT 113.135 203.925 113.305 204.115 ;
        RECT 11.335 203.115 12.705 203.925 ;
        RECT 13.635 203.115 17.305 203.925 ;
        RECT 17.315 203.115 22.825 203.925 ;
        RECT 22.845 203.055 23.275 203.840 ;
        RECT 23.295 203.115 24.665 203.925 ;
        RECT 24.675 203.115 30.185 203.925 ;
        RECT 30.195 203.115 35.705 203.925 ;
        RECT 35.725 203.055 36.155 203.840 ;
        RECT 36.175 203.115 37.545 203.925 ;
        RECT 37.555 203.115 43.065 203.925 ;
        RECT 43.075 203.115 48.585 203.925 ;
        RECT 48.605 203.055 49.035 203.840 ;
        RECT 49.055 203.115 50.425 203.925 ;
        RECT 50.435 203.115 55.945 203.925 ;
        RECT 55.955 203.115 61.465 203.925 ;
        RECT 61.485 203.055 61.915 203.840 ;
        RECT 61.935 203.115 63.305 203.925 ;
        RECT 63.315 203.115 68.825 203.925 ;
        RECT 68.835 203.115 74.345 203.925 ;
        RECT 74.365 203.055 74.795 203.840 ;
        RECT 74.815 203.115 76.185 203.925 ;
        RECT 76.195 203.115 81.705 203.925 ;
        RECT 81.715 203.115 87.225 203.925 ;
        RECT 87.245 203.055 87.675 203.840 ;
        RECT 87.695 203.115 89.065 203.925 ;
        RECT 89.075 203.115 94.585 203.925 ;
        RECT 94.595 203.115 100.105 203.925 ;
        RECT 100.125 203.055 100.555 203.840 ;
        RECT 101.035 203.115 106.545 203.925 ;
        RECT 106.555 203.115 112.065 203.925 ;
        RECT 112.075 203.115 113.445 203.925 ;
      LAYER nwell ;
        RECT 11.140 199.895 113.640 202.725 ;
      LAYER pwell ;
        RECT 11.335 198.695 12.705 199.505 ;
        RECT 13.635 198.695 19.145 199.505 ;
        RECT 19.155 198.695 24.665 199.505 ;
        RECT 24.675 198.695 30.185 199.505 ;
        RECT 30.195 198.695 35.705 199.505 ;
        RECT 35.725 198.780 36.155 199.565 ;
        RECT 36.635 198.695 39.385 199.505 ;
        RECT 39.395 198.695 44.905 199.505 ;
        RECT 44.915 198.695 50.425 199.505 ;
        RECT 50.435 198.695 55.945 199.505 ;
        RECT 55.965 198.695 57.315 199.605 ;
        RECT 58.265 198.695 59.615 199.605 ;
        RECT 59.635 199.375 60.980 199.605 ;
        RECT 59.635 198.695 61.465 199.375 ;
        RECT 61.485 198.780 61.915 199.565 ;
        RECT 61.935 199.375 62.855 199.605 ;
        RECT 65.685 199.375 66.615 199.595 ;
        RECT 61.935 198.695 71.125 199.375 ;
        RECT 71.135 198.695 72.965 199.505 ;
        RECT 72.985 198.695 74.335 199.605 ;
        RECT 74.365 198.695 75.715 199.605 ;
        RECT 76.195 198.695 81.705 199.505 ;
        RECT 81.715 198.695 87.225 199.505 ;
        RECT 87.245 198.780 87.675 199.565 ;
        RECT 88.155 198.695 89.985 199.505 ;
        RECT 89.995 198.695 95.505 199.505 ;
        RECT 95.515 198.695 101.025 199.505 ;
        RECT 101.035 198.695 106.545 199.505 ;
        RECT 106.555 198.695 112.065 199.505 ;
        RECT 112.075 198.695 113.445 199.505 ;
        RECT 11.475 198.485 11.645 198.695 ;
        RECT 13.315 198.530 13.475 198.650 ;
        RECT 16.995 198.485 17.165 198.675 ;
        RECT 18.835 198.505 19.005 198.695 ;
        RECT 22.515 198.485 22.685 198.675 ;
        RECT 23.490 198.535 23.610 198.645 ;
        RECT 24.355 198.505 24.525 198.695 ;
        RECT 26.195 198.485 26.365 198.675 ;
        RECT 29.875 198.505 30.045 198.695 ;
        RECT 31.715 198.485 31.885 198.675 ;
        RECT 35.395 198.505 35.565 198.695 ;
        RECT 36.370 198.535 36.490 198.645 ;
        RECT 37.235 198.485 37.405 198.675 ;
        RECT 39.075 198.505 39.245 198.695 ;
        RECT 42.755 198.485 42.925 198.675 ;
        RECT 44.595 198.505 44.765 198.695 ;
        RECT 48.275 198.485 48.445 198.675 ;
        RECT 49.250 198.535 49.370 198.645 ;
        RECT 50.115 198.505 50.285 198.695 ;
        RECT 51.035 198.485 51.205 198.675 ;
        RECT 51.495 198.485 51.665 198.675 ;
        RECT 55.635 198.505 55.805 198.695 ;
        RECT 57.015 198.505 57.185 198.695 ;
        RECT 57.935 198.540 58.095 198.650 ;
        RECT 58.395 198.505 58.565 198.695 ;
        RECT 61.155 198.505 61.325 198.695 ;
        RECT 62.130 198.535 62.250 198.645 ;
        RECT 65.755 198.485 65.925 198.675 ;
        RECT 67.135 198.485 67.305 198.675 ;
        RECT 67.595 198.485 67.765 198.675 ;
        RECT 70.815 198.505 70.985 198.695 ;
        RECT 71.275 198.530 71.435 198.640 ;
        RECT 71.735 198.485 71.905 198.675 ;
        RECT 72.655 198.505 72.825 198.695 ;
        RECT 73.115 198.485 73.285 198.695 ;
        RECT 74.495 198.505 74.665 198.695 ;
        RECT 75.930 198.535 76.050 198.645 ;
        RECT 81.395 198.505 81.565 198.695 ;
        RECT 83.695 198.485 83.865 198.675 ;
        RECT 86.915 198.505 87.085 198.695 ;
        RECT 87.375 198.485 87.545 198.675 ;
        RECT 87.890 198.535 88.010 198.645 ;
        RECT 89.675 198.505 89.845 198.695 ;
        RECT 92.895 198.485 93.065 198.675 ;
        RECT 95.195 198.505 95.365 198.695 ;
        RECT 98.415 198.485 98.585 198.675 ;
        RECT 98.875 198.485 99.045 198.675 ;
        RECT 100.715 198.645 100.885 198.695 ;
        RECT 100.715 198.535 100.890 198.645 ;
        RECT 100.715 198.505 100.885 198.535 ;
        RECT 106.235 198.485 106.405 198.695 ;
        RECT 111.755 198.485 111.925 198.695 ;
        RECT 113.135 198.485 113.305 198.695 ;
        RECT 11.335 197.675 12.705 198.485 ;
        RECT 13.635 197.675 17.305 198.485 ;
        RECT 17.315 197.675 22.825 198.485 ;
        RECT 22.845 197.615 23.275 198.400 ;
        RECT 23.755 197.675 26.505 198.485 ;
        RECT 26.515 197.675 32.025 198.485 ;
        RECT 32.035 197.675 37.545 198.485 ;
        RECT 37.555 197.675 43.065 198.485 ;
        RECT 43.075 197.675 48.585 198.485 ;
        RECT 48.605 197.615 49.035 198.400 ;
        RECT 49.515 197.675 51.345 198.485 ;
        RECT 51.355 197.805 61.725 198.485 ;
        RECT 55.865 197.585 56.795 197.805 ;
        RECT 59.515 197.575 61.725 197.805 ;
        RECT 62.395 197.805 66.065 198.485 ;
        RECT 62.395 197.575 63.325 197.805 ;
        RECT 66.075 197.675 67.445 198.485 ;
        RECT 67.555 197.575 70.665 198.485 ;
        RECT 71.605 197.575 72.955 198.485 ;
        RECT 72.975 197.705 74.345 198.485 ;
        RECT 74.365 197.615 74.795 198.400 ;
        RECT 74.815 197.805 84.005 198.485 ;
        RECT 74.815 197.575 75.735 197.805 ;
        RECT 78.565 197.585 79.495 197.805 ;
        RECT 84.015 197.675 87.685 198.485 ;
        RECT 87.695 197.675 93.205 198.485 ;
        RECT 93.215 197.675 98.725 198.485 ;
        RECT 98.735 197.705 100.105 198.485 ;
        RECT 100.125 197.615 100.555 198.400 ;
        RECT 101.035 197.675 106.545 198.485 ;
        RECT 106.555 197.675 112.065 198.485 ;
        RECT 112.075 197.675 113.445 198.485 ;
      LAYER nwell ;
        RECT 11.140 194.455 113.640 197.285 ;
      LAYER pwell ;
        RECT 11.335 193.255 12.705 194.065 ;
        RECT 13.635 193.255 19.145 194.065 ;
        RECT 19.155 193.255 24.665 194.065 ;
        RECT 24.675 193.255 30.185 194.065 ;
        RECT 30.195 193.255 35.705 194.065 ;
        RECT 35.725 193.340 36.155 194.125 ;
        RECT 36.635 193.255 40.305 194.065 ;
        RECT 40.315 193.255 45.825 194.065 ;
        RECT 45.835 193.255 51.345 194.065 ;
        RECT 51.355 193.255 56.865 194.065 ;
        RECT 56.875 193.255 58.245 194.035 ;
        RECT 58.545 193.255 61.465 194.165 ;
        RECT 61.485 193.340 61.915 194.125 ;
        RECT 65.355 193.935 68.355 194.165 ;
        RECT 61.935 193.255 63.765 193.935 ;
        RECT 63.775 193.845 68.355 193.935 ;
        RECT 63.775 193.485 68.365 193.845 ;
        RECT 63.775 193.255 65.345 193.485 ;
        RECT 67.435 193.295 68.365 193.485 ;
        RECT 67.435 193.255 68.355 193.295 ;
        RECT 68.375 193.255 69.725 194.165 ;
        RECT 69.755 193.935 70.675 194.165 ;
        RECT 73.505 193.935 74.435 194.155 ;
        RECT 69.755 193.255 78.945 193.935 ;
        RECT 78.955 193.255 81.705 194.065 ;
        RECT 81.715 193.255 87.225 194.065 ;
        RECT 87.245 193.340 87.675 194.125 ;
        RECT 88.155 193.255 89.985 194.065 ;
        RECT 89.995 193.255 91.365 194.035 ;
        RECT 91.375 193.255 94.125 194.065 ;
        RECT 94.135 193.935 95.055 194.165 ;
        RECT 97.885 193.935 98.815 194.155 ;
        RECT 94.135 193.255 103.325 193.935 ;
        RECT 103.795 193.255 106.545 194.065 ;
        RECT 106.555 193.255 112.065 194.065 ;
        RECT 112.075 193.255 113.445 194.065 ;
        RECT 11.475 193.045 11.645 193.255 ;
        RECT 13.315 193.090 13.475 193.210 ;
        RECT 16.995 193.045 17.165 193.235 ;
        RECT 18.835 193.065 19.005 193.255 ;
        RECT 22.515 193.045 22.685 193.235 ;
        RECT 24.355 193.045 24.525 193.255 ;
        RECT 29.875 193.045 30.045 193.255 ;
        RECT 35.395 193.065 35.565 193.255 ;
        RECT 36.370 193.095 36.490 193.205 ;
        RECT 39.075 193.045 39.245 193.235 ;
        RECT 39.995 193.065 40.165 193.255 ;
        RECT 45.515 193.065 45.685 193.255 ;
        RECT 48.275 193.045 48.445 193.235 ;
        RECT 50.575 193.045 50.745 193.235 ;
        RECT 51.035 193.065 51.205 193.255 ;
        RECT 56.095 193.045 56.265 193.235 ;
        RECT 56.555 193.065 56.725 193.255 ;
        RECT 57.475 193.045 57.645 193.235 ;
        RECT 57.935 193.205 58.105 193.255 ;
        RECT 57.935 193.095 58.110 193.205 ;
        RECT 57.935 193.065 58.105 193.095 ;
        RECT 60.695 193.045 60.865 193.235 ;
        RECT 61.150 193.065 61.320 193.255 ;
        RECT 62.995 193.045 63.165 193.235 ;
        RECT 11.335 192.235 12.705 193.045 ;
        RECT 13.635 192.235 17.305 193.045 ;
        RECT 17.315 192.235 22.825 193.045 ;
        RECT 22.845 192.175 23.275 192.960 ;
        RECT 23.295 192.235 24.665 193.045 ;
        RECT 24.675 192.235 30.185 193.045 ;
        RECT 30.195 192.365 39.385 193.045 ;
        RECT 39.395 192.365 48.585 193.045 ;
        RECT 30.195 192.135 31.115 192.365 ;
        RECT 33.945 192.145 34.875 192.365 ;
        RECT 39.395 192.135 40.315 192.365 ;
        RECT 43.145 192.145 44.075 192.365 ;
        RECT 48.605 192.175 49.035 192.960 ;
        RECT 49.055 192.235 50.885 193.045 ;
        RECT 50.895 192.235 56.405 193.045 ;
        RECT 56.425 192.135 57.775 193.045 ;
        RECT 58.255 192.235 61.005 193.045 ;
        RECT 61.015 192.365 63.305 193.045 ;
        RECT 63.455 193.015 63.625 193.255 ;
        RECT 63.915 193.065 64.085 193.255 ;
        RECT 67.595 193.045 67.765 193.235 ;
        RECT 69.440 193.065 69.610 193.255 ;
        RECT 69.895 193.065 70.065 193.235 ;
        RECT 69.895 193.045 70.060 193.065 ;
        RECT 70.355 193.045 70.525 193.235 ;
        RECT 72.250 193.095 72.370 193.205 ;
        RECT 74.035 193.045 74.205 193.235 ;
        RECT 78.635 193.065 78.805 193.255 ;
        RECT 80.015 193.045 80.185 193.235 ;
        RECT 80.475 193.045 80.645 193.235 ;
        RECT 81.395 193.065 81.565 193.255 ;
        RECT 83.235 193.045 83.405 193.235 ;
        RECT 83.695 193.045 83.865 193.235 ;
        RECT 86.915 193.065 87.085 193.255 ;
        RECT 87.890 193.095 88.010 193.205 ;
        RECT 89.675 193.065 89.845 193.255 ;
        RECT 90.135 193.065 90.305 193.255 ;
        RECT 93.815 193.045 93.985 193.255 ;
        RECT 94.275 193.045 94.445 193.235 ;
        RECT 97.955 193.045 98.125 193.235 ;
        RECT 99.795 193.090 99.955 193.200 ;
        RECT 103.015 193.065 103.185 193.255 ;
        RECT 103.530 193.095 103.650 193.205 ;
        RECT 106.235 193.065 106.405 193.255 ;
        RECT 109.455 193.045 109.625 193.235 ;
        RECT 109.970 193.095 110.090 193.205 ;
        RECT 111.755 193.045 111.925 193.255 ;
        RECT 113.135 193.045 113.305 193.255 ;
        RECT 65.580 193.015 66.525 193.045 ;
        RECT 63.455 192.815 66.525 193.015 ;
        RECT 61.015 192.135 61.935 192.365 ;
        RECT 63.315 192.335 66.525 192.815 ;
        RECT 63.315 192.135 64.245 192.335 ;
        RECT 65.580 192.135 66.525 192.335 ;
        RECT 66.535 192.235 67.905 193.045 ;
        RECT 68.225 192.365 70.060 193.045 ;
        RECT 70.215 192.365 72.045 193.045 ;
        RECT 68.225 192.135 69.155 192.365 ;
        RECT 72.515 192.235 74.345 193.045 ;
        RECT 74.365 192.175 74.795 192.960 ;
        RECT 74.815 192.235 80.325 193.045 ;
        RECT 80.335 192.265 81.705 193.045 ;
        RECT 81.715 192.235 83.545 193.045 ;
        RECT 83.565 192.135 84.915 193.045 ;
        RECT 84.935 192.365 94.125 193.045 ;
        RECT 94.245 192.365 97.710 193.045 ;
        RECT 84.935 192.135 85.855 192.365 ;
        RECT 88.685 192.145 89.615 192.365 ;
        RECT 96.790 192.135 97.710 192.365 ;
        RECT 97.825 192.135 99.175 193.045 ;
        RECT 100.125 192.175 100.555 192.960 ;
        RECT 100.575 192.365 109.765 193.045 ;
        RECT 100.575 192.135 101.495 192.365 ;
        RECT 104.325 192.145 105.255 192.365 ;
        RECT 110.235 192.235 112.065 193.045 ;
        RECT 112.075 192.235 113.445 193.045 ;
      LAYER nwell ;
        RECT 11.140 189.015 113.640 191.845 ;
      LAYER pwell ;
        RECT 11.335 187.815 12.705 188.625 ;
        RECT 13.175 187.815 16.845 188.625 ;
        RECT 16.855 187.815 22.365 188.625 ;
        RECT 26.885 188.495 27.815 188.715 ;
        RECT 30.645 188.495 31.565 188.725 ;
        RECT 34.775 188.495 35.705 188.725 ;
        RECT 22.375 187.815 31.565 188.495 ;
        RECT 31.805 187.815 35.705 188.495 ;
        RECT 35.725 187.900 36.155 188.685 ;
        RECT 36.175 187.815 38.005 188.625 ;
        RECT 38.025 187.815 39.375 188.725 ;
        RECT 42.050 188.495 42.970 188.725 ;
        RECT 39.505 187.815 42.970 188.495 ;
        RECT 43.075 187.815 44.445 188.595 ;
        RECT 44.455 188.495 45.375 188.725 ;
        RECT 48.205 188.495 49.135 188.715 ;
        RECT 44.455 187.815 53.645 188.495 ;
        RECT 54.115 187.815 57.225 188.725 ;
        RECT 57.430 188.495 58.350 188.725 ;
        RECT 57.430 187.815 60.895 188.495 ;
        RECT 61.485 187.900 61.915 188.685 ;
        RECT 61.935 188.525 62.865 188.725 ;
        RECT 64.200 188.525 65.145 188.725 ;
        RECT 61.935 188.045 65.145 188.525 ;
        RECT 62.075 187.845 65.145 188.045 ;
        RECT 11.475 187.605 11.645 187.815 ;
        RECT 12.910 187.655 13.030 187.765 ;
        RECT 13.315 187.650 13.475 187.760 ;
        RECT 16.535 187.625 16.705 187.815 ;
        RECT 16.995 187.605 17.165 187.795 ;
        RECT 22.055 187.625 22.225 187.815 ;
        RECT 22.515 187.605 22.685 187.815 ;
        RECT 23.490 187.655 23.610 187.765 ;
        RECT 24.815 187.605 24.985 187.795 ;
        RECT 25.275 187.605 25.445 187.795 ;
        RECT 35.120 187.625 35.290 187.815 ;
        RECT 37.695 187.625 37.865 187.815 ;
        RECT 38.155 187.605 38.325 187.795 ;
        RECT 39.075 187.625 39.245 187.815 ;
        RECT 39.535 187.605 39.705 187.815 ;
        RECT 40.050 187.655 40.170 187.765 ;
        RECT 43.215 187.625 43.385 187.815 ;
        RECT 43.860 187.605 44.030 187.795 ;
        RECT 48.000 187.605 48.170 187.795 ;
        RECT 49.655 187.650 49.815 187.760 ;
        RECT 50.115 187.605 50.285 187.795 ;
        RECT 52.415 187.605 52.585 187.795 ;
        RECT 52.875 187.605 53.045 187.795 ;
        RECT 53.335 187.625 53.505 187.815 ;
        RECT 53.850 187.655 53.970 187.765 ;
        RECT 57.015 187.625 57.185 187.815 ;
        RECT 60.695 187.625 60.865 187.815 ;
        RECT 61.210 187.655 61.330 187.765 ;
        RECT 62.075 187.625 62.245 187.845 ;
        RECT 64.200 187.815 65.145 187.845 ;
        RECT 65.155 187.815 67.445 188.725 ;
        RECT 68.825 188.495 69.745 188.725 ;
        RECT 67.455 187.815 69.745 188.495 ;
        RECT 69.755 187.815 75.265 188.625 ;
        RECT 75.645 188.615 76.565 188.725 ;
        RECT 75.645 188.495 77.980 188.615 ;
        RECT 82.645 188.495 83.565 188.715 ;
        RECT 75.645 187.815 84.925 188.495 ;
        RECT 85.395 187.815 87.225 188.625 ;
        RECT 87.245 187.900 87.675 188.685 ;
        RECT 90.895 188.495 91.825 188.725 ;
        RECT 87.925 187.815 91.825 188.495 ;
        RECT 91.835 187.815 93.665 188.625 ;
        RECT 93.685 187.815 95.035 188.725 ;
        RECT 98.255 188.495 99.185 188.725 ;
        RECT 102.395 188.495 103.325 188.725 ;
        RECT 95.285 187.815 99.185 188.495 ;
        RECT 99.425 187.815 103.325 188.495 ;
        RECT 103.795 187.815 105.165 188.595 ;
        RECT 105.175 187.815 106.545 188.625 ;
        RECT 106.555 187.815 112.065 188.625 ;
        RECT 112.075 187.815 113.445 188.625 ;
        RECT 65.300 187.625 65.470 187.815 ;
        RECT 67.135 187.605 67.305 187.795 ;
        RECT 67.595 187.625 67.765 187.815 ;
        RECT 72.655 187.605 72.825 187.795 ;
        RECT 73.115 187.605 73.285 187.795 ;
        RECT 74.955 187.625 75.125 187.815 ;
        RECT 75.415 187.650 75.575 187.760 ;
        RECT 79.280 187.605 79.450 187.795 ;
        RECT 80.935 187.605 81.105 187.795 ;
        RECT 81.450 187.655 81.570 187.765 ;
        RECT 84.615 187.625 84.785 187.815 ;
        RECT 85.130 187.655 85.250 187.765 ;
        RECT 86.915 187.605 87.085 187.815 ;
        RECT 87.375 187.605 87.545 187.795 ;
        RECT 91.240 187.625 91.410 187.815 ;
        RECT 91.515 187.650 91.675 187.760 ;
        RECT 91.975 187.605 92.145 187.795 ;
        RECT 93.355 187.625 93.525 187.815 ;
        RECT 93.815 187.625 93.985 187.815 ;
        RECT 96.575 187.605 96.745 187.795 ;
        RECT 98.415 187.605 98.585 187.795 ;
        RECT 98.600 187.625 98.770 187.815 ;
        RECT 98.875 187.605 99.045 187.795 ;
        RECT 100.715 187.605 100.885 187.795 ;
        RECT 102.740 187.625 102.910 187.815 ;
        RECT 103.530 187.655 103.650 187.765 ;
        RECT 103.935 187.625 104.105 187.815 ;
        RECT 106.235 187.625 106.405 187.815 ;
        RECT 107.615 187.605 107.785 187.795 ;
        RECT 108.130 187.655 108.250 187.765 ;
        RECT 111.755 187.605 111.925 187.815 ;
        RECT 113.135 187.605 113.305 187.815 ;
        RECT 11.335 186.795 12.705 187.605 ;
        RECT 13.635 186.795 17.305 187.605 ;
        RECT 17.315 186.795 22.825 187.605 ;
        RECT 22.845 186.735 23.275 187.520 ;
        RECT 23.765 186.695 25.115 187.605 ;
        RECT 25.245 186.925 28.710 187.605 ;
        RECT 27.790 186.695 28.710 186.925 ;
        RECT 29.185 186.925 38.465 187.605 ;
        RECT 29.185 186.805 31.520 186.925 ;
        RECT 29.185 186.695 30.105 186.805 ;
        RECT 36.185 186.705 37.105 186.925 ;
        RECT 38.475 186.825 39.845 187.605 ;
        RECT 40.545 186.925 44.445 187.605 ;
        RECT 44.685 186.925 48.585 187.605 ;
        RECT 43.515 186.695 44.445 186.925 ;
        RECT 47.655 186.695 48.585 186.925 ;
        RECT 48.605 186.735 49.035 187.520 ;
        RECT 49.975 186.825 51.345 187.605 ;
        RECT 51.355 186.795 52.725 187.605 ;
        RECT 52.735 186.925 61.925 187.605 ;
        RECT 57.245 186.705 58.175 186.925 ;
        RECT 61.005 186.695 61.925 186.925 ;
        RECT 61.935 186.795 67.445 187.605 ;
        RECT 67.455 186.795 72.965 187.605 ;
        RECT 72.985 186.695 74.335 187.605 ;
        RECT 74.365 186.735 74.795 187.520 ;
        RECT 75.965 186.925 79.865 187.605 ;
        RECT 78.935 186.695 79.865 186.925 ;
        RECT 79.885 186.695 81.235 187.605 ;
        RECT 81.715 186.795 87.225 187.605 ;
        RECT 87.345 186.925 90.810 187.605 ;
        RECT 89.890 186.695 90.810 186.925 ;
        RECT 91.835 186.825 93.205 187.605 ;
        RECT 93.310 186.925 96.775 187.605 ;
        RECT 93.310 186.695 94.230 186.925 ;
        RECT 96.895 186.795 98.725 187.605 ;
        RECT 98.745 186.695 100.095 187.605 ;
        RECT 100.125 186.735 100.555 187.520 ;
        RECT 100.685 186.925 104.150 187.605 ;
        RECT 103.230 186.695 104.150 186.925 ;
        RECT 104.350 186.925 107.815 187.605 ;
        RECT 104.350 186.695 105.270 186.925 ;
        RECT 108.395 186.795 112.065 187.605 ;
        RECT 112.075 186.795 113.445 187.605 ;
      LAYER nwell ;
        RECT 11.140 183.575 113.640 186.405 ;
      LAYER pwell ;
        RECT 11.335 182.375 12.705 183.185 ;
        RECT 13.635 182.375 17.305 183.185 ;
        RECT 17.315 182.375 22.825 183.185 ;
        RECT 22.835 182.375 24.205 183.155 ;
        RECT 24.225 182.375 25.575 183.285 ;
        RECT 26.515 183.055 27.445 183.285 ;
        RECT 33.310 183.055 34.230 183.285 ;
        RECT 26.515 182.375 30.415 183.055 ;
        RECT 30.765 182.375 34.230 183.055 ;
        RECT 34.345 182.375 35.695 183.285 ;
        RECT 35.725 182.460 36.155 183.245 ;
        RECT 36.185 182.375 37.535 183.285 ;
        RECT 37.555 182.375 39.385 183.185 ;
        RECT 39.395 182.375 40.765 183.155 ;
        RECT 41.235 182.375 43.065 183.185 ;
        RECT 43.085 182.375 44.435 183.285 ;
        RECT 44.465 182.375 45.815 183.285 ;
        RECT 48.490 183.055 49.410 183.285 ;
        RECT 45.945 182.375 49.410 183.055 ;
        RECT 50.435 182.375 55.945 183.185 ;
        RECT 55.955 182.375 61.465 183.185 ;
        RECT 61.485 182.460 61.915 183.245 ;
        RECT 63.095 182.605 65.850 183.285 ;
        RECT 63.095 182.375 65.365 182.605 ;
        RECT 66.535 182.375 72.045 183.185 ;
        RECT 72.425 183.175 73.345 183.285 ;
        RECT 72.425 183.055 74.760 183.175 ;
        RECT 79.425 183.055 80.345 183.275 ;
        RECT 72.425 182.375 81.705 183.055 ;
        RECT 81.715 182.375 83.085 183.155 ;
        RECT 83.095 182.375 84.465 183.185 ;
        RECT 84.485 182.375 85.835 183.285 ;
        RECT 85.865 182.375 87.215 183.285 ;
        RECT 87.245 182.460 87.675 183.245 ;
        RECT 87.695 183.055 88.615 183.285 ;
        RECT 91.445 183.055 92.375 183.275 ;
        RECT 99.550 183.055 100.470 183.285 ;
        RECT 87.695 182.375 96.885 183.055 ;
        RECT 97.005 182.375 100.470 183.055 ;
        RECT 100.585 182.375 101.935 183.285 ;
        RECT 101.955 183.055 102.875 183.285 ;
        RECT 105.705 183.055 106.635 183.275 ;
        RECT 101.955 182.375 111.145 183.055 ;
        RECT 112.075 182.375 113.445 183.185 ;
        RECT 11.475 182.165 11.645 182.375 ;
        RECT 13.315 182.210 13.475 182.330 ;
        RECT 16.995 182.185 17.165 182.375 ;
        RECT 18.835 182.165 19.005 182.355 ;
        RECT 19.295 182.165 19.465 182.355 ;
        RECT 22.515 182.185 22.685 182.375 ;
        RECT 22.975 182.185 23.145 182.375 ;
        RECT 23.895 182.210 24.055 182.320 ;
        RECT 24.355 182.165 24.525 182.375 ;
        RECT 26.195 182.220 26.355 182.330 ;
        RECT 26.930 182.185 27.100 182.375 ;
        RECT 30.795 182.185 30.965 182.375 ;
        RECT 31.250 182.165 31.420 182.355 ;
        RECT 31.715 182.165 31.885 182.355 ;
        RECT 35.395 182.185 35.565 182.375 ;
        RECT 37.235 182.185 37.405 182.375 ;
        RECT 38.800 182.165 38.970 182.355 ;
        RECT 39.075 182.185 39.245 182.375 ;
        RECT 40.455 182.185 40.625 182.375 ;
        RECT 40.970 182.215 41.090 182.325 ;
        RECT 42.755 182.185 42.925 182.375 ;
        RECT 44.135 182.185 44.305 182.375 ;
        RECT 44.595 182.185 44.765 182.375 ;
        RECT 45.975 182.185 46.145 182.375 ;
        RECT 48.275 182.165 48.445 182.355 ;
        RECT 49.250 182.215 49.370 182.325 ;
        RECT 50.115 182.220 50.275 182.330 ;
        RECT 51.035 182.165 51.205 182.355 ;
        RECT 55.635 182.185 55.805 182.375 ;
        RECT 56.555 182.165 56.725 182.355 ;
        RECT 57.015 182.185 57.185 182.355 ;
        RECT 61.155 182.185 61.325 182.375 ;
        RECT 63.095 182.355 63.165 182.375 ;
        RECT 62.535 182.220 62.695 182.330 ;
        RECT 62.995 182.185 63.165 182.355 ;
        RECT 57.115 182.165 57.185 182.185 ;
        RECT 62.995 182.165 63.065 182.185 ;
        RECT 63.455 182.165 63.625 182.355 ;
        RECT 66.270 182.215 66.390 182.325 ;
        RECT 68.110 182.215 68.230 182.325 ;
        RECT 69.435 182.165 69.605 182.355 ;
        RECT 69.950 182.215 70.070 182.325 ;
        RECT 71.735 182.185 71.905 182.375 ;
        RECT 73.760 182.165 73.930 182.355 ;
        RECT 75.010 182.215 75.130 182.325 ;
        RECT 78.820 182.165 78.990 182.355 ;
        RECT 80.935 182.165 81.105 182.355 ;
        RECT 81.395 182.185 81.565 182.375 ;
        RECT 82.775 182.185 82.945 182.375 ;
        RECT 84.155 182.185 84.325 182.375 ;
        RECT 85.535 182.185 85.705 182.375 ;
        RECT 85.995 182.185 86.165 182.375 ;
        RECT 90.135 182.165 90.305 182.355 ;
        RECT 90.650 182.215 90.770 182.325 ;
        RECT 91.330 182.165 91.500 182.355 ;
        RECT 95.655 182.210 95.815 182.320 ;
        RECT 96.575 182.185 96.745 182.375 ;
        RECT 97.035 182.185 97.205 182.375 ;
        RECT 99.520 182.165 99.690 182.355 ;
        RECT 100.715 182.185 100.885 182.375 ;
        RECT 109.455 182.165 109.625 182.355 ;
        RECT 109.970 182.215 110.090 182.325 ;
        RECT 110.835 182.185 111.005 182.375 ;
        RECT 111.755 182.165 111.925 182.355 ;
        RECT 113.135 182.165 113.305 182.375 ;
        RECT 11.335 181.355 12.705 182.165 ;
        RECT 13.635 181.355 19.145 182.165 ;
        RECT 19.265 181.485 22.730 182.165 ;
        RECT 21.810 181.255 22.730 181.485 ;
        RECT 22.845 181.295 23.275 182.080 ;
        RECT 24.325 181.485 27.790 182.165 ;
        RECT 26.870 181.255 27.790 181.485 ;
        RECT 28.090 181.255 31.565 182.165 ;
        RECT 31.685 181.485 35.150 182.165 ;
        RECT 35.485 181.485 39.385 182.165 ;
        RECT 34.230 181.255 35.150 181.485 ;
        RECT 38.455 181.255 39.385 181.485 ;
        RECT 39.395 181.485 48.585 182.165 ;
        RECT 39.395 181.255 40.315 181.485 ;
        RECT 43.145 181.265 44.075 181.485 ;
        RECT 48.605 181.295 49.035 182.080 ;
        RECT 49.515 181.355 51.345 182.165 ;
        RECT 51.355 181.355 56.865 182.165 ;
        RECT 57.115 181.935 59.385 182.165 ;
        RECT 60.795 181.935 63.065 182.165 ;
        RECT 57.115 181.255 59.870 181.935 ;
        RECT 60.310 181.255 63.065 181.935 ;
        RECT 63.315 181.935 64.885 182.165 ;
        RECT 66.975 182.125 67.895 182.165 ;
        RECT 66.975 181.935 67.905 182.125 ;
        RECT 63.315 181.575 67.905 181.935 ;
        RECT 63.315 181.485 67.895 181.575 ;
        RECT 64.895 181.255 67.895 181.485 ;
        RECT 68.385 181.255 69.735 182.165 ;
        RECT 70.445 181.485 74.345 182.165 ;
        RECT 73.415 181.255 74.345 181.485 ;
        RECT 74.365 181.295 74.795 182.080 ;
        RECT 75.505 181.485 79.405 182.165 ;
        RECT 78.475 181.255 79.405 181.485 ;
        RECT 79.415 181.355 81.245 182.165 ;
        RECT 81.255 181.485 90.445 182.165 ;
        RECT 90.915 181.485 94.815 182.165 ;
        RECT 96.205 181.485 100.105 182.165 ;
        RECT 81.255 181.255 82.175 181.485 ;
        RECT 85.005 181.265 85.935 181.485 ;
        RECT 90.915 181.255 91.845 181.485 ;
        RECT 99.175 181.255 100.105 181.485 ;
        RECT 100.125 181.295 100.555 182.080 ;
        RECT 100.575 181.485 109.765 182.165 ;
        RECT 100.575 181.255 101.495 181.485 ;
        RECT 104.325 181.265 105.255 181.485 ;
        RECT 110.235 181.355 112.065 182.165 ;
        RECT 112.075 181.355 113.445 182.165 ;
      LAYER nwell ;
        RECT 11.140 178.135 113.640 180.965 ;
      LAYER pwell ;
        RECT 11.335 176.935 12.705 177.745 ;
        RECT 13.175 176.935 15.005 177.745 ;
        RECT 15.015 176.935 20.525 177.745 ;
        RECT 25.045 177.615 25.975 177.835 ;
        RECT 28.805 177.615 29.725 177.845 ;
        RECT 20.535 176.935 29.725 177.615 ;
        RECT 30.195 176.935 32.025 177.745 ;
        RECT 32.230 176.935 35.705 177.845 ;
        RECT 35.725 177.020 36.155 177.805 ;
        RECT 36.635 176.935 39.385 177.745 ;
        RECT 39.395 176.935 42.870 177.845 ;
        RECT 45.730 177.615 46.650 177.845 ;
        RECT 43.185 176.935 46.650 177.615 ;
        RECT 46.755 176.935 48.125 177.715 ;
        RECT 48.135 176.935 50.885 177.745 ;
        RECT 50.895 176.935 52.265 177.715 ;
        RECT 52.285 176.935 55.025 177.615 ;
        RECT 55.495 176.935 57.325 177.745 ;
        RECT 57.335 176.935 59.945 177.845 ;
        RECT 60.095 176.935 61.465 177.745 ;
        RECT 61.485 177.020 61.915 177.805 ;
        RECT 61.945 176.935 63.295 177.845 ;
        RECT 63.555 177.165 66.310 177.845 ;
        RECT 72.410 177.615 73.330 177.845 ;
        RECT 63.555 176.935 65.825 177.165 ;
        RECT 66.995 176.935 69.735 177.615 ;
        RECT 69.865 176.935 73.330 177.615 ;
        RECT 73.435 177.615 74.355 177.845 ;
        RECT 77.185 177.615 78.115 177.835 ;
        RECT 83.095 177.615 84.025 177.845 ;
        RECT 73.435 176.935 82.625 177.615 ;
        RECT 83.095 176.935 86.995 177.615 ;
        RECT 87.245 177.020 87.675 177.805 ;
        RECT 90.350 177.615 91.270 177.845 ;
        RECT 87.805 176.935 91.270 177.615 ;
        RECT 91.375 176.935 92.745 177.715 ;
        RECT 92.755 176.935 96.230 177.845 ;
        RECT 96.895 176.935 99.645 177.745 ;
        RECT 102.855 177.615 103.785 177.845 ;
        RECT 99.885 176.935 103.785 177.615 ;
        RECT 104.255 176.935 105.625 177.715 ;
        RECT 106.555 176.935 107.925 177.715 ;
        RECT 108.395 176.935 112.065 177.745 ;
        RECT 112.075 176.935 113.445 177.745 ;
        RECT 11.475 176.725 11.645 176.935 ;
        RECT 12.910 176.775 13.030 176.885 ;
        RECT 13.315 176.770 13.475 176.880 ;
        RECT 14.695 176.745 14.865 176.935 ;
        RECT 16.995 176.725 17.165 176.915 ;
        RECT 20.215 176.745 20.385 176.935 ;
        RECT 20.675 176.745 20.845 176.935 ;
        RECT 22.515 176.725 22.685 176.915 ;
        RECT 23.490 176.775 23.610 176.885 ;
        RECT 24.815 176.725 24.985 176.915 ;
        RECT 25.275 176.725 25.445 176.915 ;
        RECT 26.930 176.725 27.100 176.915 ;
        RECT 29.930 176.775 30.050 176.885 ;
        RECT 31.715 176.745 31.885 176.935 ;
        RECT 34.200 176.725 34.370 176.915 ;
        RECT 34.990 176.775 35.110 176.885 ;
        RECT 35.390 176.745 35.560 176.935 ;
        RECT 36.370 176.775 36.490 176.885 ;
        RECT 38.610 176.725 38.780 176.915 ;
        RECT 39.075 176.725 39.245 176.935 ;
        RECT 39.540 176.745 39.710 176.935 ;
        RECT 43.215 176.745 43.385 176.935 ;
        RECT 46.160 176.725 46.330 176.915 ;
        RECT 46.950 176.775 47.070 176.885 ;
        RECT 47.355 176.725 47.525 176.915 ;
        RECT 47.815 176.745 47.985 176.935 ;
        RECT 50.575 176.745 50.745 176.935 ;
        RECT 51.035 176.745 51.205 176.935 ;
        RECT 54.715 176.745 54.885 176.935 ;
        RECT 55.230 176.775 55.350 176.885 ;
        RECT 57.015 176.745 57.185 176.935 ;
        RECT 57.480 176.745 57.650 176.935 ;
        RECT 57.935 176.725 58.105 176.915 ;
        RECT 58.450 176.775 58.570 176.885 ;
        RECT 58.855 176.725 59.025 176.915 ;
        RECT 61.155 176.745 61.325 176.935 ;
        RECT 62.075 176.725 62.245 176.935 ;
        RECT 63.555 176.915 63.625 176.935 ;
        RECT 62.535 176.725 62.705 176.915 ;
        RECT 63.455 176.745 63.625 176.915 ;
        RECT 64.375 176.725 64.545 176.915 ;
        RECT 66.730 176.775 66.850 176.885 ;
        RECT 67.135 176.725 67.305 176.935 ;
        RECT 69.895 176.725 70.065 176.935 ;
        RECT 70.360 176.725 70.530 176.915 ;
        RECT 74.090 176.775 74.210 176.885 ;
        RECT 75.415 176.770 75.575 176.880 ;
        RECT 75.875 176.725 76.045 176.915 ;
        RECT 79.555 176.725 79.725 176.915 ;
        RECT 80.935 176.725 81.105 176.915 ;
        RECT 82.315 176.745 82.485 176.935 ;
        RECT 82.830 176.775 82.950 176.885 ;
        RECT 83.510 176.745 83.680 176.935 ;
        RECT 84.615 176.725 84.785 176.915 ;
        RECT 87.835 176.745 88.005 176.935 ;
        RECT 92.435 176.915 92.605 176.935 ;
        RECT 88.300 176.725 88.470 176.915 ;
        RECT 92.030 176.775 92.150 176.885 ;
        RECT 92.435 176.745 92.610 176.915 ;
        RECT 92.900 176.745 93.070 176.935 ;
        RECT 99.335 176.915 99.505 176.935 ;
        RECT 96.630 176.775 96.750 176.885 ;
        RECT 99.330 176.745 99.505 176.915 ;
        RECT 99.850 176.775 99.970 176.885 ;
        RECT 101.175 176.770 101.335 176.880 ;
        RECT 103.200 176.745 103.370 176.935 ;
        RECT 103.990 176.775 104.110 176.885 ;
        RECT 104.395 176.745 104.565 176.935 ;
        RECT 106.235 176.780 106.395 176.890 ;
        RECT 92.440 176.725 92.610 176.745 ;
        RECT 99.330 176.725 99.500 176.745 ;
        RECT 106.695 176.725 106.865 176.935 ;
        RECT 107.155 176.725 107.325 176.915 ;
        RECT 108.130 176.775 108.250 176.885 ;
        RECT 111.755 176.725 111.925 176.935 ;
        RECT 113.135 176.725 113.305 176.935 ;
        RECT 11.335 175.915 12.705 176.725 ;
        RECT 13.635 175.915 17.305 176.725 ;
        RECT 17.315 175.915 22.825 176.725 ;
        RECT 22.845 175.855 23.275 176.640 ;
        RECT 23.755 175.945 25.125 176.725 ;
        RECT 25.145 175.815 26.495 176.725 ;
        RECT 26.515 176.045 30.415 176.725 ;
        RECT 30.885 176.045 34.785 176.725 ;
        RECT 26.515 175.815 27.445 176.045 ;
        RECT 33.855 175.815 34.785 176.045 ;
        RECT 35.450 175.815 38.925 176.725 ;
        RECT 39.045 176.045 42.510 176.725 ;
        RECT 42.845 176.045 46.745 176.725 ;
        RECT 41.590 175.815 42.510 176.045 ;
        RECT 45.815 175.815 46.745 176.045 ;
        RECT 47.225 175.815 48.575 176.725 ;
        RECT 48.605 175.855 49.035 176.640 ;
        RECT 49.055 176.045 58.245 176.725 ;
        RECT 58.715 176.045 60.545 176.725 ;
        RECT 49.055 175.815 49.975 176.045 ;
        RECT 52.805 175.825 53.735 176.045 ;
        RECT 59.200 175.815 60.545 176.045 ;
        RECT 60.555 176.045 62.385 176.725 ;
        RECT 62.395 176.045 64.225 176.725 ;
        RECT 60.555 175.815 61.900 176.045 ;
        RECT 62.880 175.815 64.225 176.045 ;
        RECT 64.235 175.815 66.955 176.725 ;
        RECT 66.995 176.045 68.825 176.725 ;
        RECT 67.480 175.815 68.825 176.045 ;
        RECT 68.835 175.915 70.205 176.725 ;
        RECT 70.215 175.815 73.690 176.725 ;
        RECT 74.365 175.855 74.795 176.640 ;
        RECT 75.845 176.045 79.310 176.725 ;
        RECT 78.390 175.815 79.310 176.045 ;
        RECT 79.415 175.945 80.785 176.725 ;
        RECT 80.905 176.045 84.370 176.725 ;
        RECT 84.585 176.045 88.050 176.725 ;
        RECT 83.450 175.815 84.370 176.045 ;
        RECT 87.130 175.815 88.050 176.045 ;
        RECT 88.155 175.815 91.630 176.725 ;
        RECT 92.295 175.815 95.770 176.725 ;
        RECT 96.170 175.815 99.645 176.725 ;
        RECT 100.125 175.855 100.555 176.640 ;
        RECT 101.495 175.915 107.005 176.725 ;
        RECT 107.015 175.945 108.385 176.725 ;
        RECT 108.395 175.915 112.065 176.725 ;
        RECT 112.075 175.915 113.445 176.725 ;
      LAYER nwell ;
        RECT 11.140 172.695 113.640 175.525 ;
      LAYER pwell ;
        RECT 11.335 171.495 12.705 172.305 ;
        RECT 13.175 171.495 16.845 172.305 ;
        RECT 16.855 171.495 22.365 172.305 ;
        RECT 25.030 172.175 25.950 172.405 ;
        RECT 22.485 171.495 25.950 172.175 ;
        RECT 26.055 172.175 26.975 172.405 ;
        RECT 29.805 172.175 30.735 172.395 ;
        RECT 26.055 171.495 35.245 172.175 ;
        RECT 35.725 171.580 36.155 172.365 ;
        RECT 36.175 171.495 37.545 172.275 ;
        RECT 38.670 171.495 42.145 172.405 ;
        RECT 45.355 172.175 46.285 172.405 ;
        RECT 49.495 172.175 50.425 172.405 ;
        RECT 42.385 171.495 46.285 172.175 ;
        RECT 46.525 171.495 50.425 172.175 ;
        RECT 50.435 172.175 51.355 172.405 ;
        RECT 54.185 172.175 55.115 172.395 ;
        RECT 50.435 171.495 59.625 172.175 ;
        RECT 59.635 171.495 61.465 172.305 ;
        RECT 61.485 171.580 61.915 172.365 ;
        RECT 61.935 171.495 63.305 172.305 ;
        RECT 63.315 172.175 64.660 172.405 ;
        RECT 63.315 171.495 65.145 172.175 ;
        RECT 65.810 171.495 69.285 172.405 ;
        RECT 69.295 171.495 72.770 172.405 ;
        RECT 73.445 171.495 74.795 172.405 ;
        RECT 74.815 171.495 77.425 172.405 ;
        RECT 78.035 172.175 78.955 172.405 ;
        RECT 81.785 172.175 82.715 172.395 ;
        RECT 78.035 171.495 87.225 172.175 ;
        RECT 87.245 171.580 87.675 172.365 ;
        RECT 87.890 171.495 91.365 172.405 ;
        RECT 91.570 171.495 95.045 172.405 ;
        RECT 99.175 172.175 100.105 172.405 ;
        RECT 96.205 171.495 100.105 172.175 ;
        RECT 101.045 171.495 102.395 172.405 ;
        RECT 102.415 172.175 103.335 172.405 ;
        RECT 106.165 172.175 107.095 172.395 ;
        RECT 102.415 171.495 111.605 172.175 ;
        RECT 112.075 171.495 113.445 172.305 ;
        RECT 11.475 171.285 11.645 171.495 ;
        RECT 12.910 171.335 13.030 171.445 ;
        RECT 13.315 171.330 13.475 171.440 ;
        RECT 16.535 171.305 16.705 171.495 ;
        RECT 16.995 171.285 17.165 171.475 ;
        RECT 22.055 171.305 22.225 171.495 ;
        RECT 22.515 171.285 22.685 171.495 ;
        RECT 23.490 171.335 23.610 171.445 ;
        RECT 24.815 171.285 24.985 171.475 ;
        RECT 26.195 171.285 26.365 171.475 ;
        RECT 26.660 171.285 26.830 171.475 ;
        RECT 30.340 171.285 30.510 171.475 ;
        RECT 34.935 171.305 35.105 171.495 ;
        RECT 35.450 171.335 35.570 171.445 ;
        RECT 37.235 171.285 37.405 171.495 ;
        RECT 37.700 171.285 37.870 171.475 ;
        RECT 38.155 171.340 38.315 171.450 ;
        RECT 41.380 171.285 41.550 171.475 ;
        RECT 41.830 171.305 42.000 171.495 ;
        RECT 45.060 171.285 45.230 171.475 ;
        RECT 45.700 171.305 45.870 171.495 ;
        RECT 49.195 171.285 49.365 171.475 ;
        RECT 49.840 171.305 50.010 171.495 ;
        RECT 53.335 171.330 53.495 171.440 ;
        RECT 54.715 171.285 54.885 171.475 ;
        RECT 55.175 171.285 55.345 171.475 ;
        RECT 57.015 171.330 57.175 171.440 ;
        RECT 59.315 171.305 59.485 171.495 ;
        RECT 61.155 171.305 61.325 171.495 ;
        RECT 62.535 171.285 62.705 171.475 ;
        RECT 62.995 171.305 63.165 171.495 ;
        RECT 64.375 171.285 64.545 171.475 ;
        RECT 64.835 171.305 65.005 171.495 ;
        RECT 65.350 171.335 65.470 171.445 ;
        RECT 68.970 171.305 69.140 171.495 ;
        RECT 69.440 171.305 69.610 171.495 ;
        RECT 69.895 171.285 70.065 171.475 ;
        RECT 70.360 171.285 70.530 171.475 ;
        RECT 73.170 171.335 73.290 171.445 ;
        RECT 73.575 171.305 73.745 171.495 ;
        RECT 74.090 171.335 74.210 171.445 ;
        RECT 74.960 171.305 75.130 171.495 ;
        RECT 75.415 171.330 75.575 171.440 ;
        RECT 75.875 171.285 76.045 171.475 ;
        RECT 77.770 171.335 77.890 171.445 ;
        RECT 86.455 171.285 86.625 171.475 ;
        RECT 86.915 171.285 87.085 171.495 ;
        RECT 91.050 171.305 91.220 171.495 ;
        RECT 94.730 171.305 94.900 171.495 ;
        RECT 95.655 171.340 95.815 171.450 ;
        RECT 97.035 171.285 97.205 171.475 ;
        RECT 98.415 171.285 98.585 171.475 ;
        RECT 99.520 171.305 99.690 171.495 ;
        RECT 99.795 171.285 99.965 171.475 ;
        RECT 100.715 171.340 100.875 171.450 ;
        RECT 101.175 171.305 101.345 171.495 ;
        RECT 101.635 171.285 101.805 171.475 ;
        RECT 102.150 171.335 102.270 171.445 ;
        RECT 111.295 171.285 111.465 171.495 ;
        RECT 111.810 171.335 111.930 171.445 ;
        RECT 113.135 171.285 113.305 171.495 ;
        RECT 11.335 170.475 12.705 171.285 ;
        RECT 13.635 170.475 17.305 171.285 ;
        RECT 17.315 170.475 22.825 171.285 ;
        RECT 22.845 170.415 23.275 171.200 ;
        RECT 23.765 170.375 25.115 171.285 ;
        RECT 25.135 170.475 26.505 171.285 ;
        RECT 26.515 170.375 29.990 171.285 ;
        RECT 30.195 170.375 33.670 171.285 ;
        RECT 33.875 170.475 37.545 171.285 ;
        RECT 37.555 170.375 41.030 171.285 ;
        RECT 41.235 170.375 44.710 171.285 ;
        RECT 44.915 170.375 48.390 171.285 ;
        RECT 48.605 170.415 49.035 171.200 ;
        RECT 49.165 170.605 52.630 171.285 ;
        RECT 51.710 170.375 52.630 170.605 ;
        RECT 53.665 170.375 55.015 171.285 ;
        RECT 55.035 170.505 56.405 171.285 ;
        RECT 57.335 170.475 62.845 171.285 ;
        RECT 62.855 170.605 64.685 171.285 ;
        RECT 62.855 170.375 64.200 170.605 ;
        RECT 64.695 170.475 70.205 171.285 ;
        RECT 70.215 170.375 73.690 171.285 ;
        RECT 74.365 170.415 74.795 171.200 ;
        RECT 75.735 170.605 84.840 171.285 ;
        RECT 84.935 170.475 86.765 171.285 ;
        RECT 86.785 170.375 88.135 171.285 ;
        RECT 88.155 170.605 97.345 171.285 ;
        RECT 88.155 170.375 89.075 170.605 ;
        RECT 91.905 170.385 92.835 170.605 ;
        RECT 97.355 170.505 98.725 171.285 ;
        RECT 98.735 170.475 100.105 171.285 ;
        RECT 100.125 170.415 100.555 171.200 ;
        RECT 100.585 170.375 101.935 171.285 ;
        RECT 102.415 170.605 111.605 171.285 ;
        RECT 102.415 170.375 103.335 170.605 ;
        RECT 106.165 170.385 107.095 170.605 ;
        RECT 112.075 170.475 113.445 171.285 ;
      LAYER nwell ;
        RECT 11.140 167.255 113.640 170.085 ;
      LAYER pwell ;
        RECT 11.335 166.055 12.705 166.865 ;
        RECT 13.175 166.055 14.545 166.835 ;
        RECT 14.565 166.055 15.915 166.965 ;
        RECT 16.865 166.055 18.215 166.965 ;
        RECT 19.595 166.735 20.515 166.955 ;
        RECT 26.595 166.855 27.515 166.965 ;
        RECT 25.180 166.735 27.515 166.855 ;
        RECT 18.235 166.055 27.515 166.735 ;
        RECT 28.355 166.055 32.025 166.865 ;
        RECT 32.035 166.055 35.510 166.965 ;
        RECT 35.725 166.140 36.155 166.925 ;
        RECT 36.645 166.055 39.385 166.735 ;
        RECT 39.630 166.055 44.445 166.735 ;
        RECT 44.455 166.055 45.825 166.865 ;
        RECT 45.930 166.735 46.850 166.965 ;
        RECT 45.930 166.055 49.395 166.735 ;
        RECT 49.975 166.055 51.805 166.865 ;
        RECT 51.955 166.055 54.565 166.965 ;
        RECT 54.715 166.055 57.325 166.965 ;
        RECT 57.795 166.055 59.625 166.865 ;
        RECT 59.635 166.735 60.980 166.965 ;
        RECT 59.635 166.055 61.465 166.735 ;
        RECT 61.485 166.140 61.915 166.925 ;
        RECT 62.855 166.055 65.575 166.965 ;
        RECT 65.615 166.055 69.285 166.865 ;
        RECT 69.295 166.055 70.665 166.835 ;
        RECT 72.035 166.735 72.955 166.955 ;
        RECT 79.035 166.855 79.955 166.965 ;
        RECT 77.620 166.735 79.955 166.855 ;
        RECT 70.675 166.055 79.955 166.735 ;
        RECT 80.570 166.055 85.385 166.735 ;
        RECT 85.395 166.055 86.765 166.835 ;
        RECT 87.245 166.140 87.675 166.925 ;
        RECT 97.355 166.735 98.275 166.965 ;
        RECT 101.105 166.735 102.035 166.955 ;
        RECT 87.695 166.055 96.800 166.735 ;
        RECT 97.355 166.055 106.545 166.735 ;
        RECT 106.565 166.055 107.915 166.965 ;
        RECT 107.935 166.055 109.765 166.735 ;
        RECT 109.775 166.055 111.145 166.835 ;
        RECT 112.075 166.055 113.445 166.865 ;
        RECT 11.475 165.845 11.645 166.055 ;
        RECT 12.855 166.005 13.025 166.035 ;
        RECT 12.855 165.895 13.030 166.005 ;
        RECT 12.855 165.845 13.025 165.895 ;
        RECT 13.315 165.865 13.485 166.055 ;
        RECT 14.695 165.865 14.865 166.055 ;
        RECT 16.535 165.900 16.695 166.010 ;
        RECT 16.995 165.865 17.165 166.055 ;
        RECT 18.375 165.865 18.545 166.055 ;
        RECT 22.570 165.895 22.690 166.005 ;
        RECT 23.490 165.895 23.610 166.005 ;
        RECT 24.815 165.845 24.985 166.035 ;
        RECT 25.550 165.845 25.720 166.035 ;
        RECT 28.090 165.895 28.210 166.005 ;
        RECT 29.415 165.845 29.585 166.035 ;
        RECT 31.715 165.865 31.885 166.055 ;
        RECT 32.180 165.865 32.350 166.055 ;
        RECT 36.370 165.895 36.490 166.005 ;
        RECT 39.075 165.865 39.245 166.055 ;
        RECT 44.135 165.865 44.305 166.055 ;
        RECT 45.515 165.865 45.685 166.055 ;
        RECT 47.355 165.845 47.525 166.035 ;
        RECT 48.275 165.890 48.435 166.000 ;
        RECT 49.195 165.865 49.365 166.055 ;
        RECT 49.710 165.895 49.830 166.005 ;
        RECT 50.115 165.845 50.285 166.035 ;
        RECT 51.495 165.865 51.665 166.055 ;
        RECT 52.870 165.845 53.040 166.035 ;
        RECT 54.250 165.865 54.420 166.055 ;
        RECT 55.635 165.845 55.805 166.035 ;
        RECT 56.150 165.895 56.270 166.005 ;
        RECT 57.010 165.865 57.180 166.055 ;
        RECT 57.530 165.895 57.650 166.005 ;
        RECT 59.315 165.865 59.485 166.055 ;
        RECT 61.155 165.865 61.325 166.055 ;
        RECT 61.615 165.845 61.785 166.035 ;
        RECT 62.075 165.845 62.245 166.035 ;
        RECT 62.535 165.900 62.695 166.010 ;
        RECT 62.995 165.865 63.165 166.055 ;
        RECT 68.975 165.865 69.145 166.055 ;
        RECT 69.435 165.865 69.605 166.055 ;
        RECT 70.815 165.865 70.985 166.055 ;
        RECT 74.035 165.845 74.205 166.035 ;
        RECT 75.415 165.890 75.575 166.000 ;
        RECT 75.875 165.845 76.045 166.035 ;
        RECT 85.075 165.865 85.245 166.055 ;
        RECT 86.455 165.865 86.625 166.055 ;
        RECT 86.970 165.895 87.090 166.005 ;
        RECT 87.835 165.865 88.005 166.055 ;
        RECT 96.110 165.845 96.280 166.035 ;
        RECT 96.575 165.845 96.745 166.035 ;
        RECT 97.090 165.895 97.210 166.005 ;
        RECT 104.120 165.845 104.290 166.035 ;
        RECT 104.855 165.845 105.025 166.035 ;
        RECT 106.235 165.865 106.405 166.055 ;
        RECT 106.695 165.865 106.865 166.055 ;
        RECT 109.455 165.845 109.625 166.055 ;
        RECT 109.970 165.895 110.090 166.005 ;
        RECT 110.835 165.865 111.005 166.055 ;
        RECT 111.755 165.845 111.925 166.035 ;
        RECT 113.135 165.845 113.305 166.055 ;
        RECT 11.335 165.035 12.705 165.845 ;
        RECT 12.715 165.165 21.995 165.845 ;
        RECT 14.075 164.945 14.995 165.165 ;
        RECT 19.660 165.045 21.995 165.165 ;
        RECT 21.075 164.935 21.995 165.045 ;
        RECT 22.845 164.975 23.275 165.760 ;
        RECT 23.755 165.065 25.125 165.845 ;
        RECT 25.135 165.165 29.035 165.845 ;
        RECT 29.275 165.165 38.380 165.845 ;
        RECT 38.475 165.165 47.665 165.845 ;
        RECT 25.135 164.935 26.065 165.165 ;
        RECT 38.475 164.935 39.395 165.165 ;
        RECT 42.225 164.945 43.155 165.165 ;
        RECT 48.605 164.975 49.035 165.760 ;
        RECT 49.055 165.035 50.425 165.845 ;
        RECT 50.575 164.935 53.185 165.845 ;
        RECT 53.205 165.165 55.945 165.845 ;
        RECT 56.415 165.035 61.925 165.845 ;
        RECT 61.935 165.165 64.675 165.845 ;
        RECT 65.065 165.165 74.345 165.845 ;
        RECT 65.065 165.045 67.400 165.165 ;
        RECT 65.065 164.935 65.985 165.045 ;
        RECT 72.065 164.945 72.985 165.165 ;
        RECT 74.365 164.975 74.795 165.760 ;
        RECT 75.735 165.165 85.015 165.845 ;
        RECT 77.095 164.945 78.015 165.165 ;
        RECT 82.680 165.045 85.015 165.165 ;
        RECT 84.095 164.935 85.015 165.045 ;
        RECT 85.415 164.935 96.425 165.845 ;
        RECT 96.545 165.165 100.010 165.845 ;
        RECT 99.090 164.935 100.010 165.165 ;
        RECT 100.125 164.975 100.555 165.760 ;
        RECT 100.805 165.165 104.705 165.845 ;
        RECT 104.825 165.165 108.290 165.845 ;
        RECT 103.775 164.935 104.705 165.165 ;
        RECT 107.370 164.935 108.290 165.165 ;
        RECT 108.395 165.065 109.765 165.845 ;
        RECT 110.235 165.035 112.065 165.845 ;
        RECT 112.075 165.035 113.445 165.845 ;
      LAYER nwell ;
        RECT 11.140 161.815 113.640 164.645 ;
      LAYER pwell ;
        RECT 11.335 160.615 12.705 161.425 ;
        RECT 12.725 160.615 14.075 161.525 ;
        RECT 17.315 161.295 18.245 161.525 ;
        RECT 22.375 161.295 23.305 161.525 ;
        RECT 31.025 161.295 31.955 161.515 ;
        RECT 34.785 161.295 35.705 161.525 ;
        RECT 14.475 160.615 16.900 161.295 ;
        RECT 17.315 160.615 21.215 161.295 ;
        RECT 22.375 160.615 26.275 161.295 ;
        RECT 26.515 160.615 35.705 161.295 ;
        RECT 35.725 160.700 36.155 161.485 ;
        RECT 39.375 161.295 40.305 161.525 ;
        RECT 36.405 160.615 40.305 161.295 ;
        RECT 40.315 161.295 41.235 161.525 ;
        RECT 44.065 161.295 44.995 161.515 ;
        RECT 40.315 160.615 49.505 161.295 ;
        RECT 49.515 160.615 50.885 161.395 ;
        RECT 50.895 160.615 56.405 161.425 ;
        RECT 56.425 160.615 57.775 161.525 ;
        RECT 57.795 161.295 59.140 161.525 ;
        RECT 59.635 161.295 60.980 161.525 ;
        RECT 57.795 160.615 59.625 161.295 ;
        RECT 59.635 160.615 61.465 161.295 ;
        RECT 61.485 160.700 61.915 161.485 ;
        RECT 62.420 161.295 63.765 161.525 ;
        RECT 64.260 161.295 65.605 161.525 ;
        RECT 61.935 160.615 63.765 161.295 ;
        RECT 63.775 160.615 65.605 161.295 ;
        RECT 66.075 160.615 69.745 161.425 ;
        RECT 69.755 160.615 71.125 161.395 ;
        RECT 71.135 161.295 72.065 161.525 ;
        RECT 71.135 160.615 75.035 161.295 ;
        RECT 75.285 160.615 76.635 161.525 ;
        RECT 76.665 160.615 78.015 161.525 ;
        RECT 82.155 161.295 83.085 161.525 ;
        RECT 86.295 161.295 87.225 161.525 ;
        RECT 79.185 160.615 83.085 161.295 ;
        RECT 83.325 160.615 87.225 161.295 ;
        RECT 87.245 160.700 87.675 161.485 ;
        RECT 87.790 161.295 88.710 161.525 ;
        RECT 87.790 160.615 91.255 161.295 ;
        RECT 91.375 160.615 92.745 161.395 ;
        RECT 95.955 161.295 96.885 161.525 ;
        RECT 92.985 160.615 96.885 161.295 ;
        RECT 97.450 161.295 98.370 161.525 ;
        RECT 104.235 161.295 105.165 161.525 ;
        RECT 107.830 161.295 108.750 161.525 ;
        RECT 97.450 160.615 100.915 161.295 ;
        RECT 101.265 160.615 105.165 161.295 ;
        RECT 105.285 160.615 108.750 161.295 ;
        RECT 108.855 160.615 111.465 161.525 ;
        RECT 112.075 160.615 113.445 161.425 ;
        RECT 11.475 160.405 11.645 160.615 ;
        RECT 12.910 160.455 13.030 160.565 ;
        RECT 13.315 160.405 13.485 160.595 ;
        RECT 13.775 160.425 13.945 160.615 ;
        RECT 16.995 160.425 17.165 160.595 ;
        RECT 17.730 160.425 17.900 160.615 ;
        RECT 22.055 160.460 22.215 160.570 ;
        RECT 22.790 160.425 22.960 160.615 ;
        RECT 23.435 160.405 23.605 160.595 ;
        RECT 26.655 160.425 26.825 160.615 ;
        RECT 28.035 160.405 28.205 160.595 ;
        RECT 31.710 160.405 31.880 160.595 ;
        RECT 32.175 160.405 32.345 160.595 ;
        RECT 33.555 160.405 33.725 160.595 ;
        RECT 37.235 160.405 37.405 160.595 ;
        RECT 39.720 160.425 39.890 160.615 ;
        RECT 41.190 160.405 41.360 160.595 ;
        RECT 45.110 160.455 45.230 160.565 ;
        RECT 45.515 160.405 45.685 160.595 ;
        RECT 49.195 160.425 49.365 160.615 ;
        RECT 49.655 160.450 49.815 160.560 ;
        RECT 50.115 160.405 50.285 160.595 ;
        RECT 50.575 160.425 50.745 160.615 ;
        RECT 51.500 160.405 51.670 160.595 ;
        RECT 56.095 160.425 56.265 160.615 ;
        RECT 56.555 160.425 56.725 160.615 ;
        RECT 59.315 160.425 59.485 160.615 ;
        RECT 61.155 160.425 61.325 160.615 ;
        RECT 62.075 160.425 62.245 160.615 ;
        RECT 63.915 160.425 64.085 160.615 ;
        RECT 64.375 160.405 64.545 160.595 ;
        RECT 65.755 160.565 65.925 160.595 ;
        RECT 65.755 160.455 65.930 160.565 ;
        RECT 65.755 160.405 65.925 160.455 ;
        RECT 69.435 160.425 69.605 160.615 ;
        RECT 69.620 160.405 69.790 160.595 ;
        RECT 69.895 160.425 70.065 160.615 ;
        RECT 71.550 160.425 71.720 160.615 ;
        RECT 73.760 160.405 73.930 160.595 ;
        RECT 75.010 160.455 75.130 160.565 ;
        RECT 75.415 160.405 75.585 160.595 ;
        RECT 76.335 160.425 76.505 160.615 ;
        RECT 76.850 160.455 76.970 160.565 ;
        RECT 77.715 160.425 77.885 160.615 ;
        RECT 78.635 160.460 78.795 160.570 ;
        RECT 82.500 160.425 82.670 160.615 ;
        RECT 86.455 160.405 86.625 160.595 ;
        RECT 86.640 160.425 86.810 160.615 ;
        RECT 87.375 160.450 87.535 160.560 ;
        RECT 88.755 160.405 88.925 160.595 ;
        RECT 90.595 160.405 90.765 160.595 ;
        RECT 91.055 160.425 91.225 160.615 ;
        RECT 92.435 160.425 92.605 160.615 ;
        RECT 94.270 160.405 94.440 160.595 ;
        RECT 94.740 160.405 94.910 160.595 ;
        RECT 96.300 160.425 96.470 160.615 ;
        RECT 97.090 160.455 97.210 160.565 ;
        RECT 99.795 160.405 99.965 160.595 ;
        RECT 100.715 160.425 100.885 160.615 ;
        RECT 103.015 160.405 103.185 160.595 ;
        RECT 103.480 160.405 103.650 160.595 ;
        RECT 104.580 160.425 104.750 160.615 ;
        RECT 105.315 160.425 105.485 160.615 ;
        RECT 106.290 160.455 106.410 160.565 ;
        RECT 109.000 160.425 109.170 160.615 ;
        RECT 111.755 160.565 111.925 160.595 ;
        RECT 111.755 160.455 111.930 160.565 ;
        RECT 111.755 160.405 111.925 160.455 ;
        RECT 113.135 160.405 113.305 160.615 ;
        RECT 11.335 159.595 12.705 160.405 ;
        RECT 13.175 159.725 22.455 160.405 ;
        RECT 14.535 159.505 15.455 159.725 ;
        RECT 20.120 159.605 22.455 159.725 ;
        RECT 21.535 159.495 22.455 159.605 ;
        RECT 22.845 159.535 23.275 160.320 ;
        RECT 23.295 159.625 24.665 160.405 ;
        RECT 24.770 159.725 28.235 160.405 ;
        RECT 24.770 159.495 25.690 159.725 ;
        RECT 28.550 159.495 32.025 160.405 ;
        RECT 32.045 159.495 33.395 160.405 ;
        RECT 33.525 159.725 36.990 160.405 ;
        RECT 37.205 159.725 40.670 160.405 ;
        RECT 36.070 159.495 36.990 159.725 ;
        RECT 39.750 159.495 40.670 159.725 ;
        RECT 40.775 159.725 44.675 160.405 ;
        RECT 40.775 159.495 41.705 159.725 ;
        RECT 45.375 159.495 48.585 160.405 ;
        RECT 48.605 159.535 49.035 160.320 ;
        RECT 49.985 159.495 51.335 160.405 ;
        RECT 51.355 159.495 54.830 160.405 ;
        RECT 55.405 159.725 64.685 160.405 ;
        RECT 55.405 159.605 57.740 159.725 ;
        RECT 55.405 159.495 56.325 159.605 ;
        RECT 62.405 159.505 63.325 159.725 ;
        RECT 64.695 159.595 66.065 160.405 ;
        RECT 66.305 159.725 70.205 160.405 ;
        RECT 70.445 159.725 74.345 160.405 ;
        RECT 69.275 159.495 70.205 159.725 ;
        RECT 73.415 159.495 74.345 159.725 ;
        RECT 74.365 159.535 74.795 160.320 ;
        RECT 75.275 159.625 76.645 160.405 ;
        RECT 77.485 159.725 86.765 160.405 ;
        RECT 77.485 159.605 79.820 159.725 ;
        RECT 77.485 159.495 78.405 159.605 ;
        RECT 84.485 159.505 85.405 159.725 ;
        RECT 87.705 159.495 89.055 160.405 ;
        RECT 89.075 159.595 90.905 160.405 ;
        RECT 91.110 159.495 94.585 160.405 ;
        RECT 94.595 159.495 98.070 160.405 ;
        RECT 98.275 159.595 100.105 160.405 ;
        RECT 100.125 159.535 100.555 160.320 ;
        RECT 100.575 159.595 103.325 160.405 ;
        RECT 103.335 159.495 105.945 160.405 ;
        RECT 106.555 159.595 112.065 160.405 ;
        RECT 112.075 159.595 113.445 160.405 ;
      LAYER nwell ;
        RECT 11.140 156.375 113.640 159.205 ;
      LAYER pwell ;
        RECT 11.335 155.175 12.705 155.985 ;
        RECT 12.715 155.175 14.545 155.985 ;
        RECT 14.555 155.175 15.925 155.955 ;
        RECT 15.935 155.855 16.865 156.085 ;
        RECT 29.275 155.885 30.220 156.085 ;
        RECT 15.935 155.175 19.835 155.855 ;
        RECT 20.160 155.175 29.265 155.855 ;
        RECT 29.275 155.205 32.025 155.885 ;
        RECT 34.690 155.855 35.610 156.085 ;
        RECT 29.275 155.175 30.220 155.205 ;
        RECT 11.475 154.965 11.645 155.175 ;
        RECT 13.775 154.965 13.945 155.155 ;
        RECT 14.235 154.965 14.405 155.175 ;
        RECT 15.615 154.985 15.785 155.175 ;
        RECT 16.350 154.985 16.520 155.175 ;
        RECT 16.535 154.965 16.705 155.155 ;
        RECT 17.270 154.965 17.440 155.155 ;
        RECT 22.515 154.965 22.685 155.155 ;
        RECT 24.355 154.965 24.525 155.155 ;
        RECT 24.820 154.965 24.990 155.155 ;
        RECT 28.955 154.985 29.125 155.175 ;
        RECT 31.710 154.965 31.880 155.205 ;
        RECT 32.145 155.175 35.610 155.855 ;
        RECT 35.725 155.260 36.155 156.045 ;
        RECT 36.175 155.885 37.120 156.085 ;
        RECT 36.175 155.205 38.925 155.885 ;
        RECT 36.175 155.175 37.120 155.205 ;
        RECT 32.175 154.965 32.345 155.175 ;
        RECT 36.770 154.965 36.940 155.155 ;
        RECT 38.610 154.985 38.780 155.205 ;
        RECT 38.935 155.175 42.410 156.085 ;
        RECT 43.535 155.175 44.905 155.955 ;
        RECT 45.010 155.855 45.930 156.085 ;
        RECT 45.010 155.175 48.475 155.855 ;
        RECT 48.595 155.175 49.965 155.985 ;
        RECT 50.345 155.975 51.265 156.085 ;
        RECT 50.345 155.855 52.680 155.975 ;
        RECT 57.345 155.855 58.265 156.075 ;
        RECT 50.345 155.175 59.625 155.855 ;
        RECT 60.095 155.175 61.465 155.955 ;
        RECT 61.485 155.260 61.915 156.045 ;
        RECT 61.935 155.175 63.765 155.985 ;
        RECT 63.775 155.855 65.120 156.085 ;
        RECT 63.775 155.175 65.605 155.855 ;
        RECT 65.810 155.175 69.285 156.085 ;
        RECT 69.665 155.975 70.585 156.085 ;
        RECT 69.665 155.855 72.000 155.975 ;
        RECT 76.665 155.855 77.585 156.075 ;
        RECT 69.665 155.175 78.945 155.855 ;
        RECT 79.425 155.175 80.775 156.085 ;
        RECT 83.995 155.855 84.925 156.085 ;
        RECT 81.025 155.175 84.925 155.855 ;
        RECT 84.935 155.175 86.305 155.955 ;
        RECT 87.245 155.260 87.675 156.045 ;
        RECT 88.155 155.175 90.905 155.985 ;
        RECT 91.110 155.175 94.585 156.085 ;
        RECT 94.595 155.175 96.425 155.985 ;
        RECT 96.435 155.175 99.910 156.085 ;
        RECT 100.115 155.175 103.590 156.085 ;
        RECT 104.265 155.175 105.615 156.085 ;
        RECT 105.645 155.175 106.995 156.085 ;
        RECT 107.475 155.175 108.845 155.955 ;
        RECT 109.315 155.175 112.065 155.985 ;
        RECT 112.075 155.175 113.445 155.985 ;
        RECT 39.080 154.985 39.250 155.175 ;
        RECT 40.450 154.965 40.620 155.155 ;
        RECT 40.920 154.965 41.090 155.155 ;
        RECT 43.215 155.020 43.375 155.130 ;
        RECT 43.675 154.985 43.845 155.175 ;
        RECT 44.595 154.965 44.765 155.155 ;
        RECT 48.275 155.125 48.445 155.175 ;
        RECT 48.275 155.015 48.450 155.125 ;
        RECT 48.275 154.985 48.445 155.015 ;
        RECT 49.470 154.965 49.640 155.155 ;
        RECT 49.655 154.985 49.825 155.175 ;
        RECT 59.315 154.985 59.485 155.175 ;
        RECT 59.830 155.015 59.950 155.125 ;
        RECT 60.235 154.985 60.405 155.175 ;
        RECT 62.075 154.965 62.245 155.155 ;
        RECT 63.455 154.965 63.625 155.175 ;
        RECT 63.920 154.965 64.090 155.155 ;
        RECT 65.295 154.985 65.465 155.175 ;
        RECT 68.970 154.985 69.140 155.175 ;
        RECT 70.810 154.965 70.980 155.155 ;
        RECT 72.655 154.965 72.825 155.155 ;
        RECT 74.035 154.965 74.205 155.155 ;
        RECT 75.415 155.010 75.575 155.120 ;
        RECT 78.635 154.985 78.805 155.175 ;
        RECT 79.095 155.125 79.265 155.155 ;
        RECT 79.095 155.015 79.270 155.125 ;
        RECT 79.095 154.965 79.265 155.015 ;
        RECT 79.555 154.985 79.725 155.175 ;
        RECT 84.340 154.985 84.510 155.175 ;
        RECT 84.615 154.965 84.785 155.155 ;
        RECT 85.080 154.965 85.250 155.155 ;
        RECT 85.995 154.985 86.165 155.175 ;
        RECT 86.915 155.020 87.075 155.130 ;
        RECT 87.890 155.015 88.010 155.125 ;
        RECT 89.675 154.965 89.845 155.155 ;
        RECT 90.595 154.985 90.765 155.175 ;
        RECT 11.335 154.155 12.705 154.965 ;
        RECT 12.715 154.155 14.085 154.965 ;
        RECT 14.105 154.055 15.455 154.965 ;
        RECT 15.475 154.185 16.845 154.965 ;
        RECT 16.855 154.285 20.755 154.965 ;
        RECT 16.855 154.055 17.785 154.285 ;
        RECT 20.995 154.155 22.825 154.965 ;
        RECT 22.845 154.095 23.275 154.880 ;
        RECT 23.305 154.055 24.655 154.965 ;
        RECT 24.675 154.055 28.150 154.965 ;
        RECT 28.550 154.055 32.025 154.965 ;
        RECT 32.045 154.055 33.395 154.965 ;
        RECT 33.610 154.055 37.085 154.965 ;
        RECT 37.290 154.055 40.765 154.965 ;
        RECT 40.775 154.055 44.250 154.965 ;
        RECT 44.565 154.285 48.030 154.965 ;
        RECT 47.110 154.055 48.030 154.285 ;
        RECT 48.605 154.095 49.035 154.880 ;
        RECT 49.055 154.285 52.955 154.965 ;
        RECT 53.280 154.285 62.385 154.965 ;
        RECT 49.055 154.055 49.985 154.285 ;
        RECT 62.395 154.155 63.765 154.965 ;
        RECT 63.775 154.055 67.250 154.965 ;
        RECT 67.650 154.055 71.125 154.965 ;
        RECT 71.135 154.155 72.965 154.965 ;
        RECT 72.985 154.055 74.335 154.965 ;
        RECT 74.365 154.095 74.795 154.880 ;
        RECT 75.735 154.155 79.405 154.965 ;
        RECT 79.415 154.155 84.925 154.965 ;
        RECT 84.935 154.055 88.410 154.965 ;
        RECT 88.615 154.155 89.985 154.965 ;
        RECT 89.995 154.935 90.940 154.965 ;
        RECT 92.430 154.935 92.600 155.155 ;
        RECT 94.270 154.985 94.440 155.175 ;
        RECT 96.115 155.155 96.285 155.175 ;
        RECT 96.580 155.155 96.750 155.175 ;
        RECT 96.110 154.985 96.285 155.155 ;
        RECT 96.575 154.985 96.750 155.155 ;
        RECT 100.260 154.985 100.430 155.175 ;
        RECT 96.110 154.965 96.280 154.985 ;
        RECT 96.575 154.965 96.745 154.985 ;
        RECT 102.095 154.965 102.265 155.155 ;
        RECT 103.990 155.015 104.110 155.125 ;
        RECT 104.395 154.985 104.565 155.175 ;
        RECT 105.775 154.985 105.945 155.175 ;
        RECT 107.210 155.015 107.330 155.125 ;
        RECT 107.615 154.985 107.785 155.175 ;
        RECT 109.050 155.015 109.170 155.125 ;
        RECT 111.295 154.965 111.465 155.155 ;
        RECT 111.755 155.125 111.925 155.175 ;
        RECT 111.755 155.015 111.930 155.125 ;
        RECT 111.755 154.985 111.925 155.015 ;
        RECT 113.135 154.965 113.305 155.175 ;
        RECT 89.995 154.255 92.745 154.935 ;
        RECT 89.995 154.055 90.940 154.255 ;
        RECT 92.950 154.055 96.425 154.965 ;
        RECT 96.545 154.285 100.010 154.965 ;
        RECT 99.090 154.055 100.010 154.285 ;
        RECT 100.125 154.095 100.555 154.880 ;
        RECT 100.575 154.155 102.405 154.965 ;
        RECT 102.415 154.285 111.605 154.965 ;
        RECT 102.415 154.055 103.335 154.285 ;
        RECT 106.165 154.065 107.095 154.285 ;
        RECT 112.075 154.155 113.445 154.965 ;
      LAYER nwell ;
        RECT 11.140 150.935 113.640 153.765 ;
      LAYER pwell ;
        RECT 11.335 149.735 12.705 150.545 ;
        RECT 14.075 150.415 14.995 150.635 ;
        RECT 21.075 150.535 21.995 150.645 ;
        RECT 19.660 150.415 21.995 150.535 ;
        RECT 12.715 149.735 21.995 150.415 ;
        RECT 22.835 150.415 23.755 150.645 ;
        RECT 26.585 150.415 27.515 150.635 ;
        RECT 22.835 149.735 32.025 150.415 ;
        RECT 32.230 149.735 35.705 150.645 ;
        RECT 35.725 149.820 36.155 150.605 ;
        RECT 36.185 149.735 37.535 150.645 ;
        RECT 37.555 150.415 38.485 150.645 ;
        RECT 37.555 149.735 41.455 150.415 ;
        RECT 42.155 149.735 44.905 150.545 ;
        RECT 44.915 150.415 45.835 150.645 ;
        RECT 48.665 150.415 49.595 150.635 ;
        RECT 44.915 149.735 54.105 150.415 ;
        RECT 54.115 149.735 55.945 150.545 ;
        RECT 59.155 150.415 60.085 150.645 ;
        RECT 56.185 149.735 60.085 150.415 ;
        RECT 60.095 149.735 61.465 150.545 ;
        RECT 61.485 149.820 61.915 150.605 ;
        RECT 64.695 150.415 66.040 150.645 ;
        RECT 66.535 150.415 67.880 150.645 ;
        RECT 61.945 149.735 64.685 150.415 ;
        RECT 64.695 149.735 66.525 150.415 ;
        RECT 66.535 149.735 68.365 150.415 ;
        RECT 68.375 149.735 71.850 150.645 ;
        RECT 72.540 150.415 73.885 150.645 ;
        RECT 72.055 149.735 73.885 150.415 ;
        RECT 73.895 149.735 77.565 150.545 ;
        RECT 77.575 149.735 83.085 150.545 ;
        RECT 83.105 149.735 84.455 150.645 ;
        RECT 85.395 149.735 86.765 150.515 ;
        RECT 87.245 149.820 87.675 150.605 ;
        RECT 88.155 149.735 91.825 150.545 ;
        RECT 93.640 150.445 94.585 150.645 ;
        RECT 91.835 149.765 94.585 150.445 ;
        RECT 11.475 149.525 11.645 149.735 ;
        RECT 12.855 149.685 13.025 149.735 ;
        RECT 12.855 149.575 13.030 149.685 ;
        RECT 12.855 149.545 13.025 149.575 ;
        RECT 13.315 149.525 13.485 149.715 ;
        RECT 22.570 149.575 22.690 149.685 ;
        RECT 23.895 149.570 24.055 149.680 ;
        RECT 11.335 148.715 12.705 149.525 ;
        RECT 13.175 148.845 22.455 149.525 ;
        RECT 24.215 149.495 25.160 149.525 ;
        RECT 26.650 149.495 26.820 149.715 ;
        RECT 30.520 149.525 30.690 149.715 ;
        RECT 31.255 149.525 31.425 149.715 ;
        RECT 31.715 149.545 31.885 149.735 ;
        RECT 35.390 149.545 35.560 149.735 ;
        RECT 37.235 149.545 37.405 149.735 ;
        RECT 37.970 149.545 38.140 149.735 ;
        RECT 40.510 149.575 40.630 149.685 ;
        RECT 41.890 149.575 42.010 149.685 ;
        RECT 44.130 149.525 44.300 149.715 ;
        RECT 44.595 149.545 44.765 149.735 ;
        RECT 46.895 149.525 47.065 149.715 ;
        RECT 47.355 149.525 47.525 149.715 ;
        RECT 50.115 149.525 50.285 149.715 ;
        RECT 50.575 149.525 50.745 149.715 ;
        RECT 51.960 149.525 52.130 149.715 ;
        RECT 53.795 149.545 53.965 149.735 ;
        RECT 55.635 149.545 55.805 149.735 ;
        RECT 56.095 149.570 56.255 149.680 ;
        RECT 59.500 149.545 59.670 149.735 ;
        RECT 61.155 149.545 61.325 149.735 ;
        RECT 64.375 149.545 64.545 149.735 ;
        RECT 65.755 149.525 65.925 149.715 ;
        RECT 66.215 149.525 66.385 149.735 ;
        RECT 68.055 149.545 68.225 149.735 ;
        RECT 68.520 149.545 68.690 149.735 ;
        RECT 68.975 149.525 69.145 149.715 ;
        RECT 72.195 149.545 72.365 149.735 ;
        RECT 74.035 149.525 74.205 149.715 ;
        RECT 75.875 149.525 76.045 149.715 ;
        RECT 77.255 149.545 77.425 149.735 ;
        RECT 79.740 149.525 79.910 149.715 ;
        RECT 82.775 149.545 82.945 149.735 ;
        RECT 84.155 149.545 84.325 149.735 ;
        RECT 85.075 149.580 85.235 149.690 ;
        RECT 85.535 149.545 85.705 149.735 ;
        RECT 86.970 149.575 87.090 149.685 ;
        RECT 87.890 149.575 88.010 149.685 ;
        RECT 89.215 149.525 89.385 149.715 ;
        RECT 89.675 149.525 89.845 149.715 ;
        RECT 91.515 149.545 91.685 149.735 ;
        RECT 91.980 149.545 92.150 149.765 ;
        RECT 93.640 149.735 94.585 149.765 ;
        RECT 94.790 149.735 98.265 150.645 ;
        RECT 101.475 150.415 102.405 150.645 ;
        RECT 98.505 149.735 102.405 150.415 ;
        RECT 102.785 150.535 103.705 150.645 ;
        RECT 102.785 150.415 105.120 150.535 ;
        RECT 109.785 150.415 110.705 150.635 ;
        RECT 102.785 149.735 112.065 150.415 ;
        RECT 112.075 149.735 113.445 150.545 ;
        RECT 93.410 149.575 93.530 149.685 ;
        RECT 93.820 149.525 93.990 149.715 ;
        RECT 14.535 148.625 15.455 148.845 ;
        RECT 20.120 148.725 22.455 148.845 ;
        RECT 21.535 148.615 22.455 148.725 ;
        RECT 22.845 148.655 23.275 149.440 ;
        RECT 24.215 148.815 26.965 149.495 ;
        RECT 27.205 148.845 31.105 149.525 ;
        RECT 31.115 148.845 40.305 149.525 ;
        RECT 24.215 148.615 25.160 148.815 ;
        RECT 30.175 148.615 31.105 148.845 ;
        RECT 35.625 148.625 36.555 148.845 ;
        RECT 39.385 148.615 40.305 148.845 ;
        RECT 40.970 148.615 44.445 149.525 ;
        RECT 44.455 148.715 47.205 149.525 ;
        RECT 47.225 148.615 48.575 149.525 ;
        RECT 48.605 148.655 49.035 149.440 ;
        RECT 49.055 148.715 50.425 149.525 ;
        RECT 50.435 148.745 51.805 149.525 ;
        RECT 51.815 148.615 55.290 149.525 ;
        RECT 56.785 148.845 66.065 149.525 ;
        RECT 56.785 148.725 59.120 148.845 ;
        RECT 56.785 148.615 57.705 148.725 ;
        RECT 63.785 148.625 64.705 148.845 ;
        RECT 66.075 148.615 68.795 149.525 ;
        RECT 68.835 148.845 71.575 149.525 ;
        RECT 71.595 148.715 74.345 149.525 ;
        RECT 74.365 148.655 74.795 149.440 ;
        RECT 74.815 148.715 76.185 149.525 ;
        RECT 76.425 148.845 80.325 149.525 ;
        RECT 79.395 148.615 80.325 148.845 ;
        RECT 80.335 148.845 89.525 149.525 ;
        RECT 89.645 148.845 93.110 149.525 ;
        RECT 80.335 148.615 81.255 148.845 ;
        RECT 84.085 148.625 85.015 148.845 ;
        RECT 92.190 148.615 93.110 148.845 ;
        RECT 93.675 148.615 97.150 149.525 ;
        RECT 97.500 149.495 97.670 149.715 ;
        RECT 97.950 149.545 98.120 149.735 ;
        RECT 101.820 149.545 101.990 149.735 ;
        RECT 102.095 149.525 102.265 149.715 ;
        RECT 105.960 149.525 106.130 149.715 ;
        RECT 107.615 149.525 107.785 149.715 ;
        RECT 108.075 149.525 108.245 149.715 ;
        RECT 111.755 149.525 111.925 149.735 ;
        RECT 113.135 149.525 113.305 149.735 ;
        RECT 99.160 149.495 100.105 149.525 ;
        RECT 97.355 148.815 100.105 149.495 ;
        RECT 99.160 148.615 100.105 148.815 ;
        RECT 100.125 148.655 100.555 149.440 ;
        RECT 100.575 148.715 102.405 149.525 ;
        RECT 102.645 148.845 106.545 149.525 ;
        RECT 105.615 148.615 106.545 148.845 ;
        RECT 106.555 148.715 107.925 149.525 ;
        RECT 107.935 148.745 109.305 149.525 ;
        RECT 109.315 148.715 112.065 149.525 ;
        RECT 112.075 148.715 113.445 149.525 ;
      LAYER nwell ;
        RECT 11.140 145.495 113.640 148.325 ;
      LAYER pwell ;
        RECT 11.335 144.295 12.705 145.105 ;
        RECT 13.645 144.295 14.995 145.205 ;
        RECT 15.015 144.295 16.385 145.075 ;
        RECT 19.050 144.975 19.970 145.205 ;
        RECT 16.505 144.295 19.970 144.975 ;
        RECT 20.075 144.975 21.005 145.205 ;
        RECT 20.075 144.295 23.975 144.975 ;
        RECT 24.215 144.295 26.965 145.105 ;
        RECT 29.630 144.975 30.550 145.205 ;
        RECT 27.085 144.295 30.550 144.975 ;
        RECT 30.750 144.975 31.670 145.205 ;
        RECT 30.750 144.295 34.215 144.975 ;
        RECT 34.335 144.295 35.705 145.075 ;
        RECT 35.725 144.380 36.155 145.165 ;
        RECT 37.095 144.295 38.465 145.075 ;
        RECT 38.670 144.295 42.145 145.205 ;
        RECT 42.615 144.295 45.365 145.105 ;
        RECT 45.375 144.295 50.885 145.105 ;
        RECT 50.895 144.295 54.370 145.205 ;
        RECT 54.575 144.295 55.945 145.105 ;
        RECT 59.155 144.975 60.085 145.205 ;
        RECT 56.185 144.295 60.085 144.975 ;
        RECT 60.105 144.295 61.455 145.205 ;
        RECT 61.485 144.380 61.915 145.165 ;
        RECT 62.395 144.975 63.740 145.205 ;
        RECT 64.720 144.975 66.065 145.205 ;
        RECT 66.560 144.975 67.905 145.205 ;
        RECT 62.395 144.295 64.225 144.975 ;
        RECT 64.235 144.295 66.065 144.975 ;
        RECT 66.075 144.295 67.905 144.975 ;
        RECT 68.835 144.295 72.505 145.105 ;
        RECT 72.525 144.295 73.875 145.205 ;
        RECT 74.265 145.095 75.185 145.205 ;
        RECT 74.265 144.975 76.600 145.095 ;
        RECT 81.265 144.975 82.185 145.195 ;
        RECT 74.265 144.295 83.545 144.975 ;
        RECT 83.555 144.295 87.225 145.105 ;
        RECT 87.245 144.380 87.675 145.165 ;
        RECT 87.695 144.295 91.365 145.105 ;
        RECT 91.375 145.005 92.320 145.205 ;
        RECT 91.375 144.325 94.125 145.005 ;
        RECT 91.375 144.295 92.320 144.325 ;
        RECT 11.475 144.085 11.645 144.295 ;
        RECT 13.315 144.130 13.475 144.250 ;
        RECT 13.775 144.105 13.945 144.295 ;
        RECT 16.075 144.105 16.245 144.295 ;
        RECT 16.535 144.105 16.705 144.295 ;
        RECT 16.995 144.085 17.165 144.275 ;
        RECT 20.490 144.105 20.660 144.295 ;
        RECT 22.515 144.085 22.685 144.275 ;
        RECT 23.490 144.135 23.610 144.245 ;
        RECT 26.655 144.105 26.825 144.295 ;
        RECT 27.115 144.105 27.285 144.295 ;
        RECT 28.955 144.085 29.125 144.275 ;
        RECT 11.335 143.275 12.705 144.085 ;
        RECT 13.635 143.275 17.305 144.085 ;
        RECT 17.315 143.275 22.825 144.085 ;
        RECT 22.845 143.215 23.275 144.000 ;
        RECT 23.755 143.275 29.265 144.085 ;
        RECT 29.275 144.055 30.220 144.085 ;
        RECT 31.710 144.055 31.880 144.275 ;
        RECT 32.230 144.135 32.350 144.245 ;
        RECT 34.015 144.105 34.185 144.295 ;
        RECT 35.395 144.105 35.565 144.295 ;
        RECT 36.775 144.140 36.935 144.250 ;
        RECT 37.695 144.085 37.865 144.275 ;
        RECT 38.155 144.105 38.325 144.295 ;
        RECT 41.830 144.105 42.000 144.295 ;
        RECT 42.350 144.135 42.470 144.245 ;
        RECT 43.215 144.085 43.385 144.275 ;
        RECT 43.680 144.085 43.850 144.275 ;
        RECT 45.055 144.105 45.225 144.295 ;
        RECT 48.275 144.085 48.445 144.275 ;
        RECT 50.115 144.085 50.285 144.275 ;
        RECT 50.575 144.105 50.745 144.295 ;
        RECT 51.040 144.105 51.210 144.295 ;
        RECT 53.980 144.085 54.150 144.275 ;
        RECT 54.770 144.135 54.890 144.245 ;
        RECT 55.175 144.085 55.345 144.275 ;
        RECT 55.635 144.105 55.805 144.295 ;
        RECT 57.475 144.085 57.645 144.275 ;
        RECT 59.500 144.105 59.670 144.295 ;
        RECT 61.155 144.085 61.325 144.295 ;
        RECT 61.615 144.085 61.785 144.275 ;
        RECT 62.130 144.135 62.250 144.245 ;
        RECT 63.455 144.130 63.615 144.240 ;
        RECT 63.915 144.105 64.085 144.295 ;
        RECT 64.375 144.105 64.545 144.295 ;
        RECT 66.215 144.105 66.385 144.295 ;
        RECT 67.135 144.085 67.305 144.275 ;
        RECT 68.515 144.140 68.675 144.250 ;
        RECT 29.275 143.375 32.025 144.055 ;
        RECT 29.275 143.175 30.220 143.375 ;
        RECT 32.495 143.275 38.005 144.085 ;
        RECT 38.015 143.275 43.525 144.085 ;
        RECT 43.535 143.175 47.010 144.085 ;
        RECT 47.215 143.275 48.585 144.085 ;
        RECT 48.605 143.215 49.035 144.000 ;
        RECT 49.055 143.275 50.425 144.085 ;
        RECT 50.665 143.405 54.565 144.085 ;
        RECT 53.635 143.175 54.565 143.405 ;
        RECT 55.035 143.305 56.405 144.085 ;
        RECT 56.415 143.275 57.785 144.085 ;
        RECT 57.795 143.275 61.465 144.085 ;
        RECT 61.475 143.305 62.845 144.085 ;
        RECT 63.775 143.275 67.445 144.085 ;
        RECT 67.455 144.055 68.400 144.085 ;
        RECT 69.890 144.055 70.060 144.275 ;
        RECT 70.360 144.085 70.530 144.275 ;
        RECT 72.195 144.105 72.365 144.295 ;
        RECT 73.575 144.105 73.745 144.295 ;
        RECT 74.090 144.135 74.210 144.245 ;
        RECT 75.010 144.135 75.130 144.245 ;
        RECT 78.820 144.085 78.990 144.275 ;
        RECT 79.555 144.085 79.725 144.275 ;
        RECT 80.990 144.135 81.110 144.245 ;
        RECT 83.235 144.105 83.405 144.295 ;
        RECT 84.615 144.085 84.785 144.275 ;
        RECT 86.915 144.105 87.085 144.295 ;
        RECT 67.455 143.375 70.205 144.055 ;
        RECT 67.455 143.175 68.400 143.375 ;
        RECT 70.215 143.175 73.690 144.085 ;
        RECT 74.365 143.215 74.795 144.000 ;
        RECT 75.505 143.405 79.405 144.085 ;
        RECT 78.475 143.175 79.405 143.405 ;
        RECT 79.415 143.305 80.785 144.085 ;
        RECT 81.255 143.275 84.925 144.085 ;
        RECT 84.935 144.055 85.880 144.085 ;
        RECT 87.370 144.055 87.540 144.275 ;
        RECT 87.840 144.085 88.010 144.275 ;
        RECT 91.055 144.105 91.225 144.295 ;
        RECT 93.810 144.275 93.980 144.325 ;
        RECT 94.135 144.295 96.885 145.105 ;
        RECT 97.090 144.295 100.565 145.205 ;
        RECT 100.575 144.295 102.405 145.105 ;
        RECT 105.615 144.975 106.545 145.205 ;
        RECT 102.645 144.295 106.545 144.975 ;
        RECT 106.565 144.295 107.915 145.205 ;
        RECT 107.935 144.295 109.305 145.075 ;
        RECT 109.315 144.295 112.065 145.105 ;
        RECT 112.075 144.295 113.445 145.105 ;
        RECT 91.570 144.135 91.690 144.245 ;
        RECT 93.355 144.085 93.525 144.275 ;
        RECT 93.810 144.105 93.990 144.275 ;
        RECT 96.575 144.105 96.745 144.295 ;
        RECT 93.820 144.085 93.990 144.105 ;
        RECT 84.935 143.375 87.685 144.055 ;
        RECT 84.935 143.175 85.880 143.375 ;
        RECT 87.695 143.175 91.170 144.085 ;
        RECT 91.835 143.275 93.665 144.085 ;
        RECT 93.675 143.175 97.150 144.085 ;
        RECT 97.355 144.055 98.300 144.085 ;
        RECT 99.790 144.055 99.960 144.275 ;
        RECT 100.250 144.105 100.420 144.295 ;
        RECT 100.770 144.135 100.890 144.245 ;
        RECT 101.175 144.085 101.345 144.275 ;
        RECT 102.095 144.105 102.265 144.295 ;
        RECT 105.960 144.105 106.130 144.295 ;
        RECT 107.615 144.105 107.785 144.295 ;
        RECT 108.075 144.105 108.245 144.295 ;
        RECT 111.755 144.085 111.925 144.295 ;
        RECT 113.135 144.085 113.305 144.295 ;
        RECT 97.355 143.375 100.105 144.055 ;
        RECT 97.355 143.175 98.300 143.375 ;
        RECT 100.125 143.215 100.555 144.000 ;
        RECT 101.045 143.175 102.395 144.085 ;
        RECT 102.785 143.405 112.065 144.085 ;
        RECT 102.785 143.285 105.120 143.405 ;
        RECT 102.785 143.175 103.705 143.285 ;
        RECT 109.785 143.185 110.705 143.405 ;
        RECT 112.075 143.275 113.445 144.085 ;
      LAYER nwell ;
        RECT 11.140 140.055 113.640 142.885 ;
      LAYER pwell ;
        RECT 11.335 138.855 12.705 139.665 ;
        RECT 13.175 138.855 16.845 139.665 ;
        RECT 16.865 138.855 18.215 139.765 ;
        RECT 19.155 139.535 20.085 139.765 ;
        RECT 19.155 138.855 23.055 139.535 ;
        RECT 24.225 138.855 25.575 139.765 ;
        RECT 26.255 139.675 27.205 139.765 ;
        RECT 29.495 139.675 30.445 139.765 ;
        RECT 26.255 138.855 28.185 139.675 ;
        RECT 11.475 138.645 11.645 138.855 ;
        RECT 12.910 138.695 13.030 138.805 ;
        RECT 16.535 138.665 16.705 138.855 ;
        RECT 17.915 138.665 18.085 138.855 ;
        RECT 18.835 138.700 18.995 138.810 ;
        RECT 19.570 138.665 19.740 138.855 ;
        RECT 22.515 138.645 22.685 138.835 ;
        RECT 23.895 138.700 24.055 138.810 ;
        RECT 24.355 138.665 24.525 138.855 ;
        RECT 28.035 138.835 28.185 138.855 ;
        RECT 28.515 138.855 30.445 139.675 ;
        RECT 30.655 138.855 32.025 139.665 ;
        RECT 32.035 138.855 35.705 139.665 ;
        RECT 35.725 138.940 36.155 139.725 ;
        RECT 36.635 138.855 38.465 139.665 ;
        RECT 40.280 139.565 41.225 139.765 ;
        RECT 43.040 139.565 43.985 139.765 ;
        RECT 38.475 138.885 41.225 139.565 ;
        RECT 41.235 138.885 43.985 139.565 ;
        RECT 28.515 138.835 28.665 138.855 ;
        RECT 25.790 138.695 25.910 138.805 ;
        RECT 28.035 138.665 28.205 138.835 ;
        RECT 28.495 138.665 28.665 138.835 ;
        RECT 31.715 138.665 31.885 138.855 ;
        RECT 32.635 138.645 32.805 138.835 ;
        RECT 34.935 138.665 35.105 138.835 ;
        RECT 35.395 138.665 35.565 138.855 ;
        RECT 35.855 138.690 36.015 138.800 ;
        RECT 36.370 138.695 36.490 138.805 ;
        RECT 38.155 138.665 38.325 138.855 ;
        RECT 38.620 138.835 38.790 138.885 ;
        RECT 40.280 138.855 41.225 138.885 ;
        RECT 38.610 138.665 38.790 138.835 ;
        RECT 39.130 138.695 39.250 138.805 ;
        RECT 41.380 138.665 41.550 138.885 ;
        RECT 43.040 138.855 43.985 138.885 ;
        RECT 43.995 138.855 45.365 139.665 ;
        RECT 45.375 138.855 48.850 139.765 ;
        RECT 49.425 139.655 50.345 139.765 ;
        RECT 49.425 139.535 51.760 139.655 ;
        RECT 56.425 139.535 57.345 139.755 ;
        RECT 49.425 138.855 58.705 139.535 ;
        RECT 58.715 138.855 61.465 139.665 ;
        RECT 61.485 138.940 61.915 139.725 ;
        RECT 61.935 138.855 63.765 139.665 ;
        RECT 63.775 138.855 69.285 139.665 ;
        RECT 69.295 138.855 72.770 139.765 ;
        RECT 72.975 138.855 74.805 139.665 ;
        RECT 78.015 139.535 78.945 139.765 ;
        RECT 75.045 138.855 78.945 139.535 ;
        RECT 79.415 138.855 80.785 139.635 ;
        RECT 80.795 138.855 82.165 139.635 ;
        RECT 82.175 138.855 83.545 139.665 ;
        RECT 83.555 138.855 87.225 139.665 ;
        RECT 87.245 138.940 87.675 139.725 ;
        RECT 87.695 138.855 93.205 139.665 ;
        RECT 96.415 139.535 97.345 139.765 ;
        RECT 93.445 138.855 97.345 139.535 ;
        RECT 97.815 138.855 100.565 139.665 ;
        RECT 100.945 139.655 101.865 139.765 ;
        RECT 100.945 139.535 103.280 139.655 ;
        RECT 107.945 139.535 108.865 139.755 ;
        RECT 100.945 138.855 110.225 139.535 ;
        RECT 110.235 138.855 112.065 139.665 ;
        RECT 112.075 138.855 113.445 139.665 ;
        RECT 45.055 138.835 45.225 138.855 ;
        RECT 34.935 138.645 35.085 138.665 ;
        RECT 11.335 137.835 12.705 138.645 ;
        RECT 13.545 137.965 22.825 138.645 ;
        RECT 13.545 137.845 15.880 137.965 ;
        RECT 13.545 137.735 14.465 137.845 ;
        RECT 20.545 137.745 21.465 137.965 ;
        RECT 22.845 137.775 23.275 138.560 ;
        RECT 23.665 137.965 32.945 138.645 ;
        RECT 23.665 137.845 26.000 137.965 ;
        RECT 23.665 137.735 24.585 137.845 ;
        RECT 30.665 137.745 31.585 137.965 ;
        RECT 33.155 137.825 35.085 138.645 ;
        RECT 36.175 138.615 37.120 138.645 ;
        RECT 38.610 138.615 38.780 138.665 ;
        RECT 44.595 138.645 44.765 138.835 ;
        RECT 45.055 138.665 45.230 138.835 ;
        RECT 45.520 138.665 45.690 138.855 ;
        RECT 49.250 138.695 49.370 138.805 ;
        RECT 45.060 138.645 45.230 138.665 ;
        RECT 51.035 138.645 51.205 138.835 ;
        RECT 51.495 138.645 51.665 138.835 ;
        RECT 56.280 138.645 56.450 138.835 ;
        RECT 57.475 138.690 57.635 138.800 ;
        RECT 57.935 138.645 58.105 138.835 ;
        RECT 58.395 138.665 58.565 138.855 ;
        RECT 61.155 138.665 61.325 138.855 ;
        RECT 62.535 138.645 62.705 138.835 ;
        RECT 63.455 138.665 63.625 138.855 ;
        RECT 64.375 138.645 64.545 138.835 ;
        RECT 64.890 138.695 65.010 138.805 ;
        RECT 67.595 138.645 67.765 138.835 ;
        RECT 68.975 138.665 69.145 138.855 ;
        RECT 69.440 138.665 69.610 138.855 ;
        RECT 36.175 137.935 38.925 138.615 ;
        RECT 33.155 137.735 34.105 137.825 ;
        RECT 36.175 137.735 37.120 137.935 ;
        RECT 39.395 137.835 44.905 138.645 ;
        RECT 44.915 137.735 48.390 138.645 ;
        RECT 48.605 137.775 49.035 138.560 ;
        RECT 49.515 137.835 51.345 138.645 ;
        RECT 51.365 137.735 52.715 138.645 ;
        RECT 52.965 137.965 56.865 138.645 ;
        RECT 55.935 137.735 56.865 137.965 ;
        RECT 57.795 137.865 59.165 138.645 ;
        RECT 59.175 137.835 62.845 138.645 ;
        RECT 62.855 137.965 64.685 138.645 ;
        RECT 65.155 137.835 67.905 138.645 ;
        RECT 67.915 138.615 68.860 138.645 ;
        RECT 70.350 138.615 70.520 138.835 ;
        RECT 70.870 138.695 70.990 138.805 ;
        RECT 72.655 138.645 72.825 138.835 ;
        RECT 74.035 138.645 74.205 138.835 ;
        RECT 74.495 138.665 74.665 138.855 ;
        RECT 78.360 138.665 78.530 138.855 ;
        RECT 79.150 138.695 79.270 138.805 ;
        RECT 79.555 138.665 79.725 138.855 ;
        RECT 80.935 138.665 81.105 138.855 ;
        RECT 83.235 138.665 83.405 138.855 ;
        RECT 84.155 138.645 84.325 138.835 ;
        RECT 84.670 138.695 84.790 138.805 ;
        RECT 86.915 138.665 87.085 138.855 ;
        RECT 88.480 138.645 88.650 138.835 ;
        RECT 92.895 138.665 93.065 138.855 ;
        RECT 96.760 138.665 96.930 138.855 ;
        RECT 97.550 138.695 97.670 138.805 ;
        RECT 98.415 138.645 98.585 138.835 ;
        RECT 99.795 138.645 99.965 138.835 ;
        RECT 100.255 138.665 100.425 138.855 ;
        RECT 100.770 138.695 100.890 138.805 ;
        RECT 104.580 138.645 104.750 138.835 ;
        RECT 105.775 138.690 105.935 138.800 ;
        RECT 106.235 138.645 106.405 138.835 ;
        RECT 108.075 138.690 108.235 138.800 ;
        RECT 109.915 138.665 110.085 138.855 ;
        RECT 111.755 138.645 111.925 138.855 ;
        RECT 113.135 138.645 113.305 138.855 ;
        RECT 67.915 137.935 70.665 138.615 ;
        RECT 67.915 137.735 68.860 137.935 ;
        RECT 71.135 137.835 72.965 138.645 ;
        RECT 72.985 137.735 74.335 138.645 ;
        RECT 74.365 137.775 74.795 138.560 ;
        RECT 75.185 137.965 84.465 138.645 ;
        RECT 85.165 137.965 89.065 138.645 ;
        RECT 75.185 137.845 77.520 137.965 ;
        RECT 75.185 137.735 76.105 137.845 ;
        RECT 82.185 137.745 83.105 137.965 ;
        RECT 88.135 137.735 89.065 137.965 ;
        RECT 89.445 137.965 98.725 138.645 ;
        RECT 89.445 137.845 91.780 137.965 ;
        RECT 89.445 137.735 90.365 137.845 ;
        RECT 96.445 137.745 97.365 137.965 ;
        RECT 98.735 137.835 100.105 138.645 ;
        RECT 100.125 137.775 100.555 138.560 ;
        RECT 101.265 137.965 105.165 138.645 ;
        RECT 104.235 137.735 105.165 137.965 ;
        RECT 106.095 137.865 107.465 138.645 ;
        RECT 108.395 137.835 112.065 138.645 ;
        RECT 112.075 137.835 113.445 138.645 ;
      LAYER nwell ;
        RECT 11.140 134.615 113.640 137.445 ;
      LAYER pwell ;
        RECT 11.335 133.415 12.705 134.225 ;
        RECT 12.715 133.415 16.385 134.225 ;
        RECT 19.595 134.095 20.525 134.325 ;
        RECT 16.625 133.415 20.525 134.095 ;
        RECT 20.995 133.415 22.365 134.195 ;
        RECT 22.375 133.415 25.125 134.225 ;
        RECT 25.135 133.415 26.505 134.195 ;
        RECT 26.515 134.095 27.445 134.325 ;
        RECT 34.555 134.235 35.505 134.325 ;
        RECT 26.515 133.415 30.415 134.095 ;
        RECT 30.655 133.415 33.405 134.225 ;
        RECT 33.575 133.415 35.505 134.235 ;
        RECT 35.725 133.500 36.155 134.285 ;
        RECT 37.095 134.125 38.040 134.325 ;
        RECT 37.095 133.445 39.845 134.125 ;
        RECT 37.095 133.415 38.040 133.445 ;
        RECT 11.475 133.205 11.645 133.415 ;
        RECT 16.075 133.225 16.245 133.415 ;
        RECT 19.940 133.225 20.110 133.415 ;
        RECT 20.730 133.255 20.850 133.365 ;
        RECT 22.055 133.205 22.225 133.415 ;
        RECT 22.570 133.255 22.690 133.365 ;
        RECT 23.435 133.205 23.605 133.395 ;
        RECT 24.815 133.225 24.985 133.415 ;
        RECT 25.275 133.225 25.445 133.415 ;
        RECT 26.930 133.225 27.100 133.415 ;
        RECT 28.955 133.205 29.125 133.395 ;
        RECT 29.690 133.205 29.860 133.395 ;
        RECT 33.095 133.225 33.265 133.415 ;
        RECT 33.575 133.395 33.725 133.415 ;
        RECT 33.555 133.365 33.725 133.395 ;
        RECT 33.555 133.255 33.730 133.365 ;
        RECT 33.555 133.225 33.725 133.255 ;
        RECT 34.015 133.225 34.185 133.395 ;
        RECT 36.315 133.225 36.485 133.395 ;
        RECT 36.775 133.260 36.935 133.370 ;
        RECT 39.530 133.225 39.700 133.445 ;
        RECT 39.855 133.415 43.330 134.325 ;
        RECT 43.535 133.415 47.010 134.325 ;
        RECT 47.215 133.415 50.690 134.325 ;
        RECT 52.185 134.215 53.105 134.325 ;
        RECT 52.185 134.095 54.520 134.215 ;
        RECT 59.185 134.095 60.105 134.315 ;
        RECT 52.185 133.415 61.465 134.095 ;
        RECT 61.485 133.500 61.915 134.285 ;
        RECT 61.935 133.415 63.305 134.225 ;
        RECT 63.315 134.125 64.260 134.325 ;
        RECT 63.315 133.445 66.065 134.125 ;
        RECT 63.315 133.415 64.260 133.445 ;
        RECT 40.000 133.395 40.170 133.415 ;
        RECT 39.995 133.225 40.170 133.395 ;
        RECT 34.035 133.205 34.185 133.225 ;
        RECT 36.335 133.205 36.485 133.225 ;
        RECT 39.995 133.205 40.165 133.225 ;
        RECT 11.335 132.395 12.705 133.205 ;
        RECT 13.085 132.525 22.365 133.205 ;
        RECT 13.085 132.405 15.420 132.525 ;
        RECT 13.085 132.295 14.005 132.405 ;
        RECT 20.085 132.305 21.005 132.525 ;
        RECT 22.845 132.335 23.275 133.120 ;
        RECT 23.305 132.295 24.655 133.205 ;
        RECT 25.595 132.395 29.265 133.205 ;
        RECT 29.275 132.525 33.175 133.205 ;
        RECT 29.275 132.295 30.205 132.525 ;
        RECT 34.035 132.385 35.965 133.205 ;
        RECT 36.335 132.385 38.265 133.205 ;
        RECT 38.475 132.395 40.305 133.205 ;
        RECT 40.460 133.175 40.630 133.395 ;
        RECT 43.680 133.225 43.850 133.415 ;
        RECT 42.120 133.175 43.065 133.205 ;
        RECT 40.315 132.495 43.065 133.175 ;
        RECT 35.015 132.295 35.965 132.385 ;
        RECT 37.315 132.295 38.265 132.385 ;
        RECT 42.120 132.295 43.065 132.495 ;
        RECT 43.075 133.175 44.020 133.205 ;
        RECT 45.510 133.175 45.680 133.395 ;
        RECT 47.360 133.225 47.530 133.415 ;
        RECT 48.275 133.205 48.445 133.395 ;
        RECT 50.575 133.205 50.745 133.395 ;
        RECT 51.035 133.205 51.205 133.395 ;
        RECT 51.495 133.260 51.655 133.370 ;
        RECT 55.820 133.205 55.990 133.395 ;
        RECT 57.015 133.250 57.175 133.360 ;
        RECT 57.475 133.205 57.645 133.395 ;
        RECT 61.155 133.205 61.325 133.415 ;
        RECT 62.995 133.205 63.165 133.415 ;
        RECT 65.295 133.225 65.465 133.395 ;
        RECT 65.750 133.365 65.920 133.445 ;
        RECT 66.075 133.415 69.550 134.325 ;
        RECT 69.755 133.415 73.230 134.325 ;
        RECT 76.635 134.095 77.565 134.325 ;
        RECT 73.665 133.415 77.565 134.095 ;
        RECT 77.945 134.215 78.865 134.325 ;
        RECT 77.945 134.095 80.280 134.215 ;
        RECT 84.945 134.095 85.865 134.315 ;
        RECT 77.945 133.415 87.225 134.095 ;
        RECT 87.245 133.500 87.675 134.285 ;
        RECT 87.705 133.415 89.055 134.325 ;
        RECT 89.075 133.415 90.445 134.195 ;
        RECT 90.915 133.415 92.745 134.225 ;
        RECT 92.765 133.415 94.115 134.325 ;
        RECT 94.135 133.415 95.965 134.225 ;
        RECT 95.975 133.415 97.345 134.195 ;
        RECT 97.355 133.415 101.025 134.225 ;
        RECT 101.035 133.415 106.545 134.225 ;
        RECT 106.555 133.415 112.065 134.225 ;
        RECT 112.075 133.415 113.445 134.225 ;
        RECT 65.750 133.255 65.930 133.365 ;
        RECT 65.750 133.225 65.920 133.255 ;
        RECT 66.220 133.225 66.390 133.415 ;
        RECT 65.295 133.205 65.445 133.225 ;
        RECT 67.595 133.205 67.765 133.395 ;
        RECT 43.075 132.495 45.825 133.175 ;
        RECT 43.075 132.295 44.020 132.495 ;
        RECT 45.835 132.395 48.585 133.205 ;
        RECT 48.605 132.335 49.035 133.120 ;
        RECT 49.055 132.395 50.885 133.205 ;
        RECT 50.905 132.295 52.255 133.205 ;
        RECT 52.505 132.525 56.405 133.205 ;
        RECT 55.475 132.295 56.405 132.525 ;
        RECT 57.335 132.425 58.705 133.205 ;
        RECT 58.715 132.395 61.465 133.205 ;
        RECT 61.475 132.525 63.305 133.205 ;
        RECT 63.515 132.385 65.445 133.205 ;
        RECT 66.075 132.395 67.905 133.205 ;
        RECT 68.060 133.175 68.230 133.395 ;
        RECT 69.900 133.225 70.070 133.415 ;
        RECT 72.655 133.225 72.825 133.395 ;
        RECT 72.655 133.205 72.805 133.225 ;
        RECT 74.035 133.205 74.205 133.395 ;
        RECT 76.980 133.225 77.150 133.415 ;
        RECT 84.155 133.205 84.325 133.395 ;
        RECT 86.915 133.225 87.085 133.415 ;
        RECT 88.755 133.225 88.925 133.415 ;
        RECT 89.675 133.205 89.845 133.395 ;
        RECT 90.135 133.225 90.305 133.415 ;
        RECT 90.650 133.255 90.770 133.365 ;
        RECT 92.435 133.225 92.605 133.415 ;
        RECT 92.895 133.250 93.055 133.360 ;
        RECT 93.815 133.225 93.985 133.415 ;
        RECT 95.195 133.225 95.365 133.395 ;
        RECT 95.655 133.225 95.825 133.415 ;
        RECT 97.035 133.225 97.205 133.415 ;
        RECT 99.795 133.225 99.965 133.395 ;
        RECT 100.715 133.365 100.885 133.415 ;
        RECT 100.715 133.255 100.890 133.365 ;
        RECT 100.715 133.225 100.885 133.255 ;
        RECT 90.155 133.205 90.305 133.225 ;
        RECT 95.195 133.205 95.345 133.225 ;
        RECT 69.720 133.175 70.665 133.205 ;
        RECT 67.915 132.495 70.665 133.175 ;
        RECT 63.515 132.295 64.465 132.385 ;
        RECT 69.720 132.295 70.665 132.495 ;
        RECT 70.875 132.385 72.805 133.205 ;
        RECT 72.975 132.395 74.345 133.205 ;
        RECT 70.875 132.295 71.825 132.385 ;
        RECT 74.365 132.335 74.795 133.120 ;
        RECT 75.185 132.525 84.465 133.205 ;
        RECT 75.185 132.405 77.520 132.525 ;
        RECT 75.185 132.295 76.105 132.405 ;
        RECT 82.185 132.305 83.105 132.525 ;
        RECT 84.475 132.395 89.985 133.205 ;
        RECT 90.155 132.385 92.085 133.205 ;
        RECT 91.135 132.295 92.085 132.385 ;
        RECT 93.415 132.385 95.345 133.205 ;
        RECT 95.675 133.205 95.825 133.225 ;
        RECT 99.795 133.205 99.945 133.225 ;
        RECT 104.395 133.205 104.565 133.395 ;
        RECT 104.855 133.205 105.025 133.395 ;
        RECT 106.235 133.225 106.405 133.415 ;
        RECT 106.695 133.250 106.855 133.360 ;
        RECT 107.155 133.205 107.325 133.395 ;
        RECT 111.755 133.205 111.925 133.415 ;
        RECT 113.135 133.205 113.305 133.415 ;
        RECT 95.675 132.385 97.605 133.205 ;
        RECT 93.415 132.295 94.365 132.385 ;
        RECT 96.655 132.295 97.605 132.385 ;
        RECT 98.015 132.385 99.945 133.205 ;
        RECT 98.015 132.295 98.965 132.385 ;
        RECT 100.125 132.335 100.555 133.120 ;
        RECT 101.035 132.395 104.705 133.205 ;
        RECT 104.725 132.295 106.075 133.205 ;
        RECT 107.015 132.425 108.385 133.205 ;
        RECT 108.395 132.395 112.065 133.205 ;
        RECT 112.075 132.395 113.445 133.205 ;
      LAYER nwell ;
        RECT 11.140 129.175 113.640 132.005 ;
      LAYER pwell ;
        RECT 11.335 127.975 12.705 128.785 ;
        RECT 12.715 127.975 16.385 128.785 ;
        RECT 16.405 127.975 17.755 128.885 ;
        RECT 23.975 128.795 24.925 128.885 ;
        RECT 17.775 127.975 19.145 128.785 ;
        RECT 19.155 127.975 20.525 128.755 ;
        RECT 21.455 127.975 22.825 128.755 ;
        RECT 22.995 127.975 24.925 128.795 ;
        RECT 26.495 128.655 27.415 128.875 ;
        RECT 33.495 128.775 34.415 128.885 ;
        RECT 32.080 128.655 34.415 128.775 ;
        RECT 25.135 127.975 34.415 128.655 ;
        RECT 35.725 128.060 36.155 128.845 ;
        RECT 36.185 127.975 37.535 128.885 ;
        RECT 38.695 128.795 39.645 128.885 ;
        RECT 40.995 128.795 41.945 128.885 ;
        RECT 37.715 127.975 39.645 128.795 ;
        RECT 40.015 127.975 41.945 128.795 ;
        RECT 42.165 127.975 44.905 128.655 ;
        RECT 45.055 127.975 47.665 128.885 ;
        RECT 48.135 127.975 49.965 128.785 ;
        RECT 49.985 127.975 51.335 128.885 ;
        RECT 51.725 128.775 52.645 128.885 ;
        RECT 51.725 128.655 54.060 128.775 ;
        RECT 58.725 128.655 59.645 128.875 ;
        RECT 51.725 127.975 61.005 128.655 ;
        RECT 61.485 128.060 61.915 128.845 ;
        RECT 68.595 128.795 69.545 128.885 ;
        RECT 61.935 127.975 63.305 128.785 ;
        RECT 63.315 127.975 66.055 128.655 ;
        RECT 66.075 127.975 67.445 128.785 ;
        RECT 67.615 127.975 69.545 128.795 ;
        RECT 69.955 128.795 70.905 128.885 ;
        RECT 69.955 127.975 71.885 128.795 ;
        RECT 75.255 128.655 76.185 128.885 ;
        RECT 72.285 127.975 76.185 128.655 ;
        RECT 76.195 127.975 77.565 128.785 ;
        RECT 77.585 127.975 78.935 128.885 ;
        RECT 78.965 127.975 80.315 128.885 ;
        RECT 86.075 128.795 87.025 128.885 ;
        RECT 81.255 127.975 82.620 128.655 ;
        RECT 83.095 127.975 84.925 128.785 ;
        RECT 85.095 127.975 87.025 128.795 ;
        RECT 87.245 128.060 87.675 128.845 ;
        RECT 101.015 128.655 101.945 128.885 ;
        RECT 87.695 127.975 96.800 128.655 ;
        RECT 98.045 127.975 101.945 128.655 ;
        RECT 102.325 128.775 103.245 128.885 ;
        RECT 102.325 128.655 104.660 128.775 ;
        RECT 109.325 128.655 110.245 128.875 ;
        RECT 102.325 127.975 111.605 128.655 ;
        RECT 112.075 127.975 113.445 128.785 ;
        RECT 11.475 127.765 11.645 127.975 ;
        RECT 13.775 127.765 13.945 127.955 ;
        RECT 14.235 127.765 14.405 127.955 ;
        RECT 15.615 127.765 15.785 127.955 ;
        RECT 16.075 127.785 16.245 127.975 ;
        RECT 17.270 127.765 17.440 127.955 ;
        RECT 17.455 127.785 17.625 127.975 ;
        RECT 18.835 127.785 19.005 127.975 ;
        RECT 19.295 127.785 19.465 127.975 ;
        RECT 21.135 127.925 21.295 127.930 ;
        RECT 21.135 127.820 21.310 127.925 ;
        RECT 21.190 127.815 21.310 127.820 ;
        RECT 21.595 127.765 21.765 127.975 ;
        RECT 22.995 127.955 23.145 127.975 ;
        RECT 22.975 127.785 23.145 127.955 ;
        RECT 24.355 127.785 24.525 127.955 ;
        RECT 24.815 127.765 24.985 127.955 ;
        RECT 25.275 127.785 25.445 127.975 ;
        RECT 26.470 127.765 26.640 127.955 ;
        RECT 30.390 127.815 30.510 127.925 ;
        RECT 34.200 127.765 34.370 127.955 ;
        RECT 35.395 127.820 35.555 127.930 ;
        RECT 36.315 127.785 36.485 127.975 ;
        RECT 37.715 127.955 37.865 127.975 ;
        RECT 40.015 127.955 40.165 127.975 ;
        RECT 37.695 127.785 37.865 127.955 ;
        RECT 38.340 127.765 38.510 127.955 ;
        RECT 39.995 127.785 40.165 127.955 ;
        RECT 44.595 127.785 44.765 127.975 ;
        RECT 47.350 127.785 47.520 127.975 ;
        RECT 47.815 127.925 47.985 127.955 ;
        RECT 47.815 127.815 47.990 127.925 ;
        RECT 48.330 127.815 48.450 127.925 ;
        RECT 49.250 127.815 49.370 127.925 ;
        RECT 47.815 127.765 47.985 127.815 ;
        RECT 49.655 127.765 49.825 127.975 ;
        RECT 50.115 127.785 50.285 127.975 ;
        RECT 54.440 127.765 54.610 127.955 ;
        RECT 55.175 127.765 55.345 127.955 ;
        RECT 57.015 127.810 57.175 127.920 ;
        RECT 60.695 127.765 60.865 127.975 ;
        RECT 61.210 127.815 61.330 127.925 ;
        RECT 62.995 127.785 63.165 127.975 ;
        RECT 63.455 127.785 63.625 127.975 ;
        RECT 66.215 127.765 66.385 127.955 ;
        RECT 67.135 127.785 67.305 127.975 ;
        RECT 67.615 127.955 67.765 127.975 ;
        RECT 71.735 127.955 71.885 127.975 ;
        RECT 67.595 127.785 67.765 127.955 ;
        RECT 68.515 127.785 68.685 127.955 ;
        RECT 71.735 127.785 71.905 127.955 ;
        RECT 68.515 127.765 68.665 127.785 ;
        RECT 72.380 127.765 72.550 127.955 ;
        RECT 74.035 127.765 74.205 127.955 ;
        RECT 75.600 127.785 75.770 127.975 ;
        RECT 77.255 127.785 77.425 127.975 ;
        RECT 77.715 127.785 77.885 127.975 ;
        RECT 80.015 127.785 80.185 127.975 ;
        RECT 80.935 127.820 81.095 127.930 ;
        RECT 82.775 127.785 82.945 127.955 ;
        RECT 83.695 127.765 83.865 127.955 ;
        RECT 84.615 127.785 84.785 127.975 ;
        RECT 85.095 127.955 85.245 127.975 ;
        RECT 85.075 127.785 85.245 127.955 ;
        RECT 85.535 127.765 85.705 127.955 ;
        RECT 87.835 127.785 88.005 127.975 ;
        RECT 89.400 127.765 89.570 127.955 ;
        RECT 90.135 127.765 90.305 127.955 ;
        RECT 91.515 127.785 91.685 127.955 ;
        RECT 91.535 127.765 91.685 127.785 ;
        RECT 97.220 127.765 97.390 127.955 ;
        RECT 97.495 127.820 97.655 127.930 ;
        RECT 98.415 127.810 98.575 127.920 ;
        RECT 98.875 127.765 99.045 127.955 ;
        RECT 100.770 127.815 100.890 127.925 ;
        RECT 101.360 127.785 101.530 127.975 ;
        RECT 110.375 127.765 110.545 127.955 ;
        RECT 111.295 127.785 111.465 127.975 ;
        RECT 111.755 127.925 111.925 127.955 ;
        RECT 111.755 127.815 111.930 127.925 ;
        RECT 111.755 127.765 111.925 127.815 ;
        RECT 113.135 127.765 113.305 127.975 ;
        RECT 11.335 126.955 12.705 127.765 ;
        RECT 12.725 126.855 14.075 127.765 ;
        RECT 14.105 126.855 15.455 127.765 ;
        RECT 15.475 126.985 16.845 127.765 ;
        RECT 16.855 127.085 20.755 127.765 ;
        RECT 16.855 126.855 17.785 127.085 ;
        RECT 21.465 126.855 22.815 127.765 ;
        RECT 22.845 126.895 23.275 127.680 ;
        RECT 23.295 127.085 24.250 127.765 ;
        RECT 24.675 126.985 26.045 127.765 ;
        RECT 26.055 127.085 29.955 127.765 ;
        RECT 30.885 127.085 34.785 127.765 ;
        RECT 35.025 127.085 38.925 127.765 ;
        RECT 39.020 127.085 48.125 127.765 ;
        RECT 26.055 126.855 26.985 127.085 ;
        RECT 33.855 126.855 34.785 127.085 ;
        RECT 37.995 126.855 38.925 127.085 ;
        RECT 48.605 126.895 49.035 127.680 ;
        RECT 49.525 126.855 50.875 127.765 ;
        RECT 51.125 127.085 55.025 127.765 ;
        RECT 54.095 126.855 55.025 127.085 ;
        RECT 55.035 126.985 56.405 127.765 ;
        RECT 57.335 126.955 61.005 127.765 ;
        RECT 61.015 126.955 66.525 127.765 ;
        RECT 66.735 126.945 68.665 127.765 ;
        RECT 69.065 127.085 72.965 127.765 ;
        RECT 66.735 126.855 67.685 126.945 ;
        RECT 72.035 126.855 72.965 127.085 ;
        RECT 72.975 126.955 74.345 127.765 ;
        RECT 74.365 126.895 74.795 127.680 ;
        RECT 74.900 127.085 84.005 127.765 ;
        RECT 84.015 126.955 85.845 127.765 ;
        RECT 86.085 127.085 89.985 127.765 ;
        RECT 89.055 126.855 89.985 127.085 ;
        RECT 90.005 126.855 91.355 127.765 ;
        RECT 91.535 126.945 93.465 127.765 ;
        RECT 93.905 127.085 97.805 127.765 ;
        RECT 92.515 126.855 93.465 126.945 ;
        RECT 96.875 126.855 97.805 127.085 ;
        RECT 98.745 126.855 100.095 127.765 ;
        RECT 100.125 126.895 100.555 127.680 ;
        RECT 101.405 127.085 110.685 127.765 ;
        RECT 101.405 126.965 103.740 127.085 ;
        RECT 101.405 126.855 102.325 126.965 ;
        RECT 108.405 126.865 109.325 127.085 ;
        RECT 110.695 126.955 112.065 127.765 ;
        RECT 112.075 126.955 113.445 127.765 ;
      LAYER nwell ;
        RECT 11.140 123.735 113.640 126.565 ;
      LAYER pwell ;
        RECT 11.335 122.535 12.705 123.345 ;
        RECT 13.545 123.335 14.465 123.445 ;
        RECT 13.545 123.215 15.880 123.335 ;
        RECT 20.545 123.215 21.465 123.435 ;
        RECT 34.555 123.355 35.505 123.445 ;
        RECT 13.545 122.535 22.825 123.215 ;
        RECT 23.840 122.535 32.945 123.215 ;
        RECT 33.575 122.535 35.505 123.355 ;
        RECT 35.725 122.620 36.155 123.405 ;
        RECT 37.115 122.535 48.125 123.445 ;
        RECT 48.505 123.335 49.425 123.445 ;
        RECT 48.505 123.215 50.840 123.335 ;
        RECT 55.505 123.215 56.425 123.435 ;
        RECT 48.505 122.535 57.785 123.215 ;
        RECT 57.795 122.535 61.465 123.345 ;
        RECT 61.485 122.620 61.915 123.405 ;
        RECT 61.935 122.535 64.685 123.345 ;
        RECT 64.705 122.535 66.055 123.445 ;
        RECT 69.275 123.215 70.205 123.445 ;
        RECT 66.305 122.535 70.205 123.215 ;
        RECT 70.215 122.535 72.045 123.345 ;
        RECT 72.425 123.335 73.345 123.445 ;
        RECT 72.425 123.215 74.760 123.335 ;
        RECT 79.425 123.215 80.345 123.435 ;
        RECT 84.915 123.215 85.845 123.445 ;
        RECT 72.425 122.535 81.705 123.215 ;
        RECT 81.945 122.535 85.845 123.215 ;
        RECT 85.855 122.535 87.225 123.345 ;
        RECT 87.245 122.620 87.675 123.405 ;
        RECT 88.525 123.335 89.445 123.445 ;
        RECT 88.525 123.215 90.860 123.335 ;
        RECT 95.525 123.215 96.445 123.435 ;
        RECT 88.525 122.535 97.805 123.215 ;
        RECT 97.815 122.535 99.185 123.315 ;
        RECT 99.195 122.535 100.565 123.345 ;
        RECT 103.775 123.215 104.705 123.445 ;
        RECT 100.805 122.535 104.705 123.215 ;
        RECT 104.715 122.535 106.085 123.345 ;
        RECT 106.095 122.535 107.465 123.315 ;
        RECT 108.395 122.535 112.065 123.345 ;
        RECT 112.075 122.535 113.445 123.345 ;
        RECT 11.475 122.325 11.645 122.535 ;
        RECT 12.910 122.375 13.030 122.485 ;
        RECT 22.055 122.325 22.225 122.515 ;
        RECT 22.515 122.485 22.685 122.535 ;
        RECT 22.515 122.375 22.690 122.485 ;
        RECT 22.515 122.345 22.685 122.375 ;
        RECT 23.435 122.325 23.605 122.515 ;
        RECT 32.635 122.345 32.805 122.535 ;
        RECT 33.575 122.515 33.725 122.535 ;
        RECT 33.150 122.375 33.270 122.485 ;
        RECT 33.555 122.345 33.725 122.515 ;
        RECT 36.775 122.380 36.935 122.490 ;
        RECT 42.295 122.325 42.465 122.515 ;
        RECT 46.160 122.325 46.330 122.515 ;
        RECT 46.895 122.325 47.065 122.515 ;
        RECT 47.810 122.345 47.980 122.535 ;
        RECT 48.330 122.375 48.450 122.485 ;
        RECT 50.575 122.325 50.745 122.515 ;
        RECT 51.310 122.325 51.480 122.515 ;
        RECT 57.475 122.345 57.645 122.535 ;
        RECT 58.580 122.325 58.750 122.515 ;
        RECT 59.315 122.325 59.485 122.515 ;
        RECT 60.695 122.325 60.865 122.515 ;
        RECT 61.155 122.345 61.325 122.535 ;
        RECT 64.375 122.345 64.545 122.535 ;
        RECT 64.835 122.345 65.005 122.535 ;
        RECT 69.620 122.345 69.790 122.535 ;
        RECT 71.275 122.325 71.445 122.515 ;
        RECT 71.735 122.345 71.905 122.535 ;
        RECT 72.655 122.325 72.825 122.515 ;
        RECT 74.035 122.325 74.205 122.515 ;
        RECT 74.955 122.325 75.125 122.515 ;
        RECT 81.395 122.345 81.565 122.535 ;
        RECT 85.260 122.345 85.430 122.535 ;
        RECT 85.535 122.325 85.705 122.515 ;
        RECT 85.995 122.325 86.165 122.515 ;
        RECT 86.915 122.345 87.085 122.535 ;
        RECT 87.890 122.375 88.010 122.485 ;
        RECT 88.295 122.325 88.465 122.515 ;
        RECT 89.675 122.325 89.845 122.515 ;
        RECT 90.135 122.325 90.305 122.515 ;
        RECT 94.920 122.325 95.090 122.515 ;
        RECT 95.710 122.375 95.830 122.485 ;
        RECT 97.495 122.345 97.665 122.535 ;
        RECT 98.875 122.345 99.045 122.535 ;
        RECT 99.520 122.325 99.690 122.515 ;
        RECT 100.255 122.345 100.425 122.535 ;
        RECT 104.120 122.345 104.290 122.535 ;
        RECT 105.775 122.345 105.945 122.535 ;
        RECT 106.235 122.345 106.405 122.535 ;
        RECT 108.075 122.380 108.235 122.490 ;
        RECT 109.915 122.325 110.085 122.515 ;
        RECT 111.755 122.325 111.925 122.535 ;
        RECT 113.135 122.325 113.305 122.535 ;
        RECT 11.335 121.515 12.705 122.325 ;
        RECT 13.085 121.645 22.365 122.325 ;
        RECT 13.085 121.525 15.420 121.645 ;
        RECT 13.085 121.415 14.005 121.525 ;
        RECT 20.085 121.425 21.005 121.645 ;
        RECT 22.845 121.455 23.275 122.240 ;
        RECT 23.295 121.645 32.575 122.325 ;
        RECT 24.655 121.425 25.575 121.645 ;
        RECT 30.240 121.525 32.575 121.645 ;
        RECT 31.655 121.415 32.575 121.525 ;
        RECT 33.325 121.645 42.605 122.325 ;
        RECT 42.845 121.645 46.745 122.325 ;
        RECT 33.325 121.525 35.660 121.645 ;
        RECT 33.325 121.415 34.245 121.525 ;
        RECT 40.325 121.425 41.245 121.645 ;
        RECT 45.815 121.415 46.745 121.645 ;
        RECT 46.755 121.545 48.125 122.325 ;
        RECT 48.605 121.455 49.035 122.240 ;
        RECT 49.055 121.515 50.885 122.325 ;
        RECT 50.895 121.645 54.795 122.325 ;
        RECT 55.265 121.645 59.165 122.325 ;
        RECT 50.895 121.415 51.825 121.645 ;
        RECT 58.235 121.415 59.165 121.645 ;
        RECT 59.175 121.545 60.545 122.325 ;
        RECT 60.565 121.415 61.915 122.325 ;
        RECT 62.305 121.645 71.585 122.325 ;
        RECT 62.305 121.525 64.640 121.645 ;
        RECT 62.305 121.415 63.225 121.525 ;
        RECT 69.305 121.425 70.225 121.645 ;
        RECT 71.595 121.545 72.965 122.325 ;
        RECT 72.975 121.545 74.345 122.325 ;
        RECT 74.365 121.455 74.795 122.240 ;
        RECT 74.825 121.415 76.175 122.325 ;
        RECT 76.565 121.645 85.845 122.325 ;
        RECT 76.565 121.525 78.900 121.645 ;
        RECT 76.565 121.415 77.485 121.525 ;
        RECT 83.565 121.425 84.485 121.645 ;
        RECT 85.865 121.415 87.215 122.325 ;
        RECT 87.235 121.545 88.605 122.325 ;
        RECT 88.615 121.545 89.985 122.325 ;
        RECT 90.005 121.415 91.355 122.325 ;
        RECT 91.605 121.645 95.505 122.325 ;
        RECT 96.205 121.645 100.105 122.325 ;
        RECT 94.575 121.415 95.505 121.645 ;
        RECT 99.175 121.415 100.105 121.645 ;
        RECT 100.125 121.455 100.555 122.240 ;
        RECT 100.945 121.645 110.225 122.325 ;
        RECT 100.945 121.525 103.280 121.645 ;
        RECT 100.945 121.415 101.865 121.525 ;
        RECT 107.945 121.425 108.865 121.645 ;
        RECT 110.235 121.515 112.065 122.325 ;
        RECT 112.075 121.515 113.445 122.325 ;
      LAYER nwell ;
        RECT 11.140 118.295 113.640 121.125 ;
      LAYER pwell ;
        RECT 11.335 117.095 12.705 117.905 ;
        RECT 12.915 117.775 15.125 118.005 ;
        RECT 17.845 117.775 18.775 117.995 ;
        RECT 24.655 117.775 25.575 117.995 ;
        RECT 31.655 117.895 32.575 118.005 ;
        RECT 30.240 117.775 32.575 117.895 ;
        RECT 12.915 117.095 23.285 117.775 ;
        RECT 23.295 117.095 32.575 117.775 ;
        RECT 33.875 117.095 35.245 117.875 ;
        RECT 35.725 117.180 36.155 117.965 ;
        RECT 36.175 117.095 38.005 117.905 ;
        RECT 39.765 117.895 40.685 118.005 ;
        RECT 38.015 117.095 39.385 117.875 ;
        RECT 39.765 117.775 42.100 117.895 ;
        RECT 46.765 117.775 47.685 117.995 ;
        RECT 39.765 117.095 49.045 117.775 ;
        RECT 49.055 117.095 50.425 117.905 ;
        RECT 52.185 117.895 53.105 118.005 ;
        RECT 50.435 117.095 51.805 117.875 ;
        RECT 52.185 117.775 54.520 117.895 ;
        RECT 59.185 117.775 60.105 117.995 ;
        RECT 52.185 117.095 61.465 117.775 ;
        RECT 61.485 117.180 61.915 117.965 ;
        RECT 61.945 117.095 63.295 118.005 ;
        RECT 63.315 117.095 64.685 117.905 ;
        RECT 65.065 117.895 65.985 118.005 ;
        RECT 65.065 117.775 67.400 117.895 ;
        RECT 72.065 117.775 72.985 117.995 ;
        RECT 65.065 117.095 74.345 117.775 ;
        RECT 74.355 117.095 76.185 117.905 ;
        RECT 76.195 117.095 77.565 117.875 ;
        RECT 78.935 117.775 79.855 117.995 ;
        RECT 85.935 117.895 86.855 118.005 ;
        RECT 84.520 117.775 86.855 117.895 ;
        RECT 77.575 117.095 86.855 117.775 ;
        RECT 87.245 117.180 87.675 117.965 ;
        RECT 88.155 117.095 90.905 117.905 ;
        RECT 91.285 117.895 92.205 118.005 ;
        RECT 91.285 117.775 93.620 117.895 ;
        RECT 98.285 117.775 99.205 117.995 ;
        RECT 91.285 117.095 100.565 117.775 ;
        RECT 101.035 117.095 103.785 117.905 ;
        RECT 103.805 117.095 105.155 118.005 ;
        RECT 105.175 117.095 106.545 117.875 ;
        RECT 106.555 117.095 112.065 117.905 ;
        RECT 112.075 117.095 113.445 117.905 ;
        RECT 11.475 116.885 11.645 117.095 ;
        RECT 15.155 116.885 15.325 117.075 ;
        RECT 15.615 116.885 15.785 117.075 ;
        RECT 17.270 116.885 17.440 117.075 ;
        RECT 22.515 116.885 22.685 117.075 ;
        RECT 22.975 116.905 23.145 117.095 ;
        RECT 23.435 116.905 23.605 117.095 ;
        RECT 24.355 116.885 24.525 117.075 ;
        RECT 29.875 116.885 30.045 117.075 ;
        RECT 31.255 116.885 31.425 117.075 ;
        RECT 31.770 116.935 31.890 117.045 ;
        RECT 33.555 116.940 33.715 117.050 ;
        RECT 34.935 116.905 35.105 117.095 ;
        RECT 35.450 116.935 35.570 117.045 ;
        RECT 37.235 116.885 37.405 117.075 ;
        RECT 37.695 116.905 37.865 117.095 ;
        RECT 38.155 116.905 38.325 117.095 ;
        RECT 42.755 116.885 42.925 117.075 ;
        RECT 44.135 116.885 44.305 117.075 ;
        RECT 44.650 116.935 44.770 117.045 ;
        RECT 48.275 116.885 48.445 117.075 ;
        RECT 48.735 116.905 48.905 117.095 ;
        RECT 49.195 116.885 49.365 117.075 ;
        RECT 50.115 116.905 50.285 117.095 ;
        RECT 51.495 116.905 51.665 117.095 ;
        RECT 59.315 116.930 59.475 117.040 ;
        RECT 61.155 116.905 61.325 117.095 ;
        RECT 62.995 116.885 63.165 117.095 ;
        RECT 64.375 116.905 64.545 117.095 ;
        RECT 68.515 116.885 68.685 117.075 ;
        RECT 74.035 116.885 74.205 117.095 ;
        RECT 75.415 116.930 75.575 117.040 ;
        RECT 75.875 116.905 76.045 117.095 ;
        RECT 76.335 116.905 76.505 117.095 ;
        RECT 77.715 116.905 77.885 117.095 ;
        RECT 79.095 116.885 79.265 117.075 ;
        RECT 84.615 116.885 84.785 117.075 ;
        RECT 87.890 116.935 88.010 117.045 ;
        RECT 90.135 116.885 90.305 117.075 ;
        RECT 90.595 116.905 90.765 117.095 ;
        RECT 95.655 116.885 95.825 117.075 ;
        RECT 96.115 116.885 96.285 117.075 ;
        RECT 99.795 116.885 99.965 117.075 ;
        RECT 100.255 116.905 100.425 117.095 ;
        RECT 100.770 116.935 100.890 117.045 ;
        RECT 103.475 116.905 103.645 117.095 ;
        RECT 103.935 116.885 104.105 117.095 ;
        RECT 105.315 116.885 105.485 117.095 ;
        RECT 105.775 116.885 105.945 117.075 ;
        RECT 107.615 116.930 107.775 117.040 ;
        RECT 108.995 116.885 109.165 117.075 ;
        RECT 111.755 116.885 111.925 117.095 ;
        RECT 113.135 116.885 113.305 117.095 ;
        RECT 11.335 116.075 12.705 116.885 ;
        RECT 12.715 116.075 15.465 116.885 ;
        RECT 15.475 116.105 16.845 116.885 ;
        RECT 16.855 116.205 20.755 116.885 ;
        RECT 16.855 115.975 17.785 116.205 ;
        RECT 20.995 116.075 22.825 116.885 ;
        RECT 22.845 116.015 23.275 116.800 ;
        RECT 23.295 116.075 24.665 116.885 ;
        RECT 24.675 116.075 30.185 116.885 ;
        RECT 30.205 115.975 31.555 116.885 ;
        RECT 32.035 116.075 37.545 116.885 ;
        RECT 37.555 116.075 43.065 116.885 ;
        RECT 43.085 115.975 44.435 116.885 ;
        RECT 44.915 116.075 48.585 116.885 ;
        RECT 48.605 116.015 49.035 116.800 ;
        RECT 49.055 116.205 58.335 116.885 ;
        RECT 50.415 115.985 51.335 116.205 ;
        RECT 56.000 116.085 58.335 116.205 ;
        RECT 57.415 115.975 58.335 116.085 ;
        RECT 59.635 116.075 63.305 116.885 ;
        RECT 63.315 116.075 68.825 116.885 ;
        RECT 68.835 116.075 74.345 116.885 ;
        RECT 74.365 116.015 74.795 116.800 ;
        RECT 75.735 116.075 79.405 116.885 ;
        RECT 79.415 116.075 84.925 116.885 ;
        RECT 84.935 116.075 90.445 116.885 ;
        RECT 90.455 116.075 95.965 116.885 ;
        RECT 95.975 116.105 97.345 116.885 ;
        RECT 97.355 116.075 100.105 116.885 ;
        RECT 100.125 116.015 100.555 116.800 ;
        RECT 100.575 116.075 104.245 116.885 ;
        RECT 104.255 116.105 105.625 116.885 ;
        RECT 105.645 115.975 106.995 116.885 ;
        RECT 107.935 116.105 109.305 116.885 ;
        RECT 109.315 116.075 112.065 116.885 ;
        RECT 112.075 116.075 113.445 116.885 ;
      LAYER nwell ;
        RECT 11.140 112.855 113.640 115.685 ;
      LAYER pwell ;
        RECT 11.335 111.655 12.705 112.465 ;
        RECT 12.715 111.655 14.085 112.465 ;
        RECT 14.295 112.335 16.505 112.565 ;
        RECT 19.225 112.335 20.155 112.555 ;
        RECT 14.295 111.655 24.665 112.335 ;
        RECT 24.675 111.655 27.425 112.465 ;
        RECT 27.445 111.655 28.795 112.565 ;
        RECT 28.815 111.655 30.185 112.465 ;
        RECT 30.195 111.655 35.705 112.465 ;
        RECT 35.725 111.740 36.155 112.525 ;
        RECT 36.175 111.655 37.545 112.435 ;
        RECT 38.015 111.655 39.845 112.465 ;
        RECT 39.855 111.655 41.225 112.435 ;
        RECT 41.235 111.655 43.985 112.465 ;
        RECT 43.995 111.655 45.365 112.435 ;
        RECT 46.295 111.655 49.965 112.465 ;
        RECT 49.985 111.655 51.335 112.565 ;
        RECT 51.355 111.655 53.965 112.565 ;
        RECT 54.115 111.655 56.865 112.465 ;
        RECT 56.875 111.655 58.245 112.435 ;
        RECT 58.255 111.655 60.085 112.465 ;
        RECT 60.095 111.655 61.465 112.435 ;
        RECT 61.485 111.740 61.915 112.525 ;
        RECT 62.855 111.655 66.525 112.465 ;
        RECT 66.545 111.655 67.895 112.565 ;
        RECT 67.915 111.655 69.285 112.435 ;
        RECT 69.305 111.655 70.655 112.565 ;
        RECT 70.675 111.655 73.285 112.565 ;
        RECT 73.895 111.655 77.565 112.465 ;
        RECT 77.575 111.655 83.085 112.465 ;
        RECT 83.095 111.655 84.465 112.435 ;
        RECT 84.475 111.655 87.225 112.465 ;
        RECT 87.245 111.740 87.675 112.525 ;
        RECT 88.155 111.655 89.525 112.435 ;
        RECT 89.995 111.655 93.665 112.465 ;
        RECT 93.675 111.655 95.045 112.435 ;
        RECT 95.975 111.655 97.345 112.435 ;
        RECT 97.355 111.655 98.725 112.435 ;
        RECT 98.735 111.655 101.485 112.465 ;
        RECT 106.005 112.335 106.935 112.555 ;
        RECT 109.655 112.335 111.865 112.565 ;
        RECT 101.495 111.655 111.865 112.335 ;
        RECT 112.075 111.655 113.445 112.465 ;
        RECT 11.475 111.445 11.645 111.655 ;
        RECT 13.775 111.465 13.945 111.655 ;
        RECT 17.915 111.445 18.085 111.635 ;
        RECT 19.295 111.445 19.465 111.635 ;
        RECT 21.135 111.445 21.305 111.635 ;
        RECT 22.515 111.445 22.685 111.635 ;
        RECT 24.355 111.445 24.525 111.655 ;
        RECT 25.735 111.445 25.905 111.635 ;
        RECT 26.195 111.445 26.365 111.635 ;
        RECT 27.115 111.465 27.285 111.655 ;
        RECT 28.495 111.465 28.665 111.655 ;
        RECT 29.875 111.465 30.045 111.655 ;
        RECT 35.395 111.465 35.565 111.655 ;
        RECT 37.235 111.465 37.405 111.655 ;
        RECT 37.695 111.605 37.865 111.635 ;
        RECT 37.695 111.495 37.870 111.605 ;
        RECT 37.695 111.445 37.865 111.495 ;
        RECT 39.535 111.465 39.705 111.655 ;
        RECT 40.915 111.465 41.085 111.655 ;
        RECT 43.675 111.465 43.845 111.655 ;
        RECT 44.135 111.465 44.305 111.655 ;
        RECT 45.975 111.500 46.135 111.610 ;
        RECT 48.275 111.445 48.445 111.635 ;
        RECT 49.195 111.445 49.365 111.635 ;
        RECT 49.655 111.465 49.825 111.655 ;
        RECT 50.115 111.465 50.285 111.655 ;
        RECT 51.035 111.490 51.195 111.600 ;
        RECT 51.500 111.465 51.670 111.655 ;
        RECT 56.555 111.465 56.725 111.655 ;
        RECT 57.015 111.465 57.185 111.655 ;
        RECT 59.775 111.465 59.945 111.655 ;
        RECT 60.235 111.465 60.405 111.655 ;
        RECT 61.615 111.445 61.785 111.635 ;
        RECT 62.535 111.490 62.695 111.610 ;
        RECT 66.215 111.465 66.385 111.655 ;
        RECT 67.595 111.465 67.765 111.655 ;
        RECT 68.975 111.465 69.145 111.655 ;
        RECT 70.355 111.465 70.525 111.655 ;
        RECT 70.820 111.465 70.990 111.655 ;
        RECT 73.115 111.445 73.285 111.635 ;
        RECT 73.630 111.495 73.750 111.605 ;
        RECT 74.035 111.490 74.195 111.600 ;
        RECT 75.875 111.445 76.045 111.635 ;
        RECT 76.390 111.495 76.510 111.605 ;
        RECT 76.795 111.445 76.965 111.635 ;
        RECT 77.255 111.465 77.425 111.655 ;
        RECT 82.775 111.465 82.945 111.655 ;
        RECT 83.235 111.465 83.405 111.655 ;
        RECT 86.915 111.465 87.085 111.655 ;
        RECT 87.890 111.495 88.010 111.605 ;
        RECT 88.295 111.445 88.465 111.655 ;
        RECT 89.730 111.495 89.850 111.605 ;
        RECT 93.355 111.465 93.525 111.655 ;
        RECT 93.815 111.465 93.985 111.655 ;
        RECT 95.655 111.500 95.815 111.610 ;
        RECT 96.115 111.465 96.285 111.655 ;
        RECT 98.415 111.465 98.585 111.655 ;
        RECT 98.875 111.445 99.045 111.635 ;
        RECT 99.795 111.490 99.955 111.600 ;
        RECT 101.175 111.465 101.345 111.655 ;
        RECT 101.635 111.445 101.805 111.655 ;
        RECT 113.135 111.445 113.305 111.655 ;
        RECT 11.335 110.635 12.705 111.445 ;
        RECT 12.715 110.635 18.225 111.445 ;
        RECT 18.245 110.535 19.595 111.445 ;
        RECT 19.615 110.635 21.445 111.445 ;
        RECT 21.455 110.665 22.825 111.445 ;
        RECT 22.845 110.575 23.275 111.360 ;
        RECT 23.295 110.665 24.665 111.445 ;
        RECT 24.675 110.665 26.045 111.445 ;
        RECT 26.055 110.665 27.425 111.445 ;
        RECT 27.635 110.765 38.005 111.445 ;
        RECT 38.215 110.765 48.585 111.445 ;
        RECT 27.635 110.535 29.845 110.765 ;
        RECT 32.565 110.545 33.495 110.765 ;
        RECT 38.215 110.535 40.425 110.765 ;
        RECT 43.145 110.545 44.075 110.765 ;
        RECT 48.605 110.575 49.035 111.360 ;
        RECT 49.055 110.665 50.425 111.445 ;
        RECT 51.555 110.765 61.925 111.445 ;
        RECT 63.055 110.765 73.425 111.445 ;
        RECT 51.555 110.535 53.765 110.765 ;
        RECT 56.485 110.545 57.415 110.765 ;
        RECT 63.055 110.535 65.265 110.765 ;
        RECT 67.985 110.545 68.915 110.765 ;
        RECT 74.365 110.575 74.795 111.360 ;
        RECT 74.815 110.665 76.185 111.445 ;
        RECT 76.655 110.665 78.025 111.445 ;
        RECT 78.235 110.765 88.605 111.445 ;
        RECT 88.815 110.765 99.185 111.445 ;
        RECT 78.235 110.535 80.445 110.765 ;
        RECT 83.165 110.545 84.095 110.765 ;
        RECT 88.815 110.535 91.025 110.765 ;
        RECT 93.745 110.545 94.675 110.765 ;
        RECT 100.125 110.575 100.555 111.360 ;
        RECT 101.495 110.765 111.865 111.445 ;
        RECT 106.005 110.545 106.935 110.765 ;
        RECT 109.655 110.535 111.865 110.765 ;
        RECT 112.075 110.635 113.445 111.445 ;
      LAYER nwell ;
        RECT 11.140 107.415 113.640 110.245 ;
      LAYER pwell ;
        RECT 11.335 106.215 12.705 107.025 ;
        RECT 13.185 106.215 14.535 107.125 ;
        RECT 14.755 106.895 16.965 107.125 ;
        RECT 19.685 106.895 20.615 107.115 ;
        RECT 29.645 106.895 30.575 107.115 ;
        RECT 33.295 106.895 35.505 107.125 ;
        RECT 14.755 106.215 25.125 106.895 ;
        RECT 25.135 106.215 35.505 106.895 ;
        RECT 35.725 106.300 36.155 107.085 ;
        RECT 36.185 106.215 37.535 107.125 ;
        RECT 38.025 106.215 39.375 107.125 ;
        RECT 39.855 106.215 43.525 107.025 ;
        RECT 43.545 106.215 44.895 107.125 ;
        RECT 45.115 106.895 47.325 107.125 ;
        RECT 50.045 106.895 50.975 107.115 ;
        RECT 45.115 106.215 55.485 106.895 ;
        RECT 55.505 106.215 56.855 107.125 ;
        RECT 57.345 106.215 58.695 107.125 ;
        RECT 58.715 106.215 61.465 107.025 ;
        RECT 61.485 106.300 61.915 107.085 ;
        RECT 62.135 106.895 64.345 107.125 ;
        RECT 67.065 106.895 67.995 107.115 ;
        RECT 73.635 106.895 75.845 107.125 ;
        RECT 78.565 106.895 79.495 107.115 ;
        RECT 62.135 106.215 72.505 106.895 ;
        RECT 73.635 106.215 84.005 106.895 ;
        RECT 84.025 106.215 85.375 107.125 ;
        RECT 85.865 106.215 87.215 107.125 ;
        RECT 87.245 106.300 87.675 107.085 ;
        RECT 87.895 106.895 90.105 107.125 ;
        RECT 92.825 106.895 93.755 107.115 ;
        RECT 103.705 106.895 104.635 107.115 ;
        RECT 107.355 106.895 109.565 107.125 ;
        RECT 87.895 106.215 98.265 106.895 ;
        RECT 99.195 106.215 109.565 106.895 ;
        RECT 110.695 106.215 112.065 106.995 ;
        RECT 112.075 106.215 113.445 107.025 ;
        RECT 11.475 106.005 11.645 106.215 ;
        RECT 12.910 106.055 13.030 106.165 ;
        RECT 14.235 106.025 14.405 106.215 ;
        RECT 15.615 106.005 15.785 106.195 ;
        RECT 21.135 106.005 21.305 106.195 ;
        RECT 22.515 106.005 22.685 106.195 ;
        RECT 24.815 106.025 24.985 106.215 ;
        RECT 25.275 106.025 25.445 106.215 ;
        RECT 33.555 106.005 33.725 106.195 ;
        RECT 35.395 106.005 35.565 106.195 ;
        RECT 37.235 106.005 37.405 106.215 ;
        RECT 37.750 106.055 37.870 106.165 ;
        RECT 39.075 106.025 39.245 106.215 ;
        RECT 39.590 106.055 39.710 106.165 ;
        RECT 42.755 106.005 42.925 106.195 ;
        RECT 43.215 106.025 43.385 106.215 ;
        RECT 44.595 106.025 44.765 106.215 ;
        RECT 48.275 106.005 48.445 106.195 ;
        RECT 50.115 106.005 50.285 106.195 ;
        RECT 55.175 106.025 55.345 106.215 ;
        RECT 55.635 106.005 55.805 106.195 ;
        RECT 56.555 106.025 56.725 106.215 ;
        RECT 57.070 106.055 57.190 106.165 ;
        RECT 57.475 106.025 57.645 106.215 ;
        RECT 61.155 106.005 61.325 106.215 ;
        RECT 63.455 106.005 63.625 106.195 ;
        RECT 63.915 106.005 64.085 106.195 ;
        RECT 72.195 106.025 72.365 106.215 ;
        RECT 73.115 106.060 73.275 106.170 ;
        RECT 75.875 106.005 76.045 106.195 ;
        RECT 77.255 106.005 77.425 106.195 ;
        RECT 78.635 106.005 78.805 106.195 ;
        RECT 81.395 106.005 81.565 106.195 ;
        RECT 83.695 106.025 83.865 106.215 ;
        RECT 85.075 106.025 85.245 106.215 ;
        RECT 85.590 106.055 85.710 106.165 ;
        RECT 85.995 106.025 86.165 106.215 ;
        RECT 86.915 106.005 87.085 106.195 ;
        RECT 87.890 106.055 88.010 106.165 ;
        RECT 88.295 106.005 88.465 106.195 ;
        RECT 89.675 106.005 89.845 106.195 ;
        RECT 97.955 106.025 98.125 106.215 ;
        RECT 98.875 106.060 99.035 106.170 ;
        RECT 99.335 106.025 99.505 106.215 ;
        RECT 111.745 106.195 111.915 106.215 ;
        RECT 101.635 106.005 101.805 106.195 ;
        RECT 103.015 106.005 103.185 106.195 ;
        RECT 104.395 106.005 104.565 106.195 ;
        RECT 105.315 106.050 105.475 106.160 ;
        RECT 105.775 106.005 105.945 106.195 ;
        RECT 108.075 106.005 108.245 106.195 ;
        RECT 110.375 106.060 110.535 106.170 ;
        RECT 111.745 106.025 111.925 106.195 ;
        RECT 111.755 106.005 111.925 106.025 ;
        RECT 113.135 106.005 113.305 106.215 ;
        RECT 11.335 105.195 12.705 106.005 ;
        RECT 13.175 105.195 15.925 106.005 ;
        RECT 15.935 105.195 21.445 106.005 ;
        RECT 21.465 105.095 22.815 106.005 ;
        RECT 22.845 105.135 23.275 105.920 ;
        RECT 23.495 105.325 33.865 106.005 ;
        RECT 23.495 105.095 25.705 105.325 ;
        RECT 28.425 105.105 29.355 105.325 ;
        RECT 33.875 105.195 35.705 106.005 ;
        RECT 35.725 105.135 36.155 105.920 ;
        RECT 36.175 105.195 37.545 106.005 ;
        RECT 37.555 105.195 43.065 106.005 ;
        RECT 43.075 105.195 48.585 106.005 ;
        RECT 48.605 105.135 49.035 105.920 ;
        RECT 49.065 105.095 50.415 106.005 ;
        RECT 50.435 105.195 55.945 106.005 ;
        RECT 55.955 105.195 61.465 106.005 ;
        RECT 61.485 105.135 61.915 105.920 ;
        RECT 61.935 105.195 63.765 106.005 ;
        RECT 63.775 105.325 74.145 106.005 ;
        RECT 68.285 105.105 69.215 105.325 ;
        RECT 71.935 105.095 74.145 105.325 ;
        RECT 74.365 105.135 74.795 105.920 ;
        RECT 74.825 105.095 76.175 106.005 ;
        RECT 76.195 105.195 77.565 106.005 ;
        RECT 77.585 105.095 78.935 106.005 ;
        RECT 78.955 105.195 81.705 106.005 ;
        RECT 81.715 105.195 87.225 106.005 ;
        RECT 87.245 105.135 87.675 105.920 ;
        RECT 88.165 105.095 89.515 106.005 ;
        RECT 89.535 105.325 99.905 106.005 ;
        RECT 94.045 105.105 94.975 105.325 ;
        RECT 97.695 105.095 99.905 105.325 ;
        RECT 100.125 105.135 100.555 105.920 ;
        RECT 100.585 105.095 101.935 106.005 ;
        RECT 101.955 105.195 103.325 106.005 ;
        RECT 103.345 105.095 104.695 106.005 ;
        RECT 105.645 105.095 106.995 106.005 ;
        RECT 107.015 105.195 108.385 106.005 ;
        RECT 108.395 105.195 112.065 106.005 ;
        RECT 112.075 105.195 113.445 106.005 ;
      LAYER nwell ;
        RECT 11.140 103.200 113.640 104.805 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 11.330 203.945 113.450 204.115 ;
        RECT 11.415 203.195 12.625 203.945 ;
        RECT 11.415 202.655 11.935 203.195 ;
        RECT 13.715 203.175 17.225 203.945 ;
        RECT 17.400 203.400 22.745 203.945 ;
        RECT 12.105 202.485 12.625 203.025 ;
        RECT 11.415 201.395 12.625 202.485 ;
        RECT 13.715 202.485 15.405 203.005 ;
        RECT 15.575 202.655 17.225 203.175 ;
        RECT 13.715 201.395 17.225 202.485 ;
        RECT 18.990 201.830 19.340 203.080 ;
        RECT 20.820 202.570 21.160 203.400 ;
        RECT 22.915 203.220 23.205 203.945 ;
        RECT 23.375 203.195 24.585 203.945 ;
        RECT 24.760 203.400 30.105 203.945 ;
        RECT 30.280 203.400 35.625 203.945 ;
        RECT 17.400 201.395 22.745 201.830 ;
        RECT 22.915 201.395 23.205 202.560 ;
        RECT 23.375 202.485 23.895 203.025 ;
        RECT 24.065 202.655 24.585 203.195 ;
        RECT 23.375 201.395 24.585 202.485 ;
        RECT 26.350 201.830 26.700 203.080 ;
        RECT 28.180 202.570 28.520 203.400 ;
        RECT 31.870 201.830 32.220 203.080 ;
        RECT 33.700 202.570 34.040 203.400 ;
        RECT 35.795 203.220 36.085 203.945 ;
        RECT 36.255 203.195 37.465 203.945 ;
        RECT 37.640 203.400 42.985 203.945 ;
        RECT 43.160 203.400 48.505 203.945 ;
        RECT 24.760 201.395 30.105 201.830 ;
        RECT 30.280 201.395 35.625 201.830 ;
        RECT 35.795 201.395 36.085 202.560 ;
        RECT 36.255 202.485 36.775 203.025 ;
        RECT 36.945 202.655 37.465 203.195 ;
        RECT 36.255 201.395 37.465 202.485 ;
        RECT 39.230 201.830 39.580 203.080 ;
        RECT 41.060 202.570 41.400 203.400 ;
        RECT 44.750 201.830 45.100 203.080 ;
        RECT 46.580 202.570 46.920 203.400 ;
        RECT 48.675 203.220 48.965 203.945 ;
        RECT 49.135 203.195 50.345 203.945 ;
        RECT 50.520 203.400 55.865 203.945 ;
        RECT 56.040 203.400 61.385 203.945 ;
        RECT 37.640 201.395 42.985 201.830 ;
        RECT 43.160 201.395 48.505 201.830 ;
        RECT 48.675 201.395 48.965 202.560 ;
        RECT 49.135 202.485 49.655 203.025 ;
        RECT 49.825 202.655 50.345 203.195 ;
        RECT 49.135 201.395 50.345 202.485 ;
        RECT 52.110 201.830 52.460 203.080 ;
        RECT 53.940 202.570 54.280 203.400 ;
        RECT 57.630 201.830 57.980 203.080 ;
        RECT 59.460 202.570 59.800 203.400 ;
        RECT 61.555 203.220 61.845 203.945 ;
        RECT 62.015 203.195 63.225 203.945 ;
        RECT 63.400 203.400 68.745 203.945 ;
        RECT 68.920 203.400 74.265 203.945 ;
        RECT 50.520 201.395 55.865 201.830 ;
        RECT 56.040 201.395 61.385 201.830 ;
        RECT 61.555 201.395 61.845 202.560 ;
        RECT 62.015 202.485 62.535 203.025 ;
        RECT 62.705 202.655 63.225 203.195 ;
        RECT 62.015 201.395 63.225 202.485 ;
        RECT 64.990 201.830 65.340 203.080 ;
        RECT 66.820 202.570 67.160 203.400 ;
        RECT 70.510 201.830 70.860 203.080 ;
        RECT 72.340 202.570 72.680 203.400 ;
        RECT 74.435 203.220 74.725 203.945 ;
        RECT 74.895 203.195 76.105 203.945 ;
        RECT 76.280 203.400 81.625 203.945 ;
        RECT 81.800 203.400 87.145 203.945 ;
        RECT 63.400 201.395 68.745 201.830 ;
        RECT 68.920 201.395 74.265 201.830 ;
        RECT 74.435 201.395 74.725 202.560 ;
        RECT 74.895 202.485 75.415 203.025 ;
        RECT 75.585 202.655 76.105 203.195 ;
        RECT 74.895 201.395 76.105 202.485 ;
        RECT 77.870 201.830 78.220 203.080 ;
        RECT 79.700 202.570 80.040 203.400 ;
        RECT 83.390 201.830 83.740 203.080 ;
        RECT 85.220 202.570 85.560 203.400 ;
        RECT 87.315 203.220 87.605 203.945 ;
        RECT 87.775 203.195 88.985 203.945 ;
        RECT 89.160 203.400 94.505 203.945 ;
        RECT 94.680 203.400 100.025 203.945 ;
        RECT 76.280 201.395 81.625 201.830 ;
        RECT 81.800 201.395 87.145 201.830 ;
        RECT 87.315 201.395 87.605 202.560 ;
        RECT 87.775 202.485 88.295 203.025 ;
        RECT 88.465 202.655 88.985 203.195 ;
        RECT 87.775 201.395 88.985 202.485 ;
        RECT 90.750 201.830 91.100 203.080 ;
        RECT 92.580 202.570 92.920 203.400 ;
        RECT 96.270 201.830 96.620 203.080 ;
        RECT 98.100 202.570 98.440 203.400 ;
        RECT 100.195 203.220 100.485 203.945 ;
        RECT 101.120 203.400 106.465 203.945 ;
        RECT 106.640 203.400 111.985 203.945 ;
        RECT 89.160 201.395 94.505 201.830 ;
        RECT 94.680 201.395 100.025 201.830 ;
        RECT 100.195 201.395 100.485 202.560 ;
        RECT 102.710 201.830 103.060 203.080 ;
        RECT 104.540 202.570 104.880 203.400 ;
        RECT 108.230 201.830 108.580 203.080 ;
        RECT 110.060 202.570 110.400 203.400 ;
        RECT 112.155 203.195 113.365 203.945 ;
        RECT 112.155 202.485 112.675 203.025 ;
        RECT 112.845 202.655 113.365 203.195 ;
        RECT 101.120 201.395 106.465 201.830 ;
        RECT 106.640 201.395 111.985 201.830 ;
        RECT 112.155 201.395 113.365 202.485 ;
        RECT 11.330 201.225 113.450 201.395 ;
        RECT 11.415 200.135 12.625 201.225 ;
        RECT 13.720 200.790 19.065 201.225 ;
        RECT 19.240 200.790 24.585 201.225 ;
        RECT 24.760 200.790 30.105 201.225 ;
        RECT 30.280 200.790 35.625 201.225 ;
        RECT 11.415 199.425 11.935 199.965 ;
        RECT 12.105 199.595 12.625 200.135 ;
        RECT 15.310 199.540 15.660 200.790 ;
        RECT 11.415 198.675 12.625 199.425 ;
        RECT 17.140 199.220 17.480 200.050 ;
        RECT 20.830 199.540 21.180 200.790 ;
        RECT 22.660 199.220 23.000 200.050 ;
        RECT 26.350 199.540 26.700 200.790 ;
        RECT 28.180 199.220 28.520 200.050 ;
        RECT 31.870 199.540 32.220 200.790 ;
        RECT 35.795 200.060 36.085 201.225 ;
        RECT 36.715 200.135 39.305 201.225 ;
        RECT 39.480 200.790 44.825 201.225 ;
        RECT 45.000 200.790 50.345 201.225 ;
        RECT 50.520 200.790 55.865 201.225 ;
        RECT 33.700 199.220 34.040 200.050 ;
        RECT 36.715 199.615 37.925 200.135 ;
        RECT 38.095 199.445 39.305 199.965 ;
        RECT 41.070 199.540 41.420 200.790 ;
        RECT 13.720 198.675 19.065 199.220 ;
        RECT 19.240 198.675 24.585 199.220 ;
        RECT 24.760 198.675 30.105 199.220 ;
        RECT 30.280 198.675 35.625 199.220 ;
        RECT 35.795 198.675 36.085 199.400 ;
        RECT 36.715 198.675 39.305 199.445 ;
        RECT 42.900 199.220 43.240 200.050 ;
        RECT 46.590 199.540 46.940 200.790 ;
        RECT 48.420 199.220 48.760 200.050 ;
        RECT 52.110 199.540 52.460 200.790 ;
        RECT 56.095 200.085 56.305 201.225 ;
        RECT 56.475 200.075 56.805 201.055 ;
        RECT 56.975 200.085 57.205 201.225 ;
        RECT 58.375 200.085 58.605 201.225 ;
        RECT 58.775 200.075 59.105 201.055 ;
        RECT 59.275 200.085 59.485 201.225 ;
        RECT 59.720 200.075 59.980 201.225 ;
        RECT 60.155 200.150 60.410 201.055 ;
        RECT 60.580 200.465 60.910 201.225 ;
        RECT 61.125 200.295 61.295 201.055 ;
        RECT 53.940 199.220 54.280 200.050 ;
        RECT 39.480 198.675 44.825 199.220 ;
        RECT 45.000 198.675 50.345 199.220 ;
        RECT 50.520 198.675 55.865 199.220 ;
        RECT 56.095 198.675 56.305 199.495 ;
        RECT 56.475 199.475 56.725 200.075 ;
        RECT 56.895 199.665 57.225 199.915 ;
        RECT 58.355 199.665 58.685 199.915 ;
        RECT 56.475 198.845 56.805 199.475 ;
        RECT 56.975 198.675 57.205 199.495 ;
        RECT 58.375 198.675 58.605 199.495 ;
        RECT 58.855 199.475 59.105 200.075 ;
        RECT 58.775 198.845 59.105 199.475 ;
        RECT 59.275 198.675 59.485 199.495 ;
        RECT 59.720 198.675 59.980 199.515 ;
        RECT 60.155 199.420 60.325 200.150 ;
        RECT 60.580 200.125 61.295 200.295 ;
        RECT 60.580 199.915 60.750 200.125 ;
        RECT 61.555 200.060 61.845 201.225 ;
        RECT 62.020 200.035 62.275 200.915 ;
        RECT 62.445 200.085 62.750 201.225 ;
        RECT 63.090 200.845 63.420 201.225 ;
        RECT 63.600 200.675 63.770 200.965 ;
        RECT 63.940 200.765 64.190 201.225 ;
        RECT 62.970 200.505 63.770 200.675 ;
        RECT 64.360 200.715 65.230 201.055 ;
        RECT 60.495 199.585 60.750 199.915 ;
        RECT 60.155 198.845 60.410 199.420 ;
        RECT 60.580 199.395 60.750 199.585 ;
        RECT 61.030 199.575 61.385 199.945 ;
        RECT 60.580 199.225 61.295 199.395 ;
        RECT 60.580 198.675 60.910 199.055 ;
        RECT 61.125 198.845 61.295 199.225 ;
        RECT 61.555 198.675 61.845 199.400 ;
        RECT 62.020 199.385 62.230 200.035 ;
        RECT 62.970 199.915 63.140 200.505 ;
        RECT 64.360 200.335 64.530 200.715 ;
        RECT 65.465 200.595 65.635 201.055 ;
        RECT 65.805 200.765 66.175 201.225 ;
        RECT 66.470 200.625 66.640 200.965 ;
        RECT 66.810 200.795 67.140 201.225 ;
        RECT 67.375 200.625 67.545 200.965 ;
        RECT 63.310 200.165 64.530 200.335 ;
        RECT 64.700 200.255 65.160 200.545 ;
        RECT 65.465 200.425 66.025 200.595 ;
        RECT 66.470 200.455 67.545 200.625 ;
        RECT 67.715 200.725 68.395 201.055 ;
        RECT 68.610 200.725 68.860 201.055 ;
        RECT 69.030 200.765 69.280 201.225 ;
        RECT 65.855 200.285 66.025 200.425 ;
        RECT 64.700 200.245 65.665 200.255 ;
        RECT 64.360 200.075 64.530 200.165 ;
        RECT 64.990 200.085 65.665 200.245 ;
        RECT 62.400 199.885 63.140 199.915 ;
        RECT 62.400 199.585 63.315 199.885 ;
        RECT 62.990 199.410 63.315 199.585 ;
        RECT 62.020 198.855 62.275 199.385 ;
        RECT 62.445 198.675 62.750 199.135 ;
        RECT 62.995 199.055 63.315 199.410 ;
        RECT 63.485 199.625 64.025 199.995 ;
        RECT 64.360 199.905 64.765 200.075 ;
        RECT 63.485 199.225 63.725 199.625 ;
        RECT 64.205 199.455 64.425 199.735 ;
        RECT 63.895 199.285 64.425 199.455 ;
        RECT 63.895 199.055 64.065 199.285 ;
        RECT 64.595 199.125 64.765 199.905 ;
        RECT 64.935 199.295 65.285 199.915 ;
        RECT 65.455 199.295 65.665 200.085 ;
        RECT 65.855 200.115 67.355 200.285 ;
        RECT 65.855 199.425 66.025 200.115 ;
        RECT 67.715 199.945 67.885 200.725 ;
        RECT 68.690 200.595 68.860 200.725 ;
        RECT 66.195 199.775 67.885 199.945 ;
        RECT 68.055 200.165 68.520 200.555 ;
        RECT 68.690 200.425 69.085 200.595 ;
        RECT 66.195 199.595 66.365 199.775 ;
        RECT 62.995 198.885 64.065 199.055 ;
        RECT 64.235 198.675 64.425 199.115 ;
        RECT 64.595 198.845 65.545 199.125 ;
        RECT 65.855 199.035 66.115 199.425 ;
        RECT 66.535 199.355 67.325 199.605 ;
        RECT 65.765 198.865 66.115 199.035 ;
        RECT 66.325 198.675 66.655 199.135 ;
        RECT 67.530 199.065 67.700 199.775 ;
        RECT 68.055 199.575 68.225 200.165 ;
        RECT 67.870 199.355 68.225 199.575 ;
        RECT 68.395 199.355 68.745 199.975 ;
        RECT 68.915 199.065 69.085 200.425 ;
        RECT 69.450 200.255 69.775 201.040 ;
        RECT 69.255 199.205 69.715 200.255 ;
        RECT 67.530 198.895 68.385 199.065 ;
        RECT 68.590 198.895 69.085 199.065 ;
        RECT 69.255 198.675 69.585 199.035 ;
        RECT 69.945 198.935 70.115 201.055 ;
        RECT 70.285 200.725 70.615 201.225 ;
        RECT 70.785 200.555 71.040 201.055 ;
        RECT 70.290 200.385 71.040 200.555 ;
        RECT 70.290 199.395 70.520 200.385 ;
        RECT 70.690 199.565 71.040 200.215 ;
        RECT 71.215 200.135 72.885 201.225 ;
        RECT 71.215 199.615 71.965 200.135 ;
        RECT 73.095 200.085 73.325 201.225 ;
        RECT 73.495 200.075 73.825 201.055 ;
        RECT 73.995 200.085 74.205 201.225 ;
        RECT 74.475 200.085 74.705 201.225 ;
        RECT 74.875 200.075 75.205 201.055 ;
        RECT 75.375 200.085 75.585 201.225 ;
        RECT 76.280 200.790 81.625 201.225 ;
        RECT 81.800 200.790 87.145 201.225 ;
        RECT 72.135 199.445 72.885 199.965 ;
        RECT 73.075 199.665 73.405 199.915 ;
        RECT 70.290 199.225 71.040 199.395 ;
        RECT 70.285 198.675 70.615 199.055 ;
        RECT 70.785 198.935 71.040 199.225 ;
        RECT 71.215 198.675 72.885 199.445 ;
        RECT 73.095 198.675 73.325 199.495 ;
        RECT 73.575 199.475 73.825 200.075 ;
        RECT 74.455 199.665 74.785 199.915 ;
        RECT 73.495 198.845 73.825 199.475 ;
        RECT 73.995 198.675 74.205 199.495 ;
        RECT 74.475 198.675 74.705 199.495 ;
        RECT 74.955 199.475 75.205 200.075 ;
        RECT 77.870 199.540 78.220 200.790 ;
        RECT 74.875 198.845 75.205 199.475 ;
        RECT 75.375 198.675 75.585 199.495 ;
        RECT 79.700 199.220 80.040 200.050 ;
        RECT 83.390 199.540 83.740 200.790 ;
        RECT 87.315 200.060 87.605 201.225 ;
        RECT 88.235 200.135 89.905 201.225 ;
        RECT 90.080 200.790 95.425 201.225 ;
        RECT 95.600 200.790 100.945 201.225 ;
        RECT 101.120 200.790 106.465 201.225 ;
        RECT 106.640 200.790 111.985 201.225 ;
        RECT 85.220 199.220 85.560 200.050 ;
        RECT 88.235 199.615 88.985 200.135 ;
        RECT 89.155 199.445 89.905 199.965 ;
        RECT 91.670 199.540 92.020 200.790 ;
        RECT 76.280 198.675 81.625 199.220 ;
        RECT 81.800 198.675 87.145 199.220 ;
        RECT 87.315 198.675 87.605 199.400 ;
        RECT 88.235 198.675 89.905 199.445 ;
        RECT 93.500 199.220 93.840 200.050 ;
        RECT 97.190 199.540 97.540 200.790 ;
        RECT 99.020 199.220 99.360 200.050 ;
        RECT 102.710 199.540 103.060 200.790 ;
        RECT 104.540 199.220 104.880 200.050 ;
        RECT 108.230 199.540 108.580 200.790 ;
        RECT 112.155 200.135 113.365 201.225 ;
        RECT 110.060 199.220 110.400 200.050 ;
        RECT 112.155 199.595 112.675 200.135 ;
        RECT 112.845 199.425 113.365 199.965 ;
        RECT 90.080 198.675 95.425 199.220 ;
        RECT 95.600 198.675 100.945 199.220 ;
        RECT 101.120 198.675 106.465 199.220 ;
        RECT 106.640 198.675 111.985 199.220 ;
        RECT 112.155 198.675 113.365 199.425 ;
        RECT 11.330 198.505 113.450 198.675 ;
        RECT 11.415 197.755 12.625 198.505 ;
        RECT 11.415 197.215 11.935 197.755 ;
        RECT 13.715 197.735 17.225 198.505 ;
        RECT 17.400 197.960 22.745 198.505 ;
        RECT 12.105 197.045 12.625 197.585 ;
        RECT 11.415 195.955 12.625 197.045 ;
        RECT 13.715 197.045 15.405 197.565 ;
        RECT 15.575 197.215 17.225 197.735 ;
        RECT 13.715 195.955 17.225 197.045 ;
        RECT 18.990 196.390 19.340 197.640 ;
        RECT 20.820 197.130 21.160 197.960 ;
        RECT 22.915 197.780 23.205 198.505 ;
        RECT 23.835 197.735 26.425 198.505 ;
        RECT 26.600 197.960 31.945 198.505 ;
        RECT 32.120 197.960 37.465 198.505 ;
        RECT 37.640 197.960 42.985 198.505 ;
        RECT 43.160 197.960 48.505 198.505 ;
        RECT 17.400 195.955 22.745 196.390 ;
        RECT 22.915 195.955 23.205 197.120 ;
        RECT 23.835 197.045 25.045 197.565 ;
        RECT 25.215 197.215 26.425 197.735 ;
        RECT 23.835 195.955 26.425 197.045 ;
        RECT 28.190 196.390 28.540 197.640 ;
        RECT 30.020 197.130 30.360 197.960 ;
        RECT 33.710 196.390 34.060 197.640 ;
        RECT 35.540 197.130 35.880 197.960 ;
        RECT 39.230 196.390 39.580 197.640 ;
        RECT 41.060 197.130 41.400 197.960 ;
        RECT 44.750 196.390 45.100 197.640 ;
        RECT 46.580 197.130 46.920 197.960 ;
        RECT 48.675 197.780 48.965 198.505 ;
        RECT 49.595 197.735 51.265 198.505 ;
        RECT 51.440 197.955 51.695 198.245 ;
        RECT 51.865 198.125 52.195 198.505 ;
        RECT 51.440 197.785 52.190 197.955 ;
        RECT 26.600 195.955 31.945 196.390 ;
        RECT 32.120 195.955 37.465 196.390 ;
        RECT 37.640 195.955 42.985 196.390 ;
        RECT 43.160 195.955 48.505 196.390 ;
        RECT 48.675 195.955 48.965 197.120 ;
        RECT 49.595 197.045 50.345 197.565 ;
        RECT 50.515 197.215 51.265 197.735 ;
        RECT 49.595 195.955 51.265 197.045 ;
        RECT 51.440 196.965 51.790 197.615 ;
        RECT 51.960 196.795 52.190 197.785 ;
        RECT 51.440 196.625 52.190 196.795 ;
        RECT 51.440 196.125 51.695 196.625 ;
        RECT 51.865 195.955 52.195 196.455 ;
        RECT 52.365 196.125 52.535 198.245 ;
        RECT 52.895 198.145 53.225 198.505 ;
        RECT 53.395 198.115 53.890 198.285 ;
        RECT 54.095 198.115 54.950 198.285 ;
        RECT 52.765 196.925 53.225 197.975 ;
        RECT 52.705 196.140 53.030 196.925 ;
        RECT 53.395 196.755 53.565 198.115 ;
        RECT 53.735 197.205 54.085 197.825 ;
        RECT 54.255 197.605 54.610 197.825 ;
        RECT 54.255 197.015 54.425 197.605 ;
        RECT 54.780 197.405 54.950 198.115 ;
        RECT 55.825 198.045 56.155 198.505 ;
        RECT 56.365 198.145 56.715 198.315 ;
        RECT 55.155 197.575 55.945 197.825 ;
        RECT 56.365 197.755 56.625 198.145 ;
        RECT 56.935 198.055 57.885 198.335 ;
        RECT 58.055 198.065 58.245 198.505 ;
        RECT 58.415 198.125 59.485 198.295 ;
        RECT 56.115 197.405 56.285 197.585 ;
        RECT 53.395 196.585 53.790 196.755 ;
        RECT 53.960 196.625 54.425 197.015 ;
        RECT 54.595 197.235 56.285 197.405 ;
        RECT 53.620 196.455 53.790 196.585 ;
        RECT 54.595 196.455 54.765 197.235 ;
        RECT 56.455 197.065 56.625 197.755 ;
        RECT 55.125 196.895 56.625 197.065 ;
        RECT 56.815 197.095 57.025 197.885 ;
        RECT 57.195 197.265 57.545 197.885 ;
        RECT 57.715 197.275 57.885 198.055 ;
        RECT 58.415 197.895 58.585 198.125 ;
        RECT 58.055 197.725 58.585 197.895 ;
        RECT 58.055 197.445 58.275 197.725 ;
        RECT 58.755 197.555 58.995 197.955 ;
        RECT 57.715 197.105 58.120 197.275 ;
        RECT 58.455 197.185 58.995 197.555 ;
        RECT 59.165 197.770 59.485 198.125 ;
        RECT 59.165 197.515 59.490 197.770 ;
        RECT 59.685 197.695 59.855 198.505 ;
        RECT 60.025 197.855 60.355 198.335 ;
        RECT 60.525 198.035 60.695 198.505 ;
        RECT 60.865 197.855 61.195 198.335 ;
        RECT 61.365 198.035 61.535 198.505 ;
        RECT 62.480 198.250 62.815 198.295 ;
        RECT 60.025 197.685 61.790 197.855 ;
        RECT 59.165 197.305 61.195 197.515 ;
        RECT 59.165 197.295 59.510 197.305 ;
        RECT 56.815 196.935 57.490 197.095 ;
        RECT 57.950 197.015 58.120 197.105 ;
        RECT 56.815 196.925 57.780 196.935 ;
        RECT 56.455 196.755 56.625 196.895 ;
        RECT 53.200 195.955 53.450 196.415 ;
        RECT 53.620 196.125 53.870 196.455 ;
        RECT 54.085 196.125 54.765 196.455 ;
        RECT 54.935 196.555 56.010 196.725 ;
        RECT 56.455 196.585 57.015 196.755 ;
        RECT 57.320 196.635 57.780 196.925 ;
        RECT 57.950 196.845 59.170 197.015 ;
        RECT 54.935 196.215 55.105 196.555 ;
        RECT 55.340 195.955 55.670 196.385 ;
        RECT 55.840 196.215 56.010 196.555 ;
        RECT 56.305 195.955 56.675 196.415 ;
        RECT 56.845 196.125 57.015 196.585 ;
        RECT 57.950 196.465 58.120 196.845 ;
        RECT 59.340 196.675 59.510 197.295 ;
        RECT 61.380 197.135 61.790 197.685 ;
        RECT 57.250 196.125 58.120 196.465 ;
        RECT 58.710 196.505 59.510 196.675 ;
        RECT 58.290 195.955 58.540 196.415 ;
        RECT 58.710 196.215 58.880 196.505 ;
        RECT 59.060 195.955 59.390 196.335 ;
        RECT 59.685 195.955 59.855 197.015 ;
        RECT 60.065 196.965 61.790 197.135 ;
        RECT 62.475 197.785 62.815 198.250 ;
        RECT 62.985 198.125 63.315 198.505 ;
        RECT 62.475 197.095 62.645 197.785 ;
        RECT 62.815 197.265 63.075 197.595 ;
        RECT 60.065 196.125 60.355 196.965 ;
        RECT 60.525 195.955 60.695 196.795 ;
        RECT 60.905 196.125 61.155 196.965 ;
        RECT 61.365 195.955 61.535 196.795 ;
        RECT 62.475 196.125 62.735 197.095 ;
        RECT 62.905 196.715 63.075 197.265 ;
        RECT 63.245 196.895 63.585 197.925 ;
        RECT 63.775 197.145 64.045 198.170 ;
        RECT 63.775 196.975 64.085 197.145 ;
        RECT 63.775 196.895 64.045 196.975 ;
        RECT 64.270 196.895 64.550 198.170 ;
        RECT 64.750 198.005 64.980 198.335 ;
        RECT 65.225 198.125 65.555 198.505 ;
        RECT 64.750 196.715 64.920 198.005 ;
        RECT 65.725 197.935 65.900 198.335 ;
        RECT 65.270 197.765 65.900 197.935 ;
        RECT 65.270 197.595 65.440 197.765 ;
        RECT 66.155 197.755 67.365 198.505 ;
        RECT 65.090 197.265 65.440 197.595 ;
        RECT 62.905 196.545 64.920 196.715 ;
        RECT 65.270 196.745 65.440 197.265 ;
        RECT 65.620 196.915 65.985 197.595 ;
        RECT 66.155 197.045 66.675 197.585 ;
        RECT 66.845 197.215 67.365 197.755 ;
        RECT 67.535 197.765 68.000 198.310 ;
        RECT 65.270 196.575 65.900 196.745 ;
        RECT 62.930 195.955 63.260 196.365 ;
        RECT 63.460 196.125 63.630 196.545 ;
        RECT 63.845 195.955 64.515 196.365 ;
        RECT 64.750 196.125 64.920 196.545 ;
        RECT 65.225 195.955 65.555 196.395 ;
        RECT 65.725 196.125 65.900 196.575 ;
        RECT 66.155 195.955 67.365 197.045 ;
        RECT 67.535 196.805 67.705 197.765 ;
        RECT 68.505 197.685 68.675 198.505 ;
        RECT 68.845 197.855 69.175 198.335 ;
        RECT 69.345 198.115 69.695 198.505 ;
        RECT 69.865 197.935 70.095 198.335 ;
        RECT 69.585 197.855 70.095 197.935 ;
        RECT 68.845 197.765 70.095 197.855 ;
        RECT 70.265 197.765 70.585 198.245 ;
        RECT 68.845 197.685 69.755 197.765 ;
        RECT 67.875 197.145 68.120 197.595 ;
        RECT 68.380 197.315 69.075 197.515 ;
        RECT 69.245 197.345 69.845 197.515 ;
        RECT 69.245 197.145 69.415 197.345 ;
        RECT 70.075 197.175 70.245 197.595 ;
        RECT 67.875 196.975 69.415 197.145 ;
        RECT 69.585 197.005 70.245 197.175 ;
        RECT 69.585 196.805 69.755 197.005 ;
        RECT 70.415 196.835 70.585 197.765 ;
        RECT 71.715 197.685 71.945 198.505 ;
        RECT 72.115 197.705 72.445 198.335 ;
        RECT 71.695 197.265 72.025 197.515 ;
        RECT 72.195 197.105 72.445 197.705 ;
        RECT 72.615 197.685 72.825 198.505 ;
        RECT 73.145 197.955 73.315 198.335 ;
        RECT 73.495 198.125 73.825 198.505 ;
        RECT 73.145 197.785 73.810 197.955 ;
        RECT 74.005 197.830 74.265 198.335 ;
        RECT 73.075 197.235 73.405 197.605 ;
        RECT 73.640 197.530 73.810 197.785 ;
        RECT 67.535 196.635 69.755 196.805 ;
        RECT 69.925 196.635 70.585 196.835 ;
        RECT 67.535 195.955 67.835 196.465 ;
        RECT 68.005 196.125 68.335 196.635 ;
        RECT 69.925 196.465 70.095 196.635 ;
        RECT 68.505 195.955 69.135 196.465 ;
        RECT 69.715 196.295 70.095 196.465 ;
        RECT 70.265 195.955 70.565 196.465 ;
        RECT 71.715 195.955 71.945 197.095 ;
        RECT 72.115 196.125 72.445 197.105 ;
        RECT 73.640 197.200 73.925 197.530 ;
        RECT 72.615 195.955 72.825 197.095 ;
        RECT 73.640 197.055 73.810 197.200 ;
        RECT 73.145 196.885 73.810 197.055 ;
        RECT 74.095 197.030 74.265 197.830 ;
        RECT 74.435 197.780 74.725 198.505 ;
        RECT 74.900 197.795 75.155 198.325 ;
        RECT 75.325 198.045 75.630 198.505 ;
        RECT 75.875 198.125 76.945 198.295 ;
        RECT 74.900 197.145 75.110 197.795 ;
        RECT 75.875 197.770 76.195 198.125 ;
        RECT 75.870 197.595 76.195 197.770 ;
        RECT 75.280 197.295 76.195 197.595 ;
        RECT 76.365 197.555 76.605 197.955 ;
        RECT 76.775 197.895 76.945 198.125 ;
        RECT 77.115 198.065 77.305 198.505 ;
        RECT 77.475 198.055 78.425 198.335 ;
        RECT 78.645 198.145 78.995 198.315 ;
        RECT 76.775 197.725 77.305 197.895 ;
        RECT 75.280 197.265 76.020 197.295 ;
        RECT 73.145 196.125 73.315 196.885 ;
        RECT 73.495 195.955 73.825 196.715 ;
        RECT 73.995 196.125 74.265 197.030 ;
        RECT 74.435 195.955 74.725 197.120 ;
        RECT 74.900 196.265 75.155 197.145 ;
        RECT 75.325 195.955 75.630 197.095 ;
        RECT 75.850 196.675 76.020 197.265 ;
        RECT 76.365 197.185 76.905 197.555 ;
        RECT 77.085 197.445 77.305 197.725 ;
        RECT 77.475 197.275 77.645 198.055 ;
        RECT 77.240 197.105 77.645 197.275 ;
        RECT 77.815 197.265 78.165 197.885 ;
        RECT 77.240 197.015 77.410 197.105 ;
        RECT 78.335 197.095 78.545 197.885 ;
        RECT 76.190 196.845 77.410 197.015 ;
        RECT 77.870 196.935 78.545 197.095 ;
        RECT 75.850 196.505 76.650 196.675 ;
        RECT 75.970 195.955 76.300 196.335 ;
        RECT 76.480 196.215 76.650 196.505 ;
        RECT 77.240 196.465 77.410 196.845 ;
        RECT 77.580 196.925 78.545 196.935 ;
        RECT 78.735 197.755 78.995 198.145 ;
        RECT 79.205 198.045 79.535 198.505 ;
        RECT 80.410 198.115 81.265 198.285 ;
        RECT 81.470 198.115 81.965 198.285 ;
        RECT 82.135 198.145 82.465 198.505 ;
        RECT 78.735 197.065 78.905 197.755 ;
        RECT 79.075 197.405 79.245 197.585 ;
        RECT 79.415 197.575 80.205 197.825 ;
        RECT 80.410 197.405 80.580 198.115 ;
        RECT 80.750 197.605 81.105 197.825 ;
        RECT 79.075 197.235 80.765 197.405 ;
        RECT 77.580 196.635 78.040 196.925 ;
        RECT 78.735 196.895 80.235 197.065 ;
        RECT 78.735 196.755 78.905 196.895 ;
        RECT 78.345 196.585 78.905 196.755 ;
        RECT 76.820 195.955 77.070 196.415 ;
        RECT 77.240 196.125 78.110 196.465 ;
        RECT 78.345 196.125 78.515 196.585 ;
        RECT 79.350 196.555 80.425 196.725 ;
        RECT 78.685 195.955 79.055 196.415 ;
        RECT 79.350 196.215 79.520 196.555 ;
        RECT 79.690 195.955 80.020 196.385 ;
        RECT 80.255 196.215 80.425 196.555 ;
        RECT 80.595 196.455 80.765 197.235 ;
        RECT 80.935 197.015 81.105 197.605 ;
        RECT 81.275 197.205 81.625 197.825 ;
        RECT 80.935 196.625 81.400 197.015 ;
        RECT 81.795 196.755 81.965 198.115 ;
        RECT 82.135 196.925 82.595 197.975 ;
        RECT 81.570 196.585 81.965 196.755 ;
        RECT 81.570 196.455 81.740 196.585 ;
        RECT 80.595 196.125 81.275 196.455 ;
        RECT 81.490 196.125 81.740 196.455 ;
        RECT 81.910 195.955 82.160 196.415 ;
        RECT 82.330 196.140 82.655 196.925 ;
        RECT 82.825 196.125 82.995 198.245 ;
        RECT 83.165 198.125 83.495 198.505 ;
        RECT 83.665 197.955 83.920 198.245 ;
        RECT 83.170 197.785 83.920 197.955 ;
        RECT 83.170 196.795 83.400 197.785 ;
        RECT 84.095 197.735 87.605 198.505 ;
        RECT 87.780 197.960 93.125 198.505 ;
        RECT 93.300 197.960 98.645 198.505 ;
        RECT 83.570 196.965 83.920 197.615 ;
        RECT 84.095 197.045 85.785 197.565 ;
        RECT 85.955 197.215 87.605 197.735 ;
        RECT 83.170 196.625 83.920 196.795 ;
        RECT 83.165 195.955 83.495 196.455 ;
        RECT 83.665 196.125 83.920 196.625 ;
        RECT 84.095 195.955 87.605 197.045 ;
        RECT 89.370 196.390 89.720 197.640 ;
        RECT 91.200 197.130 91.540 197.960 ;
        RECT 94.890 196.390 95.240 197.640 ;
        RECT 96.720 197.130 97.060 197.960 ;
        RECT 98.905 197.955 99.075 198.335 ;
        RECT 99.255 198.125 99.585 198.505 ;
        RECT 98.905 197.785 99.570 197.955 ;
        RECT 99.765 197.830 100.025 198.335 ;
        RECT 98.835 197.235 99.165 197.605 ;
        RECT 99.400 197.530 99.570 197.785 ;
        RECT 99.400 197.200 99.685 197.530 ;
        RECT 99.400 197.055 99.570 197.200 ;
        RECT 98.905 196.885 99.570 197.055 ;
        RECT 99.855 197.030 100.025 197.830 ;
        RECT 100.195 197.780 100.485 198.505 ;
        RECT 101.120 197.960 106.465 198.505 ;
        RECT 106.640 197.960 111.985 198.505 ;
        RECT 87.780 195.955 93.125 196.390 ;
        RECT 93.300 195.955 98.645 196.390 ;
        RECT 98.905 196.125 99.075 196.885 ;
        RECT 99.255 195.955 99.585 196.715 ;
        RECT 99.755 196.125 100.025 197.030 ;
        RECT 100.195 195.955 100.485 197.120 ;
        RECT 102.710 196.390 103.060 197.640 ;
        RECT 104.540 197.130 104.880 197.960 ;
        RECT 108.230 196.390 108.580 197.640 ;
        RECT 110.060 197.130 110.400 197.960 ;
        RECT 112.155 197.755 113.365 198.505 ;
        RECT 112.155 197.045 112.675 197.585 ;
        RECT 112.845 197.215 113.365 197.755 ;
        RECT 101.120 195.955 106.465 196.390 ;
        RECT 106.640 195.955 111.985 196.390 ;
        RECT 112.155 195.955 113.365 197.045 ;
        RECT 11.330 195.785 113.450 195.955 ;
        RECT 11.415 194.695 12.625 195.785 ;
        RECT 13.720 195.350 19.065 195.785 ;
        RECT 19.240 195.350 24.585 195.785 ;
        RECT 24.760 195.350 30.105 195.785 ;
        RECT 30.280 195.350 35.625 195.785 ;
        RECT 11.415 193.985 11.935 194.525 ;
        RECT 12.105 194.155 12.625 194.695 ;
        RECT 15.310 194.100 15.660 195.350 ;
        RECT 11.415 193.235 12.625 193.985 ;
        RECT 17.140 193.780 17.480 194.610 ;
        RECT 20.830 194.100 21.180 195.350 ;
        RECT 22.660 193.780 23.000 194.610 ;
        RECT 26.350 194.100 26.700 195.350 ;
        RECT 28.180 193.780 28.520 194.610 ;
        RECT 31.870 194.100 32.220 195.350 ;
        RECT 35.795 194.620 36.085 195.785 ;
        RECT 36.715 194.695 40.225 195.785 ;
        RECT 40.400 195.350 45.745 195.785 ;
        RECT 45.920 195.350 51.265 195.785 ;
        RECT 51.440 195.350 56.785 195.785 ;
        RECT 33.700 193.780 34.040 194.610 ;
        RECT 36.715 194.175 38.405 194.695 ;
        RECT 38.575 194.005 40.225 194.525 ;
        RECT 41.990 194.100 42.340 195.350 ;
        RECT 13.720 193.235 19.065 193.780 ;
        RECT 19.240 193.235 24.585 193.780 ;
        RECT 24.760 193.235 30.105 193.780 ;
        RECT 30.280 193.235 35.625 193.780 ;
        RECT 35.795 193.235 36.085 193.960 ;
        RECT 36.715 193.235 40.225 194.005 ;
        RECT 43.820 193.780 44.160 194.610 ;
        RECT 47.510 194.100 47.860 195.350 ;
        RECT 49.340 193.780 49.680 194.610 ;
        RECT 53.030 194.100 53.380 195.350 ;
        RECT 56.955 194.710 57.225 195.615 ;
        RECT 57.395 195.025 57.725 195.785 ;
        RECT 57.905 194.855 58.075 195.615 ;
        RECT 58.635 195.145 58.965 195.575 ;
        RECT 54.860 193.780 55.200 194.610 ;
        RECT 56.955 193.910 57.125 194.710 ;
        RECT 57.410 194.685 58.075 194.855 ;
        RECT 58.510 194.975 58.965 195.145 ;
        RECT 59.145 195.145 59.395 195.565 ;
        RECT 59.625 195.315 59.955 195.785 ;
        RECT 60.185 195.145 60.435 195.565 ;
        RECT 59.145 194.975 60.435 195.145 ;
        RECT 57.410 194.540 57.580 194.685 ;
        RECT 57.295 194.210 57.580 194.540 ;
        RECT 57.410 193.955 57.580 194.210 ;
        RECT 57.815 194.135 58.145 194.505 ;
        RECT 58.510 193.975 58.680 194.975 ;
        RECT 58.850 194.145 59.095 194.805 ;
        RECT 59.310 194.145 59.575 194.805 ;
        RECT 59.770 194.145 60.055 194.805 ;
        RECT 60.230 194.475 60.445 194.805 ;
        RECT 60.625 194.645 60.875 195.785 ;
        RECT 61.045 194.725 61.375 195.575 ;
        RECT 60.230 194.145 60.535 194.475 ;
        RECT 60.705 194.145 61.015 194.475 ;
        RECT 60.705 193.975 60.875 194.145 ;
        RECT 40.400 193.235 45.745 193.780 ;
        RECT 45.920 193.235 51.265 193.780 ;
        RECT 51.440 193.235 56.785 193.780 ;
        RECT 56.955 193.405 57.215 193.910 ;
        RECT 57.410 193.785 58.075 193.955 ;
        RECT 58.510 193.805 60.875 193.975 ;
        RECT 61.185 193.960 61.375 194.725 ;
        RECT 61.555 194.620 61.845 195.785 ;
        RECT 62.020 195.360 62.355 195.785 ;
        RECT 62.525 195.180 62.710 195.585 ;
        RECT 62.045 195.005 62.710 195.180 ;
        RECT 62.915 195.005 63.245 195.785 ;
        RECT 62.045 193.975 62.385 195.005 ;
        RECT 63.415 194.815 63.685 195.585 ;
        RECT 62.555 194.645 63.685 194.815 ;
        RECT 62.555 194.145 62.805 194.645 ;
        RECT 57.395 193.235 57.725 193.615 ;
        RECT 57.905 193.405 58.075 193.785 ;
        RECT 58.665 193.235 58.995 193.635 ;
        RECT 59.165 193.465 59.495 193.805 ;
        RECT 60.545 193.235 60.875 193.635 ;
        RECT 61.045 193.450 61.375 193.960 ;
        RECT 61.555 193.235 61.845 193.960 ;
        RECT 62.045 193.805 62.730 193.975 ;
        RECT 62.985 193.895 63.345 194.475 ;
        RECT 62.020 193.235 62.355 193.635 ;
        RECT 62.525 193.405 62.730 193.805 ;
        RECT 63.515 193.735 63.685 194.645 ;
        RECT 62.940 193.235 63.215 193.715 ;
        RECT 63.425 193.405 63.685 193.735 ;
        RECT 63.855 195.285 64.115 195.615 ;
        RECT 64.425 195.405 64.755 195.785 ;
        RECT 63.855 194.605 64.025 195.285 ;
        RECT 64.995 195.235 65.185 195.615 ;
        RECT 65.435 195.405 65.765 195.785 ;
        RECT 65.975 195.235 66.145 195.615 ;
        RECT 66.340 195.405 66.670 195.785 ;
        RECT 66.930 195.235 67.100 195.615 ;
        RECT 67.525 195.405 67.855 195.785 ;
        RECT 64.195 194.775 64.545 195.105 ;
        RECT 64.995 195.065 65.735 195.235 ;
        RECT 64.815 194.725 65.395 194.895 ;
        RECT 64.815 194.605 64.985 194.725 ;
        RECT 63.855 194.435 64.985 194.605 ;
        RECT 65.565 194.555 65.735 195.065 ;
        RECT 63.855 193.735 64.025 194.435 ;
        RECT 65.165 194.385 65.735 194.555 ;
        RECT 65.905 195.065 67.855 195.235 ;
        RECT 64.375 194.095 64.995 194.265 ;
        RECT 64.375 193.915 64.585 194.095 ;
        RECT 65.165 193.905 65.335 194.385 ;
        RECT 65.905 194.075 66.075 195.065 ;
        RECT 66.665 194.475 66.850 194.785 ;
        RECT 67.120 194.475 67.315 194.785 ;
        RECT 63.855 193.405 64.115 193.735 ;
        RECT 64.425 193.235 64.755 193.615 ;
        RECT 64.935 193.575 65.335 193.905 ;
        RECT 65.525 193.745 66.075 194.075 ;
        RECT 66.245 193.575 66.415 194.475 ;
        RECT 64.935 193.405 66.415 193.575 ;
        RECT 66.665 194.145 66.895 194.475 ;
        RECT 67.120 194.145 67.375 194.475 ;
        RECT 67.685 194.145 67.855 195.065 ;
        RECT 66.665 193.565 66.850 194.145 ;
        RECT 67.120 193.570 67.315 194.145 ;
        RECT 67.525 193.235 67.855 193.615 ;
        RECT 68.025 193.405 68.285 195.615 ;
        RECT 68.455 194.645 68.715 195.785 ;
        RECT 68.885 194.635 69.215 195.615 ;
        RECT 69.385 194.645 69.665 195.785 ;
        RECT 68.475 194.225 68.810 194.475 ;
        RECT 68.980 194.035 69.150 194.635 ;
        RECT 69.840 194.595 70.095 195.475 ;
        RECT 70.265 194.645 70.570 195.785 ;
        RECT 70.910 195.405 71.240 195.785 ;
        RECT 71.420 195.235 71.590 195.525 ;
        RECT 71.760 195.325 72.010 195.785 ;
        RECT 70.790 195.065 71.590 195.235 ;
        RECT 72.180 195.275 73.050 195.615 ;
        RECT 69.320 194.205 69.655 194.475 ;
        RECT 68.455 193.405 69.150 194.035 ;
        RECT 69.355 193.235 69.665 194.035 ;
        RECT 69.840 193.945 70.050 194.595 ;
        RECT 70.790 194.475 70.960 195.065 ;
        RECT 72.180 194.895 72.350 195.275 ;
        RECT 73.285 195.155 73.455 195.615 ;
        RECT 73.625 195.325 73.995 195.785 ;
        RECT 74.290 195.185 74.460 195.525 ;
        RECT 74.630 195.355 74.960 195.785 ;
        RECT 75.195 195.185 75.365 195.525 ;
        RECT 71.130 194.725 72.350 194.895 ;
        RECT 72.520 194.815 72.980 195.105 ;
        RECT 73.285 194.985 73.845 195.155 ;
        RECT 74.290 195.015 75.365 195.185 ;
        RECT 75.535 195.285 76.215 195.615 ;
        RECT 76.430 195.285 76.680 195.615 ;
        RECT 76.850 195.325 77.100 195.785 ;
        RECT 73.675 194.845 73.845 194.985 ;
        RECT 72.520 194.805 73.485 194.815 ;
        RECT 72.180 194.635 72.350 194.725 ;
        RECT 72.810 194.645 73.485 194.805 ;
        RECT 70.220 194.445 70.960 194.475 ;
        RECT 70.220 194.145 71.135 194.445 ;
        RECT 70.810 193.970 71.135 194.145 ;
        RECT 69.840 193.415 70.095 193.945 ;
        RECT 70.265 193.235 70.570 193.695 ;
        RECT 70.815 193.615 71.135 193.970 ;
        RECT 71.305 194.185 71.845 194.555 ;
        RECT 72.180 194.465 72.585 194.635 ;
        RECT 71.305 193.785 71.545 194.185 ;
        RECT 72.025 194.015 72.245 194.295 ;
        RECT 71.715 193.845 72.245 194.015 ;
        RECT 71.715 193.615 71.885 193.845 ;
        RECT 72.415 193.685 72.585 194.465 ;
        RECT 72.755 193.855 73.105 194.475 ;
        RECT 73.275 193.855 73.485 194.645 ;
        RECT 73.675 194.675 75.175 194.845 ;
        RECT 73.675 193.985 73.845 194.675 ;
        RECT 75.535 194.505 75.705 195.285 ;
        RECT 76.510 195.155 76.680 195.285 ;
        RECT 74.015 194.335 75.705 194.505 ;
        RECT 75.875 194.725 76.340 195.115 ;
        RECT 76.510 194.985 76.905 195.155 ;
        RECT 74.015 194.155 74.185 194.335 ;
        RECT 70.815 193.445 71.885 193.615 ;
        RECT 72.055 193.235 72.245 193.675 ;
        RECT 72.415 193.405 73.365 193.685 ;
        RECT 73.675 193.595 73.935 193.985 ;
        RECT 74.355 193.915 75.145 194.165 ;
        RECT 73.585 193.425 73.935 193.595 ;
        RECT 74.145 193.235 74.475 193.695 ;
        RECT 75.350 193.625 75.520 194.335 ;
        RECT 75.875 194.135 76.045 194.725 ;
        RECT 75.690 193.915 76.045 194.135 ;
        RECT 76.215 193.915 76.565 194.535 ;
        RECT 76.735 193.625 76.905 194.985 ;
        RECT 77.270 194.815 77.595 195.600 ;
        RECT 77.075 193.765 77.535 194.815 ;
        RECT 75.350 193.455 76.205 193.625 ;
        RECT 76.410 193.455 76.905 193.625 ;
        RECT 77.075 193.235 77.405 193.595 ;
        RECT 77.765 193.495 77.935 195.615 ;
        RECT 78.105 195.285 78.435 195.785 ;
        RECT 78.605 195.115 78.860 195.615 ;
        RECT 78.110 194.945 78.860 195.115 ;
        RECT 78.110 193.955 78.340 194.945 ;
        RECT 78.510 194.125 78.860 194.775 ;
        RECT 79.035 194.695 81.625 195.785 ;
        RECT 81.800 195.350 87.145 195.785 ;
        RECT 79.035 194.175 80.245 194.695 ;
        RECT 80.415 194.005 81.625 194.525 ;
        RECT 83.390 194.100 83.740 195.350 ;
        RECT 87.315 194.620 87.605 195.785 ;
        RECT 88.235 194.695 89.905 195.785 ;
        RECT 90.165 194.855 90.335 195.615 ;
        RECT 90.515 195.025 90.845 195.785 ;
        RECT 78.110 193.785 78.860 193.955 ;
        RECT 78.105 193.235 78.435 193.615 ;
        RECT 78.605 193.495 78.860 193.785 ;
        RECT 79.035 193.235 81.625 194.005 ;
        RECT 85.220 193.780 85.560 194.610 ;
        RECT 88.235 194.175 88.985 194.695 ;
        RECT 90.165 194.685 90.830 194.855 ;
        RECT 91.015 194.710 91.285 195.615 ;
        RECT 90.660 194.540 90.830 194.685 ;
        RECT 89.155 194.005 89.905 194.525 ;
        RECT 90.095 194.135 90.425 194.505 ;
        RECT 90.660 194.210 90.945 194.540 ;
        RECT 81.800 193.235 87.145 193.780 ;
        RECT 87.315 193.235 87.605 193.960 ;
        RECT 88.235 193.235 89.905 194.005 ;
        RECT 90.660 193.955 90.830 194.210 ;
        RECT 90.165 193.785 90.830 193.955 ;
        RECT 91.115 193.910 91.285 194.710 ;
        RECT 91.455 194.695 94.045 195.785 ;
        RECT 91.455 194.175 92.665 194.695 ;
        RECT 94.220 194.595 94.475 195.475 ;
        RECT 94.645 194.645 94.950 195.785 ;
        RECT 95.290 195.405 95.620 195.785 ;
        RECT 95.800 195.235 95.970 195.525 ;
        RECT 96.140 195.325 96.390 195.785 ;
        RECT 95.170 195.065 95.970 195.235 ;
        RECT 96.560 195.275 97.430 195.615 ;
        RECT 92.835 194.005 94.045 194.525 ;
        RECT 90.165 193.405 90.335 193.785 ;
        RECT 90.515 193.235 90.845 193.615 ;
        RECT 91.025 193.405 91.285 193.910 ;
        RECT 91.455 193.235 94.045 194.005 ;
        RECT 94.220 193.945 94.430 194.595 ;
        RECT 95.170 194.475 95.340 195.065 ;
        RECT 96.560 194.895 96.730 195.275 ;
        RECT 97.665 195.155 97.835 195.615 ;
        RECT 98.005 195.325 98.375 195.785 ;
        RECT 98.670 195.185 98.840 195.525 ;
        RECT 99.010 195.355 99.340 195.785 ;
        RECT 99.575 195.185 99.745 195.525 ;
        RECT 95.510 194.725 96.730 194.895 ;
        RECT 96.900 194.815 97.360 195.105 ;
        RECT 97.665 194.985 98.225 195.155 ;
        RECT 98.670 195.015 99.745 195.185 ;
        RECT 99.915 195.285 100.595 195.615 ;
        RECT 100.810 195.285 101.060 195.615 ;
        RECT 101.230 195.325 101.480 195.785 ;
        RECT 98.055 194.845 98.225 194.985 ;
        RECT 96.900 194.805 97.865 194.815 ;
        RECT 96.560 194.635 96.730 194.725 ;
        RECT 97.190 194.645 97.865 194.805 ;
        RECT 94.600 194.445 95.340 194.475 ;
        RECT 94.600 194.145 95.515 194.445 ;
        RECT 95.190 193.970 95.515 194.145 ;
        RECT 94.220 193.415 94.475 193.945 ;
        RECT 94.645 193.235 94.950 193.695 ;
        RECT 95.195 193.615 95.515 193.970 ;
        RECT 95.685 194.185 96.225 194.555 ;
        RECT 96.560 194.465 96.965 194.635 ;
        RECT 95.685 193.785 95.925 194.185 ;
        RECT 96.405 194.015 96.625 194.295 ;
        RECT 96.095 193.845 96.625 194.015 ;
        RECT 96.095 193.615 96.265 193.845 ;
        RECT 96.795 193.685 96.965 194.465 ;
        RECT 97.135 193.855 97.485 194.475 ;
        RECT 97.655 193.855 97.865 194.645 ;
        RECT 98.055 194.675 99.555 194.845 ;
        RECT 98.055 193.985 98.225 194.675 ;
        RECT 99.915 194.505 100.085 195.285 ;
        RECT 100.890 195.155 101.060 195.285 ;
        RECT 98.395 194.335 100.085 194.505 ;
        RECT 100.255 194.725 100.720 195.115 ;
        RECT 100.890 194.985 101.285 195.155 ;
        RECT 98.395 194.155 98.565 194.335 ;
        RECT 95.195 193.445 96.265 193.615 ;
        RECT 96.435 193.235 96.625 193.675 ;
        RECT 96.795 193.405 97.745 193.685 ;
        RECT 98.055 193.595 98.315 193.985 ;
        RECT 98.735 193.915 99.525 194.165 ;
        RECT 97.965 193.425 98.315 193.595 ;
        RECT 98.525 193.235 98.855 193.695 ;
        RECT 99.730 193.625 99.900 194.335 ;
        RECT 100.255 194.135 100.425 194.725 ;
        RECT 100.070 193.915 100.425 194.135 ;
        RECT 100.595 193.915 100.945 194.535 ;
        RECT 101.115 193.625 101.285 194.985 ;
        RECT 101.650 194.815 101.975 195.600 ;
        RECT 101.455 193.765 101.915 194.815 ;
        RECT 99.730 193.455 100.585 193.625 ;
        RECT 100.790 193.455 101.285 193.625 ;
        RECT 101.455 193.235 101.785 193.595 ;
        RECT 102.145 193.495 102.315 195.615 ;
        RECT 102.485 195.285 102.815 195.785 ;
        RECT 102.985 195.115 103.240 195.615 ;
        RECT 102.490 194.945 103.240 195.115 ;
        RECT 102.490 193.955 102.720 194.945 ;
        RECT 102.890 194.125 103.240 194.775 ;
        RECT 103.875 194.695 106.465 195.785 ;
        RECT 106.640 195.350 111.985 195.785 ;
        RECT 103.875 194.175 105.085 194.695 ;
        RECT 105.255 194.005 106.465 194.525 ;
        RECT 108.230 194.100 108.580 195.350 ;
        RECT 112.155 194.695 113.365 195.785 ;
        RECT 102.490 193.785 103.240 193.955 ;
        RECT 102.485 193.235 102.815 193.615 ;
        RECT 102.985 193.495 103.240 193.785 ;
        RECT 103.875 193.235 106.465 194.005 ;
        RECT 110.060 193.780 110.400 194.610 ;
        RECT 112.155 194.155 112.675 194.695 ;
        RECT 112.845 193.985 113.365 194.525 ;
        RECT 106.640 193.235 111.985 193.780 ;
        RECT 112.155 193.235 113.365 193.985 ;
        RECT 11.330 193.065 113.450 193.235 ;
        RECT 11.415 192.315 12.625 193.065 ;
        RECT 11.415 191.775 11.935 192.315 ;
        RECT 13.715 192.295 17.225 193.065 ;
        RECT 17.400 192.520 22.745 193.065 ;
        RECT 12.105 191.605 12.625 192.145 ;
        RECT 11.415 190.515 12.625 191.605 ;
        RECT 13.715 191.605 15.405 192.125 ;
        RECT 15.575 191.775 17.225 192.295 ;
        RECT 13.715 190.515 17.225 191.605 ;
        RECT 18.990 190.950 19.340 192.200 ;
        RECT 20.820 191.690 21.160 192.520 ;
        RECT 22.915 192.340 23.205 193.065 ;
        RECT 23.375 192.315 24.585 193.065 ;
        RECT 24.760 192.520 30.105 193.065 ;
        RECT 17.400 190.515 22.745 190.950 ;
        RECT 22.915 190.515 23.205 191.680 ;
        RECT 23.375 191.605 23.895 192.145 ;
        RECT 24.065 191.775 24.585 192.315 ;
        RECT 23.375 190.515 24.585 191.605 ;
        RECT 26.350 190.950 26.700 192.200 ;
        RECT 28.180 191.690 28.520 192.520 ;
        RECT 30.280 192.355 30.535 192.885 ;
        RECT 30.705 192.605 31.010 193.065 ;
        RECT 31.255 192.685 32.325 192.855 ;
        RECT 30.280 191.705 30.490 192.355 ;
        RECT 31.255 192.330 31.575 192.685 ;
        RECT 31.250 192.155 31.575 192.330 ;
        RECT 30.660 191.855 31.575 192.155 ;
        RECT 31.745 192.115 31.985 192.515 ;
        RECT 32.155 192.455 32.325 192.685 ;
        RECT 32.495 192.625 32.685 193.065 ;
        RECT 32.855 192.615 33.805 192.895 ;
        RECT 34.025 192.705 34.375 192.875 ;
        RECT 32.155 192.285 32.685 192.455 ;
        RECT 30.660 191.825 31.400 191.855 ;
        RECT 24.760 190.515 30.105 190.950 ;
        RECT 30.280 190.825 30.535 191.705 ;
        RECT 30.705 190.515 31.010 191.655 ;
        RECT 31.230 191.235 31.400 191.825 ;
        RECT 31.745 191.745 32.285 192.115 ;
        RECT 32.465 192.005 32.685 192.285 ;
        RECT 32.855 191.835 33.025 192.615 ;
        RECT 32.620 191.665 33.025 191.835 ;
        RECT 33.195 191.825 33.545 192.445 ;
        RECT 32.620 191.575 32.790 191.665 ;
        RECT 33.715 191.655 33.925 192.445 ;
        RECT 31.570 191.405 32.790 191.575 ;
        RECT 33.250 191.495 33.925 191.655 ;
        RECT 31.230 191.065 32.030 191.235 ;
        RECT 31.350 190.515 31.680 190.895 ;
        RECT 31.860 190.775 32.030 191.065 ;
        RECT 32.620 191.025 32.790 191.405 ;
        RECT 32.960 191.485 33.925 191.495 ;
        RECT 34.115 192.315 34.375 192.705 ;
        RECT 34.585 192.605 34.915 193.065 ;
        RECT 35.790 192.675 36.645 192.845 ;
        RECT 36.850 192.675 37.345 192.845 ;
        RECT 37.515 192.705 37.845 193.065 ;
        RECT 34.115 191.625 34.285 192.315 ;
        RECT 34.455 191.965 34.625 192.145 ;
        RECT 34.795 192.135 35.585 192.385 ;
        RECT 35.790 191.965 35.960 192.675 ;
        RECT 36.130 192.165 36.485 192.385 ;
        RECT 34.455 191.795 36.145 191.965 ;
        RECT 32.960 191.195 33.420 191.485 ;
        RECT 34.115 191.455 35.615 191.625 ;
        RECT 34.115 191.315 34.285 191.455 ;
        RECT 33.725 191.145 34.285 191.315 ;
        RECT 32.200 190.515 32.450 190.975 ;
        RECT 32.620 190.685 33.490 191.025 ;
        RECT 33.725 190.685 33.895 191.145 ;
        RECT 34.730 191.115 35.805 191.285 ;
        RECT 34.065 190.515 34.435 190.975 ;
        RECT 34.730 190.775 34.900 191.115 ;
        RECT 35.070 190.515 35.400 190.945 ;
        RECT 35.635 190.775 35.805 191.115 ;
        RECT 35.975 191.015 36.145 191.795 ;
        RECT 36.315 191.575 36.485 192.165 ;
        RECT 36.655 191.765 37.005 192.385 ;
        RECT 36.315 191.185 36.780 191.575 ;
        RECT 37.175 191.315 37.345 192.675 ;
        RECT 37.515 191.485 37.975 192.535 ;
        RECT 36.950 191.145 37.345 191.315 ;
        RECT 36.950 191.015 37.120 191.145 ;
        RECT 35.975 190.685 36.655 191.015 ;
        RECT 36.870 190.685 37.120 191.015 ;
        RECT 37.290 190.515 37.540 190.975 ;
        RECT 37.710 190.700 38.035 191.485 ;
        RECT 38.205 190.685 38.375 192.805 ;
        RECT 38.545 192.685 38.875 193.065 ;
        RECT 39.045 192.515 39.300 192.805 ;
        RECT 38.550 192.345 39.300 192.515 ;
        RECT 39.480 192.355 39.735 192.885 ;
        RECT 39.905 192.605 40.210 193.065 ;
        RECT 40.455 192.685 41.525 192.855 ;
        RECT 38.550 191.355 38.780 192.345 ;
        RECT 38.950 191.525 39.300 192.175 ;
        RECT 39.480 191.705 39.690 192.355 ;
        RECT 40.455 192.330 40.775 192.685 ;
        RECT 40.450 192.155 40.775 192.330 ;
        RECT 39.860 191.855 40.775 192.155 ;
        RECT 40.945 192.115 41.185 192.515 ;
        RECT 41.355 192.455 41.525 192.685 ;
        RECT 41.695 192.625 41.885 193.065 ;
        RECT 42.055 192.615 43.005 192.895 ;
        RECT 43.225 192.705 43.575 192.875 ;
        RECT 41.355 192.285 41.885 192.455 ;
        RECT 39.860 191.825 40.600 191.855 ;
        RECT 38.550 191.185 39.300 191.355 ;
        RECT 38.545 190.515 38.875 191.015 ;
        RECT 39.045 190.685 39.300 191.185 ;
        RECT 39.480 190.825 39.735 191.705 ;
        RECT 39.905 190.515 40.210 191.655 ;
        RECT 40.430 191.235 40.600 191.825 ;
        RECT 40.945 191.745 41.485 192.115 ;
        RECT 41.665 192.005 41.885 192.285 ;
        RECT 42.055 191.835 42.225 192.615 ;
        RECT 41.820 191.665 42.225 191.835 ;
        RECT 42.395 191.825 42.745 192.445 ;
        RECT 41.820 191.575 41.990 191.665 ;
        RECT 42.915 191.655 43.125 192.445 ;
        RECT 40.770 191.405 41.990 191.575 ;
        RECT 42.450 191.495 43.125 191.655 ;
        RECT 40.430 191.065 41.230 191.235 ;
        RECT 40.550 190.515 40.880 190.895 ;
        RECT 41.060 190.775 41.230 191.065 ;
        RECT 41.820 191.025 41.990 191.405 ;
        RECT 42.160 191.485 43.125 191.495 ;
        RECT 43.315 192.315 43.575 192.705 ;
        RECT 43.785 192.605 44.115 193.065 ;
        RECT 44.990 192.675 45.845 192.845 ;
        RECT 46.050 192.675 46.545 192.845 ;
        RECT 46.715 192.705 47.045 193.065 ;
        RECT 43.315 191.625 43.485 192.315 ;
        RECT 43.655 191.965 43.825 192.145 ;
        RECT 43.995 192.135 44.785 192.385 ;
        RECT 44.990 191.965 45.160 192.675 ;
        RECT 45.330 192.165 45.685 192.385 ;
        RECT 43.655 191.795 45.345 191.965 ;
        RECT 42.160 191.195 42.620 191.485 ;
        RECT 43.315 191.455 44.815 191.625 ;
        RECT 43.315 191.315 43.485 191.455 ;
        RECT 42.925 191.145 43.485 191.315 ;
        RECT 41.400 190.515 41.650 190.975 ;
        RECT 41.820 190.685 42.690 191.025 ;
        RECT 42.925 190.685 43.095 191.145 ;
        RECT 43.930 191.115 45.005 191.285 ;
        RECT 43.265 190.515 43.635 190.975 ;
        RECT 43.930 190.775 44.100 191.115 ;
        RECT 44.270 190.515 44.600 190.945 ;
        RECT 44.835 190.775 45.005 191.115 ;
        RECT 45.175 191.015 45.345 191.795 ;
        RECT 45.515 191.575 45.685 192.165 ;
        RECT 45.855 191.765 46.205 192.385 ;
        RECT 45.515 191.185 45.980 191.575 ;
        RECT 46.375 191.315 46.545 192.675 ;
        RECT 46.715 191.485 47.175 192.535 ;
        RECT 46.150 191.145 46.545 191.315 ;
        RECT 46.150 191.015 46.320 191.145 ;
        RECT 45.175 190.685 45.855 191.015 ;
        RECT 46.070 190.685 46.320 191.015 ;
        RECT 46.490 190.515 46.740 190.975 ;
        RECT 46.910 190.700 47.235 191.485 ;
        RECT 47.405 190.685 47.575 192.805 ;
        RECT 47.745 192.685 48.075 193.065 ;
        RECT 48.245 192.515 48.500 192.805 ;
        RECT 47.750 192.345 48.500 192.515 ;
        RECT 47.750 191.355 47.980 192.345 ;
        RECT 48.675 192.340 48.965 193.065 ;
        RECT 49.135 192.295 50.805 193.065 ;
        RECT 50.980 192.520 56.325 193.065 ;
        RECT 48.150 191.525 48.500 192.175 ;
        RECT 47.750 191.185 48.500 191.355 ;
        RECT 47.745 190.515 48.075 191.015 ;
        RECT 48.245 190.685 48.500 191.185 ;
        RECT 48.675 190.515 48.965 191.680 ;
        RECT 49.135 191.605 49.885 192.125 ;
        RECT 50.055 191.775 50.805 192.295 ;
        RECT 49.135 190.515 50.805 191.605 ;
        RECT 52.570 190.950 52.920 192.200 ;
        RECT 54.400 191.690 54.740 192.520 ;
        RECT 56.555 192.245 56.765 193.065 ;
        RECT 56.935 192.265 57.265 192.895 ;
        RECT 56.935 191.665 57.185 192.265 ;
        RECT 57.435 192.245 57.665 193.065 ;
        RECT 58.335 192.295 60.925 193.065 ;
        RECT 57.355 191.825 57.685 192.075 ;
        RECT 50.980 190.515 56.325 190.950 ;
        RECT 56.555 190.515 56.765 191.655 ;
        RECT 56.935 190.685 57.265 191.665 ;
        RECT 57.435 190.515 57.665 191.655 ;
        RECT 58.335 191.605 59.545 192.125 ;
        RECT 59.715 191.775 60.925 192.295 ;
        RECT 61.095 192.415 61.355 192.895 ;
        RECT 61.525 192.525 61.775 193.065 ;
        RECT 58.335 190.515 60.925 191.605 ;
        RECT 61.095 191.385 61.265 192.415 ;
        RECT 61.945 192.360 62.165 192.845 ;
        RECT 61.435 191.765 61.665 192.160 ;
        RECT 61.835 191.935 62.165 192.360 ;
        RECT 62.335 192.685 63.225 192.855 ;
        RECT 62.335 191.960 62.505 192.685 ;
        RECT 62.675 192.130 63.225 192.515 ;
        RECT 63.395 192.245 63.655 193.065 ;
        RECT 63.825 192.245 64.155 192.665 ;
        RECT 64.335 192.495 64.595 192.895 ;
        RECT 64.765 192.665 65.095 193.065 ;
        RECT 65.265 192.495 65.435 192.845 ;
        RECT 65.605 192.665 65.980 193.065 ;
        RECT 64.335 192.325 66.000 192.495 ;
        RECT 66.170 192.390 66.445 192.735 ;
        RECT 63.905 192.155 64.155 192.245 ;
        RECT 65.830 192.155 66.000 192.325 ;
        RECT 62.335 191.890 63.225 191.960 ;
        RECT 62.330 191.865 63.225 191.890 ;
        RECT 62.320 191.850 63.225 191.865 ;
        RECT 62.315 191.835 63.225 191.850 ;
        RECT 62.305 191.830 63.225 191.835 ;
        RECT 62.300 191.820 63.225 191.830 ;
        RECT 63.400 191.825 63.735 192.075 ;
        RECT 63.905 191.825 64.620 192.155 ;
        RECT 64.835 191.825 65.660 192.155 ;
        RECT 65.830 191.825 66.105 192.155 ;
        RECT 62.295 191.810 63.225 191.820 ;
        RECT 62.285 191.805 63.225 191.810 ;
        RECT 62.275 191.795 63.225 191.805 ;
        RECT 62.265 191.790 63.225 191.795 ;
        RECT 62.265 191.785 62.600 191.790 ;
        RECT 62.250 191.780 62.600 191.785 ;
        RECT 62.235 191.770 62.600 191.780 ;
        RECT 62.210 191.765 62.600 191.770 ;
        RECT 61.435 191.760 62.600 191.765 ;
        RECT 61.435 191.725 62.570 191.760 ;
        RECT 61.435 191.700 62.535 191.725 ;
        RECT 61.435 191.670 62.505 191.700 ;
        RECT 61.435 191.640 62.485 191.670 ;
        RECT 61.435 191.610 62.465 191.640 ;
        RECT 61.435 191.600 62.395 191.610 ;
        RECT 61.435 191.590 62.370 191.600 ;
        RECT 61.435 191.575 62.350 191.590 ;
        RECT 61.435 191.560 62.330 191.575 ;
        RECT 61.540 191.550 62.325 191.560 ;
        RECT 61.540 191.515 62.310 191.550 ;
        RECT 61.095 190.685 61.370 191.385 ;
        RECT 61.540 191.265 62.295 191.515 ;
        RECT 62.465 191.195 62.795 191.440 ;
        RECT 62.965 191.340 63.225 191.790 ;
        RECT 62.610 191.170 62.795 191.195 ;
        RECT 62.610 191.070 63.225 191.170 ;
        RECT 61.540 190.515 61.795 191.060 ;
        RECT 61.965 190.685 62.445 191.025 ;
        RECT 62.620 190.515 63.225 191.070 ;
        RECT 63.395 190.515 63.655 191.655 ;
        RECT 63.905 191.265 64.075 191.825 ;
        RECT 64.335 191.365 64.665 191.655 ;
        RECT 64.835 191.535 65.080 191.825 ;
        RECT 65.830 191.655 66.000 191.825 ;
        RECT 66.275 191.655 66.445 192.390 ;
        RECT 66.615 192.315 67.825 193.065 ;
        RECT 65.340 191.485 66.000 191.655 ;
        RECT 65.340 191.365 65.510 191.485 ;
        RECT 64.335 191.195 65.510 191.365 ;
        RECT 63.895 190.695 65.510 191.025 ;
        RECT 65.680 190.515 65.960 191.315 ;
        RECT 66.170 190.685 66.445 191.655 ;
        RECT 66.615 191.605 67.135 192.145 ;
        RECT 67.305 191.775 67.825 192.315 ;
        RECT 68.030 192.325 68.645 192.895 ;
        RECT 68.815 192.555 69.030 193.065 ;
        RECT 69.260 192.555 69.540 192.885 ;
        RECT 69.720 192.555 69.960 193.065 ;
        RECT 70.295 192.565 70.555 192.895 ;
        RECT 70.765 192.585 71.040 193.065 ;
        RECT 66.615 190.515 67.825 191.605 ;
        RECT 68.030 191.305 68.345 192.325 ;
        RECT 68.515 191.655 68.685 192.155 ;
        RECT 68.935 191.825 69.200 192.385 ;
        RECT 69.370 191.655 69.540 192.555 ;
        RECT 69.710 191.825 70.065 192.385 ;
        RECT 70.295 191.655 70.465 192.565 ;
        RECT 71.250 192.495 71.455 192.895 ;
        RECT 71.625 192.665 71.960 193.065 ;
        RECT 70.635 191.825 70.995 192.405 ;
        RECT 71.250 192.325 71.935 192.495 ;
        RECT 71.175 191.655 71.425 192.155 ;
        RECT 68.515 191.485 69.940 191.655 ;
        RECT 68.030 190.685 68.565 191.305 ;
        RECT 68.735 190.515 69.065 191.315 ;
        RECT 69.550 191.310 69.940 191.485 ;
        RECT 70.295 191.485 71.425 191.655 ;
        RECT 70.295 190.715 70.565 191.485 ;
        RECT 71.595 191.295 71.935 192.325 ;
        RECT 72.595 192.295 74.265 193.065 ;
        RECT 74.435 192.340 74.725 193.065 ;
        RECT 74.900 192.520 80.245 193.065 ;
        RECT 70.735 190.515 71.065 191.295 ;
        RECT 71.270 191.120 71.935 191.295 ;
        RECT 72.595 191.605 73.345 192.125 ;
        RECT 73.515 191.775 74.265 192.295 ;
        RECT 71.270 190.715 71.455 191.120 ;
        RECT 71.625 190.515 71.960 190.940 ;
        RECT 72.595 190.515 74.265 191.605 ;
        RECT 74.435 190.515 74.725 191.680 ;
        RECT 76.490 190.950 76.840 192.200 ;
        RECT 78.320 191.690 78.660 192.520 ;
        RECT 80.505 192.515 80.675 192.895 ;
        RECT 80.855 192.685 81.185 193.065 ;
        RECT 80.505 192.345 81.170 192.515 ;
        RECT 81.365 192.390 81.625 192.895 ;
        RECT 80.435 191.795 80.765 192.165 ;
        RECT 81.000 192.090 81.170 192.345 ;
        RECT 81.000 191.760 81.285 192.090 ;
        RECT 81.000 191.615 81.170 191.760 ;
        RECT 80.505 191.445 81.170 191.615 ;
        RECT 81.455 191.590 81.625 192.390 ;
        RECT 81.795 192.295 83.465 193.065 ;
        RECT 74.900 190.515 80.245 190.950 ;
        RECT 80.505 190.685 80.675 191.445 ;
        RECT 80.855 190.515 81.185 191.275 ;
        RECT 81.355 190.685 81.625 191.590 ;
        RECT 81.795 191.605 82.545 192.125 ;
        RECT 82.715 191.775 83.465 192.295 ;
        RECT 83.675 192.245 83.905 193.065 ;
        RECT 84.075 192.265 84.405 192.895 ;
        RECT 83.655 191.825 83.985 192.075 ;
        RECT 84.155 191.665 84.405 192.265 ;
        RECT 84.575 192.245 84.785 193.065 ;
        RECT 85.020 192.355 85.275 192.885 ;
        RECT 85.445 192.605 85.750 193.065 ;
        RECT 85.995 192.685 87.065 192.855 ;
        RECT 81.795 190.515 83.465 191.605 ;
        RECT 83.675 190.515 83.905 191.655 ;
        RECT 84.075 190.685 84.405 191.665 ;
        RECT 85.020 191.705 85.230 192.355 ;
        RECT 85.995 192.330 86.315 192.685 ;
        RECT 85.990 192.155 86.315 192.330 ;
        RECT 85.400 191.855 86.315 192.155 ;
        RECT 86.485 192.115 86.725 192.515 ;
        RECT 86.895 192.455 87.065 192.685 ;
        RECT 87.235 192.625 87.425 193.065 ;
        RECT 87.595 192.615 88.545 192.895 ;
        RECT 88.765 192.705 89.115 192.875 ;
        RECT 86.895 192.285 87.425 192.455 ;
        RECT 85.400 191.825 86.140 191.855 ;
        RECT 84.575 190.515 84.785 191.655 ;
        RECT 85.020 190.825 85.275 191.705 ;
        RECT 85.445 190.515 85.750 191.655 ;
        RECT 85.970 191.235 86.140 191.825 ;
        RECT 86.485 191.745 87.025 192.115 ;
        RECT 87.205 192.005 87.425 192.285 ;
        RECT 87.595 191.835 87.765 192.615 ;
        RECT 87.360 191.665 87.765 191.835 ;
        RECT 87.935 191.825 88.285 192.445 ;
        RECT 87.360 191.575 87.530 191.665 ;
        RECT 88.455 191.655 88.665 192.445 ;
        RECT 86.310 191.405 87.530 191.575 ;
        RECT 87.990 191.495 88.665 191.655 ;
        RECT 85.970 191.065 86.770 191.235 ;
        RECT 86.090 190.515 86.420 190.895 ;
        RECT 86.600 190.775 86.770 191.065 ;
        RECT 87.360 191.025 87.530 191.405 ;
        RECT 87.700 191.485 88.665 191.495 ;
        RECT 88.855 192.315 89.115 192.705 ;
        RECT 89.325 192.605 89.655 193.065 ;
        RECT 90.530 192.675 91.385 192.845 ;
        RECT 91.590 192.675 92.085 192.845 ;
        RECT 92.255 192.705 92.585 193.065 ;
        RECT 88.855 191.625 89.025 192.315 ;
        RECT 89.195 191.965 89.365 192.145 ;
        RECT 89.535 192.135 90.325 192.385 ;
        RECT 90.530 191.965 90.700 192.675 ;
        RECT 90.870 192.165 91.225 192.385 ;
        RECT 89.195 191.795 90.885 191.965 ;
        RECT 87.700 191.195 88.160 191.485 ;
        RECT 88.855 191.455 90.355 191.625 ;
        RECT 88.855 191.315 89.025 191.455 ;
        RECT 88.465 191.145 89.025 191.315 ;
        RECT 86.940 190.515 87.190 190.975 ;
        RECT 87.360 190.685 88.230 191.025 ;
        RECT 88.465 190.685 88.635 191.145 ;
        RECT 89.470 191.115 90.545 191.285 ;
        RECT 88.805 190.515 89.175 190.975 ;
        RECT 89.470 190.775 89.640 191.115 ;
        RECT 89.810 190.515 90.140 190.945 ;
        RECT 90.375 190.775 90.545 191.115 ;
        RECT 90.715 191.015 90.885 191.795 ;
        RECT 91.055 191.575 91.225 192.165 ;
        RECT 91.395 191.765 91.745 192.385 ;
        RECT 91.055 191.185 91.520 191.575 ;
        RECT 91.915 191.315 92.085 192.675 ;
        RECT 92.255 191.485 92.715 192.535 ;
        RECT 91.690 191.145 92.085 191.315 ;
        RECT 91.690 191.015 91.860 191.145 ;
        RECT 90.715 190.685 91.395 191.015 ;
        RECT 91.610 190.685 91.860 191.015 ;
        RECT 92.030 190.515 92.280 190.975 ;
        RECT 92.450 190.700 92.775 191.485 ;
        RECT 92.945 190.685 93.115 192.805 ;
        RECT 93.285 192.685 93.615 193.065 ;
        RECT 93.785 192.515 94.040 192.805 ;
        RECT 93.290 192.345 94.040 192.515 ;
        RECT 94.330 192.435 94.615 192.895 ;
        RECT 94.785 192.605 95.055 193.065 ;
        RECT 93.290 191.355 93.520 192.345 ;
        RECT 94.330 192.265 95.285 192.435 ;
        RECT 93.690 191.525 94.040 192.175 ;
        RECT 94.215 191.535 94.905 192.095 ;
        RECT 95.075 191.365 95.285 192.265 ;
        RECT 93.290 191.185 94.040 191.355 ;
        RECT 93.285 190.515 93.615 191.015 ;
        RECT 93.785 190.685 94.040 191.185 ;
        RECT 94.330 191.145 95.285 191.365 ;
        RECT 95.455 192.095 95.855 192.895 ;
        RECT 96.045 192.435 96.325 192.895 ;
        RECT 96.845 192.605 97.170 193.065 ;
        RECT 96.045 192.265 97.170 192.435 ;
        RECT 97.340 192.325 97.725 192.895 ;
        RECT 96.720 192.155 97.170 192.265 ;
        RECT 95.455 191.535 96.550 192.095 ;
        RECT 96.720 191.825 97.275 192.155 ;
        RECT 94.330 190.685 94.615 191.145 ;
        RECT 94.785 190.515 95.055 190.975 ;
        RECT 95.455 190.685 95.855 191.535 ;
        RECT 96.720 191.365 97.170 191.825 ;
        RECT 97.445 191.655 97.725 192.325 ;
        RECT 97.935 192.245 98.165 193.065 ;
        RECT 98.335 192.265 98.665 192.895 ;
        RECT 97.915 191.825 98.245 192.075 ;
        RECT 98.415 191.665 98.665 192.265 ;
        RECT 98.835 192.245 99.045 193.065 ;
        RECT 100.195 192.340 100.485 193.065 ;
        RECT 100.660 192.355 100.915 192.885 ;
        RECT 101.085 192.605 101.390 193.065 ;
        RECT 101.635 192.685 102.705 192.855 ;
        RECT 100.660 191.705 100.870 192.355 ;
        RECT 101.635 192.330 101.955 192.685 ;
        RECT 101.630 192.155 101.955 192.330 ;
        RECT 101.040 191.855 101.955 192.155 ;
        RECT 102.125 192.115 102.365 192.515 ;
        RECT 102.535 192.455 102.705 192.685 ;
        RECT 102.875 192.625 103.065 193.065 ;
        RECT 103.235 192.615 104.185 192.895 ;
        RECT 104.405 192.705 104.755 192.875 ;
        RECT 102.535 192.285 103.065 192.455 ;
        RECT 101.040 191.825 101.780 191.855 ;
        RECT 96.045 191.145 97.170 191.365 ;
        RECT 96.045 190.685 96.325 191.145 ;
        RECT 96.845 190.515 97.170 190.975 ;
        RECT 97.340 190.685 97.725 191.655 ;
        RECT 97.935 190.515 98.165 191.655 ;
        RECT 98.335 190.685 98.665 191.665 ;
        RECT 98.835 190.515 99.045 191.655 ;
        RECT 100.195 190.515 100.485 191.680 ;
        RECT 100.660 190.825 100.915 191.705 ;
        RECT 101.085 190.515 101.390 191.655 ;
        RECT 101.610 191.235 101.780 191.825 ;
        RECT 102.125 191.745 102.665 192.115 ;
        RECT 102.845 192.005 103.065 192.285 ;
        RECT 103.235 191.835 103.405 192.615 ;
        RECT 103.000 191.665 103.405 191.835 ;
        RECT 103.575 191.825 103.925 192.445 ;
        RECT 103.000 191.575 103.170 191.665 ;
        RECT 104.095 191.655 104.305 192.445 ;
        RECT 101.950 191.405 103.170 191.575 ;
        RECT 103.630 191.495 104.305 191.655 ;
        RECT 101.610 191.065 102.410 191.235 ;
        RECT 101.730 190.515 102.060 190.895 ;
        RECT 102.240 190.775 102.410 191.065 ;
        RECT 103.000 191.025 103.170 191.405 ;
        RECT 103.340 191.485 104.305 191.495 ;
        RECT 104.495 192.315 104.755 192.705 ;
        RECT 104.965 192.605 105.295 193.065 ;
        RECT 106.170 192.675 107.025 192.845 ;
        RECT 107.230 192.675 107.725 192.845 ;
        RECT 107.895 192.705 108.225 193.065 ;
        RECT 104.495 191.625 104.665 192.315 ;
        RECT 104.835 191.965 105.005 192.145 ;
        RECT 105.175 192.135 105.965 192.385 ;
        RECT 106.170 191.965 106.340 192.675 ;
        RECT 106.510 192.165 106.865 192.385 ;
        RECT 104.835 191.795 106.525 191.965 ;
        RECT 103.340 191.195 103.800 191.485 ;
        RECT 104.495 191.455 105.995 191.625 ;
        RECT 104.495 191.315 104.665 191.455 ;
        RECT 104.105 191.145 104.665 191.315 ;
        RECT 102.580 190.515 102.830 190.975 ;
        RECT 103.000 190.685 103.870 191.025 ;
        RECT 104.105 190.685 104.275 191.145 ;
        RECT 105.110 191.115 106.185 191.285 ;
        RECT 104.445 190.515 104.815 190.975 ;
        RECT 105.110 190.775 105.280 191.115 ;
        RECT 105.450 190.515 105.780 190.945 ;
        RECT 106.015 190.775 106.185 191.115 ;
        RECT 106.355 191.015 106.525 191.795 ;
        RECT 106.695 191.575 106.865 192.165 ;
        RECT 107.035 191.765 107.385 192.385 ;
        RECT 106.695 191.185 107.160 191.575 ;
        RECT 107.555 191.315 107.725 192.675 ;
        RECT 107.895 191.485 108.355 192.535 ;
        RECT 107.330 191.145 107.725 191.315 ;
        RECT 107.330 191.015 107.500 191.145 ;
        RECT 106.355 190.685 107.035 191.015 ;
        RECT 107.250 190.685 107.500 191.015 ;
        RECT 107.670 190.515 107.920 190.975 ;
        RECT 108.090 190.700 108.415 191.485 ;
        RECT 108.585 190.685 108.755 192.805 ;
        RECT 108.925 192.685 109.255 193.065 ;
        RECT 109.425 192.515 109.680 192.805 ;
        RECT 108.930 192.345 109.680 192.515 ;
        RECT 108.930 191.355 109.160 192.345 ;
        RECT 110.315 192.295 111.985 193.065 ;
        RECT 112.155 192.315 113.365 193.065 ;
        RECT 109.330 191.525 109.680 192.175 ;
        RECT 110.315 191.605 111.065 192.125 ;
        RECT 111.235 191.775 111.985 192.295 ;
        RECT 112.155 191.605 112.675 192.145 ;
        RECT 112.845 191.775 113.365 192.315 ;
        RECT 108.930 191.185 109.680 191.355 ;
        RECT 108.925 190.515 109.255 191.015 ;
        RECT 109.425 190.685 109.680 191.185 ;
        RECT 110.315 190.515 111.985 191.605 ;
        RECT 112.155 190.515 113.365 191.605 ;
        RECT 11.330 190.345 113.450 190.515 ;
        RECT 11.415 189.255 12.625 190.345 ;
        RECT 11.415 188.545 11.935 189.085 ;
        RECT 12.105 188.715 12.625 189.255 ;
        RECT 13.255 189.255 16.765 190.345 ;
        RECT 16.940 189.910 22.285 190.345 ;
        RECT 13.255 188.735 14.945 189.255 ;
        RECT 15.115 188.565 16.765 189.085 ;
        RECT 18.530 188.660 18.880 189.910 ;
        RECT 22.460 189.675 22.715 190.175 ;
        RECT 22.885 189.845 23.215 190.345 ;
        RECT 22.460 189.505 23.210 189.675 ;
        RECT 11.415 187.795 12.625 188.545 ;
        RECT 13.255 187.795 16.765 188.565 ;
        RECT 20.360 188.340 20.700 189.170 ;
        RECT 22.460 188.685 22.810 189.335 ;
        RECT 22.980 188.515 23.210 189.505 ;
        RECT 22.460 188.345 23.210 188.515 ;
        RECT 16.940 187.795 22.285 188.340 ;
        RECT 22.460 188.055 22.715 188.345 ;
        RECT 22.885 187.795 23.215 188.175 ;
        RECT 23.385 188.055 23.555 190.175 ;
        RECT 23.725 189.375 24.050 190.160 ;
        RECT 24.220 189.885 24.470 190.345 ;
        RECT 24.640 189.845 24.890 190.175 ;
        RECT 25.105 189.845 25.785 190.175 ;
        RECT 24.640 189.715 24.810 189.845 ;
        RECT 24.415 189.545 24.810 189.715 ;
        RECT 23.785 188.325 24.245 189.375 ;
        RECT 24.415 188.185 24.585 189.545 ;
        RECT 24.980 189.285 25.445 189.675 ;
        RECT 24.755 188.475 25.105 189.095 ;
        RECT 25.275 188.695 25.445 189.285 ;
        RECT 25.615 189.065 25.785 189.845 ;
        RECT 25.955 189.745 26.125 190.085 ;
        RECT 26.360 189.915 26.690 190.345 ;
        RECT 26.860 189.745 27.030 190.085 ;
        RECT 27.325 189.885 27.695 190.345 ;
        RECT 25.955 189.575 27.030 189.745 ;
        RECT 27.865 189.715 28.035 190.175 ;
        RECT 28.270 189.835 29.140 190.175 ;
        RECT 29.310 189.885 29.560 190.345 ;
        RECT 27.475 189.545 28.035 189.715 ;
        RECT 27.475 189.405 27.645 189.545 ;
        RECT 26.145 189.235 27.645 189.405 ;
        RECT 28.340 189.375 28.800 189.665 ;
        RECT 25.615 188.895 27.305 189.065 ;
        RECT 25.275 188.475 25.630 188.695 ;
        RECT 25.800 188.185 25.970 188.895 ;
        RECT 26.175 188.475 26.965 188.725 ;
        RECT 27.135 188.715 27.305 188.895 ;
        RECT 27.475 188.545 27.645 189.235 ;
        RECT 23.915 187.795 24.245 188.155 ;
        RECT 24.415 188.015 24.910 188.185 ;
        RECT 25.115 188.015 25.970 188.185 ;
        RECT 26.845 187.795 27.175 188.255 ;
        RECT 27.385 188.155 27.645 188.545 ;
        RECT 27.835 189.365 28.800 189.375 ;
        RECT 28.970 189.455 29.140 189.835 ;
        RECT 29.730 189.795 29.900 190.085 ;
        RECT 30.080 189.965 30.410 190.345 ;
        RECT 29.730 189.625 30.530 189.795 ;
        RECT 27.835 189.205 28.510 189.365 ;
        RECT 28.970 189.285 30.190 189.455 ;
        RECT 27.835 188.415 28.045 189.205 ;
        RECT 28.970 189.195 29.140 189.285 ;
        RECT 28.215 188.415 28.565 189.035 ;
        RECT 28.735 189.025 29.140 189.195 ;
        RECT 28.735 188.245 28.905 189.025 ;
        RECT 29.075 188.575 29.295 188.855 ;
        RECT 29.475 188.745 30.015 189.115 ;
        RECT 30.360 189.035 30.530 189.625 ;
        RECT 30.750 189.205 31.055 190.345 ;
        RECT 31.225 189.155 31.480 190.035 ;
        RECT 30.360 189.005 31.100 189.035 ;
        RECT 29.075 188.405 29.605 188.575 ;
        RECT 27.385 187.985 27.735 188.155 ;
        RECT 27.955 187.965 28.905 188.245 ;
        RECT 29.075 187.795 29.265 188.235 ;
        RECT 29.435 188.175 29.605 188.405 ;
        RECT 29.775 188.345 30.015 188.745 ;
        RECT 30.185 188.705 31.100 189.005 ;
        RECT 30.185 188.530 30.510 188.705 ;
        RECT 30.185 188.175 30.505 188.530 ;
        RECT 31.270 188.505 31.480 189.155 ;
        RECT 31.655 189.585 32.170 189.995 ;
        RECT 32.405 189.585 32.575 190.345 ;
        RECT 32.745 190.005 34.775 190.175 ;
        RECT 31.655 188.775 31.995 189.585 ;
        RECT 32.745 189.340 32.915 190.005 ;
        RECT 33.310 189.665 34.435 189.835 ;
        RECT 32.165 189.150 32.915 189.340 ;
        RECT 33.085 189.325 34.095 189.495 ;
        RECT 31.655 188.605 32.885 188.775 ;
        RECT 29.435 188.005 30.505 188.175 ;
        RECT 30.750 187.795 31.055 188.255 ;
        RECT 31.225 187.975 31.480 188.505 ;
        RECT 31.930 188.000 32.175 188.605 ;
        RECT 32.395 187.795 32.905 188.330 ;
        RECT 33.085 187.965 33.275 189.325 ;
        RECT 33.445 188.305 33.720 189.125 ;
        RECT 33.925 188.525 34.095 189.325 ;
        RECT 34.265 188.535 34.435 189.665 ;
        RECT 34.605 189.035 34.775 190.005 ;
        RECT 34.945 189.205 35.115 190.345 ;
        RECT 35.285 189.205 35.620 190.175 ;
        RECT 34.605 188.705 34.800 189.035 ;
        RECT 35.025 188.705 35.280 189.035 ;
        RECT 35.025 188.535 35.195 188.705 ;
        RECT 35.450 188.535 35.620 189.205 ;
        RECT 35.795 189.180 36.085 190.345 ;
        RECT 36.255 189.255 37.925 190.345 ;
        RECT 36.255 188.735 37.005 189.255 ;
        RECT 38.155 189.205 38.365 190.345 ;
        RECT 38.535 189.195 38.865 190.175 ;
        RECT 39.035 189.205 39.265 190.345 ;
        RECT 39.590 189.715 39.875 190.175 ;
        RECT 40.045 189.885 40.315 190.345 ;
        RECT 39.590 189.495 40.545 189.715 ;
        RECT 37.175 188.565 37.925 189.085 ;
        RECT 34.265 188.365 35.195 188.535 ;
        RECT 34.265 188.330 34.440 188.365 ;
        RECT 33.445 188.135 33.725 188.305 ;
        RECT 33.445 187.965 33.720 188.135 ;
        RECT 33.910 187.965 34.440 188.330 ;
        RECT 34.865 187.795 35.195 188.195 ;
        RECT 35.365 187.965 35.620 188.535 ;
        RECT 35.795 187.795 36.085 188.520 ;
        RECT 36.255 187.795 37.925 188.565 ;
        RECT 38.155 187.795 38.365 188.615 ;
        RECT 38.535 188.595 38.785 189.195 ;
        RECT 38.955 188.785 39.285 189.035 ;
        RECT 39.475 188.765 40.165 189.325 ;
        RECT 38.535 187.965 38.865 188.595 ;
        RECT 39.035 187.795 39.265 188.615 ;
        RECT 40.335 188.595 40.545 189.495 ;
        RECT 39.590 188.425 40.545 188.595 ;
        RECT 40.715 189.325 41.115 190.175 ;
        RECT 41.305 189.715 41.585 190.175 ;
        RECT 42.105 189.885 42.430 190.345 ;
        RECT 41.305 189.495 42.430 189.715 ;
        RECT 40.715 188.765 41.810 189.325 ;
        RECT 41.980 189.035 42.430 189.495 ;
        RECT 42.600 189.205 42.985 190.175 ;
        RECT 43.245 189.415 43.415 190.175 ;
        RECT 43.595 189.585 43.925 190.345 ;
        RECT 43.245 189.245 43.910 189.415 ;
        RECT 44.095 189.270 44.365 190.175 ;
        RECT 39.590 187.965 39.875 188.425 ;
        RECT 40.045 187.795 40.315 188.255 ;
        RECT 40.715 187.965 41.115 188.765 ;
        RECT 41.980 188.705 42.535 189.035 ;
        RECT 41.980 188.595 42.430 188.705 ;
        RECT 41.305 188.425 42.430 188.595 ;
        RECT 42.705 188.535 42.985 189.205 ;
        RECT 43.740 189.100 43.910 189.245 ;
        RECT 43.175 188.695 43.505 189.065 ;
        RECT 43.740 188.770 44.025 189.100 ;
        RECT 41.305 187.965 41.585 188.425 ;
        RECT 42.105 187.795 42.430 188.255 ;
        RECT 42.600 187.965 42.985 188.535 ;
        RECT 43.740 188.515 43.910 188.770 ;
        RECT 43.245 188.345 43.910 188.515 ;
        RECT 44.195 188.470 44.365 189.270 ;
        RECT 43.245 187.965 43.415 188.345 ;
        RECT 43.595 187.795 43.925 188.175 ;
        RECT 44.105 187.965 44.365 188.470 ;
        RECT 44.540 189.155 44.795 190.035 ;
        RECT 44.965 189.205 45.270 190.345 ;
        RECT 45.610 189.965 45.940 190.345 ;
        RECT 46.120 189.795 46.290 190.085 ;
        RECT 46.460 189.885 46.710 190.345 ;
        RECT 45.490 189.625 46.290 189.795 ;
        RECT 46.880 189.835 47.750 190.175 ;
        RECT 44.540 188.505 44.750 189.155 ;
        RECT 45.490 189.035 45.660 189.625 ;
        RECT 46.880 189.455 47.050 189.835 ;
        RECT 47.985 189.715 48.155 190.175 ;
        RECT 48.325 189.885 48.695 190.345 ;
        RECT 48.990 189.745 49.160 190.085 ;
        RECT 49.330 189.915 49.660 190.345 ;
        RECT 49.895 189.745 50.065 190.085 ;
        RECT 45.830 189.285 47.050 189.455 ;
        RECT 47.220 189.375 47.680 189.665 ;
        RECT 47.985 189.545 48.545 189.715 ;
        RECT 48.990 189.575 50.065 189.745 ;
        RECT 50.235 189.845 50.915 190.175 ;
        RECT 51.130 189.845 51.380 190.175 ;
        RECT 51.550 189.885 51.800 190.345 ;
        RECT 48.375 189.405 48.545 189.545 ;
        RECT 47.220 189.365 48.185 189.375 ;
        RECT 46.880 189.195 47.050 189.285 ;
        RECT 47.510 189.205 48.185 189.365 ;
        RECT 44.920 189.005 45.660 189.035 ;
        RECT 44.920 188.705 45.835 189.005 ;
        RECT 45.510 188.530 45.835 188.705 ;
        RECT 44.540 187.975 44.795 188.505 ;
        RECT 44.965 187.795 45.270 188.255 ;
        RECT 45.515 188.175 45.835 188.530 ;
        RECT 46.005 188.745 46.545 189.115 ;
        RECT 46.880 189.025 47.285 189.195 ;
        RECT 46.005 188.345 46.245 188.745 ;
        RECT 46.725 188.575 46.945 188.855 ;
        RECT 46.415 188.405 46.945 188.575 ;
        RECT 46.415 188.175 46.585 188.405 ;
        RECT 47.115 188.245 47.285 189.025 ;
        RECT 47.455 188.415 47.805 189.035 ;
        RECT 47.975 188.415 48.185 189.205 ;
        RECT 48.375 189.235 49.875 189.405 ;
        RECT 48.375 188.545 48.545 189.235 ;
        RECT 50.235 189.065 50.405 189.845 ;
        RECT 51.210 189.715 51.380 189.845 ;
        RECT 48.715 188.895 50.405 189.065 ;
        RECT 50.575 189.285 51.040 189.675 ;
        RECT 51.210 189.545 51.605 189.715 ;
        RECT 48.715 188.715 48.885 188.895 ;
        RECT 45.515 188.005 46.585 188.175 ;
        RECT 46.755 187.795 46.945 188.235 ;
        RECT 47.115 187.965 48.065 188.245 ;
        RECT 48.375 188.155 48.635 188.545 ;
        RECT 49.055 188.475 49.845 188.725 ;
        RECT 48.285 187.985 48.635 188.155 ;
        RECT 48.845 187.795 49.175 188.255 ;
        RECT 50.050 188.185 50.220 188.895 ;
        RECT 50.575 188.695 50.745 189.285 ;
        RECT 50.390 188.475 50.745 188.695 ;
        RECT 50.915 188.475 51.265 189.095 ;
        RECT 51.435 188.185 51.605 189.545 ;
        RECT 51.970 189.375 52.295 190.160 ;
        RECT 51.775 188.325 52.235 189.375 ;
        RECT 50.050 188.015 50.905 188.185 ;
        RECT 51.110 188.015 51.605 188.185 ;
        RECT 51.775 187.795 52.105 188.155 ;
        RECT 52.465 188.055 52.635 190.175 ;
        RECT 52.805 189.845 53.135 190.345 ;
        RECT 53.305 189.675 53.560 190.175 ;
        RECT 54.215 189.835 54.515 190.345 ;
        RECT 54.685 189.835 55.065 190.005 ;
        RECT 55.645 189.835 56.275 190.345 ;
        RECT 52.810 189.505 53.560 189.675 ;
        RECT 54.685 189.665 54.855 189.835 ;
        RECT 56.445 189.665 56.775 190.175 ;
        RECT 56.945 189.835 57.245 190.345 ;
        RECT 52.810 188.515 53.040 189.505 ;
        RECT 54.195 189.465 54.855 189.665 ;
        RECT 55.025 189.495 57.245 189.665 ;
        RECT 53.210 188.685 53.560 189.335 ;
        RECT 54.195 188.535 54.365 189.465 ;
        RECT 55.025 189.295 55.195 189.495 ;
        RECT 54.535 189.125 55.195 189.295 ;
        RECT 55.365 189.155 56.905 189.325 ;
        RECT 54.535 188.705 54.705 189.125 ;
        RECT 55.365 188.955 55.535 189.155 ;
        RECT 54.935 188.785 55.535 188.955 ;
        RECT 55.705 188.785 56.400 188.985 ;
        RECT 56.660 188.705 56.905 189.155 ;
        RECT 55.025 188.535 55.935 188.615 ;
        RECT 52.810 188.345 53.560 188.515 ;
        RECT 52.805 187.795 53.135 188.175 ;
        RECT 53.305 188.055 53.560 188.345 ;
        RECT 54.195 188.055 54.515 188.535 ;
        RECT 54.685 188.445 55.935 188.535 ;
        RECT 54.685 188.365 55.195 188.445 ;
        RECT 54.685 187.965 54.915 188.365 ;
        RECT 55.085 187.795 55.435 188.185 ;
        RECT 55.605 187.965 55.935 188.445 ;
        RECT 56.105 187.795 56.275 188.615 ;
        RECT 57.075 188.535 57.245 189.495 ;
        RECT 56.780 187.990 57.245 188.535 ;
        RECT 57.415 189.205 57.800 190.175 ;
        RECT 57.970 189.885 58.295 190.345 ;
        RECT 58.815 189.715 59.095 190.175 ;
        RECT 57.970 189.495 59.095 189.715 ;
        RECT 57.415 188.535 57.695 189.205 ;
        RECT 57.970 189.035 58.420 189.495 ;
        RECT 59.285 189.325 59.685 190.175 ;
        RECT 60.085 189.885 60.355 190.345 ;
        RECT 60.525 189.715 60.810 190.175 ;
        RECT 57.865 188.705 58.420 189.035 ;
        RECT 58.590 188.765 59.685 189.325 ;
        RECT 57.970 188.595 58.420 188.705 ;
        RECT 57.415 187.965 57.800 188.535 ;
        RECT 57.970 188.425 59.095 188.595 ;
        RECT 57.970 187.795 58.295 188.255 ;
        RECT 58.815 187.965 59.095 188.425 ;
        RECT 59.285 187.965 59.685 188.765 ;
        RECT 59.855 189.495 60.810 189.715 ;
        RECT 59.855 188.595 60.065 189.495 ;
        RECT 60.235 188.765 60.925 189.325 ;
        RECT 61.555 189.180 61.845 190.345 ;
        RECT 62.015 189.205 62.275 190.345 ;
        RECT 62.515 189.835 64.130 190.165 ;
        RECT 62.525 189.035 62.695 189.595 ;
        RECT 62.955 189.495 64.130 189.665 ;
        RECT 64.300 189.545 64.580 190.345 ;
        RECT 62.955 189.205 63.285 189.495 ;
        RECT 63.960 189.375 64.130 189.495 ;
        RECT 63.455 189.035 63.700 189.325 ;
        RECT 63.960 189.205 64.620 189.375 ;
        RECT 64.790 189.205 65.065 190.175 ;
        RECT 65.235 189.205 65.495 190.345 ;
        RECT 65.665 189.375 65.995 190.175 ;
        RECT 66.165 189.545 66.335 190.345 ;
        RECT 66.535 189.375 66.865 190.175 ;
        RECT 67.065 189.545 67.345 190.345 ;
        RECT 67.535 189.790 68.140 190.345 ;
        RECT 68.315 189.835 68.795 190.175 ;
        RECT 68.965 189.800 69.220 190.345 ;
        RECT 67.535 189.690 68.150 189.790 ;
        RECT 67.965 189.665 68.150 189.690 ;
        RECT 65.665 189.205 66.945 189.375 ;
        RECT 64.450 189.035 64.620 189.205 ;
        RECT 62.020 188.785 62.355 189.035 ;
        RECT 62.525 188.705 63.240 189.035 ;
        RECT 63.455 188.705 64.280 189.035 ;
        RECT 64.450 188.705 64.725 189.035 ;
        RECT 62.525 188.615 62.775 188.705 ;
        RECT 59.855 188.425 60.810 188.595 ;
        RECT 60.085 187.795 60.355 188.255 ;
        RECT 60.525 187.965 60.810 188.425 ;
        RECT 61.555 187.795 61.845 188.520 ;
        RECT 62.015 187.795 62.275 188.615 ;
        RECT 62.445 188.195 62.775 188.615 ;
        RECT 64.450 188.535 64.620 188.705 ;
        RECT 62.955 188.365 64.620 188.535 ;
        RECT 64.895 188.470 65.065 189.205 ;
        RECT 65.260 188.705 65.545 189.035 ;
        RECT 65.745 188.705 66.125 189.035 ;
        RECT 66.295 188.705 66.605 189.035 ;
        RECT 62.955 187.965 63.215 188.365 ;
        RECT 63.385 187.795 63.715 188.195 ;
        RECT 63.885 188.015 64.055 188.365 ;
        RECT 64.225 187.795 64.600 188.195 ;
        RECT 64.790 188.125 65.065 188.470 ;
        RECT 65.240 187.795 65.575 188.535 ;
        RECT 65.745 188.010 65.960 188.705 ;
        RECT 66.295 188.535 66.500 188.705 ;
        RECT 66.775 188.535 66.945 189.205 ;
        RECT 67.125 188.705 67.365 189.375 ;
        RECT 67.535 189.070 67.795 189.520 ;
        RECT 67.965 189.420 68.295 189.665 ;
        RECT 68.465 189.345 69.220 189.595 ;
        RECT 69.390 189.475 69.665 190.175 ;
        RECT 69.840 189.910 75.185 190.345 ;
        RECT 68.450 189.310 69.220 189.345 ;
        RECT 68.435 189.300 69.220 189.310 ;
        RECT 68.430 189.285 69.325 189.300 ;
        RECT 68.410 189.270 69.325 189.285 ;
        RECT 68.390 189.260 69.325 189.270 ;
        RECT 68.365 189.250 69.325 189.260 ;
        RECT 68.295 189.220 69.325 189.250 ;
        RECT 68.275 189.190 69.325 189.220 ;
        RECT 68.255 189.160 69.325 189.190 ;
        RECT 68.225 189.135 69.325 189.160 ;
        RECT 68.190 189.100 69.325 189.135 ;
        RECT 68.160 189.095 69.325 189.100 ;
        RECT 68.160 189.090 68.550 189.095 ;
        RECT 68.160 189.080 68.525 189.090 ;
        RECT 68.160 189.075 68.510 189.080 ;
        RECT 68.160 189.070 68.495 189.075 ;
        RECT 67.535 189.065 68.495 189.070 ;
        RECT 67.535 189.055 68.485 189.065 ;
        RECT 67.535 189.050 68.475 189.055 ;
        RECT 67.535 189.040 68.465 189.050 ;
        RECT 67.535 189.030 68.460 189.040 ;
        RECT 67.535 189.025 68.455 189.030 ;
        RECT 67.535 189.010 68.445 189.025 ;
        RECT 67.535 188.995 68.440 189.010 ;
        RECT 67.535 188.970 68.430 188.995 ;
        RECT 67.535 188.900 68.425 188.970 ;
        RECT 66.150 188.010 66.500 188.535 ;
        RECT 66.670 187.965 67.365 188.535 ;
        RECT 67.535 188.345 68.085 188.730 ;
        RECT 68.255 188.175 68.425 188.900 ;
        RECT 67.535 188.005 68.425 188.175 ;
        RECT 68.595 188.500 68.925 188.925 ;
        RECT 69.095 188.700 69.325 189.095 ;
        RECT 68.595 188.015 68.815 188.500 ;
        RECT 69.495 188.445 69.665 189.475 ;
        RECT 71.430 188.660 71.780 189.910 ;
        RECT 75.730 189.365 75.985 190.035 ;
        RECT 76.165 189.545 76.450 190.345 ;
        RECT 76.630 189.625 76.960 190.135 ;
        RECT 68.985 187.795 69.235 188.335 ;
        RECT 69.405 187.965 69.665 188.445 ;
        RECT 73.260 188.340 73.600 189.170 ;
        RECT 75.730 188.505 75.910 189.365 ;
        RECT 76.630 189.035 76.880 189.625 ;
        RECT 77.230 189.475 77.400 190.085 ;
        RECT 77.570 189.655 77.900 190.345 ;
        RECT 78.130 189.795 78.370 190.085 ;
        RECT 78.570 189.965 78.990 190.345 ;
        RECT 79.170 189.875 79.800 190.125 ;
        RECT 80.270 189.965 80.600 190.345 ;
        RECT 79.170 189.795 79.340 189.875 ;
        RECT 80.770 189.795 80.940 190.085 ;
        RECT 81.120 189.965 81.500 190.345 ;
        RECT 81.740 189.960 82.570 190.130 ;
        RECT 78.130 189.625 79.340 189.795 ;
        RECT 76.080 188.705 76.880 189.035 ;
        RECT 69.840 187.795 75.185 188.340 ;
        RECT 75.730 188.305 75.985 188.505 ;
        RECT 75.645 188.135 75.985 188.305 ;
        RECT 75.730 187.975 75.985 188.135 ;
        RECT 76.165 187.795 76.450 188.255 ;
        RECT 76.630 188.055 76.880 188.705 ;
        RECT 77.080 189.455 77.400 189.475 ;
        RECT 77.080 189.285 79.000 189.455 ;
        RECT 77.080 188.390 77.270 189.285 ;
        RECT 79.170 189.115 79.340 189.625 ;
        RECT 79.510 189.365 80.030 189.675 ;
        RECT 77.440 188.945 79.340 189.115 ;
        RECT 77.440 188.885 77.770 188.945 ;
        RECT 77.920 188.715 78.250 188.775 ;
        RECT 77.590 188.445 78.250 188.715 ;
        RECT 77.080 188.060 77.400 188.390 ;
        RECT 77.580 187.795 78.240 188.275 ;
        RECT 78.440 188.185 78.610 188.945 ;
        RECT 79.510 188.775 79.690 189.185 ;
        RECT 78.780 188.605 79.110 188.725 ;
        RECT 79.860 188.605 80.030 189.365 ;
        RECT 78.780 188.435 80.030 188.605 ;
        RECT 80.200 189.545 81.570 189.795 ;
        RECT 80.200 188.775 80.390 189.545 ;
        RECT 81.320 189.285 81.570 189.545 ;
        RECT 80.560 189.115 80.810 189.275 ;
        RECT 81.740 189.115 81.910 189.960 ;
        RECT 82.805 189.675 82.975 190.175 ;
        RECT 83.145 189.845 83.475 190.345 ;
        RECT 82.080 189.285 82.580 189.665 ;
        RECT 82.805 189.505 83.500 189.675 ;
        RECT 80.560 188.945 81.910 189.115 ;
        RECT 81.490 188.905 81.910 188.945 ;
        RECT 80.200 188.435 80.620 188.775 ;
        RECT 80.910 188.445 81.320 188.775 ;
        RECT 78.440 188.015 79.290 188.185 ;
        RECT 79.850 187.795 80.170 188.255 ;
        RECT 80.370 188.005 80.620 188.435 ;
        RECT 80.910 187.795 81.320 188.235 ;
        RECT 81.490 188.175 81.660 188.905 ;
        RECT 81.830 188.355 82.180 188.725 ;
        RECT 82.360 188.415 82.580 189.285 ;
        RECT 82.750 188.715 83.160 189.335 ;
        RECT 83.330 188.535 83.500 189.505 ;
        RECT 82.805 188.345 83.500 188.535 ;
        RECT 81.490 187.975 82.505 188.175 ;
        RECT 82.805 188.015 82.975 188.345 ;
        RECT 83.145 187.795 83.475 188.175 ;
        RECT 83.690 188.055 83.915 190.175 ;
        RECT 84.085 189.845 84.415 190.345 ;
        RECT 84.585 189.675 84.755 190.175 ;
        RECT 84.090 189.505 84.755 189.675 ;
        RECT 84.090 188.515 84.320 189.505 ;
        RECT 84.490 188.685 84.840 189.335 ;
        RECT 85.475 189.255 87.145 190.345 ;
        RECT 85.475 188.735 86.225 189.255 ;
        RECT 87.315 189.180 87.605 190.345 ;
        RECT 87.775 189.585 88.290 189.995 ;
        RECT 88.525 189.585 88.695 190.345 ;
        RECT 88.865 190.005 90.895 190.175 ;
        RECT 86.395 188.565 87.145 189.085 ;
        RECT 87.775 188.775 88.115 189.585 ;
        RECT 88.865 189.340 89.035 190.005 ;
        RECT 89.430 189.665 90.555 189.835 ;
        RECT 88.285 189.150 89.035 189.340 ;
        RECT 89.205 189.325 90.215 189.495 ;
        RECT 87.775 188.605 89.005 188.775 ;
        RECT 84.090 188.345 84.755 188.515 ;
        RECT 84.085 187.795 84.415 188.175 ;
        RECT 84.585 188.055 84.755 188.345 ;
        RECT 85.475 187.795 87.145 188.565 ;
        RECT 87.315 187.795 87.605 188.520 ;
        RECT 88.050 188.000 88.295 188.605 ;
        RECT 88.515 187.795 89.025 188.330 ;
        RECT 89.205 187.965 89.395 189.325 ;
        RECT 89.565 188.645 89.840 189.125 ;
        RECT 89.565 188.475 89.845 188.645 ;
        RECT 90.045 188.525 90.215 189.325 ;
        RECT 90.385 188.535 90.555 189.665 ;
        RECT 90.725 189.035 90.895 190.005 ;
        RECT 91.065 189.205 91.235 190.345 ;
        RECT 91.405 189.205 91.740 190.175 ;
        RECT 90.725 188.705 90.920 189.035 ;
        RECT 91.145 188.705 91.400 189.035 ;
        RECT 91.145 188.535 91.315 188.705 ;
        RECT 91.570 188.535 91.740 189.205 ;
        RECT 91.915 189.255 93.585 190.345 ;
        RECT 91.915 188.735 92.665 189.255 ;
        RECT 93.795 189.205 94.025 190.345 ;
        RECT 94.195 189.195 94.525 190.175 ;
        RECT 94.695 189.205 94.905 190.345 ;
        RECT 95.135 189.585 95.650 189.995 ;
        RECT 95.885 189.585 96.055 190.345 ;
        RECT 96.225 190.005 98.255 190.175 ;
        RECT 92.835 188.565 93.585 189.085 ;
        RECT 93.775 188.785 94.105 189.035 ;
        RECT 89.565 187.965 89.840 188.475 ;
        RECT 90.385 188.365 91.315 188.535 ;
        RECT 90.385 188.330 90.560 188.365 ;
        RECT 90.030 187.965 90.560 188.330 ;
        RECT 90.985 187.795 91.315 188.195 ;
        RECT 91.485 187.965 91.740 188.535 ;
        RECT 91.915 187.795 93.585 188.565 ;
        RECT 93.795 187.795 94.025 188.615 ;
        RECT 94.275 188.595 94.525 189.195 ;
        RECT 95.135 188.775 95.475 189.585 ;
        RECT 96.225 189.340 96.395 190.005 ;
        RECT 96.790 189.665 97.915 189.835 ;
        RECT 95.645 189.150 96.395 189.340 ;
        RECT 96.565 189.325 97.575 189.495 ;
        RECT 94.195 187.965 94.525 188.595 ;
        RECT 94.695 187.795 94.905 188.615 ;
        RECT 95.135 188.605 96.365 188.775 ;
        RECT 95.410 188.000 95.655 188.605 ;
        RECT 95.875 187.795 96.385 188.330 ;
        RECT 96.565 187.965 96.755 189.325 ;
        RECT 96.925 188.305 97.200 189.125 ;
        RECT 97.405 188.525 97.575 189.325 ;
        RECT 97.745 188.535 97.915 189.665 ;
        RECT 98.085 189.035 98.255 190.005 ;
        RECT 98.425 189.205 98.595 190.345 ;
        RECT 98.765 189.205 99.100 190.175 ;
        RECT 98.085 188.705 98.280 189.035 ;
        RECT 98.505 188.705 98.760 189.035 ;
        RECT 98.505 188.535 98.675 188.705 ;
        RECT 98.930 188.535 99.100 189.205 ;
        RECT 99.275 189.585 99.790 189.995 ;
        RECT 100.025 189.585 100.195 190.345 ;
        RECT 100.365 190.005 102.395 190.175 ;
        RECT 99.275 188.775 99.615 189.585 ;
        RECT 100.365 189.340 100.535 190.005 ;
        RECT 100.930 189.665 102.055 189.835 ;
        RECT 99.785 189.150 100.535 189.340 ;
        RECT 100.705 189.325 101.715 189.495 ;
        RECT 99.275 188.605 100.505 188.775 ;
        RECT 97.745 188.365 98.675 188.535 ;
        RECT 97.745 188.330 97.920 188.365 ;
        RECT 96.925 188.135 97.205 188.305 ;
        RECT 96.925 187.965 97.200 188.135 ;
        RECT 97.390 187.965 97.920 188.330 ;
        RECT 98.345 187.795 98.675 188.195 ;
        RECT 98.845 187.965 99.100 188.535 ;
        RECT 99.550 188.000 99.795 188.605 ;
        RECT 100.015 187.795 100.525 188.330 ;
        RECT 100.705 187.965 100.895 189.325 ;
        RECT 101.065 188.985 101.340 189.125 ;
        RECT 101.065 188.815 101.345 188.985 ;
        RECT 101.065 187.965 101.340 188.815 ;
        RECT 101.545 188.525 101.715 189.325 ;
        RECT 101.885 188.535 102.055 189.665 ;
        RECT 102.225 189.035 102.395 190.005 ;
        RECT 102.565 189.205 102.735 190.345 ;
        RECT 102.905 189.205 103.240 190.175 ;
        RECT 103.965 189.415 104.135 190.175 ;
        RECT 104.315 189.585 104.645 190.345 ;
        RECT 103.965 189.245 104.630 189.415 ;
        RECT 104.815 189.270 105.085 190.175 ;
        RECT 102.225 188.705 102.420 189.035 ;
        RECT 102.645 188.705 102.900 189.035 ;
        RECT 102.645 188.535 102.815 188.705 ;
        RECT 103.070 188.535 103.240 189.205 ;
        RECT 104.460 189.100 104.630 189.245 ;
        RECT 103.895 188.695 104.225 189.065 ;
        RECT 104.460 188.770 104.745 189.100 ;
        RECT 101.885 188.365 102.815 188.535 ;
        RECT 101.885 188.330 102.060 188.365 ;
        RECT 101.530 187.965 102.060 188.330 ;
        RECT 102.485 187.795 102.815 188.195 ;
        RECT 102.985 187.965 103.240 188.535 ;
        RECT 104.460 188.515 104.630 188.770 ;
        RECT 103.965 188.345 104.630 188.515 ;
        RECT 104.915 188.470 105.085 189.270 ;
        RECT 105.255 189.255 106.465 190.345 ;
        RECT 106.640 189.910 111.985 190.345 ;
        RECT 105.255 188.715 105.775 189.255 ;
        RECT 105.945 188.545 106.465 189.085 ;
        RECT 108.230 188.660 108.580 189.910 ;
        RECT 112.155 189.255 113.365 190.345 ;
        RECT 103.965 187.965 104.135 188.345 ;
        RECT 104.315 187.795 104.645 188.175 ;
        RECT 104.825 187.965 105.085 188.470 ;
        RECT 105.255 187.795 106.465 188.545 ;
        RECT 110.060 188.340 110.400 189.170 ;
        RECT 112.155 188.715 112.675 189.255 ;
        RECT 112.845 188.545 113.365 189.085 ;
        RECT 106.640 187.795 111.985 188.340 ;
        RECT 112.155 187.795 113.365 188.545 ;
        RECT 11.330 187.625 113.450 187.795 ;
        RECT 11.415 186.875 12.625 187.625 ;
        RECT 11.415 186.335 11.935 186.875 ;
        RECT 13.715 186.855 17.225 187.625 ;
        RECT 17.400 187.080 22.745 187.625 ;
        RECT 12.105 186.165 12.625 186.705 ;
        RECT 11.415 185.075 12.625 186.165 ;
        RECT 13.715 186.165 15.405 186.685 ;
        RECT 15.575 186.335 17.225 186.855 ;
        RECT 13.715 185.075 17.225 186.165 ;
        RECT 18.990 185.510 19.340 186.760 ;
        RECT 20.820 186.250 21.160 187.080 ;
        RECT 22.915 186.900 23.205 187.625 ;
        RECT 23.895 186.805 24.105 187.625 ;
        RECT 24.275 186.825 24.605 187.455 ;
        RECT 17.400 185.075 22.745 185.510 ;
        RECT 22.915 185.075 23.205 186.240 ;
        RECT 24.275 186.225 24.525 186.825 ;
        RECT 24.775 186.805 25.005 187.625 ;
        RECT 25.330 186.995 25.615 187.455 ;
        RECT 25.785 187.165 26.055 187.625 ;
        RECT 25.330 186.825 26.285 186.995 ;
        RECT 24.695 186.385 25.025 186.635 ;
        RECT 23.895 185.075 24.105 186.215 ;
        RECT 24.275 185.245 24.605 186.225 ;
        RECT 24.775 185.075 25.005 186.215 ;
        RECT 25.215 186.095 25.905 186.655 ;
        RECT 26.075 185.925 26.285 186.825 ;
        RECT 25.330 185.705 26.285 185.925 ;
        RECT 26.455 186.655 26.855 187.455 ;
        RECT 27.045 186.995 27.325 187.455 ;
        RECT 27.845 187.165 28.170 187.625 ;
        RECT 27.045 186.825 28.170 186.995 ;
        RECT 28.340 186.885 28.725 187.455 ;
        RECT 27.720 186.715 28.170 186.825 ;
        RECT 26.455 186.095 27.550 186.655 ;
        RECT 27.720 186.385 28.275 186.715 ;
        RECT 25.330 185.245 25.615 185.705 ;
        RECT 25.785 185.075 26.055 185.535 ;
        RECT 26.455 185.245 26.855 186.095 ;
        RECT 27.720 185.925 28.170 186.385 ;
        RECT 28.445 186.215 28.725 186.885 ;
        RECT 27.045 185.705 28.170 185.925 ;
        RECT 27.045 185.245 27.325 185.705 ;
        RECT 27.845 185.075 28.170 185.535 ;
        RECT 28.340 185.245 28.725 186.215 ;
        RECT 29.270 186.915 29.525 187.445 ;
        RECT 29.705 187.165 29.990 187.625 ;
        RECT 29.270 186.055 29.450 186.915 ;
        RECT 30.170 186.715 30.420 187.365 ;
        RECT 29.620 186.385 30.420 186.715 ;
        RECT 29.270 185.925 29.525 186.055 ;
        RECT 29.185 185.755 29.525 185.925 ;
        RECT 29.270 185.385 29.525 185.755 ;
        RECT 29.705 185.075 29.990 185.875 ;
        RECT 30.170 185.795 30.420 186.385 ;
        RECT 30.620 187.030 30.940 187.360 ;
        RECT 31.120 187.145 31.780 187.625 ;
        RECT 31.980 187.235 32.830 187.405 ;
        RECT 30.620 186.135 30.810 187.030 ;
        RECT 31.130 186.705 31.790 186.975 ;
        RECT 31.460 186.645 31.790 186.705 ;
        RECT 30.980 186.475 31.310 186.535 ;
        RECT 31.980 186.475 32.150 187.235 ;
        RECT 33.390 187.165 33.710 187.625 ;
        RECT 33.910 186.985 34.160 187.415 ;
        RECT 34.450 187.185 34.860 187.625 ;
        RECT 35.030 187.245 36.045 187.445 ;
        RECT 32.320 186.815 33.570 186.985 ;
        RECT 32.320 186.695 32.650 186.815 ;
        RECT 30.980 186.305 32.880 186.475 ;
        RECT 30.620 185.965 32.540 186.135 ;
        RECT 30.620 185.945 30.940 185.965 ;
        RECT 30.170 185.285 30.500 185.795 ;
        RECT 30.770 185.335 30.940 185.945 ;
        RECT 32.710 185.795 32.880 186.305 ;
        RECT 33.050 186.235 33.230 186.645 ;
        RECT 33.400 186.055 33.570 186.815 ;
        RECT 31.110 185.075 31.440 185.765 ;
        RECT 31.670 185.625 32.880 185.795 ;
        RECT 33.050 185.745 33.570 186.055 ;
        RECT 33.740 186.645 34.160 186.985 ;
        RECT 34.450 186.645 34.860 186.975 ;
        RECT 33.740 185.875 33.930 186.645 ;
        RECT 35.030 186.515 35.200 187.245 ;
        RECT 36.345 187.075 36.515 187.405 ;
        RECT 36.685 187.245 37.015 187.625 ;
        RECT 35.370 186.695 35.720 187.065 ;
        RECT 35.030 186.475 35.450 186.515 ;
        RECT 34.100 186.305 35.450 186.475 ;
        RECT 34.100 186.145 34.350 186.305 ;
        RECT 34.860 185.875 35.110 186.135 ;
        RECT 33.740 185.625 35.110 185.875 ;
        RECT 31.670 185.335 31.910 185.625 ;
        RECT 32.710 185.545 32.880 185.625 ;
        RECT 32.110 185.075 32.530 185.455 ;
        RECT 32.710 185.295 33.340 185.545 ;
        RECT 33.810 185.075 34.140 185.455 ;
        RECT 34.310 185.335 34.480 185.625 ;
        RECT 35.280 185.460 35.450 186.305 ;
        RECT 35.900 186.135 36.120 187.005 ;
        RECT 36.345 186.885 37.040 187.075 ;
        RECT 35.620 185.755 36.120 186.135 ;
        RECT 36.290 186.085 36.700 186.705 ;
        RECT 36.870 185.915 37.040 186.885 ;
        RECT 36.345 185.745 37.040 185.915 ;
        RECT 34.660 185.075 35.040 185.455 ;
        RECT 35.280 185.290 36.110 185.460 ;
        RECT 36.345 185.245 36.515 185.745 ;
        RECT 36.685 185.075 37.015 185.575 ;
        RECT 37.230 185.245 37.455 187.365 ;
        RECT 37.625 187.245 37.955 187.625 ;
        RECT 38.125 187.075 38.295 187.365 ;
        RECT 37.630 186.905 38.295 187.075 ;
        RECT 38.555 186.950 38.815 187.455 ;
        RECT 38.995 187.245 39.325 187.625 ;
        RECT 39.505 187.075 39.675 187.455 ;
        RECT 37.630 185.915 37.860 186.905 ;
        RECT 38.030 186.085 38.380 186.735 ;
        RECT 38.555 186.150 38.725 186.950 ;
        RECT 39.010 186.905 39.675 187.075 ;
        RECT 39.010 186.650 39.180 186.905 ;
        RECT 40.670 186.815 40.915 187.420 ;
        RECT 41.135 187.090 41.645 187.625 ;
        RECT 38.895 186.320 39.180 186.650 ;
        RECT 39.415 186.355 39.745 186.725 ;
        RECT 40.395 186.645 41.625 186.815 ;
        RECT 39.010 186.175 39.180 186.320 ;
        RECT 37.630 185.745 38.295 185.915 ;
        RECT 37.625 185.075 37.955 185.575 ;
        RECT 38.125 185.245 38.295 185.745 ;
        RECT 38.555 185.245 38.825 186.150 ;
        RECT 39.010 186.005 39.675 186.175 ;
        RECT 38.995 185.075 39.325 185.835 ;
        RECT 39.505 185.245 39.675 186.005 ;
        RECT 40.395 185.835 40.735 186.645 ;
        RECT 40.905 186.080 41.655 186.270 ;
        RECT 40.395 185.425 40.910 185.835 ;
        RECT 41.145 185.075 41.315 185.835 ;
        RECT 41.485 185.415 41.655 186.080 ;
        RECT 41.825 186.095 42.015 187.455 ;
        RECT 42.185 187.285 42.460 187.455 ;
        RECT 42.185 187.115 42.465 187.285 ;
        RECT 42.185 186.295 42.460 187.115 ;
        RECT 42.650 187.090 43.180 187.455 ;
        RECT 43.605 187.225 43.935 187.625 ;
        RECT 43.005 187.055 43.180 187.090 ;
        RECT 42.665 186.095 42.835 186.895 ;
        RECT 41.825 185.925 42.835 186.095 ;
        RECT 43.005 186.885 43.935 187.055 ;
        RECT 44.105 186.885 44.360 187.455 ;
        RECT 43.005 185.755 43.175 186.885 ;
        RECT 43.765 186.715 43.935 186.885 ;
        RECT 42.050 185.585 43.175 185.755 ;
        RECT 43.345 186.385 43.540 186.715 ;
        RECT 43.765 186.385 44.020 186.715 ;
        RECT 43.345 185.415 43.515 186.385 ;
        RECT 44.190 186.215 44.360 186.885 ;
        RECT 44.810 186.815 45.055 187.420 ;
        RECT 45.275 187.090 45.785 187.625 ;
        RECT 41.485 185.245 43.515 185.415 ;
        RECT 43.685 185.075 43.855 186.215 ;
        RECT 44.025 185.245 44.360 186.215 ;
        RECT 44.535 186.645 45.765 186.815 ;
        RECT 44.535 185.835 44.875 186.645 ;
        RECT 45.045 186.080 45.795 186.270 ;
        RECT 44.535 185.425 45.050 185.835 ;
        RECT 45.285 185.075 45.455 185.835 ;
        RECT 45.625 185.415 45.795 186.080 ;
        RECT 45.965 186.095 46.155 187.455 ;
        RECT 46.325 186.945 46.600 187.455 ;
        RECT 46.790 187.090 47.320 187.455 ;
        RECT 47.745 187.225 48.075 187.625 ;
        RECT 47.145 187.055 47.320 187.090 ;
        RECT 46.325 186.775 46.605 186.945 ;
        RECT 46.325 186.295 46.600 186.775 ;
        RECT 46.805 186.095 46.975 186.895 ;
        RECT 45.965 185.925 46.975 186.095 ;
        RECT 47.145 186.885 48.075 187.055 ;
        RECT 48.245 186.885 48.500 187.455 ;
        RECT 48.675 186.900 48.965 187.625 ;
        RECT 50.145 187.075 50.315 187.455 ;
        RECT 50.495 187.245 50.825 187.625 ;
        RECT 50.145 186.905 50.810 187.075 ;
        RECT 51.005 186.950 51.265 187.455 ;
        RECT 47.145 185.755 47.315 186.885 ;
        RECT 47.905 186.715 48.075 186.885 ;
        RECT 46.190 185.585 47.315 185.755 ;
        RECT 47.485 186.385 47.680 186.715 ;
        RECT 47.905 186.385 48.160 186.715 ;
        RECT 47.485 185.415 47.655 186.385 ;
        RECT 48.330 186.215 48.500 186.885 ;
        RECT 50.075 186.355 50.405 186.725 ;
        RECT 50.640 186.650 50.810 186.905 ;
        RECT 50.640 186.320 50.925 186.650 ;
        RECT 45.625 185.245 47.655 185.415 ;
        RECT 47.825 185.075 47.995 186.215 ;
        RECT 48.165 185.245 48.500 186.215 ;
        RECT 48.675 185.075 48.965 186.240 ;
        RECT 50.640 186.175 50.810 186.320 ;
        RECT 50.145 186.005 50.810 186.175 ;
        RECT 51.095 186.150 51.265 186.950 ;
        RECT 51.435 186.875 52.645 187.625 ;
        RECT 52.820 187.075 53.075 187.365 ;
        RECT 53.245 187.245 53.575 187.625 ;
        RECT 52.820 186.905 53.570 187.075 ;
        RECT 50.145 185.245 50.315 186.005 ;
        RECT 50.495 185.075 50.825 185.835 ;
        RECT 50.995 185.245 51.265 186.150 ;
        RECT 51.435 186.165 51.955 186.705 ;
        RECT 52.125 186.335 52.645 186.875 ;
        RECT 51.435 185.075 52.645 186.165 ;
        RECT 52.820 186.085 53.170 186.735 ;
        RECT 53.340 185.915 53.570 186.905 ;
        RECT 52.820 185.745 53.570 185.915 ;
        RECT 52.820 185.245 53.075 185.745 ;
        RECT 53.245 185.075 53.575 185.575 ;
        RECT 53.745 185.245 53.915 187.365 ;
        RECT 54.275 187.265 54.605 187.625 ;
        RECT 54.775 187.235 55.270 187.405 ;
        RECT 55.475 187.235 56.330 187.405 ;
        RECT 54.145 186.045 54.605 187.095 ;
        RECT 54.085 185.260 54.410 186.045 ;
        RECT 54.775 185.875 54.945 187.235 ;
        RECT 55.115 186.325 55.465 186.945 ;
        RECT 55.635 186.725 55.990 186.945 ;
        RECT 55.635 186.135 55.805 186.725 ;
        RECT 56.160 186.525 56.330 187.235 ;
        RECT 57.205 187.165 57.535 187.625 ;
        RECT 57.745 187.265 58.095 187.435 ;
        RECT 56.535 186.695 57.325 186.945 ;
        RECT 57.745 186.875 58.005 187.265 ;
        RECT 58.315 187.175 59.265 187.455 ;
        RECT 59.435 187.185 59.625 187.625 ;
        RECT 59.795 187.245 60.865 187.415 ;
        RECT 57.495 186.525 57.665 186.705 ;
        RECT 54.775 185.705 55.170 185.875 ;
        RECT 55.340 185.745 55.805 186.135 ;
        RECT 55.975 186.355 57.665 186.525 ;
        RECT 55.000 185.575 55.170 185.705 ;
        RECT 55.975 185.575 56.145 186.355 ;
        RECT 57.835 186.185 58.005 186.875 ;
        RECT 56.505 186.015 58.005 186.185 ;
        RECT 58.195 186.215 58.405 187.005 ;
        RECT 58.575 186.385 58.925 187.005 ;
        RECT 59.095 186.395 59.265 187.175 ;
        RECT 59.795 187.015 59.965 187.245 ;
        RECT 59.435 186.845 59.965 187.015 ;
        RECT 59.435 186.565 59.655 186.845 ;
        RECT 60.135 186.675 60.375 187.075 ;
        RECT 59.095 186.225 59.500 186.395 ;
        RECT 59.835 186.305 60.375 186.675 ;
        RECT 60.545 186.890 60.865 187.245 ;
        RECT 61.110 187.165 61.415 187.625 ;
        RECT 61.585 186.915 61.840 187.445 ;
        RECT 62.020 187.080 67.365 187.625 ;
        RECT 67.540 187.080 72.885 187.625 ;
        RECT 60.545 186.715 60.870 186.890 ;
        RECT 60.545 186.415 61.460 186.715 ;
        RECT 60.720 186.385 61.460 186.415 ;
        RECT 58.195 186.055 58.870 186.215 ;
        RECT 59.330 186.135 59.500 186.225 ;
        RECT 58.195 186.045 59.160 186.055 ;
        RECT 57.835 185.875 58.005 186.015 ;
        RECT 54.580 185.075 54.830 185.535 ;
        RECT 55.000 185.245 55.250 185.575 ;
        RECT 55.465 185.245 56.145 185.575 ;
        RECT 56.315 185.675 57.390 185.845 ;
        RECT 57.835 185.705 58.395 185.875 ;
        RECT 58.700 185.755 59.160 186.045 ;
        RECT 59.330 185.965 60.550 186.135 ;
        RECT 56.315 185.335 56.485 185.675 ;
        RECT 56.720 185.075 57.050 185.505 ;
        RECT 57.220 185.335 57.390 185.675 ;
        RECT 57.685 185.075 58.055 185.535 ;
        RECT 58.225 185.245 58.395 185.705 ;
        RECT 59.330 185.585 59.500 185.965 ;
        RECT 60.720 185.795 60.890 186.385 ;
        RECT 61.630 186.265 61.840 186.915 ;
        RECT 58.630 185.245 59.500 185.585 ;
        RECT 60.090 185.625 60.890 185.795 ;
        RECT 59.670 185.075 59.920 185.535 ;
        RECT 60.090 185.335 60.260 185.625 ;
        RECT 60.440 185.075 60.770 185.455 ;
        RECT 61.110 185.075 61.415 186.215 ;
        RECT 61.585 185.385 61.840 186.265 ;
        RECT 63.610 185.510 63.960 186.760 ;
        RECT 65.440 186.250 65.780 187.080 ;
        RECT 69.130 185.510 69.480 186.760 ;
        RECT 70.960 186.250 71.300 187.080 ;
        RECT 73.095 186.805 73.325 187.625 ;
        RECT 73.495 186.825 73.825 187.455 ;
        RECT 73.075 186.385 73.405 186.635 ;
        RECT 73.575 186.225 73.825 186.825 ;
        RECT 73.995 186.805 74.205 187.625 ;
        RECT 74.435 186.900 74.725 187.625 ;
        RECT 76.090 186.815 76.335 187.420 ;
        RECT 76.555 187.090 77.065 187.625 ;
        RECT 75.815 186.645 77.045 186.815 ;
        RECT 62.020 185.075 67.365 185.510 ;
        RECT 67.540 185.075 72.885 185.510 ;
        RECT 73.095 185.075 73.325 186.215 ;
        RECT 73.495 185.245 73.825 186.225 ;
        RECT 73.995 185.075 74.205 186.215 ;
        RECT 74.435 185.075 74.725 186.240 ;
        RECT 75.815 185.835 76.155 186.645 ;
        RECT 76.325 186.080 77.075 186.270 ;
        RECT 75.815 185.425 76.330 185.835 ;
        RECT 76.565 185.075 76.735 185.835 ;
        RECT 76.905 185.415 77.075 186.080 ;
        RECT 77.245 186.095 77.435 187.455 ;
        RECT 77.605 186.945 77.880 187.455 ;
        RECT 78.070 187.090 78.600 187.455 ;
        RECT 79.025 187.225 79.355 187.625 ;
        RECT 78.425 187.055 78.600 187.090 ;
        RECT 77.605 186.775 77.885 186.945 ;
        RECT 77.605 186.295 77.880 186.775 ;
        RECT 78.085 186.095 78.255 186.895 ;
        RECT 77.245 185.925 78.255 186.095 ;
        RECT 78.425 186.885 79.355 187.055 ;
        RECT 79.525 186.885 79.780 187.455 ;
        RECT 78.425 185.755 78.595 186.885 ;
        RECT 79.185 186.715 79.355 186.885 ;
        RECT 77.470 185.585 78.595 185.755 ;
        RECT 78.765 186.385 78.960 186.715 ;
        RECT 79.185 186.385 79.440 186.715 ;
        RECT 78.765 185.415 78.935 186.385 ;
        RECT 79.610 186.215 79.780 186.885 ;
        RECT 80.015 186.805 80.225 187.625 ;
        RECT 80.395 186.825 80.725 187.455 ;
        RECT 80.395 186.225 80.645 186.825 ;
        RECT 80.895 186.805 81.125 187.625 ;
        RECT 81.800 187.080 87.145 187.625 ;
        RECT 80.815 186.385 81.145 186.635 ;
        RECT 76.905 185.245 78.935 185.415 ;
        RECT 79.105 185.075 79.275 186.215 ;
        RECT 79.445 185.245 79.780 186.215 ;
        RECT 80.015 185.075 80.225 186.215 ;
        RECT 80.395 185.245 80.725 186.225 ;
        RECT 80.895 185.075 81.125 186.215 ;
        RECT 83.390 185.510 83.740 186.760 ;
        RECT 85.220 186.250 85.560 187.080 ;
        RECT 87.430 186.995 87.715 187.455 ;
        RECT 87.885 187.165 88.155 187.625 ;
        RECT 87.430 186.825 88.385 186.995 ;
        RECT 87.315 186.095 88.005 186.655 ;
        RECT 88.175 185.925 88.385 186.825 ;
        RECT 87.430 185.705 88.385 185.925 ;
        RECT 88.555 186.655 88.955 187.455 ;
        RECT 89.145 186.995 89.425 187.455 ;
        RECT 89.945 187.165 90.270 187.625 ;
        RECT 89.145 186.825 90.270 186.995 ;
        RECT 90.440 186.885 90.825 187.455 ;
        RECT 92.005 187.075 92.175 187.455 ;
        RECT 92.355 187.245 92.685 187.625 ;
        RECT 92.005 186.905 92.670 187.075 ;
        RECT 92.865 186.950 93.125 187.455 ;
        RECT 89.820 186.715 90.270 186.825 ;
        RECT 88.555 186.095 89.650 186.655 ;
        RECT 89.820 186.385 90.375 186.715 ;
        RECT 81.800 185.075 87.145 185.510 ;
        RECT 87.430 185.245 87.715 185.705 ;
        RECT 87.885 185.075 88.155 185.535 ;
        RECT 88.555 185.245 88.955 186.095 ;
        RECT 89.820 185.925 90.270 186.385 ;
        RECT 90.545 186.215 90.825 186.885 ;
        RECT 91.935 186.355 92.265 186.725 ;
        RECT 92.500 186.650 92.670 186.905 ;
        RECT 89.145 185.705 90.270 185.925 ;
        RECT 89.145 185.245 89.425 185.705 ;
        RECT 89.945 185.075 90.270 185.535 ;
        RECT 90.440 185.245 90.825 186.215 ;
        RECT 92.500 186.320 92.785 186.650 ;
        RECT 92.500 186.175 92.670 186.320 ;
        RECT 92.005 186.005 92.670 186.175 ;
        RECT 92.955 186.150 93.125 186.950 ;
        RECT 92.005 185.245 92.175 186.005 ;
        RECT 92.355 185.075 92.685 185.835 ;
        RECT 92.855 185.245 93.125 186.150 ;
        RECT 93.295 186.885 93.680 187.455 ;
        RECT 93.850 187.165 94.175 187.625 ;
        RECT 94.695 186.995 94.975 187.455 ;
        RECT 93.295 186.215 93.575 186.885 ;
        RECT 93.850 186.825 94.975 186.995 ;
        RECT 93.850 186.715 94.300 186.825 ;
        RECT 93.745 186.385 94.300 186.715 ;
        RECT 95.165 186.655 95.565 187.455 ;
        RECT 95.965 187.165 96.235 187.625 ;
        RECT 96.405 186.995 96.690 187.455 ;
        RECT 93.295 185.245 93.680 186.215 ;
        RECT 93.850 185.925 94.300 186.385 ;
        RECT 94.470 186.095 95.565 186.655 ;
        RECT 93.850 185.705 94.975 185.925 ;
        RECT 93.850 185.075 94.175 185.535 ;
        RECT 94.695 185.245 94.975 185.705 ;
        RECT 95.165 185.245 95.565 186.095 ;
        RECT 95.735 186.825 96.690 186.995 ;
        RECT 96.975 186.855 98.645 187.625 ;
        RECT 95.735 185.925 95.945 186.825 ;
        RECT 96.115 186.095 96.805 186.655 ;
        RECT 96.975 186.165 97.725 186.685 ;
        RECT 97.895 186.335 98.645 186.855 ;
        RECT 98.855 186.805 99.085 187.625 ;
        RECT 99.255 186.825 99.585 187.455 ;
        RECT 98.835 186.385 99.165 186.635 ;
        RECT 99.335 186.225 99.585 186.825 ;
        RECT 99.755 186.805 99.965 187.625 ;
        RECT 100.195 186.900 100.485 187.625 ;
        RECT 100.770 186.995 101.055 187.455 ;
        RECT 101.225 187.165 101.495 187.625 ;
        RECT 100.770 186.825 101.725 186.995 ;
        RECT 95.735 185.705 96.690 185.925 ;
        RECT 95.965 185.075 96.235 185.535 ;
        RECT 96.405 185.245 96.690 185.705 ;
        RECT 96.975 185.075 98.645 186.165 ;
        RECT 98.855 185.075 99.085 186.215 ;
        RECT 99.255 185.245 99.585 186.225 ;
        RECT 99.755 185.075 99.965 186.215 ;
        RECT 100.195 185.075 100.485 186.240 ;
        RECT 100.655 186.095 101.345 186.655 ;
        RECT 101.515 185.925 101.725 186.825 ;
        RECT 100.770 185.705 101.725 185.925 ;
        RECT 101.895 186.655 102.295 187.455 ;
        RECT 102.485 186.995 102.765 187.455 ;
        RECT 103.285 187.165 103.610 187.625 ;
        RECT 102.485 186.825 103.610 186.995 ;
        RECT 103.780 186.885 104.165 187.455 ;
        RECT 103.160 186.715 103.610 186.825 ;
        RECT 101.895 186.095 102.990 186.655 ;
        RECT 103.160 186.385 103.715 186.715 ;
        RECT 100.770 185.245 101.055 185.705 ;
        RECT 101.225 185.075 101.495 185.535 ;
        RECT 101.895 185.245 102.295 186.095 ;
        RECT 103.160 185.925 103.610 186.385 ;
        RECT 103.885 186.215 104.165 186.885 ;
        RECT 102.485 185.705 103.610 185.925 ;
        RECT 102.485 185.245 102.765 185.705 ;
        RECT 103.285 185.075 103.610 185.535 ;
        RECT 103.780 185.245 104.165 186.215 ;
        RECT 104.335 186.885 104.720 187.455 ;
        RECT 104.890 187.165 105.215 187.625 ;
        RECT 105.735 186.995 106.015 187.455 ;
        RECT 104.335 186.215 104.615 186.885 ;
        RECT 104.890 186.825 106.015 186.995 ;
        RECT 104.890 186.715 105.340 186.825 ;
        RECT 104.785 186.385 105.340 186.715 ;
        RECT 106.205 186.655 106.605 187.455 ;
        RECT 107.005 187.165 107.275 187.625 ;
        RECT 107.445 186.995 107.730 187.455 ;
        RECT 104.335 185.245 104.720 186.215 ;
        RECT 104.890 185.925 105.340 186.385 ;
        RECT 105.510 186.095 106.605 186.655 ;
        RECT 104.890 185.705 106.015 185.925 ;
        RECT 104.890 185.075 105.215 185.535 ;
        RECT 105.735 185.245 106.015 185.705 ;
        RECT 106.205 185.245 106.605 186.095 ;
        RECT 106.775 186.825 107.730 186.995 ;
        RECT 108.475 186.855 111.985 187.625 ;
        RECT 112.155 186.875 113.365 187.625 ;
        RECT 106.775 185.925 106.985 186.825 ;
        RECT 107.155 186.095 107.845 186.655 ;
        RECT 108.475 186.165 110.165 186.685 ;
        RECT 110.335 186.335 111.985 186.855 ;
        RECT 112.155 186.165 112.675 186.705 ;
        RECT 112.845 186.335 113.365 186.875 ;
        RECT 106.775 185.705 107.730 185.925 ;
        RECT 107.005 185.075 107.275 185.535 ;
        RECT 107.445 185.245 107.730 185.705 ;
        RECT 108.475 185.075 111.985 186.165 ;
        RECT 112.155 185.075 113.365 186.165 ;
        RECT 11.330 184.905 113.450 185.075 ;
        RECT 11.415 183.815 12.625 184.905 ;
        RECT 11.415 183.105 11.935 183.645 ;
        RECT 12.105 183.275 12.625 183.815 ;
        RECT 13.715 183.815 17.225 184.905 ;
        RECT 17.400 184.470 22.745 184.905 ;
        RECT 13.715 183.295 15.405 183.815 ;
        RECT 15.575 183.125 17.225 183.645 ;
        RECT 18.990 183.220 19.340 184.470 ;
        RECT 23.005 183.975 23.175 184.735 ;
        RECT 23.355 184.145 23.685 184.905 ;
        RECT 23.005 183.805 23.670 183.975 ;
        RECT 23.855 183.830 24.125 184.735 ;
        RECT 11.415 182.355 12.625 183.105 ;
        RECT 13.715 182.355 17.225 183.125 ;
        RECT 20.820 182.900 21.160 183.730 ;
        RECT 23.500 183.660 23.670 183.805 ;
        RECT 22.935 183.255 23.265 183.625 ;
        RECT 23.500 183.330 23.785 183.660 ;
        RECT 23.500 183.075 23.670 183.330 ;
        RECT 23.005 182.905 23.670 183.075 ;
        RECT 23.955 183.030 24.125 183.830 ;
        RECT 24.335 183.765 24.565 184.905 ;
        RECT 24.735 183.755 25.065 184.735 ;
        RECT 25.235 183.765 25.445 184.905 ;
        RECT 26.600 183.765 26.935 184.735 ;
        RECT 27.105 183.765 27.275 184.905 ;
        RECT 27.445 184.565 29.475 184.735 ;
        RECT 24.315 183.345 24.645 183.595 ;
        RECT 17.400 182.355 22.745 182.900 ;
        RECT 23.005 182.525 23.175 182.905 ;
        RECT 23.355 182.355 23.685 182.735 ;
        RECT 23.865 182.525 24.125 183.030 ;
        RECT 24.335 182.355 24.565 183.175 ;
        RECT 24.815 183.155 25.065 183.755 ;
        RECT 24.735 182.525 25.065 183.155 ;
        RECT 25.235 182.355 25.445 183.175 ;
        RECT 26.600 183.095 26.770 183.765 ;
        RECT 27.445 183.595 27.615 184.565 ;
        RECT 26.940 183.265 27.195 183.595 ;
        RECT 27.420 183.265 27.615 183.595 ;
        RECT 27.785 184.225 28.910 184.395 ;
        RECT 27.025 183.095 27.195 183.265 ;
        RECT 27.785 183.095 27.955 184.225 ;
        RECT 26.600 182.525 26.855 183.095 ;
        RECT 27.025 182.925 27.955 183.095 ;
        RECT 28.125 183.885 29.135 184.055 ;
        RECT 28.125 183.085 28.295 183.885 ;
        RECT 27.780 182.890 27.955 182.925 ;
        RECT 27.025 182.355 27.355 182.755 ;
        RECT 27.780 182.525 28.310 182.890 ;
        RECT 28.500 182.865 28.775 183.685 ;
        RECT 28.495 182.695 28.775 182.865 ;
        RECT 28.500 182.525 28.775 182.695 ;
        RECT 28.945 182.525 29.135 183.885 ;
        RECT 29.305 183.900 29.475 184.565 ;
        RECT 29.645 184.145 29.815 184.905 ;
        RECT 30.050 184.145 30.565 184.555 ;
        RECT 29.305 183.710 30.055 183.900 ;
        RECT 30.225 183.335 30.565 184.145 ;
        RECT 30.850 184.275 31.135 184.735 ;
        RECT 31.305 184.445 31.575 184.905 ;
        RECT 30.850 184.055 31.805 184.275 ;
        RECT 29.335 183.165 30.565 183.335 ;
        RECT 30.735 183.325 31.425 183.885 ;
        RECT 29.315 182.355 29.825 182.890 ;
        RECT 30.045 182.560 30.290 183.165 ;
        RECT 31.595 183.155 31.805 184.055 ;
        RECT 30.850 182.985 31.805 183.155 ;
        RECT 31.975 183.885 32.375 184.735 ;
        RECT 32.565 184.275 32.845 184.735 ;
        RECT 33.365 184.445 33.690 184.905 ;
        RECT 32.565 184.055 33.690 184.275 ;
        RECT 31.975 183.325 33.070 183.885 ;
        RECT 33.240 183.595 33.690 184.055 ;
        RECT 33.860 183.765 34.245 184.735 ;
        RECT 34.475 183.765 34.685 184.905 ;
        RECT 30.850 182.525 31.135 182.985 ;
        RECT 31.305 182.355 31.575 182.815 ;
        RECT 31.975 182.525 32.375 183.325 ;
        RECT 33.240 183.265 33.795 183.595 ;
        RECT 33.240 183.155 33.690 183.265 ;
        RECT 32.565 182.985 33.690 183.155 ;
        RECT 33.965 183.095 34.245 183.765 ;
        RECT 34.855 183.755 35.185 184.735 ;
        RECT 35.355 183.765 35.585 184.905 ;
        RECT 32.565 182.525 32.845 182.985 ;
        RECT 33.365 182.355 33.690 182.815 ;
        RECT 33.860 182.525 34.245 183.095 ;
        RECT 34.475 182.355 34.685 183.175 ;
        RECT 34.855 183.155 35.105 183.755 ;
        RECT 35.795 183.740 36.085 184.905 ;
        RECT 36.315 183.765 36.525 184.905 ;
        RECT 36.695 183.755 37.025 184.735 ;
        RECT 37.195 183.765 37.425 184.905 ;
        RECT 37.635 183.815 39.305 184.905 ;
        RECT 39.475 183.830 39.745 184.735 ;
        RECT 39.915 184.145 40.245 184.905 ;
        RECT 40.425 183.975 40.595 184.735 ;
        RECT 35.275 183.345 35.605 183.595 ;
        RECT 34.855 182.525 35.185 183.155 ;
        RECT 35.355 182.355 35.585 183.175 ;
        RECT 35.795 182.355 36.085 183.080 ;
        RECT 36.315 182.355 36.525 183.175 ;
        RECT 36.695 183.155 36.945 183.755 ;
        RECT 37.115 183.345 37.445 183.595 ;
        RECT 37.635 183.295 38.385 183.815 ;
        RECT 36.695 182.525 37.025 183.155 ;
        RECT 37.195 182.355 37.425 183.175 ;
        RECT 38.555 183.125 39.305 183.645 ;
        RECT 37.635 182.355 39.305 183.125 ;
        RECT 39.475 183.030 39.645 183.830 ;
        RECT 39.930 183.805 40.595 183.975 ;
        RECT 41.315 183.815 42.985 184.905 ;
        RECT 39.930 183.660 40.100 183.805 ;
        RECT 39.815 183.330 40.100 183.660 ;
        RECT 39.930 183.075 40.100 183.330 ;
        RECT 40.335 183.255 40.665 183.625 ;
        RECT 41.315 183.295 42.065 183.815 ;
        RECT 43.215 183.765 43.425 184.905 ;
        RECT 43.595 183.755 43.925 184.735 ;
        RECT 44.095 183.765 44.325 184.905 ;
        RECT 44.575 183.765 44.805 184.905 ;
        RECT 44.975 183.755 45.305 184.735 ;
        RECT 45.475 183.765 45.685 184.905 ;
        RECT 46.030 184.275 46.315 184.735 ;
        RECT 46.485 184.445 46.755 184.905 ;
        RECT 46.030 184.055 46.985 184.275 ;
        RECT 42.235 183.125 42.985 183.645 ;
        RECT 39.475 182.525 39.735 183.030 ;
        RECT 39.930 182.905 40.595 183.075 ;
        RECT 39.915 182.355 40.245 182.735 ;
        RECT 40.425 182.525 40.595 182.905 ;
        RECT 41.315 182.355 42.985 183.125 ;
        RECT 43.215 182.355 43.425 183.175 ;
        RECT 43.595 183.155 43.845 183.755 ;
        RECT 44.015 183.345 44.345 183.595 ;
        RECT 44.555 183.345 44.885 183.595 ;
        RECT 43.595 182.525 43.925 183.155 ;
        RECT 44.095 182.355 44.325 183.175 ;
        RECT 44.575 182.355 44.805 183.175 ;
        RECT 45.055 183.155 45.305 183.755 ;
        RECT 45.915 183.325 46.605 183.885 ;
        RECT 44.975 182.525 45.305 183.155 ;
        RECT 45.475 182.355 45.685 183.175 ;
        RECT 46.775 183.155 46.985 184.055 ;
        RECT 46.030 182.985 46.985 183.155 ;
        RECT 47.155 183.885 47.555 184.735 ;
        RECT 47.745 184.275 48.025 184.735 ;
        RECT 48.545 184.445 48.870 184.905 ;
        RECT 47.745 184.055 48.870 184.275 ;
        RECT 47.155 183.325 48.250 183.885 ;
        RECT 48.420 183.595 48.870 184.055 ;
        RECT 49.040 183.765 49.425 184.735 ;
        RECT 50.520 184.470 55.865 184.905 ;
        RECT 56.040 184.470 61.385 184.905 ;
        RECT 46.030 182.525 46.315 182.985 ;
        RECT 46.485 182.355 46.755 182.815 ;
        RECT 47.155 182.525 47.555 183.325 ;
        RECT 48.420 183.265 48.975 183.595 ;
        RECT 48.420 183.155 48.870 183.265 ;
        RECT 47.745 182.985 48.870 183.155 ;
        RECT 49.145 183.095 49.425 183.765 ;
        RECT 52.110 183.220 52.460 184.470 ;
        RECT 47.745 182.525 48.025 182.985 ;
        RECT 48.545 182.355 48.870 182.815 ;
        RECT 49.040 182.525 49.425 183.095 ;
        RECT 53.940 182.900 54.280 183.730 ;
        RECT 57.630 183.220 57.980 184.470 ;
        RECT 61.555 183.740 61.845 184.905 ;
        RECT 59.460 182.900 59.800 183.730 ;
        RECT 62.935 183.095 63.195 184.720 ;
        RECT 64.945 184.455 65.275 184.905 ;
        RECT 66.620 184.470 71.965 184.905 ;
        RECT 63.375 184.065 65.985 184.275 ;
        RECT 63.375 183.265 63.595 184.065 ;
        RECT 63.835 183.265 64.135 183.885 ;
        RECT 64.305 183.265 64.635 183.885 ;
        RECT 64.805 183.265 65.125 183.885 ;
        RECT 65.295 183.265 65.645 183.885 ;
        RECT 65.815 183.095 65.985 184.065 ;
        RECT 68.210 183.220 68.560 184.470 ;
        RECT 72.510 183.925 72.765 184.595 ;
        RECT 72.945 184.105 73.230 184.905 ;
        RECT 73.410 184.185 73.740 184.695 ;
        RECT 50.520 182.355 55.865 182.900 ;
        RECT 56.040 182.355 61.385 182.900 ;
        RECT 61.555 182.355 61.845 183.080 ;
        RECT 62.935 182.925 64.775 183.095 ;
        RECT 63.205 182.355 63.535 182.750 ;
        RECT 63.705 182.570 63.905 182.925 ;
        RECT 64.075 182.355 64.405 182.755 ;
        RECT 64.575 182.580 64.775 182.925 ;
        RECT 64.945 182.355 65.275 183.095 ;
        RECT 65.510 182.925 65.985 183.095 ;
        RECT 65.510 182.675 65.680 182.925 ;
        RECT 70.040 182.900 70.380 183.730 ;
        RECT 72.510 183.065 72.690 183.925 ;
        RECT 73.410 183.595 73.660 184.185 ;
        RECT 74.010 184.035 74.180 184.645 ;
        RECT 74.350 184.215 74.680 184.905 ;
        RECT 74.910 184.355 75.150 184.645 ;
        RECT 75.350 184.525 75.770 184.905 ;
        RECT 75.950 184.435 76.580 184.685 ;
        RECT 77.050 184.525 77.380 184.905 ;
        RECT 75.950 184.355 76.120 184.435 ;
        RECT 77.550 184.355 77.720 184.645 ;
        RECT 77.900 184.525 78.280 184.905 ;
        RECT 78.520 184.520 79.350 184.690 ;
        RECT 74.910 184.185 76.120 184.355 ;
        RECT 72.860 183.265 73.660 183.595 ;
        RECT 66.620 182.355 71.965 182.900 ;
        RECT 72.510 182.865 72.765 183.065 ;
        RECT 72.425 182.695 72.765 182.865 ;
        RECT 72.510 182.535 72.765 182.695 ;
        RECT 72.945 182.355 73.230 182.815 ;
        RECT 73.410 182.615 73.660 183.265 ;
        RECT 73.860 184.015 74.180 184.035 ;
        RECT 73.860 183.845 75.780 184.015 ;
        RECT 73.860 182.950 74.050 183.845 ;
        RECT 75.950 183.675 76.120 184.185 ;
        RECT 76.290 183.925 76.810 184.235 ;
        RECT 74.220 183.505 76.120 183.675 ;
        RECT 74.220 183.445 74.550 183.505 ;
        RECT 74.700 183.275 75.030 183.335 ;
        RECT 74.370 183.005 75.030 183.275 ;
        RECT 73.860 182.620 74.180 182.950 ;
        RECT 74.360 182.355 75.020 182.835 ;
        RECT 75.220 182.745 75.390 183.505 ;
        RECT 76.290 183.335 76.470 183.745 ;
        RECT 75.560 183.165 75.890 183.285 ;
        RECT 76.640 183.165 76.810 183.925 ;
        RECT 75.560 182.995 76.810 183.165 ;
        RECT 76.980 184.105 78.350 184.355 ;
        RECT 76.980 183.335 77.170 184.105 ;
        RECT 78.100 183.845 78.350 184.105 ;
        RECT 77.340 183.675 77.590 183.835 ;
        RECT 78.520 183.675 78.690 184.520 ;
        RECT 79.585 184.235 79.755 184.735 ;
        RECT 79.925 184.405 80.255 184.905 ;
        RECT 78.860 183.845 79.360 184.225 ;
        RECT 79.585 184.065 80.280 184.235 ;
        RECT 77.340 183.505 78.690 183.675 ;
        RECT 78.270 183.465 78.690 183.505 ;
        RECT 76.980 182.995 77.400 183.335 ;
        RECT 77.690 183.005 78.100 183.335 ;
        RECT 75.220 182.575 76.070 182.745 ;
        RECT 76.630 182.355 76.950 182.815 ;
        RECT 77.150 182.565 77.400 182.995 ;
        RECT 77.690 182.355 78.100 182.795 ;
        RECT 78.270 182.735 78.440 183.465 ;
        RECT 78.610 182.915 78.960 183.285 ;
        RECT 79.140 182.975 79.360 183.845 ;
        RECT 79.530 183.275 79.940 183.895 ;
        RECT 80.110 183.095 80.280 184.065 ;
        RECT 79.585 182.905 80.280 183.095 ;
        RECT 78.270 182.535 79.285 182.735 ;
        RECT 79.585 182.575 79.755 182.905 ;
        RECT 79.925 182.355 80.255 182.735 ;
        RECT 80.470 182.615 80.695 184.735 ;
        RECT 80.865 184.405 81.195 184.905 ;
        RECT 81.365 184.235 81.535 184.735 ;
        RECT 80.870 184.065 81.535 184.235 ;
        RECT 80.870 183.075 81.100 184.065 ;
        RECT 81.270 183.245 81.620 183.895 ;
        RECT 81.795 183.830 82.065 184.735 ;
        RECT 82.235 184.145 82.565 184.905 ;
        RECT 82.745 183.975 82.915 184.735 ;
        RECT 80.870 182.905 81.535 183.075 ;
        RECT 80.865 182.355 81.195 182.735 ;
        RECT 81.365 182.615 81.535 182.905 ;
        RECT 81.795 183.030 81.965 183.830 ;
        RECT 82.250 183.805 82.915 183.975 ;
        RECT 83.175 183.815 84.385 184.905 ;
        RECT 82.250 183.660 82.420 183.805 ;
        RECT 82.135 183.330 82.420 183.660 ;
        RECT 82.250 183.075 82.420 183.330 ;
        RECT 82.655 183.255 82.985 183.625 ;
        RECT 83.175 183.275 83.695 183.815 ;
        RECT 84.615 183.765 84.825 184.905 ;
        RECT 84.995 183.755 85.325 184.735 ;
        RECT 85.495 183.765 85.725 184.905 ;
        RECT 85.975 183.765 86.205 184.905 ;
        RECT 86.375 183.755 86.705 184.735 ;
        RECT 86.875 183.765 87.085 184.905 ;
        RECT 83.865 183.105 84.385 183.645 ;
        RECT 81.795 182.525 82.055 183.030 ;
        RECT 82.250 182.905 82.915 183.075 ;
        RECT 82.235 182.355 82.565 182.735 ;
        RECT 82.745 182.525 82.915 182.905 ;
        RECT 83.175 182.355 84.385 183.105 ;
        RECT 84.615 182.355 84.825 183.175 ;
        RECT 84.995 183.155 85.245 183.755 ;
        RECT 85.415 183.345 85.745 183.595 ;
        RECT 85.955 183.345 86.285 183.595 ;
        RECT 84.995 182.525 85.325 183.155 ;
        RECT 85.495 182.355 85.725 183.175 ;
        RECT 85.975 182.355 86.205 183.175 ;
        RECT 86.455 183.155 86.705 183.755 ;
        RECT 87.315 183.740 87.605 184.905 ;
        RECT 87.780 183.715 88.035 184.595 ;
        RECT 88.205 183.765 88.510 184.905 ;
        RECT 88.850 184.525 89.180 184.905 ;
        RECT 89.360 184.355 89.530 184.645 ;
        RECT 89.700 184.445 89.950 184.905 ;
        RECT 88.730 184.185 89.530 184.355 ;
        RECT 90.120 184.395 90.990 184.735 ;
        RECT 86.375 182.525 86.705 183.155 ;
        RECT 86.875 182.355 87.085 183.175 ;
        RECT 87.315 182.355 87.605 183.080 ;
        RECT 87.780 183.065 87.990 183.715 ;
        RECT 88.730 183.595 88.900 184.185 ;
        RECT 90.120 184.015 90.290 184.395 ;
        RECT 91.225 184.275 91.395 184.735 ;
        RECT 91.565 184.445 91.935 184.905 ;
        RECT 92.230 184.305 92.400 184.645 ;
        RECT 92.570 184.475 92.900 184.905 ;
        RECT 93.135 184.305 93.305 184.645 ;
        RECT 89.070 183.845 90.290 184.015 ;
        RECT 90.460 183.935 90.920 184.225 ;
        RECT 91.225 184.105 91.785 184.275 ;
        RECT 92.230 184.135 93.305 184.305 ;
        RECT 93.475 184.405 94.155 184.735 ;
        RECT 94.370 184.405 94.620 184.735 ;
        RECT 94.790 184.445 95.040 184.905 ;
        RECT 91.615 183.965 91.785 184.105 ;
        RECT 90.460 183.925 91.425 183.935 ;
        RECT 90.120 183.755 90.290 183.845 ;
        RECT 90.750 183.765 91.425 183.925 ;
        RECT 88.160 183.565 88.900 183.595 ;
        RECT 88.160 183.265 89.075 183.565 ;
        RECT 88.750 183.090 89.075 183.265 ;
        RECT 87.780 182.535 88.035 183.065 ;
        RECT 88.205 182.355 88.510 182.815 ;
        RECT 88.755 182.735 89.075 183.090 ;
        RECT 89.245 183.305 89.785 183.675 ;
        RECT 90.120 183.585 90.525 183.755 ;
        RECT 89.245 182.905 89.485 183.305 ;
        RECT 89.965 183.135 90.185 183.415 ;
        RECT 89.655 182.965 90.185 183.135 ;
        RECT 89.655 182.735 89.825 182.965 ;
        RECT 90.355 182.805 90.525 183.585 ;
        RECT 90.695 182.975 91.045 183.595 ;
        RECT 91.215 182.975 91.425 183.765 ;
        RECT 91.615 183.795 93.115 183.965 ;
        RECT 91.615 183.105 91.785 183.795 ;
        RECT 93.475 183.625 93.645 184.405 ;
        RECT 94.450 184.275 94.620 184.405 ;
        RECT 91.955 183.455 93.645 183.625 ;
        RECT 93.815 183.845 94.280 184.235 ;
        RECT 94.450 184.105 94.845 184.275 ;
        RECT 91.955 183.275 92.125 183.455 ;
        RECT 88.755 182.565 89.825 182.735 ;
        RECT 89.995 182.355 90.185 182.795 ;
        RECT 90.355 182.525 91.305 182.805 ;
        RECT 91.615 182.715 91.875 183.105 ;
        RECT 92.295 183.035 93.085 183.285 ;
        RECT 91.525 182.545 91.875 182.715 ;
        RECT 92.085 182.355 92.415 182.815 ;
        RECT 93.290 182.745 93.460 183.455 ;
        RECT 93.815 183.255 93.985 183.845 ;
        RECT 93.630 183.035 93.985 183.255 ;
        RECT 94.155 183.035 94.505 183.655 ;
        RECT 94.675 182.745 94.845 184.105 ;
        RECT 95.210 183.935 95.535 184.720 ;
        RECT 95.015 182.885 95.475 183.935 ;
        RECT 93.290 182.575 94.145 182.745 ;
        RECT 94.350 182.575 94.845 182.745 ;
        RECT 95.015 182.355 95.345 182.715 ;
        RECT 95.705 182.615 95.875 184.735 ;
        RECT 96.045 184.405 96.375 184.905 ;
        RECT 96.545 184.235 96.800 184.735 ;
        RECT 96.050 184.065 96.800 184.235 ;
        RECT 97.090 184.275 97.375 184.735 ;
        RECT 97.545 184.445 97.815 184.905 ;
        RECT 96.050 183.075 96.280 184.065 ;
        RECT 97.090 184.055 98.045 184.275 ;
        RECT 96.450 183.245 96.800 183.895 ;
        RECT 96.975 183.325 97.665 183.885 ;
        RECT 97.835 183.155 98.045 184.055 ;
        RECT 96.050 182.905 96.800 183.075 ;
        RECT 96.045 182.355 96.375 182.735 ;
        RECT 96.545 182.615 96.800 182.905 ;
        RECT 97.090 182.985 98.045 183.155 ;
        RECT 98.215 183.885 98.615 184.735 ;
        RECT 98.805 184.275 99.085 184.735 ;
        RECT 99.605 184.445 99.930 184.905 ;
        RECT 98.805 184.055 99.930 184.275 ;
        RECT 98.215 183.325 99.310 183.885 ;
        RECT 99.480 183.595 99.930 184.055 ;
        RECT 100.100 183.765 100.485 184.735 ;
        RECT 100.695 183.765 100.925 184.905 ;
        RECT 97.090 182.525 97.375 182.985 ;
        RECT 97.545 182.355 97.815 182.815 ;
        RECT 98.215 182.525 98.615 183.325 ;
        RECT 99.480 183.265 100.035 183.595 ;
        RECT 99.480 183.155 99.930 183.265 ;
        RECT 98.805 182.985 99.930 183.155 ;
        RECT 100.205 183.095 100.485 183.765 ;
        RECT 101.095 183.755 101.425 184.735 ;
        RECT 101.595 183.765 101.805 184.905 ;
        RECT 100.675 183.345 101.005 183.595 ;
        RECT 98.805 182.525 99.085 182.985 ;
        RECT 99.605 182.355 99.930 182.815 ;
        RECT 100.100 182.525 100.485 183.095 ;
        RECT 100.695 182.355 100.925 183.175 ;
        RECT 101.175 183.155 101.425 183.755 ;
        RECT 102.040 183.715 102.295 184.595 ;
        RECT 102.465 183.765 102.770 184.905 ;
        RECT 103.110 184.525 103.440 184.905 ;
        RECT 103.620 184.355 103.790 184.645 ;
        RECT 103.960 184.445 104.210 184.905 ;
        RECT 102.990 184.185 103.790 184.355 ;
        RECT 104.380 184.395 105.250 184.735 ;
        RECT 101.095 182.525 101.425 183.155 ;
        RECT 101.595 182.355 101.805 183.175 ;
        RECT 102.040 183.065 102.250 183.715 ;
        RECT 102.990 183.595 103.160 184.185 ;
        RECT 104.380 184.015 104.550 184.395 ;
        RECT 105.485 184.275 105.655 184.735 ;
        RECT 105.825 184.445 106.195 184.905 ;
        RECT 106.490 184.305 106.660 184.645 ;
        RECT 106.830 184.475 107.160 184.905 ;
        RECT 107.395 184.305 107.565 184.645 ;
        RECT 103.330 183.845 104.550 184.015 ;
        RECT 104.720 183.935 105.180 184.225 ;
        RECT 105.485 184.105 106.045 184.275 ;
        RECT 106.490 184.135 107.565 184.305 ;
        RECT 107.735 184.405 108.415 184.735 ;
        RECT 108.630 184.405 108.880 184.735 ;
        RECT 109.050 184.445 109.300 184.905 ;
        RECT 105.875 183.965 106.045 184.105 ;
        RECT 104.720 183.925 105.685 183.935 ;
        RECT 104.380 183.755 104.550 183.845 ;
        RECT 105.010 183.765 105.685 183.925 ;
        RECT 102.420 183.565 103.160 183.595 ;
        RECT 102.420 183.265 103.335 183.565 ;
        RECT 103.010 183.090 103.335 183.265 ;
        RECT 102.040 182.535 102.295 183.065 ;
        RECT 102.465 182.355 102.770 182.815 ;
        RECT 103.015 182.735 103.335 183.090 ;
        RECT 103.505 183.305 104.045 183.675 ;
        RECT 104.380 183.585 104.785 183.755 ;
        RECT 103.505 182.905 103.745 183.305 ;
        RECT 104.225 183.135 104.445 183.415 ;
        RECT 103.915 182.965 104.445 183.135 ;
        RECT 103.915 182.735 104.085 182.965 ;
        RECT 104.615 182.805 104.785 183.585 ;
        RECT 104.955 182.975 105.305 183.595 ;
        RECT 105.475 182.975 105.685 183.765 ;
        RECT 105.875 183.795 107.375 183.965 ;
        RECT 105.875 183.105 106.045 183.795 ;
        RECT 107.735 183.625 107.905 184.405 ;
        RECT 108.710 184.275 108.880 184.405 ;
        RECT 106.215 183.455 107.905 183.625 ;
        RECT 108.075 183.845 108.540 184.235 ;
        RECT 108.710 184.105 109.105 184.275 ;
        RECT 106.215 183.275 106.385 183.455 ;
        RECT 103.015 182.565 104.085 182.735 ;
        RECT 104.255 182.355 104.445 182.795 ;
        RECT 104.615 182.525 105.565 182.805 ;
        RECT 105.875 182.715 106.135 183.105 ;
        RECT 106.555 183.035 107.345 183.285 ;
        RECT 105.785 182.545 106.135 182.715 ;
        RECT 106.345 182.355 106.675 182.815 ;
        RECT 107.550 182.745 107.720 183.455 ;
        RECT 108.075 183.255 108.245 183.845 ;
        RECT 107.890 183.035 108.245 183.255 ;
        RECT 108.415 183.035 108.765 183.655 ;
        RECT 108.935 182.745 109.105 184.105 ;
        RECT 109.470 183.935 109.795 184.720 ;
        RECT 109.275 182.885 109.735 183.935 ;
        RECT 107.550 182.575 108.405 182.745 ;
        RECT 108.610 182.575 109.105 182.745 ;
        RECT 109.275 182.355 109.605 182.715 ;
        RECT 109.965 182.615 110.135 184.735 ;
        RECT 110.305 184.405 110.635 184.905 ;
        RECT 110.805 184.235 111.060 184.735 ;
        RECT 110.310 184.065 111.060 184.235 ;
        RECT 110.310 183.075 110.540 184.065 ;
        RECT 110.710 183.245 111.060 183.895 ;
        RECT 112.155 183.815 113.365 184.905 ;
        RECT 112.155 183.275 112.675 183.815 ;
        RECT 112.845 183.105 113.365 183.645 ;
        RECT 110.310 182.905 111.060 183.075 ;
        RECT 110.305 182.355 110.635 182.735 ;
        RECT 110.805 182.615 111.060 182.905 ;
        RECT 112.155 182.355 113.365 183.105 ;
        RECT 11.330 182.185 113.450 182.355 ;
        RECT 11.415 181.435 12.625 182.185 ;
        RECT 13.720 181.640 19.065 182.185 ;
        RECT 11.415 180.895 11.935 181.435 ;
        RECT 12.105 180.725 12.625 181.265 ;
        RECT 11.415 179.635 12.625 180.725 ;
        RECT 15.310 180.070 15.660 181.320 ;
        RECT 17.140 180.810 17.480 181.640 ;
        RECT 19.350 181.555 19.635 182.015 ;
        RECT 19.805 181.725 20.075 182.185 ;
        RECT 19.350 181.385 20.305 181.555 ;
        RECT 19.235 180.655 19.925 181.215 ;
        RECT 20.095 180.485 20.305 181.385 ;
        RECT 19.350 180.265 20.305 180.485 ;
        RECT 20.475 181.215 20.875 182.015 ;
        RECT 21.065 181.555 21.345 182.015 ;
        RECT 21.865 181.725 22.190 182.185 ;
        RECT 21.065 181.385 22.190 181.555 ;
        RECT 22.360 181.445 22.745 182.015 ;
        RECT 22.915 181.460 23.205 182.185 ;
        RECT 24.410 181.555 24.695 182.015 ;
        RECT 24.865 181.725 25.135 182.185 ;
        RECT 21.740 181.275 22.190 181.385 ;
        RECT 20.475 180.655 21.570 181.215 ;
        RECT 21.740 180.945 22.295 181.275 ;
        RECT 13.720 179.635 19.065 180.070 ;
        RECT 19.350 179.805 19.635 180.265 ;
        RECT 19.805 179.635 20.075 180.095 ;
        RECT 20.475 179.805 20.875 180.655 ;
        RECT 21.740 180.485 22.190 180.945 ;
        RECT 22.465 180.775 22.745 181.445 ;
        RECT 24.410 181.385 25.365 181.555 ;
        RECT 21.065 180.265 22.190 180.485 ;
        RECT 21.065 179.805 21.345 180.265 ;
        RECT 21.865 179.635 22.190 180.095 ;
        RECT 22.360 179.805 22.745 180.775 ;
        RECT 22.915 179.635 23.205 180.800 ;
        RECT 24.295 180.655 24.985 181.215 ;
        RECT 25.155 180.485 25.365 181.385 ;
        RECT 24.410 180.265 25.365 180.485 ;
        RECT 25.535 181.215 25.935 182.015 ;
        RECT 26.125 181.555 26.405 182.015 ;
        RECT 26.925 181.725 27.250 182.185 ;
        RECT 26.125 181.385 27.250 181.555 ;
        RECT 27.420 181.445 27.805 182.015 ;
        RECT 26.800 181.275 27.250 181.385 ;
        RECT 25.535 180.655 26.630 181.215 ;
        RECT 26.800 180.945 27.355 181.275 ;
        RECT 24.410 179.805 24.695 180.265 ;
        RECT 24.865 179.635 25.135 180.095 ;
        RECT 25.535 179.805 25.935 180.655 ;
        RECT 26.800 180.485 27.250 180.945 ;
        RECT 27.525 180.775 27.805 181.445 ;
        RECT 28.180 181.405 28.680 182.015 ;
        RECT 27.975 180.945 28.325 181.195 ;
        RECT 28.510 180.775 28.680 181.405 ;
        RECT 29.310 181.535 29.640 182.015 ;
        RECT 29.810 181.725 30.035 182.185 ;
        RECT 30.205 181.535 30.535 182.015 ;
        RECT 29.310 181.365 30.535 181.535 ;
        RECT 30.725 181.385 30.975 182.185 ;
        RECT 31.145 181.385 31.485 182.015 ;
        RECT 31.770 181.555 32.055 182.015 ;
        RECT 32.225 181.725 32.495 182.185 ;
        RECT 31.770 181.385 32.725 181.555 ;
        RECT 28.850 180.995 29.180 181.195 ;
        RECT 29.350 180.995 29.680 181.195 ;
        RECT 29.850 181.165 30.270 181.195 ;
        RECT 29.850 180.995 30.275 181.165 ;
        RECT 30.445 181.025 31.140 181.195 ;
        RECT 30.445 180.775 30.615 181.025 ;
        RECT 31.310 180.775 31.485 181.385 ;
        RECT 26.125 180.265 27.250 180.485 ;
        RECT 26.125 179.805 26.405 180.265 ;
        RECT 26.925 179.635 27.250 180.095 ;
        RECT 27.420 179.805 27.805 180.775 ;
        RECT 28.180 180.605 30.615 180.775 ;
        RECT 28.180 179.805 28.510 180.605 ;
        RECT 28.680 179.635 29.010 180.435 ;
        RECT 29.310 179.805 29.640 180.605 ;
        RECT 30.285 179.635 30.535 180.435 ;
        RECT 30.805 179.635 30.975 180.775 ;
        RECT 31.145 179.805 31.485 180.775 ;
        RECT 31.655 180.655 32.345 181.215 ;
        RECT 32.515 180.485 32.725 181.385 ;
        RECT 31.770 180.265 32.725 180.485 ;
        RECT 32.895 181.215 33.295 182.015 ;
        RECT 33.485 181.555 33.765 182.015 ;
        RECT 34.285 181.725 34.610 182.185 ;
        RECT 33.485 181.385 34.610 181.555 ;
        RECT 34.780 181.445 35.165 182.015 ;
        RECT 34.160 181.275 34.610 181.385 ;
        RECT 32.895 180.655 33.990 181.215 ;
        RECT 34.160 180.945 34.715 181.275 ;
        RECT 31.770 179.805 32.055 180.265 ;
        RECT 32.225 179.635 32.495 180.095 ;
        RECT 32.895 179.805 33.295 180.655 ;
        RECT 34.160 180.485 34.610 180.945 ;
        RECT 34.885 180.775 35.165 181.445 ;
        RECT 35.610 181.375 35.855 181.980 ;
        RECT 36.075 181.650 36.585 182.185 ;
        RECT 33.485 180.265 34.610 180.485 ;
        RECT 33.485 179.805 33.765 180.265 ;
        RECT 34.285 179.635 34.610 180.095 ;
        RECT 34.780 179.805 35.165 180.775 ;
        RECT 35.335 181.205 36.565 181.375 ;
        RECT 35.335 180.395 35.675 181.205 ;
        RECT 35.845 180.640 36.595 180.830 ;
        RECT 35.335 179.985 35.850 180.395 ;
        RECT 36.085 179.635 36.255 180.395 ;
        RECT 36.425 179.975 36.595 180.640 ;
        RECT 36.765 180.655 36.955 182.015 ;
        RECT 37.125 181.505 37.400 182.015 ;
        RECT 37.590 181.650 38.120 182.015 ;
        RECT 38.545 181.785 38.875 182.185 ;
        RECT 37.945 181.615 38.120 181.650 ;
        RECT 37.125 181.335 37.405 181.505 ;
        RECT 37.125 180.855 37.400 181.335 ;
        RECT 37.605 180.655 37.775 181.455 ;
        RECT 36.765 180.485 37.775 180.655 ;
        RECT 37.945 181.445 38.875 181.615 ;
        RECT 39.045 181.445 39.300 182.015 ;
        RECT 37.945 180.315 38.115 181.445 ;
        RECT 38.705 181.275 38.875 181.445 ;
        RECT 36.990 180.145 38.115 180.315 ;
        RECT 38.285 180.945 38.480 181.275 ;
        RECT 38.705 180.945 38.960 181.275 ;
        RECT 38.285 179.975 38.455 180.945 ;
        RECT 39.130 180.775 39.300 181.445 ;
        RECT 36.425 179.805 38.455 179.975 ;
        RECT 38.625 179.635 38.795 180.775 ;
        RECT 38.965 179.805 39.300 180.775 ;
        RECT 39.480 181.475 39.735 182.005 ;
        RECT 39.905 181.725 40.210 182.185 ;
        RECT 40.455 181.805 41.525 181.975 ;
        RECT 39.480 180.825 39.690 181.475 ;
        RECT 40.455 181.450 40.775 181.805 ;
        RECT 40.450 181.275 40.775 181.450 ;
        RECT 39.860 180.975 40.775 181.275 ;
        RECT 40.945 181.235 41.185 181.635 ;
        RECT 41.355 181.575 41.525 181.805 ;
        RECT 41.695 181.745 41.885 182.185 ;
        RECT 42.055 181.735 43.005 182.015 ;
        RECT 43.225 181.825 43.575 181.995 ;
        RECT 41.355 181.405 41.885 181.575 ;
        RECT 39.860 180.945 40.600 180.975 ;
        RECT 39.480 179.945 39.735 180.825 ;
        RECT 39.905 179.635 40.210 180.775 ;
        RECT 40.430 180.355 40.600 180.945 ;
        RECT 40.945 180.865 41.485 181.235 ;
        RECT 41.665 181.125 41.885 181.405 ;
        RECT 42.055 180.955 42.225 181.735 ;
        RECT 41.820 180.785 42.225 180.955 ;
        RECT 42.395 180.945 42.745 181.565 ;
        RECT 41.820 180.695 41.990 180.785 ;
        RECT 42.915 180.775 43.125 181.565 ;
        RECT 40.770 180.525 41.990 180.695 ;
        RECT 42.450 180.615 43.125 180.775 ;
        RECT 40.430 180.185 41.230 180.355 ;
        RECT 40.550 179.635 40.880 180.015 ;
        RECT 41.060 179.895 41.230 180.185 ;
        RECT 41.820 180.145 41.990 180.525 ;
        RECT 42.160 180.605 43.125 180.615 ;
        RECT 43.315 181.435 43.575 181.825 ;
        RECT 43.785 181.725 44.115 182.185 ;
        RECT 44.990 181.795 45.845 181.965 ;
        RECT 46.050 181.795 46.545 181.965 ;
        RECT 46.715 181.825 47.045 182.185 ;
        RECT 43.315 180.745 43.485 181.435 ;
        RECT 43.655 181.085 43.825 181.265 ;
        RECT 43.995 181.255 44.785 181.505 ;
        RECT 44.990 181.085 45.160 181.795 ;
        RECT 45.330 181.285 45.685 181.505 ;
        RECT 43.655 180.915 45.345 181.085 ;
        RECT 42.160 180.315 42.620 180.605 ;
        RECT 43.315 180.575 44.815 180.745 ;
        RECT 43.315 180.435 43.485 180.575 ;
        RECT 42.925 180.265 43.485 180.435 ;
        RECT 41.400 179.635 41.650 180.095 ;
        RECT 41.820 179.805 42.690 180.145 ;
        RECT 42.925 179.805 43.095 180.265 ;
        RECT 43.930 180.235 45.005 180.405 ;
        RECT 43.265 179.635 43.635 180.095 ;
        RECT 43.930 179.895 44.100 180.235 ;
        RECT 44.270 179.635 44.600 180.065 ;
        RECT 44.835 179.895 45.005 180.235 ;
        RECT 45.175 180.135 45.345 180.915 ;
        RECT 45.515 180.695 45.685 181.285 ;
        RECT 45.855 180.885 46.205 181.505 ;
        RECT 45.515 180.305 45.980 180.695 ;
        RECT 46.375 180.435 46.545 181.795 ;
        RECT 46.715 180.605 47.175 181.655 ;
        RECT 46.150 180.265 46.545 180.435 ;
        RECT 46.150 180.135 46.320 180.265 ;
        RECT 45.175 179.805 45.855 180.135 ;
        RECT 46.070 179.805 46.320 180.135 ;
        RECT 46.490 179.635 46.740 180.095 ;
        RECT 46.910 179.820 47.235 180.605 ;
        RECT 47.405 179.805 47.575 181.925 ;
        RECT 47.745 181.805 48.075 182.185 ;
        RECT 48.245 181.635 48.500 181.925 ;
        RECT 47.750 181.465 48.500 181.635 ;
        RECT 47.750 180.475 47.980 181.465 ;
        RECT 48.675 181.460 48.965 182.185 ;
        RECT 49.595 181.415 51.265 182.185 ;
        RECT 51.440 181.640 56.785 182.185 ;
        RECT 57.225 181.790 57.555 182.185 ;
        RECT 48.150 180.645 48.500 181.295 ;
        RECT 47.750 180.305 48.500 180.475 ;
        RECT 47.745 179.635 48.075 180.135 ;
        RECT 48.245 179.805 48.500 180.305 ;
        RECT 48.675 179.635 48.965 180.800 ;
        RECT 49.595 180.725 50.345 181.245 ;
        RECT 50.515 180.895 51.265 181.415 ;
        RECT 49.595 179.635 51.265 180.725 ;
        RECT 53.030 180.070 53.380 181.320 ;
        RECT 54.860 180.810 55.200 181.640 ;
        RECT 57.725 181.615 57.925 181.970 ;
        RECT 58.095 181.785 58.425 182.185 ;
        RECT 58.595 181.615 58.795 181.960 ;
        RECT 56.955 181.445 58.795 181.615 ;
        RECT 58.965 181.445 59.295 182.185 ;
        RECT 59.530 181.615 59.700 181.865 ;
        RECT 60.480 181.615 60.650 181.865 ;
        RECT 59.530 181.445 60.005 181.615 ;
        RECT 51.440 179.635 56.785 180.070 ;
        RECT 56.955 179.820 57.215 181.445 ;
        RECT 57.395 180.475 57.615 181.275 ;
        RECT 57.855 180.655 58.155 181.275 ;
        RECT 58.325 180.655 58.655 181.275 ;
        RECT 58.825 180.655 59.145 181.275 ;
        RECT 59.315 180.655 59.665 181.275 ;
        RECT 59.835 180.475 60.005 181.445 ;
        RECT 57.395 180.265 60.005 180.475 ;
        RECT 60.175 181.445 60.650 181.615 ;
        RECT 60.885 181.445 61.215 182.185 ;
        RECT 61.385 181.615 61.585 181.960 ;
        RECT 61.755 181.785 62.085 182.185 ;
        RECT 62.255 181.615 62.455 181.970 ;
        RECT 62.625 181.790 62.955 182.185 ;
        RECT 63.395 181.685 63.655 182.015 ;
        RECT 63.965 181.805 64.295 182.185 ;
        RECT 64.475 181.845 65.955 182.015 ;
        RECT 61.385 181.445 63.225 181.615 ;
        RECT 60.175 180.475 60.345 181.445 ;
        RECT 60.515 180.655 60.865 181.275 ;
        RECT 61.035 180.655 61.355 181.275 ;
        RECT 61.525 180.655 61.855 181.275 ;
        RECT 62.025 180.655 62.325 181.275 ;
        RECT 62.565 180.475 62.785 181.275 ;
        RECT 60.175 180.265 62.785 180.475 ;
        RECT 58.965 179.635 59.295 180.085 ;
        RECT 60.885 179.635 61.215 180.085 ;
        RECT 62.965 179.820 63.225 181.445 ;
        RECT 63.395 180.985 63.565 181.685 ;
        RECT 64.475 181.515 64.875 181.845 ;
        RECT 63.915 181.325 64.125 181.505 ;
        RECT 63.915 181.155 64.535 181.325 ;
        RECT 64.705 181.035 64.875 181.515 ;
        RECT 65.065 181.345 65.615 181.675 ;
        RECT 63.395 180.815 64.525 180.985 ;
        RECT 64.705 180.865 65.275 181.035 ;
        RECT 63.395 180.135 63.565 180.815 ;
        RECT 64.355 180.695 64.525 180.815 ;
        RECT 63.735 180.315 64.085 180.645 ;
        RECT 64.355 180.525 64.935 180.695 ;
        RECT 65.105 180.355 65.275 180.865 ;
        RECT 64.535 180.185 65.275 180.355 ;
        RECT 65.445 180.355 65.615 181.345 ;
        RECT 65.785 180.945 65.955 181.845 ;
        RECT 66.205 181.275 66.390 181.855 ;
        RECT 66.660 181.275 66.855 181.850 ;
        RECT 67.065 181.805 67.395 182.185 ;
        RECT 66.205 180.945 66.435 181.275 ;
        RECT 66.660 180.945 66.915 181.275 ;
        RECT 66.205 180.635 66.390 180.945 ;
        RECT 66.660 180.635 66.855 180.945 ;
        RECT 67.225 180.355 67.395 181.275 ;
        RECT 65.445 180.185 67.395 180.355 ;
        RECT 63.395 179.805 63.655 180.135 ;
        RECT 63.965 179.635 64.295 180.015 ;
        RECT 64.535 179.805 64.725 180.185 ;
        RECT 64.975 179.635 65.305 180.015 ;
        RECT 65.515 179.805 65.685 180.185 ;
        RECT 65.880 179.635 66.210 180.015 ;
        RECT 66.470 179.805 66.640 180.185 ;
        RECT 67.065 179.635 67.395 180.015 ;
        RECT 67.565 179.805 67.825 182.015 ;
        RECT 68.515 181.365 68.725 182.185 ;
        RECT 68.895 181.385 69.225 182.015 ;
        RECT 68.895 180.785 69.145 181.385 ;
        RECT 69.395 181.365 69.625 182.185 ;
        RECT 70.570 181.375 70.815 181.980 ;
        RECT 71.035 181.650 71.545 182.185 ;
        RECT 70.295 181.205 71.525 181.375 ;
        RECT 69.315 180.945 69.645 181.195 ;
        RECT 68.515 179.635 68.725 180.775 ;
        RECT 68.895 179.805 69.225 180.785 ;
        RECT 69.395 179.635 69.625 180.775 ;
        RECT 70.295 180.395 70.635 181.205 ;
        RECT 70.805 180.640 71.555 180.830 ;
        RECT 70.295 179.985 70.810 180.395 ;
        RECT 71.045 179.635 71.215 180.395 ;
        RECT 71.385 179.975 71.555 180.640 ;
        RECT 71.725 180.655 71.915 182.015 ;
        RECT 72.085 181.165 72.360 182.015 ;
        RECT 72.550 181.650 73.080 182.015 ;
        RECT 73.505 181.785 73.835 182.185 ;
        RECT 72.905 181.615 73.080 181.650 ;
        RECT 72.085 180.995 72.365 181.165 ;
        RECT 72.085 180.855 72.360 180.995 ;
        RECT 72.565 180.655 72.735 181.455 ;
        RECT 71.725 180.485 72.735 180.655 ;
        RECT 72.905 181.445 73.835 181.615 ;
        RECT 74.005 181.445 74.260 182.015 ;
        RECT 74.435 181.460 74.725 182.185 ;
        RECT 72.905 180.315 73.075 181.445 ;
        RECT 73.665 181.275 73.835 181.445 ;
        RECT 71.950 180.145 73.075 180.315 ;
        RECT 73.245 180.945 73.440 181.275 ;
        RECT 73.665 180.945 73.920 181.275 ;
        RECT 73.245 179.975 73.415 180.945 ;
        RECT 74.090 180.775 74.260 181.445 ;
        RECT 75.630 181.375 75.875 181.980 ;
        RECT 76.095 181.650 76.605 182.185 ;
        RECT 75.355 181.205 76.585 181.375 ;
        RECT 71.385 179.805 73.415 179.975 ;
        RECT 73.585 179.635 73.755 180.775 ;
        RECT 73.925 179.805 74.260 180.775 ;
        RECT 74.435 179.635 74.725 180.800 ;
        RECT 75.355 180.395 75.695 181.205 ;
        RECT 75.865 180.640 76.615 180.830 ;
        RECT 75.355 179.985 75.870 180.395 ;
        RECT 76.105 179.635 76.275 180.395 ;
        RECT 76.445 179.975 76.615 180.640 ;
        RECT 76.785 180.655 76.975 182.015 ;
        RECT 77.145 181.165 77.420 182.015 ;
        RECT 77.610 181.650 78.140 182.015 ;
        RECT 78.565 181.785 78.895 182.185 ;
        RECT 77.965 181.615 78.140 181.650 ;
        RECT 77.145 180.995 77.425 181.165 ;
        RECT 77.145 180.855 77.420 180.995 ;
        RECT 77.625 180.655 77.795 181.455 ;
        RECT 76.785 180.485 77.795 180.655 ;
        RECT 77.965 181.445 78.895 181.615 ;
        RECT 79.065 181.445 79.320 182.015 ;
        RECT 77.965 180.315 78.135 181.445 ;
        RECT 78.725 181.275 78.895 181.445 ;
        RECT 77.010 180.145 78.135 180.315 ;
        RECT 78.305 180.945 78.500 181.275 ;
        RECT 78.725 180.945 78.980 181.275 ;
        RECT 78.305 179.975 78.475 180.945 ;
        RECT 79.150 180.775 79.320 181.445 ;
        RECT 79.495 181.415 81.165 182.185 ;
        RECT 76.445 179.805 78.475 179.975 ;
        RECT 78.645 179.635 78.815 180.775 ;
        RECT 78.985 179.805 79.320 180.775 ;
        RECT 79.495 180.725 80.245 181.245 ;
        RECT 80.415 180.895 81.165 181.415 ;
        RECT 81.340 181.475 81.595 182.005 ;
        RECT 81.765 181.725 82.070 182.185 ;
        RECT 82.315 181.805 83.385 181.975 ;
        RECT 81.340 180.825 81.550 181.475 ;
        RECT 82.315 181.450 82.635 181.805 ;
        RECT 82.310 181.275 82.635 181.450 ;
        RECT 81.720 180.975 82.635 181.275 ;
        RECT 82.805 181.235 83.045 181.635 ;
        RECT 83.215 181.575 83.385 181.805 ;
        RECT 83.555 181.745 83.745 182.185 ;
        RECT 83.915 181.735 84.865 182.015 ;
        RECT 85.085 181.825 85.435 181.995 ;
        RECT 83.215 181.405 83.745 181.575 ;
        RECT 81.720 180.945 82.460 180.975 ;
        RECT 79.495 179.635 81.165 180.725 ;
        RECT 81.340 179.945 81.595 180.825 ;
        RECT 81.765 179.635 82.070 180.775 ;
        RECT 82.290 180.355 82.460 180.945 ;
        RECT 82.805 180.865 83.345 181.235 ;
        RECT 83.525 181.125 83.745 181.405 ;
        RECT 83.915 180.955 84.085 181.735 ;
        RECT 83.680 180.785 84.085 180.955 ;
        RECT 84.255 180.945 84.605 181.565 ;
        RECT 83.680 180.695 83.850 180.785 ;
        RECT 84.775 180.775 84.985 181.565 ;
        RECT 82.630 180.525 83.850 180.695 ;
        RECT 84.310 180.615 84.985 180.775 ;
        RECT 82.290 180.185 83.090 180.355 ;
        RECT 82.410 179.635 82.740 180.015 ;
        RECT 82.920 179.895 83.090 180.185 ;
        RECT 83.680 180.145 83.850 180.525 ;
        RECT 84.020 180.605 84.985 180.615 ;
        RECT 85.175 181.435 85.435 181.825 ;
        RECT 85.645 181.725 85.975 182.185 ;
        RECT 86.850 181.795 87.705 181.965 ;
        RECT 87.910 181.795 88.405 181.965 ;
        RECT 88.575 181.825 88.905 182.185 ;
        RECT 85.175 180.745 85.345 181.435 ;
        RECT 85.515 181.085 85.685 181.265 ;
        RECT 85.855 181.255 86.645 181.505 ;
        RECT 86.850 181.085 87.020 181.795 ;
        RECT 87.190 181.285 87.545 181.505 ;
        RECT 85.515 180.915 87.205 181.085 ;
        RECT 84.020 180.315 84.480 180.605 ;
        RECT 85.175 180.575 86.675 180.745 ;
        RECT 85.175 180.435 85.345 180.575 ;
        RECT 84.785 180.265 85.345 180.435 ;
        RECT 83.260 179.635 83.510 180.095 ;
        RECT 83.680 179.805 84.550 180.145 ;
        RECT 84.785 179.805 84.955 180.265 ;
        RECT 85.790 180.235 86.865 180.405 ;
        RECT 85.125 179.635 85.495 180.095 ;
        RECT 85.790 179.895 85.960 180.235 ;
        RECT 86.130 179.635 86.460 180.065 ;
        RECT 86.695 179.895 86.865 180.235 ;
        RECT 87.035 180.135 87.205 180.915 ;
        RECT 87.375 180.695 87.545 181.285 ;
        RECT 87.715 180.885 88.065 181.505 ;
        RECT 87.375 180.305 87.840 180.695 ;
        RECT 88.235 180.435 88.405 181.795 ;
        RECT 88.575 180.605 89.035 181.655 ;
        RECT 88.010 180.265 88.405 180.435 ;
        RECT 88.010 180.135 88.180 180.265 ;
        RECT 87.035 179.805 87.715 180.135 ;
        RECT 87.930 179.805 88.180 180.135 ;
        RECT 88.350 179.635 88.600 180.095 ;
        RECT 88.770 179.820 89.095 180.605 ;
        RECT 89.265 179.805 89.435 181.925 ;
        RECT 89.605 181.805 89.935 182.185 ;
        RECT 90.105 181.635 90.360 181.925 ;
        RECT 89.610 181.465 90.360 181.635 ;
        RECT 89.610 180.475 89.840 181.465 ;
        RECT 91.000 181.445 91.255 182.015 ;
        RECT 91.425 181.785 91.755 182.185 ;
        RECT 92.180 181.650 92.710 182.015 ;
        RECT 92.180 181.615 92.355 181.650 ;
        RECT 91.425 181.445 92.355 181.615 ;
        RECT 92.900 181.505 93.175 182.015 ;
        RECT 90.010 180.645 90.360 181.295 ;
        RECT 91.000 180.775 91.170 181.445 ;
        RECT 91.425 181.275 91.595 181.445 ;
        RECT 91.340 180.945 91.595 181.275 ;
        RECT 91.820 180.945 92.015 181.275 ;
        RECT 89.610 180.305 90.360 180.475 ;
        RECT 89.605 179.635 89.935 180.135 ;
        RECT 90.105 179.805 90.360 180.305 ;
        RECT 91.000 179.805 91.335 180.775 ;
        RECT 91.505 179.635 91.675 180.775 ;
        RECT 91.845 179.975 92.015 180.945 ;
        RECT 92.185 180.315 92.355 181.445 ;
        RECT 92.525 180.655 92.695 181.455 ;
        RECT 92.895 181.335 93.175 181.505 ;
        RECT 92.900 180.855 93.175 181.335 ;
        RECT 93.345 180.655 93.535 182.015 ;
        RECT 93.715 181.650 94.225 182.185 ;
        RECT 94.445 181.375 94.690 181.980 ;
        RECT 96.330 181.375 96.575 181.980 ;
        RECT 96.795 181.650 97.305 182.185 ;
        RECT 93.735 181.205 94.965 181.375 ;
        RECT 92.525 180.485 93.535 180.655 ;
        RECT 93.705 180.640 94.455 180.830 ;
        RECT 92.185 180.145 93.310 180.315 ;
        RECT 93.705 179.975 93.875 180.640 ;
        RECT 94.625 180.395 94.965 181.205 ;
        RECT 91.845 179.805 93.875 179.975 ;
        RECT 94.045 179.635 94.215 180.395 ;
        RECT 94.450 179.985 94.965 180.395 ;
        RECT 96.055 181.205 97.285 181.375 ;
        RECT 96.055 180.395 96.395 181.205 ;
        RECT 96.565 180.640 97.315 180.830 ;
        RECT 96.055 179.985 96.570 180.395 ;
        RECT 96.805 179.635 96.975 180.395 ;
        RECT 97.145 179.975 97.315 180.640 ;
        RECT 97.485 180.655 97.675 182.015 ;
        RECT 97.845 181.505 98.120 182.015 ;
        RECT 98.310 181.650 98.840 182.015 ;
        RECT 99.265 181.785 99.595 182.185 ;
        RECT 98.665 181.615 98.840 181.650 ;
        RECT 97.845 181.335 98.125 181.505 ;
        RECT 97.845 180.855 98.120 181.335 ;
        RECT 98.325 180.655 98.495 181.455 ;
        RECT 97.485 180.485 98.495 180.655 ;
        RECT 98.665 181.445 99.595 181.615 ;
        RECT 99.765 181.445 100.020 182.015 ;
        RECT 100.195 181.460 100.485 182.185 ;
        RECT 100.660 181.475 100.915 182.005 ;
        RECT 101.085 181.725 101.390 182.185 ;
        RECT 101.635 181.805 102.705 181.975 ;
        RECT 98.665 180.315 98.835 181.445 ;
        RECT 99.425 181.275 99.595 181.445 ;
        RECT 97.710 180.145 98.835 180.315 ;
        RECT 99.005 180.945 99.200 181.275 ;
        RECT 99.425 180.945 99.680 181.275 ;
        RECT 99.005 179.975 99.175 180.945 ;
        RECT 99.850 180.775 100.020 181.445 ;
        RECT 100.660 180.825 100.870 181.475 ;
        RECT 101.635 181.450 101.955 181.805 ;
        RECT 101.630 181.275 101.955 181.450 ;
        RECT 101.040 180.975 101.955 181.275 ;
        RECT 102.125 181.235 102.365 181.635 ;
        RECT 102.535 181.575 102.705 181.805 ;
        RECT 102.875 181.745 103.065 182.185 ;
        RECT 103.235 181.735 104.185 182.015 ;
        RECT 104.405 181.825 104.755 181.995 ;
        RECT 102.535 181.405 103.065 181.575 ;
        RECT 101.040 180.945 101.780 180.975 ;
        RECT 97.145 179.805 99.175 179.975 ;
        RECT 99.345 179.635 99.515 180.775 ;
        RECT 99.685 179.805 100.020 180.775 ;
        RECT 100.195 179.635 100.485 180.800 ;
        RECT 100.660 179.945 100.915 180.825 ;
        RECT 101.085 179.635 101.390 180.775 ;
        RECT 101.610 180.355 101.780 180.945 ;
        RECT 102.125 180.865 102.665 181.235 ;
        RECT 102.845 181.125 103.065 181.405 ;
        RECT 103.235 180.955 103.405 181.735 ;
        RECT 103.000 180.785 103.405 180.955 ;
        RECT 103.575 180.945 103.925 181.565 ;
        RECT 103.000 180.695 103.170 180.785 ;
        RECT 104.095 180.775 104.305 181.565 ;
        RECT 101.950 180.525 103.170 180.695 ;
        RECT 103.630 180.615 104.305 180.775 ;
        RECT 101.610 180.185 102.410 180.355 ;
        RECT 101.730 179.635 102.060 180.015 ;
        RECT 102.240 179.895 102.410 180.185 ;
        RECT 103.000 180.145 103.170 180.525 ;
        RECT 103.340 180.605 104.305 180.615 ;
        RECT 104.495 181.435 104.755 181.825 ;
        RECT 104.965 181.725 105.295 182.185 ;
        RECT 106.170 181.795 107.025 181.965 ;
        RECT 107.230 181.795 107.725 181.965 ;
        RECT 107.895 181.825 108.225 182.185 ;
        RECT 104.495 180.745 104.665 181.435 ;
        RECT 104.835 181.085 105.005 181.265 ;
        RECT 105.175 181.255 105.965 181.505 ;
        RECT 106.170 181.085 106.340 181.795 ;
        RECT 106.510 181.285 106.865 181.505 ;
        RECT 104.835 180.915 106.525 181.085 ;
        RECT 103.340 180.315 103.800 180.605 ;
        RECT 104.495 180.575 105.995 180.745 ;
        RECT 104.495 180.435 104.665 180.575 ;
        RECT 104.105 180.265 104.665 180.435 ;
        RECT 102.580 179.635 102.830 180.095 ;
        RECT 103.000 179.805 103.870 180.145 ;
        RECT 104.105 179.805 104.275 180.265 ;
        RECT 105.110 180.235 106.185 180.405 ;
        RECT 104.445 179.635 104.815 180.095 ;
        RECT 105.110 179.895 105.280 180.235 ;
        RECT 105.450 179.635 105.780 180.065 ;
        RECT 106.015 179.895 106.185 180.235 ;
        RECT 106.355 180.135 106.525 180.915 ;
        RECT 106.695 180.695 106.865 181.285 ;
        RECT 107.035 180.885 107.385 181.505 ;
        RECT 106.695 180.305 107.160 180.695 ;
        RECT 107.555 180.435 107.725 181.795 ;
        RECT 107.895 180.605 108.355 181.655 ;
        RECT 107.330 180.265 107.725 180.435 ;
        RECT 107.330 180.135 107.500 180.265 ;
        RECT 106.355 179.805 107.035 180.135 ;
        RECT 107.250 179.805 107.500 180.135 ;
        RECT 107.670 179.635 107.920 180.095 ;
        RECT 108.090 179.820 108.415 180.605 ;
        RECT 108.585 179.805 108.755 181.925 ;
        RECT 108.925 181.805 109.255 182.185 ;
        RECT 109.425 181.635 109.680 181.925 ;
        RECT 108.930 181.465 109.680 181.635 ;
        RECT 108.930 180.475 109.160 181.465 ;
        RECT 110.315 181.415 111.985 182.185 ;
        RECT 112.155 181.435 113.365 182.185 ;
        RECT 109.330 180.645 109.680 181.295 ;
        RECT 110.315 180.725 111.065 181.245 ;
        RECT 111.235 180.895 111.985 181.415 ;
        RECT 112.155 180.725 112.675 181.265 ;
        RECT 112.845 180.895 113.365 181.435 ;
        RECT 108.930 180.305 109.680 180.475 ;
        RECT 108.925 179.635 109.255 180.135 ;
        RECT 109.425 179.805 109.680 180.305 ;
        RECT 110.315 179.635 111.985 180.725 ;
        RECT 112.155 179.635 113.365 180.725 ;
        RECT 11.330 179.465 113.450 179.635 ;
        RECT 11.415 178.375 12.625 179.465 ;
        RECT 11.415 177.665 11.935 178.205 ;
        RECT 12.105 177.835 12.625 178.375 ;
        RECT 13.255 178.375 14.925 179.465 ;
        RECT 15.100 179.030 20.445 179.465 ;
        RECT 13.255 177.855 14.005 178.375 ;
        RECT 14.175 177.685 14.925 178.205 ;
        RECT 16.690 177.780 17.040 179.030 ;
        RECT 20.620 178.795 20.875 179.295 ;
        RECT 21.045 178.965 21.375 179.465 ;
        RECT 20.620 178.625 21.370 178.795 ;
        RECT 11.415 176.915 12.625 177.665 ;
        RECT 13.255 176.915 14.925 177.685 ;
        RECT 18.520 177.460 18.860 178.290 ;
        RECT 20.620 177.805 20.970 178.455 ;
        RECT 21.140 177.635 21.370 178.625 ;
        RECT 20.620 177.465 21.370 177.635 ;
        RECT 15.100 176.915 20.445 177.460 ;
        RECT 20.620 177.175 20.875 177.465 ;
        RECT 21.045 176.915 21.375 177.295 ;
        RECT 21.545 177.175 21.715 179.295 ;
        RECT 21.885 178.495 22.210 179.280 ;
        RECT 22.380 179.005 22.630 179.465 ;
        RECT 22.800 178.965 23.050 179.295 ;
        RECT 23.265 178.965 23.945 179.295 ;
        RECT 22.800 178.835 22.970 178.965 ;
        RECT 22.575 178.665 22.970 178.835 ;
        RECT 21.945 177.445 22.405 178.495 ;
        RECT 22.575 177.305 22.745 178.665 ;
        RECT 23.140 178.405 23.605 178.795 ;
        RECT 22.915 177.595 23.265 178.215 ;
        RECT 23.435 177.815 23.605 178.405 ;
        RECT 23.775 178.185 23.945 178.965 ;
        RECT 24.115 178.865 24.285 179.205 ;
        RECT 24.520 179.035 24.850 179.465 ;
        RECT 25.020 178.865 25.190 179.205 ;
        RECT 25.485 179.005 25.855 179.465 ;
        RECT 24.115 178.695 25.190 178.865 ;
        RECT 26.025 178.835 26.195 179.295 ;
        RECT 26.430 178.955 27.300 179.295 ;
        RECT 27.470 179.005 27.720 179.465 ;
        RECT 25.635 178.665 26.195 178.835 ;
        RECT 25.635 178.525 25.805 178.665 ;
        RECT 24.305 178.355 25.805 178.525 ;
        RECT 26.500 178.495 26.960 178.785 ;
        RECT 23.775 178.015 25.465 178.185 ;
        RECT 23.435 177.595 23.790 177.815 ;
        RECT 23.960 177.305 24.130 178.015 ;
        RECT 24.335 177.595 25.125 177.845 ;
        RECT 25.295 177.835 25.465 178.015 ;
        RECT 25.635 177.665 25.805 178.355 ;
        RECT 22.075 176.915 22.405 177.275 ;
        RECT 22.575 177.135 23.070 177.305 ;
        RECT 23.275 177.135 24.130 177.305 ;
        RECT 25.005 176.915 25.335 177.375 ;
        RECT 25.545 177.275 25.805 177.665 ;
        RECT 25.995 178.485 26.960 178.495 ;
        RECT 27.130 178.575 27.300 178.955 ;
        RECT 27.890 178.915 28.060 179.205 ;
        RECT 28.240 179.085 28.570 179.465 ;
        RECT 27.890 178.745 28.690 178.915 ;
        RECT 25.995 178.325 26.670 178.485 ;
        RECT 27.130 178.405 28.350 178.575 ;
        RECT 25.995 177.535 26.205 178.325 ;
        RECT 27.130 178.315 27.300 178.405 ;
        RECT 26.375 177.535 26.725 178.155 ;
        RECT 26.895 178.145 27.300 178.315 ;
        RECT 26.895 177.365 27.065 178.145 ;
        RECT 27.235 177.695 27.455 177.975 ;
        RECT 27.635 177.865 28.175 178.235 ;
        RECT 28.520 178.155 28.690 178.745 ;
        RECT 28.910 178.325 29.215 179.465 ;
        RECT 29.385 178.275 29.640 179.155 ;
        RECT 28.520 178.125 29.260 178.155 ;
        RECT 27.235 177.525 27.765 177.695 ;
        RECT 25.545 177.105 25.895 177.275 ;
        RECT 26.115 177.085 27.065 177.365 ;
        RECT 27.235 176.915 27.425 177.355 ;
        RECT 27.595 177.295 27.765 177.525 ;
        RECT 27.935 177.465 28.175 177.865 ;
        RECT 28.345 177.825 29.260 178.125 ;
        RECT 28.345 177.650 28.670 177.825 ;
        RECT 28.345 177.295 28.665 177.650 ;
        RECT 29.430 177.625 29.640 178.275 ;
        RECT 30.275 178.375 31.945 179.465 ;
        RECT 32.320 178.495 32.650 179.295 ;
        RECT 32.820 178.665 33.150 179.465 ;
        RECT 33.450 178.495 33.780 179.295 ;
        RECT 34.425 178.665 34.675 179.465 ;
        RECT 30.275 177.855 31.025 178.375 ;
        RECT 32.320 178.325 34.755 178.495 ;
        RECT 34.945 178.325 35.115 179.465 ;
        RECT 35.285 178.325 35.625 179.295 ;
        RECT 31.195 177.685 31.945 178.205 ;
        RECT 32.115 177.905 32.465 178.155 ;
        RECT 32.650 177.695 32.820 178.325 ;
        RECT 32.990 177.905 33.320 178.105 ;
        RECT 33.490 177.905 33.820 178.105 ;
        RECT 33.990 177.905 34.410 178.105 ;
        RECT 34.585 178.075 34.755 178.325 ;
        RECT 34.585 177.905 35.280 178.075 ;
        RECT 27.595 177.125 28.665 177.295 ;
        RECT 28.910 176.915 29.215 177.375 ;
        RECT 29.385 177.095 29.640 177.625 ;
        RECT 30.275 176.915 31.945 177.685 ;
        RECT 32.320 177.085 32.820 177.695 ;
        RECT 33.450 177.565 34.675 177.735 ;
        RECT 35.450 177.715 35.625 178.325 ;
        RECT 35.795 178.300 36.085 179.465 ;
        RECT 36.715 178.375 39.305 179.465 ;
        RECT 36.715 177.855 37.925 178.375 ;
        RECT 39.475 178.325 39.815 179.295 ;
        RECT 39.985 178.325 40.155 179.465 ;
        RECT 40.425 178.665 40.675 179.465 ;
        RECT 41.320 178.495 41.650 179.295 ;
        RECT 41.950 178.665 42.280 179.465 ;
        RECT 42.450 178.495 42.780 179.295 ;
        RECT 43.270 178.835 43.555 179.295 ;
        RECT 43.725 179.005 43.995 179.465 ;
        RECT 43.270 178.615 44.225 178.835 ;
        RECT 40.345 178.325 42.780 178.495 ;
        RECT 33.450 177.085 33.780 177.565 ;
        RECT 33.950 176.915 34.175 177.375 ;
        RECT 34.345 177.085 34.675 177.565 ;
        RECT 34.865 176.915 35.115 177.715 ;
        RECT 35.285 177.085 35.625 177.715 ;
        RECT 38.095 177.685 39.305 178.205 ;
        RECT 35.795 176.915 36.085 177.640 ;
        RECT 36.715 176.915 39.305 177.685 ;
        RECT 39.475 177.715 39.650 178.325 ;
        RECT 40.345 178.075 40.515 178.325 ;
        RECT 39.820 177.905 40.515 178.075 ;
        RECT 40.690 177.905 41.110 178.105 ;
        RECT 41.280 177.905 41.610 178.105 ;
        RECT 41.780 177.905 42.110 178.105 ;
        RECT 39.475 177.085 39.815 177.715 ;
        RECT 39.985 176.915 40.235 177.715 ;
        RECT 40.425 177.565 41.650 177.735 ;
        RECT 40.425 177.085 40.755 177.565 ;
        RECT 40.925 176.915 41.150 177.375 ;
        RECT 41.320 177.085 41.650 177.565 ;
        RECT 42.280 177.695 42.450 178.325 ;
        RECT 42.635 177.905 42.985 178.155 ;
        RECT 43.155 177.885 43.845 178.445 ;
        RECT 44.015 177.715 44.225 178.615 ;
        RECT 42.280 177.085 42.780 177.695 ;
        RECT 43.270 177.545 44.225 177.715 ;
        RECT 44.395 178.445 44.795 179.295 ;
        RECT 44.985 178.835 45.265 179.295 ;
        RECT 45.785 179.005 46.110 179.465 ;
        RECT 44.985 178.615 46.110 178.835 ;
        RECT 44.395 177.885 45.490 178.445 ;
        RECT 45.660 178.155 46.110 178.615 ;
        RECT 46.280 178.325 46.665 179.295 ;
        RECT 43.270 177.085 43.555 177.545 ;
        RECT 43.725 176.915 43.995 177.375 ;
        RECT 44.395 177.085 44.795 177.885 ;
        RECT 45.660 177.825 46.215 178.155 ;
        RECT 45.660 177.715 46.110 177.825 ;
        RECT 44.985 177.545 46.110 177.715 ;
        RECT 46.385 177.655 46.665 178.325 ;
        RECT 44.985 177.085 45.265 177.545 ;
        RECT 45.785 176.915 46.110 177.375 ;
        RECT 46.280 177.085 46.665 177.655 ;
        RECT 46.835 178.390 47.105 179.295 ;
        RECT 47.275 178.705 47.605 179.465 ;
        RECT 47.785 178.535 47.955 179.295 ;
        RECT 46.835 177.590 47.005 178.390 ;
        RECT 47.290 178.365 47.955 178.535 ;
        RECT 48.215 178.375 50.805 179.465 ;
        RECT 51.065 178.535 51.235 179.295 ;
        RECT 51.415 178.705 51.745 179.465 ;
        RECT 47.290 178.220 47.460 178.365 ;
        RECT 47.175 177.890 47.460 178.220 ;
        RECT 47.290 177.635 47.460 177.890 ;
        RECT 47.695 177.815 48.025 178.185 ;
        RECT 48.215 177.855 49.425 178.375 ;
        RECT 51.065 178.365 51.730 178.535 ;
        RECT 51.915 178.390 52.185 179.295 ;
        RECT 52.410 178.595 52.695 179.465 ;
        RECT 52.865 178.835 53.125 179.295 ;
        RECT 53.300 179.005 53.555 179.465 ;
        RECT 53.725 178.835 53.985 179.295 ;
        RECT 52.865 178.665 53.985 178.835 ;
        RECT 54.155 178.665 54.465 179.465 ;
        RECT 52.865 178.415 53.125 178.665 ;
        RECT 54.635 178.495 54.945 179.295 ;
        RECT 51.560 178.220 51.730 178.365 ;
        RECT 49.595 177.685 50.805 178.205 ;
        RECT 50.995 177.815 51.325 178.185 ;
        RECT 51.560 177.890 51.845 178.220 ;
        RECT 46.835 177.085 47.095 177.590 ;
        RECT 47.290 177.465 47.955 177.635 ;
        RECT 47.275 176.915 47.605 177.295 ;
        RECT 47.785 177.085 47.955 177.465 ;
        RECT 48.215 176.915 50.805 177.685 ;
        RECT 51.560 177.635 51.730 177.890 ;
        RECT 51.065 177.465 51.730 177.635 ;
        RECT 52.015 177.590 52.185 178.390 ;
        RECT 51.065 177.085 51.235 177.465 ;
        RECT 51.415 176.915 51.745 177.295 ;
        RECT 51.925 177.085 52.185 177.590 ;
        RECT 52.370 178.245 53.125 178.415 ;
        RECT 53.915 178.325 54.945 178.495 ;
        RECT 52.370 177.735 52.775 178.245 ;
        RECT 53.915 178.075 54.085 178.325 ;
        RECT 52.945 177.905 54.085 178.075 ;
        RECT 52.370 177.565 54.020 177.735 ;
        RECT 54.255 177.585 54.605 178.155 ;
        RECT 52.415 176.915 52.695 177.395 ;
        RECT 52.865 177.175 53.125 177.565 ;
        RECT 53.300 176.915 53.555 177.395 ;
        RECT 53.725 177.175 54.020 177.565 ;
        RECT 54.775 177.415 54.945 178.325 ;
        RECT 55.575 178.375 57.245 179.465 ;
        RECT 57.425 178.485 57.755 179.295 ;
        RECT 57.925 178.665 58.165 179.465 ;
        RECT 55.575 177.855 56.325 178.375 ;
        RECT 57.425 178.315 58.140 178.485 ;
        RECT 56.495 177.685 57.245 178.205 ;
        RECT 57.420 177.905 57.800 178.145 ;
        RECT 57.970 178.075 58.140 178.315 ;
        RECT 58.345 178.445 58.515 179.295 ;
        RECT 58.685 178.665 59.015 179.465 ;
        RECT 59.185 178.445 59.355 179.295 ;
        RECT 58.345 178.275 59.355 178.445 ;
        RECT 59.525 178.315 59.855 179.465 ;
        RECT 60.175 178.375 61.385 179.465 ;
        RECT 57.970 177.905 58.470 178.075 ;
        RECT 57.970 177.735 58.140 177.905 ;
        RECT 58.860 177.735 59.355 178.275 ;
        RECT 60.175 177.835 60.695 178.375 ;
        RECT 61.555 178.300 61.845 179.465 ;
        RECT 62.055 178.325 62.285 179.465 ;
        RECT 62.455 178.315 62.785 179.295 ;
        RECT 62.955 178.325 63.165 179.465 ;
        RECT 54.200 176.915 54.475 177.395 ;
        RECT 54.645 177.085 54.945 177.415 ;
        RECT 55.575 176.915 57.245 177.685 ;
        RECT 57.505 177.565 58.140 177.735 ;
        RECT 58.345 177.565 59.355 177.735 ;
        RECT 57.505 177.085 57.675 177.565 ;
        RECT 57.855 176.915 58.095 177.395 ;
        RECT 58.345 177.085 58.515 177.565 ;
        RECT 58.685 176.915 59.015 177.395 ;
        RECT 59.185 177.085 59.355 177.565 ;
        RECT 59.525 176.915 59.855 177.715 ;
        RECT 60.865 177.665 61.385 178.205 ;
        RECT 62.035 177.905 62.365 178.155 ;
        RECT 60.175 176.915 61.385 177.665 ;
        RECT 61.555 176.915 61.845 177.640 ;
        RECT 62.055 176.915 62.285 177.735 ;
        RECT 62.535 177.715 62.785 178.315 ;
        RECT 62.455 177.085 62.785 177.715 ;
        RECT 62.955 176.915 63.165 177.735 ;
        RECT 63.395 177.655 63.655 179.280 ;
        RECT 65.405 179.015 65.735 179.465 ;
        RECT 63.835 178.625 66.445 178.835 ;
        RECT 63.835 177.825 64.055 178.625 ;
        RECT 64.295 177.825 64.595 178.445 ;
        RECT 64.765 177.825 65.095 178.445 ;
        RECT 65.265 177.825 65.585 178.445 ;
        RECT 65.755 177.825 66.105 178.445 ;
        RECT 66.275 177.655 66.445 178.625 ;
        RECT 63.395 177.485 65.235 177.655 ;
        RECT 63.665 176.915 63.995 177.310 ;
        RECT 64.165 177.130 64.365 177.485 ;
        RECT 64.535 176.915 64.865 177.315 ;
        RECT 65.035 177.140 65.235 177.485 ;
        RECT 65.405 176.915 65.735 177.655 ;
        RECT 65.970 177.485 66.445 177.655 ;
        RECT 67.075 178.495 67.385 179.295 ;
        RECT 67.555 178.665 67.865 179.465 ;
        RECT 68.035 178.835 68.295 179.295 ;
        RECT 68.465 179.005 68.720 179.465 ;
        RECT 68.895 178.835 69.155 179.295 ;
        RECT 68.035 178.665 69.155 178.835 ;
        RECT 67.075 178.325 68.105 178.495 ;
        RECT 65.970 177.235 66.140 177.485 ;
        RECT 67.075 177.415 67.245 178.325 ;
        RECT 67.415 177.585 67.765 178.155 ;
        RECT 67.935 178.075 68.105 178.325 ;
        RECT 68.895 178.415 69.155 178.665 ;
        RECT 69.325 178.595 69.610 179.465 ;
        RECT 69.950 178.835 70.235 179.295 ;
        RECT 70.405 179.005 70.675 179.465 ;
        RECT 69.950 178.615 70.905 178.835 ;
        RECT 68.895 178.245 69.650 178.415 ;
        RECT 67.935 177.905 69.075 178.075 ;
        RECT 69.245 177.735 69.650 178.245 ;
        RECT 69.835 177.885 70.525 178.445 ;
        RECT 68.000 177.565 69.650 177.735 ;
        RECT 70.695 177.715 70.905 178.615 ;
        RECT 67.075 177.085 67.375 177.415 ;
        RECT 67.545 176.915 67.820 177.395 ;
        RECT 68.000 177.175 68.295 177.565 ;
        RECT 68.465 176.915 68.720 177.395 ;
        RECT 68.895 177.175 69.155 177.565 ;
        RECT 69.950 177.545 70.905 177.715 ;
        RECT 71.075 178.445 71.475 179.295 ;
        RECT 71.665 178.835 71.945 179.295 ;
        RECT 72.465 179.005 72.790 179.465 ;
        RECT 71.665 178.615 72.790 178.835 ;
        RECT 71.075 177.885 72.170 178.445 ;
        RECT 72.340 178.155 72.790 178.615 ;
        RECT 72.960 178.325 73.345 179.295 ;
        RECT 69.325 176.915 69.605 177.395 ;
        RECT 69.950 177.085 70.235 177.545 ;
        RECT 70.405 176.915 70.675 177.375 ;
        RECT 71.075 177.085 71.475 177.885 ;
        RECT 72.340 177.825 72.895 178.155 ;
        RECT 72.340 177.715 72.790 177.825 ;
        RECT 71.665 177.545 72.790 177.715 ;
        RECT 73.065 177.655 73.345 178.325 ;
        RECT 71.665 177.085 71.945 177.545 ;
        RECT 72.465 176.915 72.790 177.375 ;
        RECT 72.960 177.085 73.345 177.655 ;
        RECT 73.520 178.275 73.775 179.155 ;
        RECT 73.945 178.325 74.250 179.465 ;
        RECT 74.590 179.085 74.920 179.465 ;
        RECT 75.100 178.915 75.270 179.205 ;
        RECT 75.440 179.005 75.690 179.465 ;
        RECT 74.470 178.745 75.270 178.915 ;
        RECT 75.860 178.955 76.730 179.295 ;
        RECT 73.520 177.625 73.730 178.275 ;
        RECT 74.470 178.155 74.640 178.745 ;
        RECT 75.860 178.575 76.030 178.955 ;
        RECT 76.965 178.835 77.135 179.295 ;
        RECT 77.305 179.005 77.675 179.465 ;
        RECT 77.970 178.865 78.140 179.205 ;
        RECT 78.310 179.035 78.640 179.465 ;
        RECT 78.875 178.865 79.045 179.205 ;
        RECT 74.810 178.405 76.030 178.575 ;
        RECT 76.200 178.495 76.660 178.785 ;
        RECT 76.965 178.665 77.525 178.835 ;
        RECT 77.970 178.695 79.045 178.865 ;
        RECT 79.215 178.965 79.895 179.295 ;
        RECT 80.110 178.965 80.360 179.295 ;
        RECT 80.530 179.005 80.780 179.465 ;
        RECT 77.355 178.525 77.525 178.665 ;
        RECT 76.200 178.485 77.165 178.495 ;
        RECT 75.860 178.315 76.030 178.405 ;
        RECT 76.490 178.325 77.165 178.485 ;
        RECT 73.900 178.125 74.640 178.155 ;
        RECT 73.900 177.825 74.815 178.125 ;
        RECT 74.490 177.650 74.815 177.825 ;
        RECT 73.520 177.095 73.775 177.625 ;
        RECT 73.945 176.915 74.250 177.375 ;
        RECT 74.495 177.295 74.815 177.650 ;
        RECT 74.985 177.865 75.525 178.235 ;
        RECT 75.860 178.145 76.265 178.315 ;
        RECT 74.985 177.465 75.225 177.865 ;
        RECT 75.705 177.695 75.925 177.975 ;
        RECT 75.395 177.525 75.925 177.695 ;
        RECT 75.395 177.295 75.565 177.525 ;
        RECT 76.095 177.365 76.265 178.145 ;
        RECT 76.435 177.535 76.785 178.155 ;
        RECT 76.955 177.535 77.165 178.325 ;
        RECT 77.355 178.355 78.855 178.525 ;
        RECT 77.355 177.665 77.525 178.355 ;
        RECT 79.215 178.185 79.385 178.965 ;
        RECT 80.190 178.835 80.360 178.965 ;
        RECT 77.695 178.015 79.385 178.185 ;
        RECT 79.555 178.405 80.020 178.795 ;
        RECT 80.190 178.665 80.585 178.835 ;
        RECT 77.695 177.835 77.865 178.015 ;
        RECT 74.495 177.125 75.565 177.295 ;
        RECT 75.735 176.915 75.925 177.355 ;
        RECT 76.095 177.085 77.045 177.365 ;
        RECT 77.355 177.275 77.615 177.665 ;
        RECT 78.035 177.595 78.825 177.845 ;
        RECT 77.265 177.105 77.615 177.275 ;
        RECT 77.825 176.915 78.155 177.375 ;
        RECT 79.030 177.305 79.200 178.015 ;
        RECT 79.555 177.815 79.725 178.405 ;
        RECT 79.370 177.595 79.725 177.815 ;
        RECT 79.895 177.595 80.245 178.215 ;
        RECT 80.415 177.305 80.585 178.665 ;
        RECT 80.950 178.495 81.275 179.280 ;
        RECT 80.755 177.445 81.215 178.495 ;
        RECT 79.030 177.135 79.885 177.305 ;
        RECT 80.090 177.135 80.585 177.305 ;
        RECT 80.755 176.915 81.085 177.275 ;
        RECT 81.445 177.175 81.615 179.295 ;
        RECT 81.785 178.965 82.115 179.465 ;
        RECT 82.285 178.795 82.540 179.295 ;
        RECT 81.790 178.625 82.540 178.795 ;
        RECT 81.790 177.635 82.020 178.625 ;
        RECT 82.190 177.805 82.540 178.455 ;
        RECT 83.180 178.325 83.515 179.295 ;
        RECT 83.685 178.325 83.855 179.465 ;
        RECT 84.025 179.125 86.055 179.295 ;
        RECT 83.180 177.655 83.350 178.325 ;
        RECT 84.025 178.155 84.195 179.125 ;
        RECT 83.520 177.825 83.775 178.155 ;
        RECT 84.000 177.825 84.195 178.155 ;
        RECT 84.365 178.785 85.490 178.955 ;
        RECT 83.605 177.655 83.775 177.825 ;
        RECT 84.365 177.655 84.535 178.785 ;
        RECT 81.790 177.465 82.540 177.635 ;
        RECT 81.785 176.915 82.115 177.295 ;
        RECT 82.285 177.175 82.540 177.465 ;
        RECT 83.180 177.085 83.435 177.655 ;
        RECT 83.605 177.485 84.535 177.655 ;
        RECT 84.705 178.445 85.715 178.615 ;
        RECT 84.705 177.645 84.875 178.445 ;
        RECT 85.080 177.765 85.355 178.245 ;
        RECT 85.075 177.595 85.355 177.765 ;
        RECT 84.360 177.450 84.535 177.485 ;
        RECT 83.605 176.915 83.935 177.315 ;
        RECT 84.360 177.085 84.890 177.450 ;
        RECT 85.080 177.085 85.355 177.595 ;
        RECT 85.525 177.085 85.715 178.445 ;
        RECT 85.885 178.460 86.055 179.125 ;
        RECT 86.225 178.705 86.395 179.465 ;
        RECT 86.630 178.705 87.145 179.115 ;
        RECT 85.885 178.270 86.635 178.460 ;
        RECT 86.805 177.895 87.145 178.705 ;
        RECT 87.315 178.300 87.605 179.465 ;
        RECT 87.890 178.835 88.175 179.295 ;
        RECT 88.345 179.005 88.615 179.465 ;
        RECT 87.890 178.615 88.845 178.835 ;
        RECT 85.915 177.725 87.145 177.895 ;
        RECT 87.775 177.885 88.465 178.445 ;
        RECT 85.895 176.915 86.405 177.450 ;
        RECT 86.625 177.120 86.870 177.725 ;
        RECT 88.635 177.715 88.845 178.615 ;
        RECT 87.315 176.915 87.605 177.640 ;
        RECT 87.890 177.545 88.845 177.715 ;
        RECT 89.015 178.445 89.415 179.295 ;
        RECT 89.605 178.835 89.885 179.295 ;
        RECT 90.405 179.005 90.730 179.465 ;
        RECT 89.605 178.615 90.730 178.835 ;
        RECT 89.015 177.885 90.110 178.445 ;
        RECT 90.280 178.155 90.730 178.615 ;
        RECT 90.900 178.325 91.285 179.295 ;
        RECT 87.890 177.085 88.175 177.545 ;
        RECT 88.345 176.915 88.615 177.375 ;
        RECT 89.015 177.085 89.415 177.885 ;
        RECT 90.280 177.825 90.835 178.155 ;
        RECT 90.280 177.715 90.730 177.825 ;
        RECT 89.605 177.545 90.730 177.715 ;
        RECT 91.005 177.655 91.285 178.325 ;
        RECT 89.605 177.085 89.885 177.545 ;
        RECT 90.405 176.915 90.730 177.375 ;
        RECT 90.900 177.085 91.285 177.655 ;
        RECT 91.455 178.390 91.725 179.295 ;
        RECT 91.895 178.705 92.225 179.465 ;
        RECT 92.405 178.535 92.575 179.295 ;
        RECT 91.455 177.590 91.625 178.390 ;
        RECT 91.910 178.365 92.575 178.535 ;
        RECT 91.910 178.220 92.080 178.365 ;
        RECT 91.795 177.890 92.080 178.220 ;
        RECT 92.835 178.325 93.175 179.295 ;
        RECT 93.345 178.325 93.515 179.465 ;
        RECT 93.785 178.665 94.035 179.465 ;
        RECT 94.680 178.495 95.010 179.295 ;
        RECT 95.310 178.665 95.640 179.465 ;
        RECT 95.810 178.495 96.140 179.295 ;
        RECT 93.705 178.325 96.140 178.495 ;
        RECT 96.975 178.375 99.565 179.465 ;
        RECT 99.735 178.705 100.250 179.115 ;
        RECT 100.485 178.705 100.655 179.465 ;
        RECT 100.825 179.125 102.855 179.295 ;
        RECT 91.910 177.635 92.080 177.890 ;
        RECT 92.315 177.815 92.645 178.185 ;
        RECT 92.835 177.715 93.010 178.325 ;
        RECT 93.705 178.075 93.875 178.325 ;
        RECT 93.180 177.905 93.875 178.075 ;
        RECT 94.050 177.905 94.470 178.105 ;
        RECT 94.640 177.905 94.970 178.105 ;
        RECT 95.140 177.905 95.470 178.105 ;
        RECT 91.455 177.085 91.715 177.590 ;
        RECT 91.910 177.465 92.575 177.635 ;
        RECT 91.895 176.915 92.225 177.295 ;
        RECT 92.405 177.085 92.575 177.465 ;
        RECT 92.835 177.085 93.175 177.715 ;
        RECT 93.345 176.915 93.595 177.715 ;
        RECT 93.785 177.565 95.010 177.735 ;
        RECT 93.785 177.085 94.115 177.565 ;
        RECT 94.285 176.915 94.510 177.375 ;
        RECT 94.680 177.085 95.010 177.565 ;
        RECT 95.640 177.695 95.810 178.325 ;
        RECT 95.995 177.905 96.345 178.155 ;
        RECT 96.975 177.855 98.185 178.375 ;
        RECT 95.640 177.085 96.140 177.695 ;
        RECT 98.355 177.685 99.565 178.205 ;
        RECT 99.735 177.895 100.075 178.705 ;
        RECT 100.825 178.460 100.995 179.125 ;
        RECT 101.390 178.785 102.515 178.955 ;
        RECT 100.245 178.270 100.995 178.460 ;
        RECT 101.165 178.445 102.175 178.615 ;
        RECT 99.735 177.725 100.965 177.895 ;
        RECT 96.975 176.915 99.565 177.685 ;
        RECT 100.010 177.120 100.255 177.725 ;
        RECT 100.475 176.915 100.985 177.450 ;
        RECT 101.165 177.085 101.355 178.445 ;
        RECT 101.525 178.105 101.800 178.245 ;
        RECT 101.525 177.935 101.805 178.105 ;
        RECT 101.525 177.085 101.800 177.935 ;
        RECT 102.005 177.645 102.175 178.445 ;
        RECT 102.345 177.655 102.515 178.785 ;
        RECT 102.685 178.155 102.855 179.125 ;
        RECT 103.025 178.325 103.195 179.465 ;
        RECT 103.365 178.325 103.700 179.295 ;
        RECT 104.425 178.535 104.595 179.295 ;
        RECT 104.775 178.705 105.105 179.465 ;
        RECT 104.425 178.365 105.090 178.535 ;
        RECT 105.275 178.390 105.545 179.295 ;
        RECT 102.685 177.825 102.880 178.155 ;
        RECT 103.105 177.825 103.360 178.155 ;
        RECT 103.105 177.655 103.275 177.825 ;
        RECT 103.530 177.655 103.700 178.325 ;
        RECT 104.920 178.220 105.090 178.365 ;
        RECT 104.355 177.815 104.685 178.185 ;
        RECT 104.920 177.890 105.205 178.220 ;
        RECT 102.345 177.485 103.275 177.655 ;
        RECT 102.345 177.450 102.520 177.485 ;
        RECT 101.990 177.085 102.520 177.450 ;
        RECT 102.945 176.915 103.275 177.315 ;
        RECT 103.445 177.085 103.700 177.655 ;
        RECT 104.920 177.635 105.090 177.890 ;
        RECT 104.425 177.465 105.090 177.635 ;
        RECT 105.375 177.590 105.545 178.390 ;
        RECT 106.725 178.535 106.895 179.295 ;
        RECT 107.075 178.705 107.405 179.465 ;
        RECT 106.725 178.365 107.390 178.535 ;
        RECT 107.575 178.390 107.845 179.295 ;
        RECT 107.220 178.220 107.390 178.365 ;
        RECT 106.655 177.815 106.985 178.185 ;
        RECT 107.220 177.890 107.505 178.220 ;
        RECT 107.220 177.635 107.390 177.890 ;
        RECT 104.425 177.085 104.595 177.465 ;
        RECT 104.775 176.915 105.105 177.295 ;
        RECT 105.285 177.085 105.545 177.590 ;
        RECT 106.725 177.465 107.390 177.635 ;
        RECT 107.675 177.590 107.845 178.390 ;
        RECT 108.475 178.375 111.985 179.465 ;
        RECT 112.155 178.375 113.365 179.465 ;
        RECT 108.475 177.855 110.165 178.375 ;
        RECT 110.335 177.685 111.985 178.205 ;
        RECT 112.155 177.835 112.675 178.375 ;
        RECT 106.725 177.085 106.895 177.465 ;
        RECT 107.075 176.915 107.405 177.295 ;
        RECT 107.585 177.085 107.845 177.590 ;
        RECT 108.475 176.915 111.985 177.685 ;
        RECT 112.845 177.665 113.365 178.205 ;
        RECT 112.155 176.915 113.365 177.665 ;
        RECT 11.330 176.745 113.450 176.915 ;
        RECT 11.415 175.995 12.625 176.745 ;
        RECT 11.415 175.455 11.935 175.995 ;
        RECT 13.715 175.975 17.225 176.745 ;
        RECT 17.400 176.200 22.745 176.745 ;
        RECT 12.105 175.285 12.625 175.825 ;
        RECT 11.415 174.195 12.625 175.285 ;
        RECT 13.715 175.285 15.405 175.805 ;
        RECT 15.575 175.455 17.225 175.975 ;
        RECT 13.715 174.195 17.225 175.285 ;
        RECT 18.990 174.630 19.340 175.880 ;
        RECT 20.820 175.370 21.160 176.200 ;
        RECT 22.915 176.020 23.205 176.745 ;
        RECT 23.835 176.070 24.095 176.575 ;
        RECT 24.275 176.365 24.605 176.745 ;
        RECT 24.785 176.195 24.955 176.575 ;
        RECT 17.400 174.195 22.745 174.630 ;
        RECT 22.915 174.195 23.205 175.360 ;
        RECT 23.835 175.270 24.005 176.070 ;
        RECT 24.290 176.025 24.955 176.195 ;
        RECT 24.290 175.770 24.460 176.025 ;
        RECT 25.255 175.925 25.485 176.745 ;
        RECT 25.655 175.945 25.985 176.575 ;
        RECT 24.175 175.440 24.460 175.770 ;
        RECT 24.695 175.475 25.025 175.845 ;
        RECT 25.235 175.505 25.565 175.755 ;
        RECT 24.290 175.295 24.460 175.440 ;
        RECT 25.735 175.345 25.985 175.945 ;
        RECT 26.155 175.925 26.365 176.745 ;
        RECT 26.600 176.005 26.855 176.575 ;
        RECT 27.025 176.345 27.355 176.745 ;
        RECT 27.780 176.210 28.310 176.575 ;
        RECT 27.780 176.175 27.955 176.210 ;
        RECT 27.025 176.005 27.955 176.175 ;
        RECT 23.835 174.365 24.105 175.270 ;
        RECT 24.290 175.125 24.955 175.295 ;
        RECT 24.275 174.195 24.605 174.955 ;
        RECT 24.785 174.365 24.955 175.125 ;
        RECT 25.255 174.195 25.485 175.335 ;
        RECT 25.655 174.365 25.985 175.345 ;
        RECT 26.600 175.335 26.770 176.005 ;
        RECT 27.025 175.835 27.195 176.005 ;
        RECT 26.940 175.505 27.195 175.835 ;
        RECT 27.420 175.505 27.615 175.835 ;
        RECT 26.155 174.195 26.365 175.335 ;
        RECT 26.600 174.365 26.935 175.335 ;
        RECT 27.105 174.195 27.275 175.335 ;
        RECT 27.445 174.535 27.615 175.505 ;
        RECT 27.785 174.875 27.955 176.005 ;
        RECT 28.125 175.215 28.295 176.015 ;
        RECT 28.500 175.725 28.775 176.575 ;
        RECT 28.495 175.555 28.775 175.725 ;
        RECT 28.500 175.415 28.775 175.555 ;
        RECT 28.945 175.215 29.135 176.575 ;
        RECT 29.315 176.210 29.825 176.745 ;
        RECT 30.045 175.935 30.290 176.540 ;
        RECT 31.010 175.935 31.255 176.540 ;
        RECT 31.475 176.210 31.985 176.745 ;
        RECT 29.335 175.765 30.565 175.935 ;
        RECT 28.125 175.045 29.135 175.215 ;
        RECT 29.305 175.200 30.055 175.390 ;
        RECT 27.785 174.705 28.910 174.875 ;
        RECT 29.305 174.535 29.475 175.200 ;
        RECT 30.225 174.955 30.565 175.765 ;
        RECT 27.445 174.365 29.475 174.535 ;
        RECT 29.645 174.195 29.815 174.955 ;
        RECT 30.050 174.545 30.565 174.955 ;
        RECT 30.735 175.765 31.965 175.935 ;
        RECT 30.735 174.955 31.075 175.765 ;
        RECT 31.245 175.200 31.995 175.390 ;
        RECT 30.735 174.545 31.250 174.955 ;
        RECT 31.485 174.195 31.655 174.955 ;
        RECT 31.825 174.535 31.995 175.200 ;
        RECT 32.165 175.215 32.355 176.575 ;
        RECT 32.525 176.405 32.800 176.575 ;
        RECT 32.525 176.235 32.805 176.405 ;
        RECT 32.525 175.415 32.800 176.235 ;
        RECT 32.990 176.210 33.520 176.575 ;
        RECT 33.945 176.345 34.275 176.745 ;
        RECT 33.345 176.175 33.520 176.210 ;
        RECT 33.005 175.215 33.175 176.015 ;
        RECT 32.165 175.045 33.175 175.215 ;
        RECT 33.345 176.005 34.275 176.175 ;
        RECT 34.445 176.005 34.700 176.575 ;
        RECT 33.345 174.875 33.515 176.005 ;
        RECT 34.105 175.835 34.275 176.005 ;
        RECT 32.390 174.705 33.515 174.875 ;
        RECT 33.685 175.505 33.880 175.835 ;
        RECT 34.105 175.505 34.360 175.835 ;
        RECT 33.685 174.535 33.855 175.505 ;
        RECT 34.530 175.335 34.700 176.005 ;
        RECT 35.540 175.965 36.040 176.575 ;
        RECT 35.335 175.505 35.685 175.755 ;
        RECT 35.870 175.335 36.040 175.965 ;
        RECT 36.670 176.095 37.000 176.575 ;
        RECT 37.170 176.285 37.395 176.745 ;
        RECT 37.565 176.095 37.895 176.575 ;
        RECT 36.670 175.925 37.895 176.095 ;
        RECT 38.085 175.945 38.335 176.745 ;
        RECT 38.505 175.945 38.845 176.575 ;
        RECT 39.130 176.115 39.415 176.575 ;
        RECT 39.585 176.285 39.855 176.745 ;
        RECT 39.130 175.945 40.085 176.115 ;
        RECT 36.210 175.555 36.540 175.755 ;
        RECT 36.710 175.555 37.040 175.755 ;
        RECT 37.210 175.555 37.630 175.755 ;
        RECT 37.805 175.585 38.500 175.755 ;
        RECT 37.805 175.335 37.975 175.585 ;
        RECT 38.670 175.335 38.845 175.945 ;
        RECT 31.825 174.365 33.855 174.535 ;
        RECT 34.025 174.195 34.195 175.335 ;
        RECT 34.365 174.365 34.700 175.335 ;
        RECT 35.540 175.165 37.975 175.335 ;
        RECT 35.540 174.365 35.870 175.165 ;
        RECT 36.040 174.195 36.370 174.995 ;
        RECT 36.670 174.365 37.000 175.165 ;
        RECT 37.645 174.195 37.895 174.995 ;
        RECT 38.165 174.195 38.335 175.335 ;
        RECT 38.505 174.365 38.845 175.335 ;
        RECT 39.015 175.215 39.705 175.775 ;
        RECT 39.875 175.045 40.085 175.945 ;
        RECT 39.130 174.825 40.085 175.045 ;
        RECT 40.255 175.775 40.655 176.575 ;
        RECT 40.845 176.115 41.125 176.575 ;
        RECT 41.645 176.285 41.970 176.745 ;
        RECT 40.845 175.945 41.970 176.115 ;
        RECT 42.140 176.005 42.525 176.575 ;
        RECT 41.520 175.835 41.970 175.945 ;
        RECT 40.255 175.215 41.350 175.775 ;
        RECT 41.520 175.505 42.075 175.835 ;
        RECT 39.130 174.365 39.415 174.825 ;
        RECT 39.585 174.195 39.855 174.655 ;
        RECT 40.255 174.365 40.655 175.215 ;
        RECT 41.520 175.045 41.970 175.505 ;
        RECT 42.245 175.335 42.525 176.005 ;
        RECT 42.970 175.935 43.215 176.540 ;
        RECT 43.435 176.210 43.945 176.745 ;
        RECT 40.845 174.825 41.970 175.045 ;
        RECT 40.845 174.365 41.125 174.825 ;
        RECT 41.645 174.195 41.970 174.655 ;
        RECT 42.140 174.365 42.525 175.335 ;
        RECT 42.695 175.765 43.925 175.935 ;
        RECT 42.695 174.955 43.035 175.765 ;
        RECT 43.205 175.200 43.955 175.390 ;
        RECT 42.695 174.545 43.210 174.955 ;
        RECT 43.445 174.195 43.615 174.955 ;
        RECT 43.785 174.535 43.955 175.200 ;
        RECT 44.125 175.215 44.315 176.575 ;
        RECT 44.485 175.725 44.760 176.575 ;
        RECT 44.950 176.210 45.480 176.575 ;
        RECT 45.905 176.345 46.235 176.745 ;
        RECT 45.305 176.175 45.480 176.210 ;
        RECT 44.485 175.555 44.765 175.725 ;
        RECT 44.485 175.415 44.760 175.555 ;
        RECT 44.965 175.215 45.135 176.015 ;
        RECT 44.125 175.045 45.135 175.215 ;
        RECT 45.305 176.005 46.235 176.175 ;
        RECT 46.405 176.005 46.660 176.575 ;
        RECT 45.305 174.875 45.475 176.005 ;
        RECT 46.065 175.835 46.235 176.005 ;
        RECT 44.350 174.705 45.475 174.875 ;
        RECT 45.645 175.505 45.840 175.835 ;
        RECT 46.065 175.505 46.320 175.835 ;
        RECT 45.645 174.535 45.815 175.505 ;
        RECT 46.490 175.335 46.660 176.005 ;
        RECT 47.335 175.925 47.565 176.745 ;
        RECT 47.735 175.945 48.065 176.575 ;
        RECT 47.315 175.505 47.645 175.755 ;
        RECT 47.815 175.345 48.065 175.945 ;
        RECT 48.235 175.925 48.445 176.745 ;
        RECT 48.675 176.020 48.965 176.745 ;
        RECT 49.140 176.035 49.395 176.565 ;
        RECT 49.565 176.285 49.870 176.745 ;
        RECT 50.115 176.365 51.185 176.535 ;
        RECT 49.140 175.385 49.350 176.035 ;
        RECT 50.115 176.010 50.435 176.365 ;
        RECT 50.110 175.835 50.435 176.010 ;
        RECT 49.520 175.535 50.435 175.835 ;
        RECT 50.605 175.795 50.845 176.195 ;
        RECT 51.015 176.135 51.185 176.365 ;
        RECT 51.355 176.305 51.545 176.745 ;
        RECT 51.715 176.295 52.665 176.575 ;
        RECT 52.885 176.385 53.235 176.555 ;
        RECT 51.015 175.965 51.545 176.135 ;
        RECT 49.520 175.505 50.260 175.535 ;
        RECT 43.785 174.365 45.815 174.535 ;
        RECT 45.985 174.195 46.155 175.335 ;
        RECT 46.325 174.365 46.660 175.335 ;
        RECT 47.335 174.195 47.565 175.335 ;
        RECT 47.735 174.365 48.065 175.345 ;
        RECT 48.235 174.195 48.445 175.335 ;
        RECT 48.675 174.195 48.965 175.360 ;
        RECT 49.140 174.505 49.395 175.385 ;
        RECT 49.565 174.195 49.870 175.335 ;
        RECT 50.090 174.915 50.260 175.505 ;
        RECT 50.605 175.425 51.145 175.795 ;
        RECT 51.325 175.685 51.545 175.965 ;
        RECT 51.715 175.515 51.885 176.295 ;
        RECT 51.480 175.345 51.885 175.515 ;
        RECT 52.055 175.505 52.405 176.125 ;
        RECT 51.480 175.255 51.650 175.345 ;
        RECT 52.575 175.335 52.785 176.125 ;
        RECT 50.430 175.085 51.650 175.255 ;
        RECT 52.110 175.175 52.785 175.335 ;
        RECT 50.090 174.745 50.890 174.915 ;
        RECT 50.210 174.195 50.540 174.575 ;
        RECT 50.720 174.455 50.890 174.745 ;
        RECT 51.480 174.705 51.650 175.085 ;
        RECT 51.820 175.165 52.785 175.175 ;
        RECT 52.975 175.995 53.235 176.385 ;
        RECT 53.445 176.285 53.775 176.745 ;
        RECT 54.650 176.355 55.505 176.525 ;
        RECT 55.710 176.355 56.205 176.525 ;
        RECT 56.375 176.385 56.705 176.745 ;
        RECT 52.975 175.305 53.145 175.995 ;
        RECT 53.315 175.645 53.485 175.825 ;
        RECT 53.655 175.815 54.445 176.065 ;
        RECT 54.650 175.645 54.820 176.355 ;
        RECT 54.990 175.845 55.345 176.065 ;
        RECT 53.315 175.475 55.005 175.645 ;
        RECT 51.820 174.875 52.280 175.165 ;
        RECT 52.975 175.135 54.475 175.305 ;
        RECT 52.975 174.995 53.145 175.135 ;
        RECT 52.585 174.825 53.145 174.995 ;
        RECT 51.060 174.195 51.310 174.655 ;
        RECT 51.480 174.365 52.350 174.705 ;
        RECT 52.585 174.365 52.755 174.825 ;
        RECT 53.590 174.795 54.665 174.965 ;
        RECT 52.925 174.195 53.295 174.655 ;
        RECT 53.590 174.455 53.760 174.795 ;
        RECT 53.930 174.195 54.260 174.625 ;
        RECT 54.495 174.455 54.665 174.795 ;
        RECT 54.835 174.695 55.005 175.475 ;
        RECT 55.175 175.255 55.345 175.845 ;
        RECT 55.515 175.445 55.865 176.065 ;
        RECT 55.175 174.865 55.640 175.255 ;
        RECT 56.035 174.995 56.205 176.355 ;
        RECT 56.375 175.165 56.835 176.215 ;
        RECT 55.810 174.825 56.205 174.995 ;
        RECT 55.810 174.695 55.980 174.825 ;
        RECT 54.835 174.365 55.515 174.695 ;
        RECT 55.730 174.365 55.980 174.695 ;
        RECT 56.150 174.195 56.400 174.655 ;
        RECT 56.570 174.380 56.895 175.165 ;
        RECT 57.065 174.365 57.235 176.485 ;
        RECT 57.405 176.365 57.735 176.745 ;
        RECT 57.905 176.195 58.160 176.485 ;
        RECT 57.410 176.025 58.160 176.195 ;
        RECT 58.885 176.195 59.055 176.575 ;
        RECT 59.270 176.365 59.600 176.745 ;
        RECT 58.885 176.025 59.600 176.195 ;
        RECT 57.410 175.035 57.640 176.025 ;
        RECT 57.810 175.205 58.160 175.855 ;
        RECT 58.795 175.475 59.150 175.845 ;
        RECT 59.430 175.835 59.600 176.025 ;
        RECT 59.770 176.000 60.025 176.575 ;
        RECT 59.430 175.505 59.685 175.835 ;
        RECT 59.430 175.295 59.600 175.505 ;
        RECT 58.885 175.125 59.600 175.295 ;
        RECT 59.855 175.270 60.025 176.000 ;
        RECT 60.200 175.905 60.460 176.745 ;
        RECT 60.640 175.905 60.900 176.745 ;
        RECT 61.075 176.000 61.330 176.575 ;
        RECT 61.500 176.365 61.830 176.745 ;
        RECT 62.045 176.195 62.215 176.575 ;
        RECT 61.500 176.025 62.215 176.195 ;
        RECT 62.565 176.195 62.735 176.575 ;
        RECT 62.950 176.365 63.280 176.745 ;
        RECT 62.565 176.025 63.280 176.195 ;
        RECT 57.410 174.865 58.160 175.035 ;
        RECT 57.405 174.195 57.735 174.695 ;
        RECT 57.905 174.365 58.160 174.865 ;
        RECT 58.885 174.365 59.055 175.125 ;
        RECT 59.270 174.195 59.600 174.955 ;
        RECT 59.770 174.365 60.025 175.270 ;
        RECT 60.200 174.195 60.460 175.345 ;
        RECT 60.640 174.195 60.900 175.345 ;
        RECT 61.075 175.270 61.245 176.000 ;
        RECT 61.500 175.835 61.670 176.025 ;
        RECT 61.415 175.505 61.670 175.835 ;
        RECT 61.500 175.295 61.670 175.505 ;
        RECT 61.950 175.475 62.305 175.845 ;
        RECT 62.475 175.475 62.830 175.845 ;
        RECT 63.110 175.835 63.280 176.025 ;
        RECT 63.450 176.000 63.705 176.575 ;
        RECT 63.110 175.505 63.365 175.835 ;
        RECT 63.110 175.295 63.280 175.505 ;
        RECT 61.075 174.365 61.330 175.270 ;
        RECT 61.500 175.125 62.215 175.295 ;
        RECT 61.500 174.195 61.830 174.955 ;
        RECT 62.045 174.365 62.215 175.125 ;
        RECT 62.565 175.125 63.280 175.295 ;
        RECT 63.535 175.270 63.705 176.000 ;
        RECT 63.880 175.905 64.140 176.745 ;
        RECT 64.325 176.215 64.655 176.575 ;
        RECT 64.825 176.385 65.155 176.745 ;
        RECT 65.355 176.215 65.685 176.575 ;
        RECT 64.325 176.005 65.685 176.215 ;
        RECT 66.195 175.985 66.905 176.575 ;
        RECT 67.165 176.195 67.335 176.575 ;
        RECT 67.550 176.365 67.880 176.745 ;
        RECT 67.165 176.025 67.880 176.195 ;
        RECT 66.675 175.895 66.905 175.985 ;
        RECT 64.315 175.505 64.625 175.835 ;
        RECT 64.835 175.505 65.210 175.835 ;
        RECT 65.530 175.505 66.025 175.835 ;
        RECT 62.565 174.365 62.735 175.125 ;
        RECT 62.950 174.195 63.280 174.955 ;
        RECT 63.450 174.365 63.705 175.270 ;
        RECT 63.880 174.195 64.140 175.345 ;
        RECT 64.325 174.195 64.655 175.255 ;
        RECT 64.835 174.580 65.005 175.505 ;
        RECT 65.175 175.015 65.505 175.235 ;
        RECT 65.700 175.215 66.025 175.505 ;
        RECT 66.200 175.215 66.530 175.755 ;
        RECT 66.700 175.015 66.905 175.895 ;
        RECT 67.075 175.475 67.430 175.845 ;
        RECT 67.710 175.835 67.880 176.025 ;
        RECT 68.050 176.000 68.305 176.575 ;
        RECT 67.710 175.505 67.965 175.835 ;
        RECT 67.710 175.295 67.880 175.505 ;
        RECT 65.175 174.785 66.905 175.015 ;
        RECT 65.175 174.385 65.505 174.785 ;
        RECT 65.675 174.195 66.005 174.555 ;
        RECT 66.205 174.365 66.905 174.785 ;
        RECT 67.165 175.125 67.880 175.295 ;
        RECT 68.135 175.270 68.305 176.000 ;
        RECT 68.480 175.905 68.740 176.745 ;
        RECT 68.915 175.995 70.125 176.745 ;
        RECT 67.165 174.365 67.335 175.125 ;
        RECT 67.550 174.195 67.880 174.955 ;
        RECT 68.050 174.365 68.305 175.270 ;
        RECT 68.480 174.195 68.740 175.345 ;
        RECT 68.915 175.285 69.435 175.825 ;
        RECT 69.605 175.455 70.125 175.995 ;
        RECT 70.295 175.945 70.635 176.575 ;
        RECT 70.805 175.945 71.055 176.745 ;
        RECT 71.245 176.095 71.575 176.575 ;
        RECT 71.745 176.285 71.970 176.745 ;
        RECT 72.140 176.095 72.470 176.575 ;
        RECT 70.295 175.335 70.470 175.945 ;
        RECT 71.245 175.925 72.470 176.095 ;
        RECT 73.100 175.965 73.600 176.575 ;
        RECT 74.435 176.020 74.725 176.745 ;
        RECT 75.930 176.115 76.215 176.575 ;
        RECT 76.385 176.285 76.655 176.745 ;
        RECT 70.640 175.585 71.335 175.755 ;
        RECT 71.165 175.335 71.335 175.585 ;
        RECT 71.510 175.555 71.930 175.755 ;
        RECT 72.100 175.555 72.430 175.755 ;
        RECT 72.600 175.555 72.930 175.755 ;
        RECT 73.100 175.335 73.270 175.965 ;
        RECT 75.930 175.945 76.885 176.115 ;
        RECT 73.455 175.505 73.805 175.755 ;
        RECT 68.915 174.195 70.125 175.285 ;
        RECT 70.295 174.365 70.635 175.335 ;
        RECT 70.805 174.195 70.975 175.335 ;
        RECT 71.165 175.165 73.600 175.335 ;
        RECT 71.245 174.195 71.495 174.995 ;
        RECT 72.140 174.365 72.470 175.165 ;
        RECT 72.770 174.195 73.100 174.995 ;
        RECT 73.270 174.365 73.600 175.165 ;
        RECT 74.435 174.195 74.725 175.360 ;
        RECT 75.815 175.215 76.505 175.775 ;
        RECT 76.675 175.045 76.885 175.945 ;
        RECT 75.930 174.825 76.885 175.045 ;
        RECT 77.055 175.775 77.455 176.575 ;
        RECT 77.645 176.115 77.925 176.575 ;
        RECT 78.445 176.285 78.770 176.745 ;
        RECT 77.645 175.945 78.770 176.115 ;
        RECT 78.940 176.005 79.325 176.575 ;
        RECT 79.585 176.195 79.755 176.575 ;
        RECT 79.935 176.365 80.265 176.745 ;
        RECT 79.585 176.025 80.250 176.195 ;
        RECT 80.445 176.070 80.705 176.575 ;
        RECT 78.320 175.835 78.770 175.945 ;
        RECT 77.055 175.215 78.150 175.775 ;
        RECT 78.320 175.505 78.875 175.835 ;
        RECT 75.930 174.365 76.215 174.825 ;
        RECT 76.385 174.195 76.655 174.655 ;
        RECT 77.055 174.365 77.455 175.215 ;
        RECT 78.320 175.045 78.770 175.505 ;
        RECT 79.045 175.335 79.325 176.005 ;
        RECT 79.515 175.475 79.845 175.845 ;
        RECT 80.080 175.770 80.250 176.025 ;
        RECT 77.645 174.825 78.770 175.045 ;
        RECT 77.645 174.365 77.925 174.825 ;
        RECT 78.445 174.195 78.770 174.655 ;
        RECT 78.940 174.365 79.325 175.335 ;
        RECT 80.080 175.440 80.365 175.770 ;
        RECT 80.080 175.295 80.250 175.440 ;
        RECT 79.585 175.125 80.250 175.295 ;
        RECT 80.535 175.270 80.705 176.070 ;
        RECT 80.990 176.115 81.275 176.575 ;
        RECT 81.445 176.285 81.715 176.745 ;
        RECT 80.990 175.945 81.945 176.115 ;
        RECT 79.585 174.365 79.755 175.125 ;
        RECT 79.935 174.195 80.265 174.955 ;
        RECT 80.435 174.365 80.705 175.270 ;
        RECT 80.875 175.215 81.565 175.775 ;
        RECT 81.735 175.045 81.945 175.945 ;
        RECT 80.990 174.825 81.945 175.045 ;
        RECT 82.115 175.775 82.515 176.575 ;
        RECT 82.705 176.115 82.985 176.575 ;
        RECT 83.505 176.285 83.830 176.745 ;
        RECT 82.705 175.945 83.830 176.115 ;
        RECT 84.000 176.005 84.385 176.575 ;
        RECT 83.380 175.835 83.830 175.945 ;
        RECT 82.115 175.215 83.210 175.775 ;
        RECT 83.380 175.505 83.935 175.835 ;
        RECT 80.990 174.365 81.275 174.825 ;
        RECT 81.445 174.195 81.715 174.655 ;
        RECT 82.115 174.365 82.515 175.215 ;
        RECT 83.380 175.045 83.830 175.505 ;
        RECT 84.105 175.335 84.385 176.005 ;
        RECT 84.670 176.115 84.955 176.575 ;
        RECT 85.125 176.285 85.395 176.745 ;
        RECT 84.670 175.945 85.625 176.115 ;
        RECT 82.705 174.825 83.830 175.045 ;
        RECT 82.705 174.365 82.985 174.825 ;
        RECT 83.505 174.195 83.830 174.655 ;
        RECT 84.000 174.365 84.385 175.335 ;
        RECT 84.555 175.215 85.245 175.775 ;
        RECT 85.415 175.045 85.625 175.945 ;
        RECT 84.670 174.825 85.625 175.045 ;
        RECT 85.795 175.775 86.195 176.575 ;
        RECT 86.385 176.115 86.665 176.575 ;
        RECT 87.185 176.285 87.510 176.745 ;
        RECT 86.385 175.945 87.510 176.115 ;
        RECT 87.680 176.005 88.065 176.575 ;
        RECT 87.060 175.835 87.510 175.945 ;
        RECT 85.795 175.215 86.890 175.775 ;
        RECT 87.060 175.505 87.615 175.835 ;
        RECT 84.670 174.365 84.955 174.825 ;
        RECT 85.125 174.195 85.395 174.655 ;
        RECT 85.795 174.365 86.195 175.215 ;
        RECT 87.060 175.045 87.510 175.505 ;
        RECT 87.785 175.335 88.065 176.005 ;
        RECT 86.385 174.825 87.510 175.045 ;
        RECT 86.385 174.365 86.665 174.825 ;
        RECT 87.185 174.195 87.510 174.655 ;
        RECT 87.680 174.365 88.065 175.335 ;
        RECT 88.235 175.945 88.575 176.575 ;
        RECT 88.745 175.945 88.995 176.745 ;
        RECT 89.185 176.095 89.515 176.575 ;
        RECT 89.685 176.285 89.910 176.745 ;
        RECT 90.080 176.095 90.410 176.575 ;
        RECT 88.235 175.335 88.410 175.945 ;
        RECT 89.185 175.925 90.410 176.095 ;
        RECT 91.040 175.965 91.540 176.575 ;
        RECT 88.580 175.585 89.275 175.755 ;
        RECT 89.105 175.335 89.275 175.585 ;
        RECT 89.450 175.555 89.870 175.755 ;
        RECT 90.040 175.555 90.370 175.755 ;
        RECT 90.540 175.555 90.870 175.755 ;
        RECT 91.040 175.335 91.210 175.965 ;
        RECT 92.375 175.945 92.715 176.575 ;
        RECT 92.885 175.945 93.135 176.745 ;
        RECT 93.325 176.095 93.655 176.575 ;
        RECT 93.825 176.285 94.050 176.745 ;
        RECT 94.220 176.095 94.550 176.575 ;
        RECT 91.395 175.505 91.745 175.755 ;
        RECT 92.375 175.335 92.550 175.945 ;
        RECT 93.325 175.925 94.550 176.095 ;
        RECT 95.180 175.965 95.680 176.575 ;
        RECT 96.260 175.965 96.760 176.575 ;
        RECT 92.720 175.585 93.415 175.755 ;
        RECT 93.245 175.335 93.415 175.585 ;
        RECT 93.590 175.555 94.010 175.755 ;
        RECT 94.180 175.555 94.510 175.755 ;
        RECT 94.680 175.555 95.010 175.755 ;
        RECT 95.180 175.335 95.350 175.965 ;
        RECT 95.535 175.505 95.885 175.755 ;
        RECT 96.055 175.505 96.405 175.755 ;
        RECT 96.590 175.335 96.760 175.965 ;
        RECT 97.390 176.095 97.720 176.575 ;
        RECT 97.890 176.285 98.115 176.745 ;
        RECT 98.285 176.095 98.615 176.575 ;
        RECT 97.390 175.925 98.615 176.095 ;
        RECT 98.805 175.945 99.055 176.745 ;
        RECT 99.225 175.945 99.565 176.575 ;
        RECT 100.195 176.020 100.485 176.745 ;
        RECT 101.580 176.200 106.925 176.745 ;
        RECT 96.930 175.555 97.260 175.755 ;
        RECT 97.430 175.555 97.760 175.755 ;
        RECT 97.930 175.555 98.350 175.755 ;
        RECT 98.525 175.585 99.220 175.755 ;
        RECT 98.525 175.335 98.695 175.585 ;
        RECT 99.390 175.335 99.565 175.945 ;
        RECT 88.235 174.365 88.575 175.335 ;
        RECT 88.745 174.195 88.915 175.335 ;
        RECT 89.105 175.165 91.540 175.335 ;
        RECT 89.185 174.195 89.435 174.995 ;
        RECT 90.080 174.365 90.410 175.165 ;
        RECT 90.710 174.195 91.040 174.995 ;
        RECT 91.210 174.365 91.540 175.165 ;
        RECT 92.375 174.365 92.715 175.335 ;
        RECT 92.885 174.195 93.055 175.335 ;
        RECT 93.245 175.165 95.680 175.335 ;
        RECT 93.325 174.195 93.575 174.995 ;
        RECT 94.220 174.365 94.550 175.165 ;
        RECT 94.850 174.195 95.180 174.995 ;
        RECT 95.350 174.365 95.680 175.165 ;
        RECT 96.260 175.165 98.695 175.335 ;
        RECT 96.260 174.365 96.590 175.165 ;
        RECT 96.760 174.195 97.090 174.995 ;
        RECT 97.390 174.365 97.720 175.165 ;
        RECT 98.365 174.195 98.615 174.995 ;
        RECT 98.885 174.195 99.055 175.335 ;
        RECT 99.225 174.365 99.565 175.335 ;
        RECT 100.195 174.195 100.485 175.360 ;
        RECT 103.170 174.630 103.520 175.880 ;
        RECT 105.000 175.370 105.340 176.200 ;
        RECT 107.185 176.195 107.355 176.575 ;
        RECT 107.535 176.365 107.865 176.745 ;
        RECT 107.185 176.025 107.850 176.195 ;
        RECT 108.045 176.070 108.305 176.575 ;
        RECT 107.115 175.475 107.445 175.845 ;
        RECT 107.680 175.770 107.850 176.025 ;
        RECT 107.680 175.440 107.965 175.770 ;
        RECT 107.680 175.295 107.850 175.440 ;
        RECT 107.185 175.125 107.850 175.295 ;
        RECT 108.135 175.270 108.305 176.070 ;
        RECT 108.475 175.975 111.985 176.745 ;
        RECT 112.155 175.995 113.365 176.745 ;
        RECT 101.580 174.195 106.925 174.630 ;
        RECT 107.185 174.365 107.355 175.125 ;
        RECT 107.535 174.195 107.865 174.955 ;
        RECT 108.035 174.365 108.305 175.270 ;
        RECT 108.475 175.285 110.165 175.805 ;
        RECT 110.335 175.455 111.985 175.975 ;
        RECT 112.155 175.285 112.675 175.825 ;
        RECT 112.845 175.455 113.365 175.995 ;
        RECT 108.475 174.195 111.985 175.285 ;
        RECT 112.155 174.195 113.365 175.285 ;
        RECT 11.330 174.025 113.450 174.195 ;
        RECT 11.415 172.935 12.625 174.025 ;
        RECT 11.415 172.225 11.935 172.765 ;
        RECT 12.105 172.395 12.625 172.935 ;
        RECT 13.255 172.935 16.765 174.025 ;
        RECT 16.940 173.590 22.285 174.025 ;
        RECT 13.255 172.415 14.945 172.935 ;
        RECT 15.115 172.245 16.765 172.765 ;
        RECT 18.530 172.340 18.880 173.590 ;
        RECT 22.570 173.395 22.855 173.855 ;
        RECT 23.025 173.565 23.295 174.025 ;
        RECT 22.570 173.175 23.525 173.395 ;
        RECT 11.415 171.475 12.625 172.225 ;
        RECT 13.255 171.475 16.765 172.245 ;
        RECT 20.360 172.020 20.700 172.850 ;
        RECT 22.455 172.445 23.145 173.005 ;
        RECT 23.315 172.275 23.525 173.175 ;
        RECT 22.570 172.105 23.525 172.275 ;
        RECT 23.695 173.005 24.095 173.855 ;
        RECT 24.285 173.395 24.565 173.855 ;
        RECT 25.085 173.565 25.410 174.025 ;
        RECT 24.285 173.175 25.410 173.395 ;
        RECT 23.695 172.445 24.790 173.005 ;
        RECT 24.960 172.715 25.410 173.175 ;
        RECT 25.580 172.885 25.965 173.855 ;
        RECT 16.940 171.475 22.285 172.020 ;
        RECT 22.570 171.645 22.855 172.105 ;
        RECT 23.025 171.475 23.295 171.935 ;
        RECT 23.695 171.645 24.095 172.445 ;
        RECT 24.960 172.385 25.515 172.715 ;
        RECT 24.960 172.275 25.410 172.385 ;
        RECT 24.285 172.105 25.410 172.275 ;
        RECT 25.685 172.215 25.965 172.885 ;
        RECT 24.285 171.645 24.565 172.105 ;
        RECT 25.085 171.475 25.410 171.935 ;
        RECT 25.580 171.645 25.965 172.215 ;
        RECT 26.140 172.835 26.395 173.715 ;
        RECT 26.565 172.885 26.870 174.025 ;
        RECT 27.210 173.645 27.540 174.025 ;
        RECT 27.720 173.475 27.890 173.765 ;
        RECT 28.060 173.565 28.310 174.025 ;
        RECT 27.090 173.305 27.890 173.475 ;
        RECT 28.480 173.515 29.350 173.855 ;
        RECT 26.140 172.185 26.350 172.835 ;
        RECT 27.090 172.715 27.260 173.305 ;
        RECT 28.480 173.135 28.650 173.515 ;
        RECT 29.585 173.395 29.755 173.855 ;
        RECT 29.925 173.565 30.295 174.025 ;
        RECT 30.590 173.425 30.760 173.765 ;
        RECT 30.930 173.595 31.260 174.025 ;
        RECT 31.495 173.425 31.665 173.765 ;
        RECT 27.430 172.965 28.650 173.135 ;
        RECT 28.820 173.055 29.280 173.345 ;
        RECT 29.585 173.225 30.145 173.395 ;
        RECT 30.590 173.255 31.665 173.425 ;
        RECT 31.835 173.525 32.515 173.855 ;
        RECT 32.730 173.525 32.980 173.855 ;
        RECT 33.150 173.565 33.400 174.025 ;
        RECT 29.975 173.085 30.145 173.225 ;
        RECT 28.820 173.045 29.785 173.055 ;
        RECT 28.480 172.875 28.650 172.965 ;
        RECT 29.110 172.885 29.785 173.045 ;
        RECT 26.520 172.685 27.260 172.715 ;
        RECT 26.520 172.385 27.435 172.685 ;
        RECT 27.110 172.210 27.435 172.385 ;
        RECT 26.140 171.655 26.395 172.185 ;
        RECT 26.565 171.475 26.870 171.935 ;
        RECT 27.115 171.855 27.435 172.210 ;
        RECT 27.605 172.425 28.145 172.795 ;
        RECT 28.480 172.705 28.885 172.875 ;
        RECT 27.605 172.025 27.845 172.425 ;
        RECT 28.325 172.255 28.545 172.535 ;
        RECT 28.015 172.085 28.545 172.255 ;
        RECT 28.015 171.855 28.185 172.085 ;
        RECT 28.715 171.925 28.885 172.705 ;
        RECT 29.055 172.095 29.405 172.715 ;
        RECT 29.575 172.095 29.785 172.885 ;
        RECT 29.975 172.915 31.475 173.085 ;
        RECT 29.975 172.225 30.145 172.915 ;
        RECT 31.835 172.745 32.005 173.525 ;
        RECT 32.810 173.395 32.980 173.525 ;
        RECT 30.315 172.575 32.005 172.745 ;
        RECT 32.175 172.965 32.640 173.355 ;
        RECT 32.810 173.225 33.205 173.395 ;
        RECT 30.315 172.395 30.485 172.575 ;
        RECT 27.115 171.685 28.185 171.855 ;
        RECT 28.355 171.475 28.545 171.915 ;
        RECT 28.715 171.645 29.665 171.925 ;
        RECT 29.975 171.835 30.235 172.225 ;
        RECT 30.655 172.155 31.445 172.405 ;
        RECT 29.885 171.665 30.235 171.835 ;
        RECT 30.445 171.475 30.775 171.935 ;
        RECT 31.650 171.865 31.820 172.575 ;
        RECT 32.175 172.375 32.345 172.965 ;
        RECT 31.990 172.155 32.345 172.375 ;
        RECT 32.515 172.155 32.865 172.775 ;
        RECT 33.035 171.865 33.205 173.225 ;
        RECT 33.570 173.055 33.895 173.840 ;
        RECT 33.375 172.005 33.835 173.055 ;
        RECT 31.650 171.695 32.505 171.865 ;
        RECT 32.710 171.695 33.205 171.865 ;
        RECT 33.375 171.475 33.705 171.835 ;
        RECT 34.065 171.735 34.235 173.855 ;
        RECT 34.405 173.525 34.735 174.025 ;
        RECT 34.905 173.355 35.160 173.855 ;
        RECT 34.410 173.185 35.160 173.355 ;
        RECT 34.410 172.195 34.640 173.185 ;
        RECT 34.810 172.365 35.160 173.015 ;
        RECT 35.795 172.860 36.085 174.025 ;
        RECT 36.255 172.950 36.525 173.855 ;
        RECT 36.695 173.265 37.025 174.025 ;
        RECT 37.205 173.095 37.375 173.855 ;
        RECT 34.410 172.025 35.160 172.195 ;
        RECT 34.405 171.475 34.735 171.855 ;
        RECT 34.905 171.735 35.160 172.025 ;
        RECT 35.795 171.475 36.085 172.200 ;
        RECT 36.255 172.150 36.425 172.950 ;
        RECT 36.710 172.925 37.375 173.095 ;
        RECT 38.760 173.055 39.090 173.855 ;
        RECT 39.260 173.225 39.590 174.025 ;
        RECT 39.890 173.055 40.220 173.855 ;
        RECT 40.865 173.225 41.115 174.025 ;
        RECT 36.710 172.780 36.880 172.925 ;
        RECT 38.760 172.885 41.195 173.055 ;
        RECT 41.385 172.885 41.555 174.025 ;
        RECT 41.725 172.885 42.065 173.855 ;
        RECT 36.595 172.450 36.880 172.780 ;
        RECT 36.710 172.195 36.880 172.450 ;
        RECT 37.115 172.375 37.445 172.745 ;
        RECT 38.555 172.465 38.905 172.715 ;
        RECT 39.090 172.255 39.260 172.885 ;
        RECT 39.430 172.465 39.760 172.665 ;
        RECT 39.930 172.465 40.260 172.665 ;
        RECT 40.430 172.465 40.850 172.665 ;
        RECT 41.025 172.635 41.195 172.885 ;
        RECT 41.025 172.465 41.720 172.635 ;
        RECT 36.255 171.645 36.515 172.150 ;
        RECT 36.710 172.025 37.375 172.195 ;
        RECT 36.695 171.475 37.025 171.855 ;
        RECT 37.205 171.645 37.375 172.025 ;
        RECT 38.760 171.645 39.260 172.255 ;
        RECT 39.890 172.125 41.115 172.295 ;
        RECT 41.890 172.275 42.065 172.885 ;
        RECT 42.235 173.265 42.750 173.675 ;
        RECT 42.985 173.265 43.155 174.025 ;
        RECT 43.325 173.685 45.355 173.855 ;
        RECT 42.235 172.455 42.575 173.265 ;
        RECT 43.325 173.020 43.495 173.685 ;
        RECT 43.890 173.345 45.015 173.515 ;
        RECT 42.745 172.830 43.495 173.020 ;
        RECT 43.665 173.005 44.675 173.175 ;
        RECT 42.235 172.285 43.465 172.455 ;
        RECT 39.890 171.645 40.220 172.125 ;
        RECT 40.390 171.475 40.615 171.935 ;
        RECT 40.785 171.645 41.115 172.125 ;
        RECT 41.305 171.475 41.555 172.275 ;
        RECT 41.725 171.645 42.065 172.275 ;
        RECT 42.510 171.680 42.755 172.285 ;
        RECT 42.975 171.475 43.485 172.010 ;
        RECT 43.665 171.645 43.855 173.005 ;
        RECT 44.025 171.985 44.300 172.805 ;
        RECT 44.505 172.205 44.675 173.005 ;
        RECT 44.845 172.215 45.015 173.345 ;
        RECT 45.185 172.715 45.355 173.685 ;
        RECT 45.525 172.885 45.695 174.025 ;
        RECT 45.865 172.885 46.200 173.855 ;
        RECT 45.185 172.385 45.380 172.715 ;
        RECT 45.605 172.385 45.860 172.715 ;
        RECT 45.605 172.215 45.775 172.385 ;
        RECT 46.030 172.215 46.200 172.885 ;
        RECT 46.375 173.265 46.890 173.675 ;
        RECT 47.125 173.265 47.295 174.025 ;
        RECT 47.465 173.685 49.495 173.855 ;
        RECT 46.375 172.455 46.715 173.265 ;
        RECT 47.465 173.020 47.635 173.685 ;
        RECT 48.030 173.345 49.155 173.515 ;
        RECT 46.885 172.830 47.635 173.020 ;
        RECT 47.805 173.005 48.815 173.175 ;
        RECT 46.375 172.285 47.605 172.455 ;
        RECT 44.845 172.045 45.775 172.215 ;
        RECT 44.845 172.010 45.020 172.045 ;
        RECT 44.025 171.815 44.305 171.985 ;
        RECT 44.025 171.645 44.300 171.815 ;
        RECT 44.490 171.645 45.020 172.010 ;
        RECT 45.445 171.475 45.775 171.875 ;
        RECT 45.945 171.645 46.200 172.215 ;
        RECT 46.650 171.680 46.895 172.285 ;
        RECT 47.115 171.475 47.625 172.010 ;
        RECT 47.805 171.645 47.995 173.005 ;
        RECT 48.165 172.325 48.440 172.805 ;
        RECT 48.165 172.155 48.445 172.325 ;
        RECT 48.645 172.205 48.815 173.005 ;
        RECT 48.985 172.215 49.155 173.345 ;
        RECT 49.325 172.715 49.495 173.685 ;
        RECT 49.665 172.885 49.835 174.025 ;
        RECT 50.005 172.885 50.340 173.855 ;
        RECT 49.325 172.385 49.520 172.715 ;
        RECT 49.745 172.385 50.000 172.715 ;
        RECT 49.745 172.215 49.915 172.385 ;
        RECT 50.170 172.215 50.340 172.885 ;
        RECT 48.165 171.645 48.440 172.155 ;
        RECT 48.985 172.045 49.915 172.215 ;
        RECT 48.985 172.010 49.160 172.045 ;
        RECT 48.630 171.645 49.160 172.010 ;
        RECT 49.585 171.475 49.915 171.875 ;
        RECT 50.085 171.645 50.340 172.215 ;
        RECT 50.520 172.835 50.775 173.715 ;
        RECT 50.945 172.885 51.250 174.025 ;
        RECT 51.590 173.645 51.920 174.025 ;
        RECT 52.100 173.475 52.270 173.765 ;
        RECT 52.440 173.565 52.690 174.025 ;
        RECT 51.470 173.305 52.270 173.475 ;
        RECT 52.860 173.515 53.730 173.855 ;
        RECT 50.520 172.185 50.730 172.835 ;
        RECT 51.470 172.715 51.640 173.305 ;
        RECT 52.860 173.135 53.030 173.515 ;
        RECT 53.965 173.395 54.135 173.855 ;
        RECT 54.305 173.565 54.675 174.025 ;
        RECT 54.970 173.425 55.140 173.765 ;
        RECT 55.310 173.595 55.640 174.025 ;
        RECT 55.875 173.425 56.045 173.765 ;
        RECT 51.810 172.965 53.030 173.135 ;
        RECT 53.200 173.055 53.660 173.345 ;
        RECT 53.965 173.225 54.525 173.395 ;
        RECT 54.970 173.255 56.045 173.425 ;
        RECT 56.215 173.525 56.895 173.855 ;
        RECT 57.110 173.525 57.360 173.855 ;
        RECT 57.530 173.565 57.780 174.025 ;
        RECT 54.355 173.085 54.525 173.225 ;
        RECT 53.200 173.045 54.165 173.055 ;
        RECT 52.860 172.875 53.030 172.965 ;
        RECT 53.490 172.885 54.165 173.045 ;
        RECT 50.900 172.685 51.640 172.715 ;
        RECT 50.900 172.385 51.815 172.685 ;
        RECT 51.490 172.210 51.815 172.385 ;
        RECT 50.520 171.655 50.775 172.185 ;
        RECT 50.945 171.475 51.250 171.935 ;
        RECT 51.495 171.855 51.815 172.210 ;
        RECT 51.985 172.425 52.525 172.795 ;
        RECT 52.860 172.705 53.265 172.875 ;
        RECT 51.985 172.025 52.225 172.425 ;
        RECT 52.705 172.255 52.925 172.535 ;
        RECT 52.395 172.085 52.925 172.255 ;
        RECT 52.395 171.855 52.565 172.085 ;
        RECT 53.095 171.925 53.265 172.705 ;
        RECT 53.435 172.095 53.785 172.715 ;
        RECT 53.955 172.095 54.165 172.885 ;
        RECT 54.355 172.915 55.855 173.085 ;
        RECT 54.355 172.225 54.525 172.915 ;
        RECT 56.215 172.745 56.385 173.525 ;
        RECT 57.190 173.395 57.360 173.525 ;
        RECT 54.695 172.575 56.385 172.745 ;
        RECT 56.555 172.965 57.020 173.355 ;
        RECT 57.190 173.225 57.585 173.395 ;
        RECT 54.695 172.395 54.865 172.575 ;
        RECT 51.495 171.685 52.565 171.855 ;
        RECT 52.735 171.475 52.925 171.915 ;
        RECT 53.095 171.645 54.045 171.925 ;
        RECT 54.355 171.835 54.615 172.225 ;
        RECT 55.035 172.155 55.825 172.405 ;
        RECT 54.265 171.665 54.615 171.835 ;
        RECT 54.825 171.475 55.155 171.935 ;
        RECT 56.030 171.865 56.200 172.575 ;
        RECT 56.555 172.375 56.725 172.965 ;
        RECT 56.370 172.155 56.725 172.375 ;
        RECT 56.895 172.155 57.245 172.775 ;
        RECT 57.415 171.865 57.585 173.225 ;
        RECT 57.950 173.055 58.275 173.840 ;
        RECT 57.755 172.005 58.215 173.055 ;
        RECT 56.030 171.695 56.885 171.865 ;
        RECT 57.090 171.695 57.585 171.865 ;
        RECT 57.755 171.475 58.085 171.835 ;
        RECT 58.445 171.735 58.615 173.855 ;
        RECT 58.785 173.525 59.115 174.025 ;
        RECT 59.285 173.355 59.540 173.855 ;
        RECT 58.790 173.185 59.540 173.355 ;
        RECT 58.790 172.195 59.020 173.185 ;
        RECT 59.190 172.365 59.540 173.015 ;
        RECT 59.715 172.935 61.385 174.025 ;
        RECT 59.715 172.415 60.465 172.935 ;
        RECT 61.555 172.860 61.845 174.025 ;
        RECT 62.015 172.935 63.225 174.025 ;
        RECT 60.635 172.245 61.385 172.765 ;
        RECT 62.015 172.395 62.535 172.935 ;
        RECT 63.400 172.875 63.660 174.025 ;
        RECT 63.835 172.950 64.090 173.855 ;
        RECT 64.260 173.265 64.590 174.025 ;
        RECT 64.805 173.095 64.975 173.855 ;
        RECT 58.790 172.025 59.540 172.195 ;
        RECT 58.785 171.475 59.115 171.855 ;
        RECT 59.285 171.735 59.540 172.025 ;
        RECT 59.715 171.475 61.385 172.245 ;
        RECT 62.705 172.225 63.225 172.765 ;
        RECT 61.555 171.475 61.845 172.200 ;
        RECT 62.015 171.475 63.225 172.225 ;
        RECT 63.400 171.475 63.660 172.315 ;
        RECT 63.835 172.220 64.005 172.950 ;
        RECT 64.260 172.925 64.975 173.095 ;
        RECT 65.900 173.055 66.230 173.855 ;
        RECT 66.400 173.225 66.730 174.025 ;
        RECT 67.030 173.055 67.360 173.855 ;
        RECT 68.005 173.225 68.255 174.025 ;
        RECT 64.260 172.715 64.430 172.925 ;
        RECT 65.900 172.885 68.335 173.055 ;
        RECT 68.525 172.885 68.695 174.025 ;
        RECT 68.865 172.885 69.205 173.855 ;
        RECT 64.175 172.385 64.430 172.715 ;
        RECT 63.835 171.645 64.090 172.220 ;
        RECT 64.260 172.195 64.430 172.385 ;
        RECT 64.710 172.375 65.065 172.745 ;
        RECT 65.695 172.465 66.045 172.715 ;
        RECT 66.230 172.255 66.400 172.885 ;
        RECT 66.570 172.465 66.900 172.665 ;
        RECT 67.070 172.465 67.400 172.665 ;
        RECT 67.570 172.465 67.990 172.665 ;
        RECT 68.165 172.635 68.335 172.885 ;
        RECT 68.165 172.465 68.860 172.635 ;
        RECT 64.260 172.025 64.975 172.195 ;
        RECT 64.260 171.475 64.590 171.855 ;
        RECT 64.805 171.645 64.975 172.025 ;
        RECT 65.900 171.645 66.400 172.255 ;
        RECT 67.030 172.125 68.255 172.295 ;
        RECT 69.030 172.275 69.205 172.885 ;
        RECT 67.030 171.645 67.360 172.125 ;
        RECT 67.530 171.475 67.755 171.935 ;
        RECT 67.925 171.645 68.255 172.125 ;
        RECT 68.445 171.475 68.695 172.275 ;
        RECT 68.865 171.645 69.205 172.275 ;
        RECT 69.375 172.885 69.715 173.855 ;
        RECT 69.885 172.885 70.055 174.025 ;
        RECT 70.325 173.225 70.575 174.025 ;
        RECT 71.220 173.055 71.550 173.855 ;
        RECT 71.850 173.225 72.180 174.025 ;
        RECT 72.350 173.055 72.680 173.855 ;
        RECT 70.245 172.885 72.680 173.055 ;
        RECT 73.555 172.885 73.785 174.025 ;
        RECT 69.375 172.275 69.550 172.885 ;
        RECT 70.245 172.635 70.415 172.885 ;
        RECT 69.720 172.465 70.415 172.635 ;
        RECT 70.590 172.465 71.010 172.665 ;
        RECT 71.180 172.465 71.510 172.665 ;
        RECT 71.680 172.465 72.010 172.665 ;
        RECT 69.375 171.645 69.715 172.275 ;
        RECT 69.885 171.475 70.135 172.275 ;
        RECT 70.325 172.125 71.550 172.295 ;
        RECT 70.325 171.645 70.655 172.125 ;
        RECT 70.825 171.475 71.050 171.935 ;
        RECT 71.220 171.645 71.550 172.125 ;
        RECT 72.180 172.255 72.350 172.885 ;
        RECT 73.955 172.875 74.285 173.855 ;
        RECT 74.455 172.885 74.665 174.025 ;
        RECT 74.905 173.045 75.235 173.855 ;
        RECT 75.405 173.225 75.645 174.025 ;
        RECT 74.905 172.875 75.620 173.045 ;
        RECT 72.535 172.465 72.885 172.715 ;
        RECT 73.535 172.465 73.865 172.715 ;
        RECT 72.180 171.645 72.680 172.255 ;
        RECT 73.555 171.475 73.785 172.295 ;
        RECT 74.035 172.275 74.285 172.875 ;
        RECT 74.900 172.465 75.280 172.705 ;
        RECT 75.450 172.635 75.620 172.875 ;
        RECT 75.825 173.005 75.995 173.855 ;
        RECT 76.165 173.225 76.495 174.025 ;
        RECT 76.665 173.005 76.835 173.855 ;
        RECT 75.825 172.835 76.835 173.005 ;
        RECT 77.005 172.875 77.335 174.025 ;
        RECT 76.340 172.665 76.835 172.835 ;
        RECT 75.450 172.465 75.950 172.635 ;
        RECT 76.335 172.495 76.835 172.665 ;
        RECT 75.450 172.295 75.620 172.465 ;
        RECT 76.340 172.295 76.835 172.495 ;
        RECT 73.955 171.645 74.285 172.275 ;
        RECT 74.455 171.475 74.665 172.295 ;
        RECT 74.985 172.125 75.620 172.295 ;
        RECT 75.825 172.125 76.835 172.295 ;
        RECT 78.120 172.835 78.375 173.715 ;
        RECT 78.545 172.885 78.850 174.025 ;
        RECT 79.190 173.645 79.520 174.025 ;
        RECT 79.700 173.475 79.870 173.765 ;
        RECT 80.040 173.565 80.290 174.025 ;
        RECT 79.070 173.305 79.870 173.475 ;
        RECT 80.460 173.515 81.330 173.855 ;
        RECT 74.985 171.645 75.155 172.125 ;
        RECT 75.335 171.475 75.575 171.955 ;
        RECT 75.825 171.645 75.995 172.125 ;
        RECT 76.165 171.475 76.495 171.955 ;
        RECT 76.665 171.645 76.835 172.125 ;
        RECT 77.005 171.475 77.335 172.275 ;
        RECT 78.120 172.185 78.330 172.835 ;
        RECT 79.070 172.715 79.240 173.305 ;
        RECT 80.460 173.135 80.630 173.515 ;
        RECT 81.565 173.395 81.735 173.855 ;
        RECT 81.905 173.565 82.275 174.025 ;
        RECT 82.570 173.425 82.740 173.765 ;
        RECT 82.910 173.595 83.240 174.025 ;
        RECT 83.475 173.425 83.645 173.765 ;
        RECT 79.410 172.965 80.630 173.135 ;
        RECT 80.800 173.055 81.260 173.345 ;
        RECT 81.565 173.225 82.125 173.395 ;
        RECT 82.570 173.255 83.645 173.425 ;
        RECT 83.815 173.525 84.495 173.855 ;
        RECT 84.710 173.525 84.960 173.855 ;
        RECT 85.130 173.565 85.380 174.025 ;
        RECT 81.955 173.085 82.125 173.225 ;
        RECT 80.800 173.045 81.765 173.055 ;
        RECT 80.460 172.875 80.630 172.965 ;
        RECT 81.090 172.885 81.765 173.045 ;
        RECT 78.500 172.685 79.240 172.715 ;
        RECT 78.500 172.385 79.415 172.685 ;
        RECT 79.090 172.210 79.415 172.385 ;
        RECT 78.120 171.655 78.375 172.185 ;
        RECT 78.545 171.475 78.850 171.935 ;
        RECT 79.095 171.855 79.415 172.210 ;
        RECT 79.585 172.425 80.125 172.795 ;
        RECT 80.460 172.705 80.865 172.875 ;
        RECT 79.585 172.025 79.825 172.425 ;
        RECT 80.305 172.255 80.525 172.535 ;
        RECT 79.995 172.085 80.525 172.255 ;
        RECT 79.995 171.855 80.165 172.085 ;
        RECT 80.695 171.925 80.865 172.705 ;
        RECT 81.035 172.095 81.385 172.715 ;
        RECT 81.555 172.095 81.765 172.885 ;
        RECT 81.955 172.915 83.455 173.085 ;
        RECT 81.955 172.225 82.125 172.915 ;
        RECT 83.815 172.745 83.985 173.525 ;
        RECT 84.790 173.395 84.960 173.525 ;
        RECT 82.295 172.575 83.985 172.745 ;
        RECT 84.155 172.965 84.620 173.355 ;
        RECT 84.790 173.225 85.185 173.395 ;
        RECT 82.295 172.395 82.465 172.575 ;
        RECT 79.095 171.685 80.165 171.855 ;
        RECT 80.335 171.475 80.525 171.915 ;
        RECT 80.695 171.645 81.645 171.925 ;
        RECT 81.955 171.835 82.215 172.225 ;
        RECT 82.635 172.155 83.425 172.405 ;
        RECT 81.865 171.665 82.215 171.835 ;
        RECT 82.425 171.475 82.755 171.935 ;
        RECT 83.630 171.865 83.800 172.575 ;
        RECT 84.155 172.375 84.325 172.965 ;
        RECT 83.970 172.155 84.325 172.375 ;
        RECT 84.495 172.155 84.845 172.775 ;
        RECT 85.015 171.865 85.185 173.225 ;
        RECT 85.550 173.055 85.875 173.840 ;
        RECT 85.355 172.005 85.815 173.055 ;
        RECT 83.630 171.695 84.485 171.865 ;
        RECT 84.690 171.695 85.185 171.865 ;
        RECT 85.355 171.475 85.685 171.835 ;
        RECT 86.045 171.735 86.215 173.855 ;
        RECT 86.385 173.525 86.715 174.025 ;
        RECT 86.885 173.355 87.140 173.855 ;
        RECT 86.390 173.185 87.140 173.355 ;
        RECT 86.390 172.195 86.620 173.185 ;
        RECT 86.790 172.365 87.140 173.015 ;
        RECT 87.315 172.860 87.605 174.025 ;
        RECT 87.980 173.055 88.310 173.855 ;
        RECT 88.480 173.225 88.810 174.025 ;
        RECT 89.110 173.055 89.440 173.855 ;
        RECT 90.085 173.225 90.335 174.025 ;
        RECT 87.980 172.885 90.415 173.055 ;
        RECT 90.605 172.885 90.775 174.025 ;
        RECT 90.945 172.885 91.285 173.855 ;
        RECT 91.660 173.055 91.990 173.855 ;
        RECT 92.160 173.225 92.490 174.025 ;
        RECT 92.790 173.055 93.120 173.855 ;
        RECT 93.765 173.225 94.015 174.025 ;
        RECT 91.660 172.885 94.095 173.055 ;
        RECT 94.285 172.885 94.455 174.025 ;
        RECT 94.625 172.885 94.965 173.855 ;
        RECT 87.775 172.465 88.125 172.715 ;
        RECT 88.310 172.255 88.480 172.885 ;
        RECT 88.650 172.465 88.980 172.665 ;
        RECT 89.150 172.465 89.480 172.665 ;
        RECT 89.650 172.465 90.070 172.665 ;
        RECT 90.245 172.635 90.415 172.885 ;
        RECT 90.245 172.465 90.940 172.635 ;
        RECT 86.390 172.025 87.140 172.195 ;
        RECT 86.385 171.475 86.715 171.855 ;
        RECT 86.885 171.735 87.140 172.025 ;
        RECT 87.315 171.475 87.605 172.200 ;
        RECT 87.980 171.645 88.480 172.255 ;
        RECT 89.110 172.125 90.335 172.295 ;
        RECT 91.110 172.275 91.285 172.885 ;
        RECT 91.455 172.465 91.805 172.715 ;
        RECT 89.110 171.645 89.440 172.125 ;
        RECT 89.610 171.475 89.835 171.935 ;
        RECT 90.005 171.645 90.335 172.125 ;
        RECT 90.525 171.475 90.775 172.275 ;
        RECT 90.945 171.645 91.285 172.275 ;
        RECT 91.990 172.255 92.160 172.885 ;
        RECT 92.330 172.465 92.660 172.665 ;
        RECT 92.830 172.465 93.160 172.665 ;
        RECT 93.330 172.465 93.750 172.665 ;
        RECT 93.925 172.635 94.095 172.885 ;
        RECT 93.925 172.465 94.620 172.635 ;
        RECT 91.660 171.645 92.160 172.255 ;
        RECT 92.790 172.125 94.015 172.295 ;
        RECT 94.790 172.275 94.965 172.885 ;
        RECT 96.055 173.265 96.570 173.675 ;
        RECT 96.805 173.265 96.975 174.025 ;
        RECT 97.145 173.685 99.175 173.855 ;
        RECT 96.055 172.455 96.395 173.265 ;
        RECT 97.145 173.020 97.315 173.685 ;
        RECT 97.710 173.345 98.835 173.515 ;
        RECT 96.565 172.830 97.315 173.020 ;
        RECT 97.485 173.005 98.495 173.175 ;
        RECT 96.055 172.285 97.285 172.455 ;
        RECT 92.790 171.645 93.120 172.125 ;
        RECT 93.290 171.475 93.515 171.935 ;
        RECT 93.685 171.645 94.015 172.125 ;
        RECT 94.205 171.475 94.455 172.275 ;
        RECT 94.625 171.645 94.965 172.275 ;
        RECT 96.330 171.680 96.575 172.285 ;
        RECT 96.795 171.475 97.305 172.010 ;
        RECT 97.485 171.645 97.675 173.005 ;
        RECT 97.845 172.665 98.120 172.805 ;
        RECT 97.845 172.495 98.125 172.665 ;
        RECT 97.845 171.645 98.120 172.495 ;
        RECT 98.325 172.205 98.495 173.005 ;
        RECT 98.665 172.215 98.835 173.345 ;
        RECT 99.005 172.715 99.175 173.685 ;
        RECT 99.345 172.885 99.515 174.025 ;
        RECT 99.685 172.885 100.020 173.855 ;
        RECT 101.155 172.885 101.385 174.025 ;
        RECT 99.005 172.385 99.200 172.715 ;
        RECT 99.425 172.385 99.680 172.715 ;
        RECT 99.425 172.215 99.595 172.385 ;
        RECT 99.850 172.215 100.020 172.885 ;
        RECT 101.555 172.875 101.885 173.855 ;
        RECT 102.055 172.885 102.265 174.025 ;
        RECT 101.135 172.465 101.465 172.715 ;
        RECT 98.665 172.045 99.595 172.215 ;
        RECT 98.665 172.010 98.840 172.045 ;
        RECT 98.310 171.645 98.840 172.010 ;
        RECT 99.265 171.475 99.595 171.875 ;
        RECT 99.765 171.645 100.020 172.215 ;
        RECT 101.155 171.475 101.385 172.295 ;
        RECT 101.635 172.275 101.885 172.875 ;
        RECT 102.500 172.835 102.755 173.715 ;
        RECT 102.925 172.885 103.230 174.025 ;
        RECT 103.570 173.645 103.900 174.025 ;
        RECT 104.080 173.475 104.250 173.765 ;
        RECT 104.420 173.565 104.670 174.025 ;
        RECT 103.450 173.305 104.250 173.475 ;
        RECT 104.840 173.515 105.710 173.855 ;
        RECT 101.555 171.645 101.885 172.275 ;
        RECT 102.055 171.475 102.265 172.295 ;
        RECT 102.500 172.185 102.710 172.835 ;
        RECT 103.450 172.715 103.620 173.305 ;
        RECT 104.840 173.135 105.010 173.515 ;
        RECT 105.945 173.395 106.115 173.855 ;
        RECT 106.285 173.565 106.655 174.025 ;
        RECT 106.950 173.425 107.120 173.765 ;
        RECT 107.290 173.595 107.620 174.025 ;
        RECT 107.855 173.425 108.025 173.765 ;
        RECT 103.790 172.965 105.010 173.135 ;
        RECT 105.180 173.055 105.640 173.345 ;
        RECT 105.945 173.225 106.505 173.395 ;
        RECT 106.950 173.255 108.025 173.425 ;
        RECT 108.195 173.525 108.875 173.855 ;
        RECT 109.090 173.525 109.340 173.855 ;
        RECT 109.510 173.565 109.760 174.025 ;
        RECT 106.335 173.085 106.505 173.225 ;
        RECT 105.180 173.045 106.145 173.055 ;
        RECT 104.840 172.875 105.010 172.965 ;
        RECT 105.470 172.885 106.145 173.045 ;
        RECT 102.880 172.685 103.620 172.715 ;
        RECT 102.880 172.385 103.795 172.685 ;
        RECT 103.470 172.210 103.795 172.385 ;
        RECT 102.500 171.655 102.755 172.185 ;
        RECT 102.925 171.475 103.230 171.935 ;
        RECT 103.475 171.855 103.795 172.210 ;
        RECT 103.965 172.425 104.505 172.795 ;
        RECT 104.840 172.705 105.245 172.875 ;
        RECT 103.965 172.025 104.205 172.425 ;
        RECT 104.685 172.255 104.905 172.535 ;
        RECT 104.375 172.085 104.905 172.255 ;
        RECT 104.375 171.855 104.545 172.085 ;
        RECT 105.075 171.925 105.245 172.705 ;
        RECT 105.415 172.095 105.765 172.715 ;
        RECT 105.935 172.095 106.145 172.885 ;
        RECT 106.335 172.915 107.835 173.085 ;
        RECT 106.335 172.225 106.505 172.915 ;
        RECT 108.195 172.745 108.365 173.525 ;
        RECT 109.170 173.395 109.340 173.525 ;
        RECT 106.675 172.575 108.365 172.745 ;
        RECT 108.535 172.965 109.000 173.355 ;
        RECT 109.170 173.225 109.565 173.395 ;
        RECT 106.675 172.395 106.845 172.575 ;
        RECT 103.475 171.685 104.545 171.855 ;
        RECT 104.715 171.475 104.905 171.915 ;
        RECT 105.075 171.645 106.025 171.925 ;
        RECT 106.335 171.835 106.595 172.225 ;
        RECT 107.015 172.155 107.805 172.405 ;
        RECT 106.245 171.665 106.595 171.835 ;
        RECT 106.805 171.475 107.135 171.935 ;
        RECT 108.010 171.865 108.180 172.575 ;
        RECT 108.535 172.375 108.705 172.965 ;
        RECT 108.350 172.155 108.705 172.375 ;
        RECT 108.875 172.155 109.225 172.775 ;
        RECT 109.395 171.865 109.565 173.225 ;
        RECT 109.930 173.055 110.255 173.840 ;
        RECT 109.735 172.005 110.195 173.055 ;
        RECT 108.010 171.695 108.865 171.865 ;
        RECT 109.070 171.695 109.565 171.865 ;
        RECT 109.735 171.475 110.065 171.835 ;
        RECT 110.425 171.735 110.595 173.855 ;
        RECT 110.765 173.525 111.095 174.025 ;
        RECT 111.265 173.355 111.520 173.855 ;
        RECT 110.770 173.185 111.520 173.355 ;
        RECT 110.770 172.195 111.000 173.185 ;
        RECT 111.170 172.365 111.520 173.015 ;
        RECT 112.155 172.935 113.365 174.025 ;
        RECT 112.155 172.395 112.675 172.935 ;
        RECT 112.845 172.225 113.365 172.765 ;
        RECT 110.770 172.025 111.520 172.195 ;
        RECT 110.765 171.475 111.095 171.855 ;
        RECT 111.265 171.735 111.520 172.025 ;
        RECT 112.155 171.475 113.365 172.225 ;
        RECT 11.330 171.305 113.450 171.475 ;
        RECT 11.415 170.555 12.625 171.305 ;
        RECT 11.415 170.015 11.935 170.555 ;
        RECT 13.715 170.535 17.225 171.305 ;
        RECT 17.400 170.760 22.745 171.305 ;
        RECT 12.105 169.845 12.625 170.385 ;
        RECT 11.415 168.755 12.625 169.845 ;
        RECT 13.715 169.845 15.405 170.365 ;
        RECT 15.575 170.015 17.225 170.535 ;
        RECT 13.715 168.755 17.225 169.845 ;
        RECT 18.990 169.190 19.340 170.440 ;
        RECT 20.820 169.930 21.160 170.760 ;
        RECT 22.915 170.580 23.205 171.305 ;
        RECT 23.895 170.485 24.105 171.305 ;
        RECT 24.275 170.505 24.605 171.135 ;
        RECT 17.400 168.755 22.745 169.190 ;
        RECT 22.915 168.755 23.205 169.920 ;
        RECT 24.275 169.905 24.525 170.505 ;
        RECT 24.775 170.485 25.005 171.305 ;
        RECT 25.215 170.555 26.425 171.305 ;
        RECT 24.695 170.065 25.025 170.315 ;
        RECT 23.895 168.755 24.105 169.895 ;
        RECT 24.275 168.925 24.605 169.905 ;
        RECT 24.775 168.755 25.005 169.895 ;
        RECT 25.215 169.845 25.735 170.385 ;
        RECT 25.905 170.015 26.425 170.555 ;
        RECT 26.595 170.505 26.935 171.135 ;
        RECT 27.105 170.505 27.355 171.305 ;
        RECT 27.545 170.655 27.875 171.135 ;
        RECT 28.045 170.845 28.270 171.305 ;
        RECT 28.440 170.655 28.770 171.135 ;
        RECT 26.595 169.895 26.770 170.505 ;
        RECT 27.545 170.485 28.770 170.655 ;
        RECT 29.400 170.525 29.900 171.135 ;
        RECT 26.940 170.145 27.635 170.315 ;
        RECT 27.465 169.895 27.635 170.145 ;
        RECT 27.810 170.115 28.230 170.315 ;
        RECT 28.400 170.115 28.730 170.315 ;
        RECT 28.900 170.115 29.230 170.315 ;
        RECT 29.400 169.895 29.570 170.525 ;
        RECT 30.275 170.505 30.615 171.135 ;
        RECT 30.785 170.505 31.035 171.305 ;
        RECT 31.225 170.655 31.555 171.135 ;
        RECT 31.725 170.845 31.950 171.305 ;
        RECT 32.120 170.655 32.450 171.135 ;
        RECT 29.755 170.065 30.105 170.315 ;
        RECT 30.275 169.895 30.450 170.505 ;
        RECT 31.225 170.485 32.450 170.655 ;
        RECT 33.080 170.525 33.580 171.135 ;
        RECT 33.955 170.535 37.465 171.305 ;
        RECT 30.620 170.145 31.315 170.315 ;
        RECT 31.145 169.895 31.315 170.145 ;
        RECT 31.490 170.115 31.910 170.315 ;
        RECT 32.080 170.115 32.410 170.315 ;
        RECT 32.580 170.115 32.910 170.315 ;
        RECT 33.080 169.895 33.250 170.525 ;
        RECT 33.435 170.065 33.785 170.315 ;
        RECT 25.215 168.755 26.425 169.845 ;
        RECT 26.595 168.925 26.935 169.895 ;
        RECT 27.105 168.755 27.275 169.895 ;
        RECT 27.465 169.725 29.900 169.895 ;
        RECT 27.545 168.755 27.795 169.555 ;
        RECT 28.440 168.925 28.770 169.725 ;
        RECT 29.070 168.755 29.400 169.555 ;
        RECT 29.570 168.925 29.900 169.725 ;
        RECT 30.275 168.925 30.615 169.895 ;
        RECT 30.785 168.755 30.955 169.895 ;
        RECT 31.145 169.725 33.580 169.895 ;
        RECT 31.225 168.755 31.475 169.555 ;
        RECT 32.120 168.925 32.450 169.725 ;
        RECT 32.750 168.755 33.080 169.555 ;
        RECT 33.250 168.925 33.580 169.725 ;
        RECT 33.955 169.845 35.645 170.365 ;
        RECT 35.815 170.015 37.465 170.535 ;
        RECT 37.635 170.505 37.975 171.135 ;
        RECT 38.145 170.505 38.395 171.305 ;
        RECT 38.585 170.655 38.915 171.135 ;
        RECT 39.085 170.845 39.310 171.305 ;
        RECT 39.480 170.655 39.810 171.135 ;
        RECT 37.635 169.895 37.810 170.505 ;
        RECT 38.585 170.485 39.810 170.655 ;
        RECT 40.440 170.525 40.940 171.135 ;
        RECT 37.980 170.145 38.675 170.315 ;
        RECT 38.505 169.895 38.675 170.145 ;
        RECT 38.850 170.115 39.270 170.315 ;
        RECT 39.440 170.115 39.770 170.315 ;
        RECT 39.940 170.115 40.270 170.315 ;
        RECT 40.440 169.895 40.610 170.525 ;
        RECT 41.315 170.505 41.655 171.135 ;
        RECT 41.825 170.505 42.075 171.305 ;
        RECT 42.265 170.655 42.595 171.135 ;
        RECT 42.765 170.845 42.990 171.305 ;
        RECT 43.160 170.655 43.490 171.135 ;
        RECT 40.795 170.065 41.145 170.315 ;
        RECT 41.315 169.895 41.490 170.505 ;
        RECT 42.265 170.485 43.490 170.655 ;
        RECT 44.120 170.525 44.620 171.135 ;
        RECT 41.660 170.145 42.355 170.315 ;
        RECT 42.185 169.895 42.355 170.145 ;
        RECT 42.530 170.115 42.950 170.315 ;
        RECT 43.120 170.115 43.450 170.315 ;
        RECT 43.620 170.115 43.950 170.315 ;
        RECT 44.120 169.895 44.290 170.525 ;
        RECT 44.995 170.505 45.335 171.135 ;
        RECT 45.505 170.505 45.755 171.305 ;
        RECT 45.945 170.655 46.275 171.135 ;
        RECT 46.445 170.845 46.670 171.305 ;
        RECT 46.840 170.655 47.170 171.135 ;
        RECT 44.475 170.065 44.825 170.315 ;
        RECT 44.995 169.895 45.170 170.505 ;
        RECT 45.945 170.485 47.170 170.655 ;
        RECT 47.800 170.525 48.300 171.135 ;
        RECT 48.675 170.580 48.965 171.305 ;
        RECT 49.250 170.675 49.535 171.135 ;
        RECT 49.705 170.845 49.975 171.305 ;
        RECT 45.340 170.145 46.035 170.315 ;
        RECT 45.865 169.895 46.035 170.145 ;
        RECT 46.210 170.115 46.630 170.315 ;
        RECT 46.800 170.115 47.130 170.315 ;
        RECT 47.300 170.115 47.630 170.315 ;
        RECT 47.800 169.895 47.970 170.525 ;
        RECT 49.250 170.505 50.205 170.675 ;
        RECT 48.155 170.065 48.505 170.315 ;
        RECT 33.955 168.755 37.465 169.845 ;
        RECT 37.635 168.925 37.975 169.895 ;
        RECT 38.145 168.755 38.315 169.895 ;
        RECT 38.505 169.725 40.940 169.895 ;
        RECT 38.585 168.755 38.835 169.555 ;
        RECT 39.480 168.925 39.810 169.725 ;
        RECT 40.110 168.755 40.440 169.555 ;
        RECT 40.610 168.925 40.940 169.725 ;
        RECT 41.315 168.925 41.655 169.895 ;
        RECT 41.825 168.755 41.995 169.895 ;
        RECT 42.185 169.725 44.620 169.895 ;
        RECT 42.265 168.755 42.515 169.555 ;
        RECT 43.160 168.925 43.490 169.725 ;
        RECT 43.790 168.755 44.120 169.555 ;
        RECT 44.290 168.925 44.620 169.725 ;
        RECT 44.995 168.925 45.335 169.895 ;
        RECT 45.505 168.755 45.675 169.895 ;
        RECT 45.865 169.725 48.300 169.895 ;
        RECT 45.945 168.755 46.195 169.555 ;
        RECT 46.840 168.925 47.170 169.725 ;
        RECT 47.470 168.755 47.800 169.555 ;
        RECT 47.970 168.925 48.300 169.725 ;
        RECT 48.675 168.755 48.965 169.920 ;
        RECT 49.135 169.775 49.825 170.335 ;
        RECT 49.995 169.605 50.205 170.505 ;
        RECT 49.250 169.385 50.205 169.605 ;
        RECT 50.375 170.335 50.775 171.135 ;
        RECT 50.965 170.675 51.245 171.135 ;
        RECT 51.765 170.845 52.090 171.305 ;
        RECT 50.965 170.505 52.090 170.675 ;
        RECT 52.260 170.565 52.645 171.135 ;
        RECT 51.640 170.395 52.090 170.505 ;
        RECT 50.375 169.775 51.470 170.335 ;
        RECT 51.640 170.065 52.195 170.395 ;
        RECT 49.250 168.925 49.535 169.385 ;
        RECT 49.705 168.755 49.975 169.215 ;
        RECT 50.375 168.925 50.775 169.775 ;
        RECT 51.640 169.605 52.090 170.065 ;
        RECT 52.365 169.895 52.645 170.565 ;
        RECT 53.795 170.485 54.005 171.305 ;
        RECT 54.175 170.505 54.505 171.135 ;
        RECT 54.175 169.905 54.425 170.505 ;
        RECT 54.675 170.485 54.905 171.305 ;
        RECT 55.205 170.755 55.375 171.135 ;
        RECT 55.555 170.925 55.885 171.305 ;
        RECT 55.205 170.585 55.870 170.755 ;
        RECT 56.065 170.630 56.325 171.135 ;
        RECT 57.420 170.760 62.765 171.305 ;
        RECT 54.595 170.065 54.925 170.315 ;
        RECT 55.135 170.035 55.465 170.405 ;
        RECT 55.700 170.330 55.870 170.585 ;
        RECT 55.700 170.000 55.985 170.330 ;
        RECT 50.965 169.385 52.090 169.605 ;
        RECT 50.965 168.925 51.245 169.385 ;
        RECT 51.765 168.755 52.090 169.215 ;
        RECT 52.260 168.925 52.645 169.895 ;
        RECT 53.795 168.755 54.005 169.895 ;
        RECT 54.175 168.925 54.505 169.905 ;
        RECT 54.675 168.755 54.905 169.895 ;
        RECT 55.700 169.855 55.870 170.000 ;
        RECT 55.205 169.685 55.870 169.855 ;
        RECT 56.155 169.830 56.325 170.630 ;
        RECT 55.205 168.925 55.375 169.685 ;
        RECT 55.555 168.755 55.885 169.515 ;
        RECT 56.055 168.925 56.325 169.830 ;
        RECT 59.010 169.190 59.360 170.440 ;
        RECT 60.840 169.930 61.180 170.760 ;
        RECT 62.940 170.465 63.200 171.305 ;
        RECT 63.375 170.560 63.630 171.135 ;
        RECT 63.800 170.925 64.130 171.305 ;
        RECT 64.345 170.755 64.515 171.135 ;
        RECT 64.780 170.760 70.125 171.305 ;
        RECT 63.800 170.585 64.515 170.755 ;
        RECT 57.420 168.755 62.765 169.190 ;
        RECT 62.940 168.755 63.200 169.905 ;
        RECT 63.375 169.830 63.545 170.560 ;
        RECT 63.800 170.395 63.970 170.585 ;
        RECT 63.715 170.065 63.970 170.395 ;
        RECT 63.800 169.855 63.970 170.065 ;
        RECT 64.250 170.035 64.605 170.405 ;
        RECT 63.375 168.925 63.630 169.830 ;
        RECT 63.800 169.685 64.515 169.855 ;
        RECT 63.800 168.755 64.130 169.515 ;
        RECT 64.345 168.925 64.515 169.685 ;
        RECT 66.370 169.190 66.720 170.440 ;
        RECT 68.200 169.930 68.540 170.760 ;
        RECT 70.295 170.505 70.635 171.135 ;
        RECT 70.805 170.505 71.055 171.305 ;
        RECT 71.245 170.655 71.575 171.135 ;
        RECT 71.745 170.845 71.970 171.305 ;
        RECT 72.140 170.655 72.470 171.135 ;
        RECT 70.295 169.895 70.470 170.505 ;
        RECT 71.245 170.485 72.470 170.655 ;
        RECT 73.100 170.525 73.600 171.135 ;
        RECT 74.435 170.580 74.725 171.305 ;
        RECT 75.815 170.795 76.120 171.305 ;
        RECT 70.640 170.145 71.335 170.315 ;
        RECT 71.165 169.895 71.335 170.145 ;
        RECT 71.510 170.115 71.930 170.315 ;
        RECT 72.100 170.115 72.430 170.315 ;
        RECT 72.600 170.115 72.930 170.315 ;
        RECT 73.100 169.895 73.270 170.525 ;
        RECT 73.455 170.065 73.805 170.315 ;
        RECT 75.815 170.065 76.130 170.625 ;
        RECT 76.300 170.315 76.550 171.125 ;
        RECT 76.720 170.780 76.980 171.305 ;
        RECT 77.160 170.315 77.410 171.125 ;
        RECT 77.580 170.745 77.840 171.305 ;
        RECT 78.010 170.655 78.270 171.110 ;
        RECT 78.440 170.825 78.700 171.305 ;
        RECT 78.870 170.655 79.130 171.110 ;
        RECT 79.300 170.825 79.560 171.305 ;
        RECT 79.730 170.655 79.990 171.110 ;
        RECT 80.160 170.825 80.405 171.305 ;
        RECT 80.575 170.655 80.850 171.110 ;
        RECT 81.020 170.825 81.265 171.305 ;
        RECT 81.435 170.655 81.695 171.110 ;
        RECT 81.875 170.825 82.125 171.305 ;
        RECT 82.295 170.655 82.555 171.110 ;
        RECT 82.735 170.825 82.985 171.305 ;
        RECT 83.155 170.655 83.415 171.110 ;
        RECT 83.595 170.825 83.855 171.305 ;
        RECT 84.025 170.655 84.285 171.110 ;
        RECT 84.455 170.825 84.755 171.305 ;
        RECT 78.010 170.485 84.755 170.655 ;
        RECT 85.015 170.535 86.685 171.305 ;
        RECT 76.300 170.065 83.420 170.315 ;
        RECT 64.780 168.755 70.125 169.190 ;
        RECT 70.295 168.925 70.635 169.895 ;
        RECT 70.805 168.755 70.975 169.895 ;
        RECT 71.165 169.725 73.600 169.895 ;
        RECT 71.245 168.755 71.495 169.555 ;
        RECT 72.140 168.925 72.470 169.725 ;
        RECT 72.770 168.755 73.100 169.555 ;
        RECT 73.270 168.925 73.600 169.725 ;
        RECT 74.435 168.755 74.725 169.920 ;
        RECT 75.825 168.755 76.120 169.565 ;
        RECT 76.300 168.925 76.545 170.065 ;
        RECT 76.720 168.755 76.980 169.565 ;
        RECT 77.160 168.930 77.410 170.065 ;
        RECT 83.590 169.895 84.755 170.485 ;
        RECT 78.010 169.670 84.755 169.895 ;
        RECT 85.015 169.845 85.765 170.365 ;
        RECT 85.935 170.015 86.685 170.535 ;
        RECT 86.895 170.485 87.125 171.305 ;
        RECT 87.295 170.505 87.625 171.135 ;
        RECT 86.875 170.065 87.205 170.315 ;
        RECT 87.375 169.905 87.625 170.505 ;
        RECT 87.795 170.485 88.005 171.305 ;
        RECT 88.240 170.595 88.495 171.125 ;
        RECT 88.665 170.845 88.970 171.305 ;
        RECT 89.215 170.925 90.285 171.095 ;
        RECT 78.010 169.655 83.415 169.670 ;
        RECT 77.580 168.760 77.840 169.555 ;
        RECT 78.010 168.930 78.270 169.655 ;
        RECT 78.440 168.760 78.700 169.485 ;
        RECT 78.870 168.930 79.130 169.655 ;
        RECT 79.300 168.760 79.560 169.485 ;
        RECT 79.730 168.930 79.990 169.655 ;
        RECT 80.160 168.760 80.420 169.485 ;
        RECT 80.590 168.930 80.850 169.655 ;
        RECT 81.020 168.760 81.265 169.485 ;
        RECT 81.435 168.930 81.695 169.655 ;
        RECT 81.880 168.760 82.125 169.485 ;
        RECT 82.295 168.930 82.555 169.655 ;
        RECT 82.740 168.760 82.985 169.485 ;
        RECT 83.155 168.930 83.415 169.655 ;
        RECT 83.600 168.760 83.855 169.485 ;
        RECT 84.025 168.930 84.315 169.670 ;
        RECT 77.580 168.755 83.855 168.760 ;
        RECT 84.485 168.755 84.755 169.500 ;
        RECT 85.015 168.755 86.685 169.845 ;
        RECT 86.895 168.755 87.125 169.895 ;
        RECT 87.295 168.925 87.625 169.905 ;
        RECT 88.240 169.945 88.450 170.595 ;
        RECT 89.215 170.570 89.535 170.925 ;
        RECT 89.210 170.395 89.535 170.570 ;
        RECT 88.620 170.095 89.535 170.395 ;
        RECT 89.705 170.355 89.945 170.755 ;
        RECT 90.115 170.695 90.285 170.925 ;
        RECT 90.455 170.865 90.645 171.305 ;
        RECT 90.815 170.855 91.765 171.135 ;
        RECT 91.985 170.945 92.335 171.115 ;
        RECT 90.115 170.525 90.645 170.695 ;
        RECT 88.620 170.065 89.360 170.095 ;
        RECT 87.795 168.755 88.005 169.895 ;
        RECT 88.240 169.065 88.495 169.945 ;
        RECT 88.665 168.755 88.970 169.895 ;
        RECT 89.190 169.475 89.360 170.065 ;
        RECT 89.705 169.985 90.245 170.355 ;
        RECT 90.425 170.245 90.645 170.525 ;
        RECT 90.815 170.075 90.985 170.855 ;
        RECT 90.580 169.905 90.985 170.075 ;
        RECT 91.155 170.065 91.505 170.685 ;
        RECT 90.580 169.815 90.750 169.905 ;
        RECT 91.675 169.895 91.885 170.685 ;
        RECT 89.530 169.645 90.750 169.815 ;
        RECT 91.210 169.735 91.885 169.895 ;
        RECT 89.190 169.305 89.990 169.475 ;
        RECT 89.310 168.755 89.640 169.135 ;
        RECT 89.820 169.015 89.990 169.305 ;
        RECT 90.580 169.265 90.750 169.645 ;
        RECT 90.920 169.725 91.885 169.735 ;
        RECT 92.075 170.555 92.335 170.945 ;
        RECT 92.545 170.845 92.875 171.305 ;
        RECT 93.750 170.915 94.605 171.085 ;
        RECT 94.810 170.915 95.305 171.085 ;
        RECT 95.475 170.945 95.805 171.305 ;
        RECT 92.075 169.865 92.245 170.555 ;
        RECT 92.415 170.205 92.585 170.385 ;
        RECT 92.755 170.375 93.545 170.625 ;
        RECT 93.750 170.205 93.920 170.915 ;
        RECT 94.090 170.405 94.445 170.625 ;
        RECT 92.415 170.035 94.105 170.205 ;
        RECT 90.920 169.435 91.380 169.725 ;
        RECT 92.075 169.695 93.575 169.865 ;
        RECT 92.075 169.555 92.245 169.695 ;
        RECT 91.685 169.385 92.245 169.555 ;
        RECT 90.160 168.755 90.410 169.215 ;
        RECT 90.580 168.925 91.450 169.265 ;
        RECT 91.685 168.925 91.855 169.385 ;
        RECT 92.690 169.355 93.765 169.525 ;
        RECT 92.025 168.755 92.395 169.215 ;
        RECT 92.690 169.015 92.860 169.355 ;
        RECT 93.030 168.755 93.360 169.185 ;
        RECT 93.595 169.015 93.765 169.355 ;
        RECT 93.935 169.255 94.105 170.035 ;
        RECT 94.275 169.815 94.445 170.405 ;
        RECT 94.615 170.005 94.965 170.625 ;
        RECT 94.275 169.425 94.740 169.815 ;
        RECT 95.135 169.555 95.305 170.915 ;
        RECT 95.475 169.725 95.935 170.775 ;
        RECT 94.910 169.385 95.305 169.555 ;
        RECT 94.910 169.255 95.080 169.385 ;
        RECT 93.935 168.925 94.615 169.255 ;
        RECT 94.830 168.925 95.080 169.255 ;
        RECT 95.250 168.755 95.500 169.215 ;
        RECT 95.670 168.940 95.995 169.725 ;
        RECT 96.165 168.925 96.335 171.045 ;
        RECT 96.505 170.925 96.835 171.305 ;
        RECT 97.005 170.755 97.260 171.045 ;
        RECT 96.510 170.585 97.260 170.755 ;
        RECT 97.435 170.630 97.695 171.135 ;
        RECT 97.875 170.925 98.205 171.305 ;
        RECT 98.385 170.755 98.555 171.135 ;
        RECT 96.510 169.595 96.740 170.585 ;
        RECT 96.910 169.765 97.260 170.415 ;
        RECT 97.435 169.830 97.605 170.630 ;
        RECT 97.890 170.585 98.555 170.755 ;
        RECT 97.890 170.330 98.060 170.585 ;
        RECT 98.815 170.555 100.025 171.305 ;
        RECT 100.195 170.580 100.485 171.305 ;
        RECT 97.775 170.000 98.060 170.330 ;
        RECT 98.295 170.035 98.625 170.405 ;
        RECT 97.890 169.855 98.060 170.000 ;
        RECT 96.510 169.425 97.260 169.595 ;
        RECT 96.505 168.755 96.835 169.255 ;
        RECT 97.005 168.925 97.260 169.425 ;
        RECT 97.435 168.925 97.705 169.830 ;
        RECT 97.890 169.685 98.555 169.855 ;
        RECT 97.875 168.755 98.205 169.515 ;
        RECT 98.385 168.925 98.555 169.685 ;
        RECT 98.815 169.845 99.335 170.385 ;
        RECT 99.505 170.015 100.025 170.555 ;
        RECT 100.715 170.485 100.925 171.305 ;
        RECT 101.095 170.505 101.425 171.135 ;
        RECT 98.815 168.755 100.025 169.845 ;
        RECT 100.195 168.755 100.485 169.920 ;
        RECT 101.095 169.905 101.345 170.505 ;
        RECT 101.595 170.485 101.825 171.305 ;
        RECT 102.500 170.595 102.755 171.125 ;
        RECT 102.925 170.845 103.230 171.305 ;
        RECT 103.475 170.925 104.545 171.095 ;
        RECT 101.515 170.065 101.845 170.315 ;
        RECT 102.500 169.945 102.710 170.595 ;
        RECT 103.475 170.570 103.795 170.925 ;
        RECT 103.470 170.395 103.795 170.570 ;
        RECT 102.880 170.095 103.795 170.395 ;
        RECT 103.965 170.355 104.205 170.755 ;
        RECT 104.375 170.695 104.545 170.925 ;
        RECT 104.715 170.865 104.905 171.305 ;
        RECT 105.075 170.855 106.025 171.135 ;
        RECT 106.245 170.945 106.595 171.115 ;
        RECT 104.375 170.525 104.905 170.695 ;
        RECT 102.880 170.065 103.620 170.095 ;
        RECT 100.715 168.755 100.925 169.895 ;
        RECT 101.095 168.925 101.425 169.905 ;
        RECT 101.595 168.755 101.825 169.895 ;
        RECT 102.500 169.065 102.755 169.945 ;
        RECT 102.925 168.755 103.230 169.895 ;
        RECT 103.450 169.475 103.620 170.065 ;
        RECT 103.965 169.985 104.505 170.355 ;
        RECT 104.685 170.245 104.905 170.525 ;
        RECT 105.075 170.075 105.245 170.855 ;
        RECT 104.840 169.905 105.245 170.075 ;
        RECT 105.415 170.065 105.765 170.685 ;
        RECT 104.840 169.815 105.010 169.905 ;
        RECT 105.935 169.895 106.145 170.685 ;
        RECT 103.790 169.645 105.010 169.815 ;
        RECT 105.470 169.735 106.145 169.895 ;
        RECT 103.450 169.305 104.250 169.475 ;
        RECT 103.570 168.755 103.900 169.135 ;
        RECT 104.080 169.015 104.250 169.305 ;
        RECT 104.840 169.265 105.010 169.645 ;
        RECT 105.180 169.725 106.145 169.735 ;
        RECT 106.335 170.555 106.595 170.945 ;
        RECT 106.805 170.845 107.135 171.305 ;
        RECT 108.010 170.915 108.865 171.085 ;
        RECT 109.070 170.915 109.565 171.085 ;
        RECT 109.735 170.945 110.065 171.305 ;
        RECT 106.335 169.865 106.505 170.555 ;
        RECT 106.675 170.205 106.845 170.385 ;
        RECT 107.015 170.375 107.805 170.625 ;
        RECT 108.010 170.205 108.180 170.915 ;
        RECT 108.350 170.405 108.705 170.625 ;
        RECT 106.675 170.035 108.365 170.205 ;
        RECT 105.180 169.435 105.640 169.725 ;
        RECT 106.335 169.695 107.835 169.865 ;
        RECT 106.335 169.555 106.505 169.695 ;
        RECT 105.945 169.385 106.505 169.555 ;
        RECT 104.420 168.755 104.670 169.215 ;
        RECT 104.840 168.925 105.710 169.265 ;
        RECT 105.945 168.925 106.115 169.385 ;
        RECT 106.950 169.355 108.025 169.525 ;
        RECT 106.285 168.755 106.655 169.215 ;
        RECT 106.950 169.015 107.120 169.355 ;
        RECT 107.290 168.755 107.620 169.185 ;
        RECT 107.855 169.015 108.025 169.355 ;
        RECT 108.195 169.255 108.365 170.035 ;
        RECT 108.535 169.815 108.705 170.405 ;
        RECT 108.875 170.005 109.225 170.625 ;
        RECT 108.535 169.425 109.000 169.815 ;
        RECT 109.395 169.555 109.565 170.915 ;
        RECT 109.735 169.725 110.195 170.775 ;
        RECT 109.170 169.385 109.565 169.555 ;
        RECT 109.170 169.255 109.340 169.385 ;
        RECT 108.195 168.925 108.875 169.255 ;
        RECT 109.090 168.925 109.340 169.255 ;
        RECT 109.510 168.755 109.760 169.215 ;
        RECT 109.930 168.940 110.255 169.725 ;
        RECT 110.425 168.925 110.595 171.045 ;
        RECT 110.765 170.925 111.095 171.305 ;
        RECT 111.265 170.755 111.520 171.045 ;
        RECT 110.770 170.585 111.520 170.755 ;
        RECT 110.770 169.595 111.000 170.585 ;
        RECT 112.155 170.555 113.365 171.305 ;
        RECT 111.170 169.765 111.520 170.415 ;
        RECT 112.155 169.845 112.675 170.385 ;
        RECT 112.845 170.015 113.365 170.555 ;
        RECT 110.770 169.425 111.520 169.595 ;
        RECT 110.765 168.755 111.095 169.255 ;
        RECT 111.265 168.925 111.520 169.425 ;
        RECT 112.155 168.755 113.365 169.845 ;
        RECT 11.330 168.585 113.450 168.755 ;
        RECT 11.415 167.495 12.625 168.585 ;
        RECT 11.415 166.785 11.935 167.325 ;
        RECT 12.105 166.955 12.625 167.495 ;
        RECT 13.345 167.655 13.515 168.415 ;
        RECT 13.695 167.825 14.025 168.585 ;
        RECT 13.345 167.485 14.010 167.655 ;
        RECT 14.195 167.510 14.465 168.415 ;
        RECT 13.840 167.340 14.010 167.485 ;
        RECT 13.275 166.935 13.605 167.305 ;
        RECT 13.840 167.010 14.125 167.340 ;
        RECT 11.415 166.035 12.625 166.785 ;
        RECT 13.840 166.755 14.010 167.010 ;
        RECT 13.345 166.585 14.010 166.755 ;
        RECT 14.295 166.710 14.465 167.510 ;
        RECT 14.675 167.445 14.905 168.585 ;
        RECT 15.075 167.435 15.405 168.415 ;
        RECT 15.575 167.445 15.785 168.585 ;
        RECT 16.975 167.445 17.205 168.585 ;
        RECT 17.375 167.435 17.705 168.415 ;
        RECT 17.875 167.445 18.085 168.585 ;
        RECT 18.405 167.915 18.575 168.415 ;
        RECT 18.745 168.085 19.075 168.585 ;
        RECT 18.405 167.745 19.070 167.915 ;
        RECT 14.655 167.025 14.985 167.275 ;
        RECT 13.345 166.205 13.515 166.585 ;
        RECT 13.695 166.035 14.025 166.415 ;
        RECT 14.205 166.205 14.465 166.710 ;
        RECT 14.675 166.035 14.905 166.855 ;
        RECT 15.155 166.835 15.405 167.435 ;
        RECT 16.955 167.025 17.285 167.275 ;
        RECT 15.075 166.205 15.405 166.835 ;
        RECT 15.575 166.035 15.785 166.855 ;
        RECT 16.975 166.035 17.205 166.855 ;
        RECT 17.455 166.835 17.705 167.435 ;
        RECT 18.320 166.925 18.670 167.575 ;
        RECT 17.375 166.205 17.705 166.835 ;
        RECT 17.875 166.035 18.085 166.855 ;
        RECT 18.840 166.755 19.070 167.745 ;
        RECT 18.405 166.585 19.070 166.755 ;
        RECT 18.405 166.295 18.575 166.585 ;
        RECT 18.745 166.035 19.075 166.415 ;
        RECT 19.245 166.295 19.470 168.415 ;
        RECT 19.685 168.085 20.015 168.585 ;
        RECT 20.185 167.915 20.355 168.415 ;
        RECT 20.590 168.200 21.420 168.370 ;
        RECT 21.660 168.205 22.040 168.585 ;
        RECT 19.660 167.745 20.355 167.915 ;
        RECT 19.660 166.775 19.830 167.745 ;
        RECT 20.000 166.955 20.410 167.575 ;
        RECT 20.580 167.525 21.080 167.905 ;
        RECT 19.660 166.585 20.355 166.775 ;
        RECT 20.580 166.655 20.800 167.525 ;
        RECT 21.250 167.355 21.420 168.200 ;
        RECT 22.220 168.035 22.390 168.325 ;
        RECT 22.560 168.205 22.890 168.585 ;
        RECT 23.360 168.115 23.990 168.365 ;
        RECT 24.170 168.205 24.590 168.585 ;
        RECT 23.820 168.035 23.990 168.115 ;
        RECT 24.790 168.035 25.030 168.325 ;
        RECT 21.590 167.785 22.960 168.035 ;
        RECT 21.590 167.525 21.840 167.785 ;
        RECT 22.350 167.355 22.600 167.515 ;
        RECT 21.250 167.185 22.600 167.355 ;
        RECT 21.250 167.145 21.670 167.185 ;
        RECT 20.980 166.595 21.330 166.965 ;
        RECT 19.685 166.035 20.015 166.415 ;
        RECT 20.185 166.255 20.355 166.585 ;
        RECT 21.500 166.415 21.670 167.145 ;
        RECT 22.770 167.015 22.960 167.785 ;
        RECT 21.840 166.685 22.250 167.015 ;
        RECT 22.540 166.675 22.960 167.015 ;
        RECT 23.130 167.605 23.650 167.915 ;
        RECT 23.820 167.865 25.030 168.035 ;
        RECT 25.260 167.895 25.590 168.585 ;
        RECT 23.130 166.845 23.300 167.605 ;
        RECT 23.470 167.015 23.650 167.425 ;
        RECT 23.820 167.355 23.990 167.865 ;
        RECT 25.760 167.715 25.930 168.325 ;
        RECT 26.200 167.865 26.530 168.375 ;
        RECT 25.760 167.695 26.080 167.715 ;
        RECT 24.160 167.525 26.080 167.695 ;
        RECT 23.820 167.185 25.720 167.355 ;
        RECT 24.050 166.845 24.380 166.965 ;
        RECT 23.130 166.675 24.380 166.845 ;
        RECT 20.655 166.215 21.670 166.415 ;
        RECT 21.840 166.035 22.250 166.475 ;
        RECT 22.540 166.245 22.790 166.675 ;
        RECT 22.990 166.035 23.310 166.495 ;
        RECT 24.550 166.425 24.720 167.185 ;
        RECT 25.390 167.125 25.720 167.185 ;
        RECT 24.910 166.955 25.240 167.015 ;
        RECT 24.910 166.685 25.570 166.955 ;
        RECT 25.890 166.630 26.080 167.525 ;
        RECT 23.870 166.255 24.720 166.425 ;
        RECT 24.920 166.035 25.580 166.515 ;
        RECT 25.760 166.300 26.080 166.630 ;
        RECT 26.280 167.275 26.530 167.865 ;
        RECT 26.710 167.785 26.995 168.585 ;
        RECT 27.175 167.605 27.430 168.275 ;
        RECT 27.250 167.565 27.430 167.605 ;
        RECT 27.250 167.395 27.515 167.565 ;
        RECT 28.435 167.495 31.945 168.585 ;
        RECT 26.280 166.945 27.080 167.275 ;
        RECT 26.280 166.295 26.530 166.945 ;
        RECT 27.250 166.745 27.430 167.395 ;
        RECT 28.435 166.975 30.125 167.495 ;
        RECT 32.115 167.445 32.455 168.415 ;
        RECT 32.625 167.445 32.795 168.585 ;
        RECT 33.065 167.785 33.315 168.585 ;
        RECT 33.960 167.615 34.290 168.415 ;
        RECT 34.590 167.785 34.920 168.585 ;
        RECT 35.090 167.615 35.420 168.415 ;
        RECT 32.985 167.445 35.420 167.615 ;
        RECT 30.295 166.805 31.945 167.325 ;
        RECT 26.710 166.035 26.995 166.495 ;
        RECT 27.175 166.215 27.430 166.745 ;
        RECT 28.435 166.035 31.945 166.805 ;
        RECT 32.115 166.885 32.290 167.445 ;
        RECT 32.985 167.195 33.155 167.445 ;
        RECT 32.460 167.025 33.155 167.195 ;
        RECT 33.330 167.025 33.750 167.225 ;
        RECT 33.920 167.025 34.250 167.225 ;
        RECT 34.420 167.025 34.750 167.225 ;
        RECT 32.115 166.835 32.345 166.885 ;
        RECT 32.115 166.205 32.455 166.835 ;
        RECT 32.625 166.035 32.875 166.835 ;
        RECT 33.065 166.685 34.290 166.855 ;
        RECT 33.065 166.205 33.395 166.685 ;
        RECT 33.565 166.035 33.790 166.495 ;
        RECT 33.960 166.205 34.290 166.685 ;
        RECT 34.920 166.815 35.090 167.445 ;
        RECT 35.795 167.420 36.085 168.585 ;
        RECT 36.770 167.715 37.055 168.585 ;
        RECT 37.225 167.955 37.485 168.415 ;
        RECT 37.660 168.125 37.915 168.585 ;
        RECT 38.085 167.955 38.345 168.415 ;
        RECT 37.225 167.785 38.345 167.955 ;
        RECT 38.515 167.785 38.825 168.585 ;
        RECT 37.225 167.535 37.485 167.785 ;
        RECT 38.995 167.615 39.305 168.415 ;
        RECT 39.725 167.855 40.020 168.585 ;
        RECT 40.190 167.685 40.450 168.410 ;
        RECT 40.620 167.855 40.880 168.585 ;
        RECT 41.050 167.685 41.310 168.410 ;
        RECT 41.480 167.855 41.740 168.585 ;
        RECT 41.910 167.685 42.170 168.410 ;
        RECT 42.340 167.855 42.600 168.585 ;
        RECT 42.770 167.685 43.030 168.410 ;
        RECT 36.730 167.365 37.485 167.535 ;
        RECT 38.275 167.445 39.305 167.615 ;
        RECT 35.275 167.025 35.625 167.275 ;
        RECT 36.730 166.855 37.135 167.365 ;
        RECT 38.275 167.195 38.445 167.445 ;
        RECT 37.305 167.025 38.445 167.195 ;
        RECT 34.920 166.205 35.420 166.815 ;
        RECT 35.795 166.035 36.085 166.760 ;
        RECT 36.730 166.685 38.380 166.855 ;
        RECT 38.615 166.705 38.965 167.275 ;
        RECT 36.775 166.035 37.055 166.515 ;
        RECT 37.225 166.295 37.485 166.685 ;
        RECT 37.660 166.035 37.915 166.515 ;
        RECT 38.085 166.295 38.380 166.685 ;
        RECT 39.135 166.535 39.305 167.445 ;
        RECT 39.720 167.445 43.030 167.685 ;
        RECT 43.200 167.475 43.460 168.585 ;
        RECT 39.720 166.855 40.690 167.445 ;
        RECT 43.630 167.275 43.880 168.410 ;
        RECT 44.060 167.475 44.355 168.585 ;
        RECT 44.535 167.495 45.745 168.585 ;
        RECT 40.860 167.025 43.880 167.275 ;
        RECT 39.720 166.685 43.030 166.855 ;
        RECT 38.560 166.035 38.835 166.515 ;
        RECT 39.005 166.205 39.305 166.535 ;
        RECT 39.720 166.035 40.020 166.515 ;
        RECT 40.190 166.230 40.450 166.685 ;
        RECT 40.620 166.035 40.880 166.515 ;
        RECT 41.050 166.230 41.310 166.685 ;
        RECT 41.480 166.035 41.740 166.515 ;
        RECT 41.910 166.230 42.170 166.685 ;
        RECT 42.340 166.035 42.600 166.515 ;
        RECT 42.770 166.230 43.030 166.685 ;
        RECT 43.200 166.035 43.460 166.560 ;
        RECT 43.630 166.215 43.880 167.025 ;
        RECT 44.050 166.665 44.365 167.275 ;
        RECT 44.535 166.955 45.055 167.495 ;
        RECT 45.915 167.445 46.300 168.415 ;
        RECT 46.470 168.125 46.795 168.585 ;
        RECT 47.315 167.955 47.595 168.415 ;
        RECT 46.470 167.735 47.595 167.955 ;
        RECT 45.225 166.785 45.745 167.325 ;
        RECT 44.060 166.035 44.305 166.495 ;
        RECT 44.535 166.035 45.745 166.785 ;
        RECT 45.915 166.775 46.195 167.445 ;
        RECT 46.470 167.275 46.920 167.735 ;
        RECT 47.785 167.565 48.185 168.415 ;
        RECT 48.585 168.125 48.855 168.585 ;
        RECT 49.025 167.955 49.310 168.415 ;
        RECT 46.365 166.945 46.920 167.275 ;
        RECT 47.090 167.005 48.185 167.565 ;
        RECT 46.470 166.835 46.920 166.945 ;
        RECT 45.915 166.205 46.300 166.775 ;
        RECT 46.470 166.665 47.595 166.835 ;
        RECT 46.470 166.035 46.795 166.495 ;
        RECT 47.315 166.205 47.595 166.665 ;
        RECT 47.785 166.205 48.185 167.005 ;
        RECT 48.355 167.735 49.310 167.955 ;
        RECT 48.355 166.835 48.565 167.735 ;
        RECT 48.735 167.005 49.425 167.565 ;
        RECT 50.055 167.495 51.725 168.585 ;
        RECT 50.055 166.975 50.805 167.495 ;
        RECT 52.045 167.435 52.375 168.585 ;
        RECT 52.545 167.565 52.715 168.415 ;
        RECT 52.885 167.785 53.215 168.585 ;
        RECT 53.385 167.565 53.555 168.415 ;
        RECT 53.735 167.785 53.975 168.585 ;
        RECT 54.145 167.605 54.475 168.415 ;
        RECT 52.545 167.395 53.555 167.565 ;
        RECT 53.760 167.435 54.475 167.605 ;
        RECT 54.805 167.435 55.135 168.585 ;
        RECT 55.305 167.565 55.475 168.415 ;
        RECT 55.645 167.785 55.975 168.585 ;
        RECT 56.145 167.565 56.315 168.415 ;
        RECT 56.495 167.785 56.735 168.585 ;
        RECT 56.905 167.605 57.235 168.415 ;
        RECT 48.355 166.665 49.310 166.835 ;
        RECT 50.975 166.805 51.725 167.325 ;
        RECT 52.545 167.225 53.040 167.395 ;
        RECT 52.545 167.055 53.045 167.225 ;
        RECT 53.760 167.195 53.930 167.435 ;
        RECT 55.305 167.395 56.315 167.565 ;
        RECT 56.520 167.435 57.235 167.605 ;
        RECT 57.875 167.495 59.545 168.585 ;
        RECT 52.545 166.855 53.040 167.055 ;
        RECT 53.430 167.025 53.930 167.195 ;
        RECT 54.100 167.025 54.480 167.265 ;
        RECT 53.760 166.855 53.930 167.025 ;
        RECT 55.305 166.855 55.800 167.395 ;
        RECT 56.520 167.195 56.690 167.435 ;
        RECT 56.190 167.025 56.690 167.195 ;
        RECT 56.860 167.025 57.240 167.265 ;
        RECT 56.520 166.855 56.690 167.025 ;
        RECT 57.875 166.975 58.625 167.495 ;
        RECT 59.720 167.435 59.980 168.585 ;
        RECT 60.155 167.510 60.410 168.415 ;
        RECT 60.580 167.825 60.910 168.585 ;
        RECT 61.125 167.655 61.295 168.415 ;
        RECT 48.585 166.035 48.855 166.495 ;
        RECT 49.025 166.205 49.310 166.665 ;
        RECT 50.055 166.035 51.725 166.805 ;
        RECT 52.045 166.035 52.375 166.835 ;
        RECT 52.545 166.685 53.555 166.855 ;
        RECT 53.760 166.685 54.395 166.855 ;
        RECT 52.545 166.205 52.715 166.685 ;
        RECT 52.885 166.035 53.215 166.515 ;
        RECT 53.385 166.205 53.555 166.685 ;
        RECT 53.805 166.035 54.045 166.515 ;
        RECT 54.225 166.205 54.395 166.685 ;
        RECT 54.805 166.035 55.135 166.835 ;
        RECT 55.305 166.685 56.315 166.855 ;
        RECT 56.520 166.685 57.155 166.855 ;
        RECT 58.795 166.805 59.545 167.325 ;
        RECT 55.305 166.205 55.475 166.685 ;
        RECT 55.645 166.035 55.975 166.515 ;
        RECT 56.145 166.205 56.315 166.685 ;
        RECT 56.565 166.035 56.805 166.515 ;
        RECT 56.985 166.205 57.155 166.685 ;
        RECT 57.875 166.035 59.545 166.805 ;
        RECT 59.720 166.035 59.980 166.875 ;
        RECT 60.155 166.780 60.325 167.510 ;
        RECT 60.580 167.485 61.295 167.655 ;
        RECT 60.580 167.275 60.750 167.485 ;
        RECT 61.555 167.420 61.845 168.585 ;
        RECT 62.945 167.525 63.275 168.585 ;
        RECT 60.495 166.945 60.750 167.275 ;
        RECT 60.155 166.205 60.410 166.780 ;
        RECT 60.580 166.755 60.750 166.945 ;
        RECT 61.030 166.935 61.385 167.305 ;
        RECT 63.455 167.275 63.625 168.200 ;
        RECT 63.795 167.995 64.125 168.395 ;
        RECT 64.295 168.225 64.625 168.585 ;
        RECT 64.825 167.995 65.525 168.415 ;
        RECT 63.795 167.765 65.525 167.995 ;
        RECT 63.795 167.545 64.125 167.765 ;
        RECT 64.320 167.275 64.645 167.565 ;
        RECT 62.935 166.945 63.245 167.275 ;
        RECT 63.455 166.945 63.830 167.275 ;
        RECT 64.150 166.945 64.645 167.275 ;
        RECT 64.820 167.025 65.150 167.565 ;
        RECT 65.320 166.885 65.525 167.765 ;
        RECT 65.695 167.495 69.205 168.585 ;
        RECT 69.465 167.655 69.635 168.415 ;
        RECT 69.815 167.825 70.145 168.585 ;
        RECT 65.695 166.975 67.385 167.495 ;
        RECT 69.465 167.485 70.130 167.655 ;
        RECT 70.315 167.510 70.585 168.415 ;
        RECT 70.845 167.915 71.015 168.415 ;
        RECT 71.185 168.085 71.515 168.585 ;
        RECT 70.845 167.745 71.510 167.915 ;
        RECT 69.960 167.340 70.130 167.485 ;
        RECT 65.295 166.795 65.525 166.885 ;
        RECT 67.555 166.805 69.205 167.325 ;
        RECT 69.395 166.935 69.725 167.305 ;
        RECT 69.960 167.010 70.245 167.340 ;
        RECT 60.580 166.585 61.295 166.755 ;
        RECT 60.580 166.035 60.910 166.415 ;
        RECT 61.125 166.205 61.295 166.585 ;
        RECT 61.555 166.035 61.845 166.760 ;
        RECT 62.945 166.565 64.305 166.775 ;
        RECT 62.945 166.205 63.275 166.565 ;
        RECT 63.445 166.035 63.775 166.395 ;
        RECT 63.975 166.205 64.305 166.565 ;
        RECT 64.815 166.205 65.525 166.795 ;
        RECT 65.695 166.035 69.205 166.805 ;
        RECT 69.960 166.755 70.130 167.010 ;
        RECT 69.465 166.585 70.130 166.755 ;
        RECT 70.415 166.710 70.585 167.510 ;
        RECT 70.760 166.925 71.110 167.575 ;
        RECT 71.280 166.755 71.510 167.745 ;
        RECT 69.465 166.205 69.635 166.585 ;
        RECT 69.815 166.035 70.145 166.415 ;
        RECT 70.325 166.205 70.585 166.710 ;
        RECT 70.845 166.585 71.510 166.755 ;
        RECT 70.845 166.295 71.015 166.585 ;
        RECT 71.185 166.035 71.515 166.415 ;
        RECT 71.685 166.295 71.910 168.415 ;
        RECT 72.125 168.085 72.455 168.585 ;
        RECT 72.625 167.915 72.795 168.415 ;
        RECT 73.030 168.200 73.860 168.370 ;
        RECT 74.100 168.205 74.480 168.585 ;
        RECT 72.100 167.745 72.795 167.915 ;
        RECT 72.100 166.775 72.270 167.745 ;
        RECT 72.440 166.955 72.850 167.575 ;
        RECT 73.020 167.525 73.520 167.905 ;
        RECT 72.100 166.585 72.795 166.775 ;
        RECT 73.020 166.655 73.240 167.525 ;
        RECT 73.690 167.355 73.860 168.200 ;
        RECT 74.660 168.035 74.830 168.325 ;
        RECT 75.000 168.205 75.330 168.585 ;
        RECT 75.800 168.115 76.430 168.365 ;
        RECT 76.610 168.205 77.030 168.585 ;
        RECT 76.260 168.035 76.430 168.115 ;
        RECT 77.230 168.035 77.470 168.325 ;
        RECT 74.030 167.785 75.400 168.035 ;
        RECT 74.030 167.525 74.280 167.785 ;
        RECT 74.790 167.355 75.040 167.515 ;
        RECT 73.690 167.185 75.040 167.355 ;
        RECT 73.690 167.145 74.110 167.185 ;
        RECT 73.420 166.595 73.770 166.965 ;
        RECT 72.125 166.035 72.455 166.415 ;
        RECT 72.625 166.255 72.795 166.585 ;
        RECT 73.940 166.415 74.110 167.145 ;
        RECT 75.210 167.015 75.400 167.785 ;
        RECT 74.280 166.685 74.690 167.015 ;
        RECT 74.980 166.675 75.400 167.015 ;
        RECT 75.570 167.605 76.090 167.915 ;
        RECT 76.260 167.865 77.470 168.035 ;
        RECT 77.700 167.895 78.030 168.585 ;
        RECT 75.570 166.845 75.740 167.605 ;
        RECT 75.910 167.015 76.090 167.425 ;
        RECT 76.260 167.355 76.430 167.865 ;
        RECT 78.200 167.715 78.370 168.325 ;
        RECT 78.640 167.865 78.970 168.375 ;
        RECT 78.200 167.695 78.520 167.715 ;
        RECT 76.600 167.525 78.520 167.695 ;
        RECT 76.260 167.185 78.160 167.355 ;
        RECT 76.490 166.845 76.820 166.965 ;
        RECT 75.570 166.675 76.820 166.845 ;
        RECT 73.095 166.215 74.110 166.415 ;
        RECT 74.280 166.035 74.690 166.475 ;
        RECT 74.980 166.245 75.230 166.675 ;
        RECT 75.430 166.035 75.750 166.495 ;
        RECT 76.990 166.425 77.160 167.185 ;
        RECT 77.830 167.125 78.160 167.185 ;
        RECT 77.350 166.955 77.680 167.015 ;
        RECT 77.350 166.685 78.010 166.955 ;
        RECT 78.330 166.630 78.520 167.525 ;
        RECT 76.310 166.255 77.160 166.425 ;
        RECT 77.360 166.035 78.020 166.515 ;
        RECT 78.200 166.300 78.520 166.630 ;
        RECT 78.720 167.275 78.970 167.865 ;
        RECT 79.150 167.785 79.435 168.585 ;
        RECT 79.615 167.605 79.870 168.275 ;
        RECT 80.665 167.855 80.960 168.585 ;
        RECT 81.130 167.685 81.390 168.410 ;
        RECT 81.560 167.855 81.820 168.585 ;
        RECT 81.990 167.685 82.250 168.410 ;
        RECT 82.420 167.855 82.680 168.585 ;
        RECT 82.850 167.685 83.110 168.410 ;
        RECT 83.280 167.855 83.540 168.585 ;
        RECT 83.710 167.685 83.970 168.410 ;
        RECT 78.720 166.945 79.520 167.275 ;
        RECT 78.720 166.295 78.970 166.945 ;
        RECT 79.690 166.745 79.870 167.605 ;
        RECT 79.615 166.545 79.870 166.745 ;
        RECT 80.660 167.445 83.970 167.685 ;
        RECT 84.140 167.475 84.400 168.585 ;
        RECT 80.660 166.855 81.630 167.445 ;
        RECT 84.570 167.275 84.820 168.410 ;
        RECT 85.000 167.475 85.295 168.585 ;
        RECT 85.475 167.510 85.745 168.415 ;
        RECT 85.915 167.825 86.245 168.585 ;
        RECT 86.425 167.655 86.595 168.415 ;
        RECT 81.800 167.025 84.820 167.275 ;
        RECT 80.660 166.685 83.970 166.855 ;
        RECT 79.150 166.035 79.435 166.495 ;
        RECT 79.615 166.375 79.955 166.545 ;
        RECT 79.615 166.215 79.870 166.375 ;
        RECT 80.660 166.035 80.960 166.515 ;
        RECT 81.130 166.230 81.390 166.685 ;
        RECT 81.560 166.035 81.820 166.515 ;
        RECT 81.990 166.230 82.250 166.685 ;
        RECT 82.420 166.035 82.680 166.515 ;
        RECT 82.850 166.230 83.110 166.685 ;
        RECT 83.280 166.035 83.540 166.515 ;
        RECT 83.710 166.230 83.970 166.685 ;
        RECT 84.140 166.035 84.400 166.560 ;
        RECT 84.570 166.215 84.820 167.025 ;
        RECT 84.990 166.665 85.305 167.275 ;
        RECT 85.475 166.710 85.645 167.510 ;
        RECT 85.930 167.485 86.595 167.655 ;
        RECT 85.930 167.340 86.100 167.485 ;
        RECT 87.315 167.420 87.605 168.585 ;
        RECT 87.785 167.775 88.080 168.585 ;
        RECT 85.815 167.010 86.100 167.340 ;
        RECT 85.930 166.755 86.100 167.010 ;
        RECT 86.335 166.935 86.665 167.305 ;
        RECT 88.260 167.275 88.505 168.415 ;
        RECT 88.680 167.775 88.940 168.585 ;
        RECT 89.540 168.580 95.815 168.585 ;
        RECT 89.120 167.275 89.370 168.410 ;
        RECT 89.540 167.785 89.800 168.580 ;
        RECT 89.970 167.685 90.230 168.410 ;
        RECT 90.400 167.855 90.660 168.580 ;
        RECT 90.830 167.685 91.090 168.410 ;
        RECT 91.260 167.855 91.520 168.580 ;
        RECT 91.690 167.685 91.950 168.410 ;
        RECT 92.120 167.855 92.380 168.580 ;
        RECT 92.550 167.685 92.810 168.410 ;
        RECT 92.980 167.855 93.225 168.580 ;
        RECT 93.395 167.685 93.655 168.410 ;
        RECT 93.840 167.855 94.085 168.580 ;
        RECT 94.255 167.685 94.515 168.410 ;
        RECT 94.700 167.855 94.945 168.580 ;
        RECT 95.115 167.685 95.375 168.410 ;
        RECT 95.560 167.855 95.815 168.580 ;
        RECT 89.970 167.670 95.375 167.685 ;
        RECT 95.985 167.670 96.275 168.410 ;
        RECT 96.445 167.840 96.715 168.585 ;
        RECT 89.970 167.565 96.715 167.670 ;
        RECT 89.970 167.445 96.745 167.565 ;
        RECT 95.550 167.395 96.745 167.445 ;
        RECT 97.440 167.395 97.695 168.275 ;
        RECT 97.865 167.445 98.170 168.585 ;
        RECT 98.510 168.205 98.840 168.585 ;
        RECT 99.020 168.035 99.190 168.325 ;
        RECT 99.360 168.125 99.610 168.585 ;
        RECT 98.390 167.865 99.190 168.035 ;
        RECT 99.780 168.075 100.650 168.415 ;
        RECT 85.000 166.035 85.245 166.495 ;
        RECT 85.475 166.205 85.735 166.710 ;
        RECT 85.930 166.585 86.595 166.755 ;
        RECT 85.915 166.035 86.245 166.415 ;
        RECT 86.425 166.205 86.595 166.585 ;
        RECT 87.315 166.035 87.605 166.760 ;
        RECT 87.775 166.715 88.090 167.275 ;
        RECT 88.260 167.025 95.380 167.275 ;
        RECT 87.775 166.035 88.080 166.545 ;
        RECT 88.260 166.215 88.510 167.025 ;
        RECT 88.680 166.035 88.940 166.560 ;
        RECT 89.120 166.215 89.370 167.025 ;
        RECT 95.550 166.855 96.715 167.395 ;
        RECT 89.970 166.685 96.715 166.855 ;
        RECT 97.440 166.745 97.650 167.395 ;
        RECT 98.390 167.275 98.560 167.865 ;
        RECT 99.780 167.695 99.950 168.075 ;
        RECT 100.885 167.955 101.055 168.415 ;
        RECT 101.225 168.125 101.595 168.585 ;
        RECT 101.890 167.985 102.060 168.325 ;
        RECT 102.230 168.155 102.560 168.585 ;
        RECT 102.795 167.985 102.965 168.325 ;
        RECT 98.730 167.525 99.950 167.695 ;
        RECT 100.120 167.615 100.580 167.905 ;
        RECT 100.885 167.785 101.445 167.955 ;
        RECT 101.890 167.815 102.965 167.985 ;
        RECT 103.135 168.085 103.815 168.415 ;
        RECT 104.030 168.085 104.280 168.415 ;
        RECT 104.450 168.125 104.700 168.585 ;
        RECT 101.275 167.645 101.445 167.785 ;
        RECT 100.120 167.605 101.085 167.615 ;
        RECT 99.780 167.435 99.950 167.525 ;
        RECT 100.410 167.445 101.085 167.605 ;
        RECT 97.820 167.245 98.560 167.275 ;
        RECT 97.820 166.945 98.735 167.245 ;
        RECT 98.410 166.770 98.735 166.945 ;
        RECT 89.540 166.035 89.800 166.595 ;
        RECT 89.970 166.230 90.230 166.685 ;
        RECT 90.400 166.035 90.660 166.515 ;
        RECT 90.830 166.230 91.090 166.685 ;
        RECT 91.260 166.035 91.520 166.515 ;
        RECT 91.690 166.230 91.950 166.685 ;
        RECT 92.120 166.035 92.365 166.515 ;
        RECT 92.535 166.230 92.810 166.685 ;
        RECT 92.980 166.035 93.225 166.515 ;
        RECT 93.395 166.230 93.655 166.685 ;
        RECT 93.835 166.035 94.085 166.515 ;
        RECT 94.255 166.230 94.515 166.685 ;
        RECT 94.695 166.035 94.945 166.515 ;
        RECT 95.115 166.230 95.375 166.685 ;
        RECT 95.555 166.035 95.815 166.515 ;
        RECT 95.985 166.230 96.245 166.685 ;
        RECT 96.415 166.035 96.715 166.515 ;
        RECT 97.440 166.215 97.695 166.745 ;
        RECT 97.865 166.035 98.170 166.495 ;
        RECT 98.415 166.415 98.735 166.770 ;
        RECT 98.905 166.985 99.445 167.355 ;
        RECT 99.780 167.265 100.185 167.435 ;
        RECT 98.905 166.585 99.145 166.985 ;
        RECT 99.625 166.815 99.845 167.095 ;
        RECT 99.315 166.645 99.845 166.815 ;
        RECT 99.315 166.415 99.485 166.645 ;
        RECT 100.015 166.485 100.185 167.265 ;
        RECT 100.355 166.655 100.705 167.275 ;
        RECT 100.875 166.655 101.085 167.445 ;
        RECT 101.275 167.475 102.775 167.645 ;
        RECT 101.275 166.785 101.445 167.475 ;
        RECT 103.135 167.305 103.305 168.085 ;
        RECT 104.110 167.955 104.280 168.085 ;
        RECT 101.615 167.135 103.305 167.305 ;
        RECT 103.475 167.525 103.940 167.915 ;
        RECT 104.110 167.785 104.505 167.955 ;
        RECT 101.615 166.955 101.785 167.135 ;
        RECT 98.415 166.245 99.485 166.415 ;
        RECT 99.655 166.035 99.845 166.475 ;
        RECT 100.015 166.205 100.965 166.485 ;
        RECT 101.275 166.395 101.535 166.785 ;
        RECT 101.955 166.715 102.745 166.965 ;
        RECT 101.185 166.225 101.535 166.395 ;
        RECT 101.745 166.035 102.075 166.495 ;
        RECT 102.950 166.425 103.120 167.135 ;
        RECT 103.475 166.935 103.645 167.525 ;
        RECT 103.290 166.715 103.645 166.935 ;
        RECT 103.815 166.715 104.165 167.335 ;
        RECT 104.335 166.425 104.505 167.785 ;
        RECT 104.870 167.615 105.195 168.400 ;
        RECT 104.675 166.565 105.135 167.615 ;
        RECT 102.950 166.255 103.805 166.425 ;
        RECT 104.010 166.255 104.505 166.425 ;
        RECT 104.675 166.035 105.005 166.395 ;
        RECT 105.365 166.295 105.535 168.415 ;
        RECT 105.705 168.085 106.035 168.585 ;
        RECT 106.205 167.915 106.460 168.415 ;
        RECT 105.710 167.745 106.460 167.915 ;
        RECT 105.710 166.755 105.940 167.745 ;
        RECT 106.110 166.925 106.460 167.575 ;
        RECT 106.675 167.445 106.905 168.585 ;
        RECT 107.075 167.435 107.405 168.415 ;
        RECT 107.575 167.445 107.785 168.585 ;
        RECT 108.020 168.160 108.355 168.585 ;
        RECT 108.525 167.980 108.710 168.385 ;
        RECT 108.045 167.805 108.710 167.980 ;
        RECT 108.915 167.805 109.245 168.585 ;
        RECT 106.655 167.025 106.985 167.275 ;
        RECT 105.710 166.585 106.460 166.755 ;
        RECT 105.705 166.035 106.035 166.415 ;
        RECT 106.205 166.295 106.460 166.585 ;
        RECT 106.675 166.035 106.905 166.855 ;
        RECT 107.155 166.835 107.405 167.435 ;
        RECT 107.075 166.205 107.405 166.835 ;
        RECT 107.575 166.035 107.785 166.855 ;
        RECT 108.045 166.775 108.385 167.805 ;
        RECT 109.415 167.615 109.685 168.385 ;
        RECT 108.555 167.445 109.685 167.615 ;
        RECT 108.555 166.945 108.805 167.445 ;
        RECT 108.045 166.605 108.730 166.775 ;
        RECT 108.985 166.695 109.345 167.275 ;
        RECT 108.020 166.035 108.355 166.435 ;
        RECT 108.525 166.205 108.730 166.605 ;
        RECT 109.515 166.535 109.685 167.445 ;
        RECT 108.940 166.035 109.215 166.515 ;
        RECT 109.425 166.205 109.685 166.535 ;
        RECT 109.855 167.510 110.125 168.415 ;
        RECT 110.295 167.825 110.625 168.585 ;
        RECT 110.805 167.655 110.975 168.415 ;
        RECT 109.855 166.710 110.025 167.510 ;
        RECT 110.310 167.485 110.975 167.655 ;
        RECT 112.155 167.495 113.365 168.585 ;
        RECT 110.310 167.340 110.480 167.485 ;
        RECT 110.195 167.010 110.480 167.340 ;
        RECT 110.310 166.755 110.480 167.010 ;
        RECT 110.715 166.935 111.045 167.305 ;
        RECT 112.155 166.955 112.675 167.495 ;
        RECT 112.845 166.785 113.365 167.325 ;
        RECT 109.855 166.205 110.115 166.710 ;
        RECT 110.310 166.585 110.975 166.755 ;
        RECT 110.295 166.035 110.625 166.415 ;
        RECT 110.805 166.205 110.975 166.585 ;
        RECT 112.155 166.035 113.365 166.785 ;
        RECT 11.330 165.865 113.450 166.035 ;
        RECT 11.415 165.115 12.625 165.865 ;
        RECT 12.885 165.315 13.055 165.605 ;
        RECT 13.225 165.485 13.555 165.865 ;
        RECT 12.885 165.145 13.550 165.315 ;
        RECT 11.415 164.575 11.935 165.115 ;
        RECT 12.105 164.405 12.625 164.945 ;
        RECT 11.415 163.315 12.625 164.405 ;
        RECT 12.800 164.325 13.150 164.975 ;
        RECT 13.320 164.155 13.550 165.145 ;
        RECT 12.885 163.985 13.550 164.155 ;
        RECT 12.885 163.485 13.055 163.985 ;
        RECT 13.225 163.315 13.555 163.815 ;
        RECT 13.725 163.485 13.950 165.605 ;
        RECT 14.165 165.485 14.495 165.865 ;
        RECT 14.665 165.315 14.835 165.645 ;
        RECT 15.135 165.485 16.150 165.685 ;
        RECT 14.140 165.125 14.835 165.315 ;
        RECT 14.140 164.155 14.310 165.125 ;
        RECT 14.480 164.325 14.890 164.945 ;
        RECT 15.060 164.375 15.280 165.245 ;
        RECT 15.460 164.935 15.810 165.305 ;
        RECT 15.980 164.755 16.150 165.485 ;
        RECT 16.320 165.425 16.730 165.865 ;
        RECT 17.020 165.225 17.270 165.655 ;
        RECT 17.470 165.405 17.790 165.865 ;
        RECT 18.350 165.475 19.200 165.645 ;
        RECT 16.320 164.885 16.730 165.215 ;
        RECT 17.020 164.885 17.440 165.225 ;
        RECT 15.730 164.715 16.150 164.755 ;
        RECT 15.730 164.545 17.080 164.715 ;
        RECT 14.140 163.985 14.835 164.155 ;
        RECT 15.060 163.995 15.560 164.375 ;
        RECT 14.165 163.315 14.495 163.815 ;
        RECT 14.665 163.485 14.835 163.985 ;
        RECT 15.730 163.700 15.900 164.545 ;
        RECT 16.830 164.385 17.080 164.545 ;
        RECT 16.070 164.115 16.320 164.375 ;
        RECT 17.250 164.115 17.440 164.885 ;
        RECT 16.070 163.865 17.440 164.115 ;
        RECT 17.610 165.055 18.860 165.225 ;
        RECT 17.610 164.295 17.780 165.055 ;
        RECT 18.530 164.935 18.860 165.055 ;
        RECT 17.950 164.475 18.130 164.885 ;
        RECT 19.030 164.715 19.200 165.475 ;
        RECT 19.400 165.385 20.060 165.865 ;
        RECT 20.240 165.270 20.560 165.600 ;
        RECT 19.390 164.945 20.050 165.215 ;
        RECT 19.390 164.885 19.720 164.945 ;
        RECT 19.870 164.715 20.200 164.775 ;
        RECT 18.300 164.545 20.200 164.715 ;
        RECT 17.610 163.985 18.130 164.295 ;
        RECT 18.300 164.035 18.470 164.545 ;
        RECT 20.370 164.375 20.560 165.270 ;
        RECT 18.640 164.205 20.560 164.375 ;
        RECT 20.240 164.185 20.560 164.205 ;
        RECT 20.760 164.955 21.010 165.605 ;
        RECT 21.190 165.405 21.475 165.865 ;
        RECT 21.655 165.525 21.910 165.685 ;
        RECT 21.655 165.355 21.995 165.525 ;
        RECT 21.655 165.155 21.910 165.355 ;
        RECT 20.760 164.625 21.560 164.955 ;
        RECT 18.300 163.865 19.510 164.035 ;
        RECT 15.070 163.530 15.900 163.700 ;
        RECT 16.140 163.315 16.520 163.695 ;
        RECT 16.700 163.575 16.870 163.865 ;
        RECT 18.300 163.785 18.470 163.865 ;
        RECT 17.040 163.315 17.370 163.695 ;
        RECT 17.840 163.535 18.470 163.785 ;
        RECT 18.650 163.315 19.070 163.695 ;
        RECT 19.270 163.575 19.510 163.865 ;
        RECT 19.740 163.315 20.070 164.005 ;
        RECT 20.240 163.575 20.410 164.185 ;
        RECT 20.760 164.035 21.010 164.625 ;
        RECT 21.730 164.295 21.910 165.155 ;
        RECT 22.915 165.140 23.205 165.865 ;
        RECT 23.835 165.190 24.095 165.695 ;
        RECT 24.275 165.485 24.605 165.865 ;
        RECT 24.785 165.315 24.955 165.695 ;
        RECT 20.680 163.525 21.010 164.035 ;
        RECT 21.190 163.315 21.475 164.115 ;
        RECT 21.655 163.625 21.910 164.295 ;
        RECT 22.915 163.315 23.205 164.480 ;
        RECT 23.835 164.390 24.005 165.190 ;
        RECT 24.290 165.145 24.955 165.315 ;
        RECT 24.290 164.890 24.460 165.145 ;
        RECT 25.220 165.125 25.475 165.695 ;
        RECT 25.645 165.465 25.975 165.865 ;
        RECT 26.400 165.330 26.930 165.695 ;
        RECT 26.400 165.295 26.575 165.330 ;
        RECT 25.645 165.125 26.575 165.295 ;
        RECT 24.175 164.560 24.460 164.890 ;
        RECT 24.695 164.595 25.025 164.965 ;
        RECT 24.290 164.415 24.460 164.560 ;
        RECT 25.220 164.455 25.390 165.125 ;
        RECT 25.645 164.955 25.815 165.125 ;
        RECT 25.560 164.625 25.815 164.955 ;
        RECT 26.040 164.625 26.235 164.955 ;
        RECT 23.835 163.485 24.105 164.390 ;
        RECT 24.290 164.245 24.955 164.415 ;
        RECT 24.275 163.315 24.605 164.075 ;
        RECT 24.785 163.485 24.955 164.245 ;
        RECT 25.220 163.485 25.555 164.455 ;
        RECT 25.725 163.315 25.895 164.455 ;
        RECT 26.065 163.655 26.235 164.625 ;
        RECT 26.405 163.995 26.575 165.125 ;
        RECT 26.745 164.335 26.915 165.135 ;
        RECT 27.120 164.845 27.395 165.695 ;
        RECT 27.115 164.675 27.395 164.845 ;
        RECT 27.120 164.535 27.395 164.675 ;
        RECT 27.565 164.335 27.755 165.695 ;
        RECT 27.935 165.330 28.445 165.865 ;
        RECT 28.665 165.055 28.910 165.660 ;
        RECT 29.355 165.355 29.660 165.865 ;
        RECT 27.955 164.885 29.185 165.055 ;
        RECT 26.745 164.165 27.755 164.335 ;
        RECT 27.925 164.320 28.675 164.510 ;
        RECT 26.405 163.825 27.530 163.995 ;
        RECT 27.925 163.655 28.095 164.320 ;
        RECT 28.845 164.075 29.185 164.885 ;
        RECT 29.355 164.625 29.670 165.185 ;
        RECT 29.840 164.875 30.090 165.685 ;
        RECT 30.260 165.340 30.520 165.865 ;
        RECT 30.700 164.875 30.950 165.685 ;
        RECT 31.120 165.305 31.380 165.865 ;
        RECT 31.550 165.215 31.810 165.670 ;
        RECT 31.980 165.385 32.240 165.865 ;
        RECT 32.410 165.215 32.670 165.670 ;
        RECT 32.840 165.385 33.100 165.865 ;
        RECT 33.270 165.215 33.530 165.670 ;
        RECT 33.700 165.385 33.945 165.865 ;
        RECT 34.115 165.215 34.390 165.670 ;
        RECT 34.560 165.385 34.805 165.865 ;
        RECT 34.975 165.215 35.235 165.670 ;
        RECT 35.415 165.385 35.665 165.865 ;
        RECT 35.835 165.215 36.095 165.670 ;
        RECT 36.275 165.385 36.525 165.865 ;
        RECT 36.695 165.215 36.955 165.670 ;
        RECT 37.135 165.385 37.395 165.865 ;
        RECT 37.565 165.215 37.825 165.670 ;
        RECT 37.995 165.385 38.295 165.865 ;
        RECT 31.550 165.045 38.295 165.215 ;
        RECT 29.840 164.625 36.960 164.875 ;
        RECT 26.065 163.485 28.095 163.655 ;
        RECT 28.265 163.315 28.435 164.075 ;
        RECT 28.670 163.665 29.185 164.075 ;
        RECT 29.365 163.315 29.660 164.125 ;
        RECT 29.840 163.485 30.085 164.625 ;
        RECT 30.260 163.315 30.520 164.125 ;
        RECT 30.700 163.490 30.950 164.625 ;
        RECT 37.130 164.455 38.295 165.045 ;
        RECT 31.550 164.230 38.295 164.455 ;
        RECT 38.560 165.155 38.815 165.685 ;
        RECT 38.985 165.405 39.290 165.865 ;
        RECT 39.535 165.485 40.605 165.655 ;
        RECT 38.560 164.505 38.770 165.155 ;
        RECT 39.535 165.130 39.855 165.485 ;
        RECT 39.530 164.955 39.855 165.130 ;
        RECT 38.940 164.655 39.855 164.955 ;
        RECT 40.025 164.915 40.265 165.315 ;
        RECT 40.435 165.255 40.605 165.485 ;
        RECT 40.775 165.425 40.965 165.865 ;
        RECT 41.135 165.415 42.085 165.695 ;
        RECT 42.305 165.505 42.655 165.675 ;
        RECT 40.435 165.085 40.965 165.255 ;
        RECT 38.940 164.625 39.680 164.655 ;
        RECT 31.550 164.215 36.955 164.230 ;
        RECT 31.120 163.320 31.380 164.115 ;
        RECT 31.550 163.490 31.810 164.215 ;
        RECT 31.980 163.320 32.240 164.045 ;
        RECT 32.410 163.490 32.670 164.215 ;
        RECT 32.840 163.320 33.100 164.045 ;
        RECT 33.270 163.490 33.530 164.215 ;
        RECT 33.700 163.320 33.960 164.045 ;
        RECT 34.130 163.490 34.390 164.215 ;
        RECT 34.560 163.320 34.805 164.045 ;
        RECT 34.975 163.490 35.235 164.215 ;
        RECT 35.420 163.320 35.665 164.045 ;
        RECT 35.835 163.490 36.095 164.215 ;
        RECT 36.280 163.320 36.525 164.045 ;
        RECT 36.695 163.490 36.955 164.215 ;
        RECT 37.140 163.320 37.395 164.045 ;
        RECT 37.565 163.490 37.855 164.230 ;
        RECT 31.120 163.315 37.395 163.320 ;
        RECT 38.025 163.315 38.295 164.060 ;
        RECT 38.560 163.625 38.815 164.505 ;
        RECT 38.985 163.315 39.290 164.455 ;
        RECT 39.510 164.035 39.680 164.625 ;
        RECT 40.025 164.545 40.565 164.915 ;
        RECT 40.745 164.805 40.965 165.085 ;
        RECT 41.135 164.635 41.305 165.415 ;
        RECT 40.900 164.465 41.305 164.635 ;
        RECT 41.475 164.625 41.825 165.245 ;
        RECT 40.900 164.375 41.070 164.465 ;
        RECT 41.995 164.455 42.205 165.245 ;
        RECT 39.850 164.205 41.070 164.375 ;
        RECT 41.530 164.295 42.205 164.455 ;
        RECT 39.510 163.865 40.310 164.035 ;
        RECT 39.630 163.315 39.960 163.695 ;
        RECT 40.140 163.575 40.310 163.865 ;
        RECT 40.900 163.825 41.070 164.205 ;
        RECT 41.240 164.285 42.205 164.295 ;
        RECT 42.395 165.115 42.655 165.505 ;
        RECT 42.865 165.405 43.195 165.865 ;
        RECT 44.070 165.475 44.925 165.645 ;
        RECT 45.130 165.475 45.625 165.645 ;
        RECT 45.795 165.505 46.125 165.865 ;
        RECT 42.395 164.425 42.565 165.115 ;
        RECT 42.735 164.765 42.905 164.945 ;
        RECT 43.075 164.935 43.865 165.185 ;
        RECT 44.070 164.765 44.240 165.475 ;
        RECT 44.410 164.965 44.765 165.185 ;
        RECT 42.735 164.595 44.425 164.765 ;
        RECT 41.240 163.995 41.700 164.285 ;
        RECT 42.395 164.255 43.895 164.425 ;
        RECT 42.395 164.115 42.565 164.255 ;
        RECT 42.005 163.945 42.565 164.115 ;
        RECT 40.480 163.315 40.730 163.775 ;
        RECT 40.900 163.485 41.770 163.825 ;
        RECT 42.005 163.485 42.175 163.945 ;
        RECT 43.010 163.915 44.085 164.085 ;
        RECT 42.345 163.315 42.715 163.775 ;
        RECT 43.010 163.575 43.180 163.915 ;
        RECT 43.350 163.315 43.680 163.745 ;
        RECT 43.915 163.575 44.085 163.915 ;
        RECT 44.255 163.815 44.425 164.595 ;
        RECT 44.595 164.375 44.765 164.965 ;
        RECT 44.935 164.565 45.285 165.185 ;
        RECT 44.595 163.985 45.060 164.375 ;
        RECT 45.455 164.115 45.625 165.475 ;
        RECT 45.795 164.285 46.255 165.335 ;
        RECT 45.230 163.945 45.625 164.115 ;
        RECT 45.230 163.815 45.400 163.945 ;
        RECT 44.255 163.485 44.935 163.815 ;
        RECT 45.150 163.485 45.400 163.815 ;
        RECT 45.570 163.315 45.820 163.775 ;
        RECT 45.990 163.500 46.315 164.285 ;
        RECT 46.485 163.485 46.655 165.605 ;
        RECT 46.825 165.485 47.155 165.865 ;
        RECT 47.325 165.315 47.580 165.605 ;
        RECT 46.830 165.145 47.580 165.315 ;
        RECT 46.830 164.155 47.060 165.145 ;
        RECT 48.675 165.140 48.965 165.865 ;
        RECT 49.135 165.115 50.345 165.865 ;
        RECT 47.230 164.325 47.580 164.975 ;
        RECT 46.830 163.985 47.580 164.155 ;
        RECT 46.825 163.315 47.155 163.815 ;
        RECT 47.325 163.485 47.580 163.985 ;
        RECT 48.675 163.315 48.965 164.480 ;
        RECT 49.135 164.405 49.655 164.945 ;
        RECT 49.825 164.575 50.345 165.115 ;
        RECT 50.665 165.065 50.995 165.865 ;
        RECT 51.165 165.215 51.335 165.695 ;
        RECT 51.505 165.385 51.835 165.865 ;
        RECT 52.005 165.215 52.175 165.695 ;
        RECT 52.425 165.385 52.665 165.865 ;
        RECT 52.845 165.215 53.015 165.695 ;
        RECT 53.335 165.385 53.615 165.865 ;
        RECT 53.785 165.215 54.045 165.605 ;
        RECT 54.220 165.385 54.475 165.865 ;
        RECT 54.645 165.215 54.940 165.605 ;
        RECT 55.120 165.385 55.395 165.865 ;
        RECT 55.565 165.365 55.865 165.695 ;
        RECT 51.165 165.045 52.175 165.215 ;
        RECT 52.380 165.045 53.015 165.215 ;
        RECT 53.290 165.045 54.940 165.215 ;
        RECT 51.165 164.505 51.660 165.045 ;
        RECT 52.380 164.875 52.550 165.045 ;
        RECT 52.050 164.705 52.550 164.875 ;
        RECT 49.135 163.315 50.345 164.405 ;
        RECT 50.665 163.315 50.995 164.465 ;
        RECT 51.165 164.335 52.175 164.505 ;
        RECT 51.165 163.485 51.335 164.335 ;
        RECT 51.505 163.315 51.835 164.115 ;
        RECT 52.005 163.485 52.175 164.335 ;
        RECT 52.380 164.465 52.550 164.705 ;
        RECT 52.720 164.635 53.100 164.875 ;
        RECT 53.290 164.535 53.695 165.045 ;
        RECT 53.865 164.705 55.005 164.875 ;
        RECT 52.380 164.295 53.095 164.465 ;
        RECT 53.290 164.365 54.045 164.535 ;
        RECT 52.355 163.315 52.595 164.115 ;
        RECT 52.765 163.485 53.095 164.295 ;
        RECT 53.330 163.315 53.615 164.185 ;
        RECT 53.785 164.115 54.045 164.365 ;
        RECT 54.835 164.455 55.005 164.705 ;
        RECT 55.175 164.625 55.525 165.195 ;
        RECT 55.695 164.455 55.865 165.365 ;
        RECT 56.500 165.320 61.845 165.865 ;
        RECT 62.015 165.365 62.315 165.695 ;
        RECT 62.485 165.385 62.760 165.865 ;
        RECT 54.835 164.285 55.865 164.455 ;
        RECT 53.785 163.945 54.905 164.115 ;
        RECT 53.785 163.485 54.045 163.945 ;
        RECT 54.220 163.315 54.475 163.775 ;
        RECT 54.645 163.485 54.905 163.945 ;
        RECT 55.075 163.315 55.385 164.115 ;
        RECT 55.555 163.485 55.865 164.285 ;
        RECT 58.090 163.750 58.440 165.000 ;
        RECT 59.920 164.490 60.260 165.320 ;
        RECT 62.015 164.455 62.185 165.365 ;
        RECT 62.940 165.215 63.235 165.605 ;
        RECT 63.405 165.385 63.660 165.865 ;
        RECT 63.835 165.215 64.095 165.605 ;
        RECT 64.265 165.385 64.545 165.865 ;
        RECT 62.355 164.625 62.705 165.195 ;
        RECT 62.940 165.045 64.590 165.215 ;
        RECT 62.875 164.705 64.015 164.875 ;
        RECT 62.875 164.455 63.045 164.705 ;
        RECT 64.185 164.535 64.590 165.045 ;
        RECT 62.015 164.285 63.045 164.455 ;
        RECT 63.835 164.365 64.590 164.535 ;
        RECT 65.150 165.155 65.405 165.685 ;
        RECT 65.585 165.405 65.870 165.865 ;
        RECT 56.500 163.315 61.845 163.750 ;
        RECT 62.015 163.485 62.325 164.285 ;
        RECT 63.835 164.115 64.095 164.365 ;
        RECT 65.150 164.295 65.330 165.155 ;
        RECT 66.050 164.955 66.300 165.605 ;
        RECT 65.500 164.625 66.300 164.955 ;
        RECT 62.495 163.315 62.805 164.115 ;
        RECT 62.975 163.945 64.095 164.115 ;
        RECT 62.975 163.485 63.235 163.945 ;
        RECT 63.405 163.315 63.660 163.775 ;
        RECT 63.835 163.485 64.095 163.945 ;
        RECT 64.265 163.315 64.550 164.185 ;
        RECT 65.150 163.825 65.405 164.295 ;
        RECT 65.065 163.655 65.405 163.825 ;
        RECT 65.150 163.625 65.405 163.655 ;
        RECT 65.585 163.315 65.870 164.115 ;
        RECT 66.050 164.035 66.300 164.625 ;
        RECT 66.500 165.270 66.820 165.600 ;
        RECT 67.000 165.385 67.660 165.865 ;
        RECT 67.860 165.475 68.710 165.645 ;
        RECT 66.500 164.375 66.690 165.270 ;
        RECT 67.010 164.945 67.670 165.215 ;
        RECT 67.340 164.885 67.670 164.945 ;
        RECT 66.860 164.715 67.190 164.775 ;
        RECT 67.860 164.715 68.030 165.475 ;
        RECT 69.270 165.405 69.590 165.865 ;
        RECT 69.790 165.225 70.040 165.655 ;
        RECT 70.330 165.425 70.740 165.865 ;
        RECT 70.910 165.485 71.925 165.685 ;
        RECT 68.200 165.055 69.450 165.225 ;
        RECT 68.200 164.935 68.530 165.055 ;
        RECT 66.860 164.545 68.760 164.715 ;
        RECT 66.500 164.205 68.420 164.375 ;
        RECT 66.500 164.185 66.820 164.205 ;
        RECT 66.050 163.525 66.380 164.035 ;
        RECT 66.650 163.575 66.820 164.185 ;
        RECT 68.590 164.035 68.760 164.545 ;
        RECT 68.930 164.475 69.110 164.885 ;
        RECT 69.280 164.295 69.450 165.055 ;
        RECT 66.990 163.315 67.320 164.005 ;
        RECT 67.550 163.865 68.760 164.035 ;
        RECT 68.930 163.985 69.450 164.295 ;
        RECT 69.620 164.885 70.040 165.225 ;
        RECT 70.330 164.885 70.740 165.215 ;
        RECT 69.620 164.115 69.810 164.885 ;
        RECT 70.910 164.755 71.080 165.485 ;
        RECT 72.225 165.315 72.395 165.645 ;
        RECT 72.565 165.485 72.895 165.865 ;
        RECT 71.250 164.935 71.600 165.305 ;
        RECT 70.910 164.715 71.330 164.755 ;
        RECT 69.980 164.545 71.330 164.715 ;
        RECT 69.980 164.385 70.230 164.545 ;
        RECT 70.740 164.115 70.990 164.375 ;
        RECT 69.620 163.865 70.990 164.115 ;
        RECT 67.550 163.575 67.790 163.865 ;
        RECT 68.590 163.785 68.760 163.865 ;
        RECT 67.990 163.315 68.410 163.695 ;
        RECT 68.590 163.535 69.220 163.785 ;
        RECT 69.690 163.315 70.020 163.695 ;
        RECT 70.190 163.575 70.360 163.865 ;
        RECT 71.160 163.700 71.330 164.545 ;
        RECT 71.780 164.375 72.000 165.245 ;
        RECT 72.225 165.125 72.920 165.315 ;
        RECT 71.500 163.995 72.000 164.375 ;
        RECT 72.170 164.325 72.580 164.945 ;
        RECT 72.750 164.155 72.920 165.125 ;
        RECT 72.225 163.985 72.920 164.155 ;
        RECT 70.540 163.315 70.920 163.695 ;
        RECT 71.160 163.530 71.990 163.700 ;
        RECT 72.225 163.485 72.395 163.985 ;
        RECT 72.565 163.315 72.895 163.815 ;
        RECT 73.110 163.485 73.335 165.605 ;
        RECT 73.505 165.485 73.835 165.865 ;
        RECT 74.005 165.315 74.175 165.605 ;
        RECT 73.510 165.145 74.175 165.315 ;
        RECT 73.510 164.155 73.740 165.145 ;
        RECT 74.435 165.140 74.725 165.865 ;
        RECT 75.905 165.315 76.075 165.605 ;
        RECT 76.245 165.485 76.575 165.865 ;
        RECT 75.905 165.145 76.570 165.315 ;
        RECT 73.910 164.325 74.260 164.975 ;
        RECT 73.510 163.985 74.175 164.155 ;
        RECT 73.505 163.315 73.835 163.815 ;
        RECT 74.005 163.485 74.175 163.985 ;
        RECT 74.435 163.315 74.725 164.480 ;
        RECT 75.820 164.325 76.170 164.975 ;
        RECT 76.340 164.155 76.570 165.145 ;
        RECT 75.905 163.985 76.570 164.155 ;
        RECT 75.905 163.485 76.075 163.985 ;
        RECT 76.245 163.315 76.575 163.815 ;
        RECT 76.745 163.485 76.970 165.605 ;
        RECT 77.185 165.485 77.515 165.865 ;
        RECT 77.685 165.315 77.855 165.645 ;
        RECT 78.155 165.485 79.170 165.685 ;
        RECT 77.160 165.125 77.855 165.315 ;
        RECT 77.160 164.155 77.330 165.125 ;
        RECT 77.500 164.325 77.910 164.945 ;
        RECT 78.080 164.375 78.300 165.245 ;
        RECT 78.480 164.935 78.830 165.305 ;
        RECT 79.000 164.755 79.170 165.485 ;
        RECT 79.340 165.425 79.750 165.865 ;
        RECT 80.040 165.225 80.290 165.655 ;
        RECT 80.490 165.405 80.810 165.865 ;
        RECT 81.370 165.475 82.220 165.645 ;
        RECT 79.340 164.885 79.750 165.215 ;
        RECT 80.040 164.885 80.460 165.225 ;
        RECT 78.750 164.715 79.170 164.755 ;
        RECT 78.750 164.545 80.100 164.715 ;
        RECT 77.160 163.985 77.855 164.155 ;
        RECT 78.080 163.995 78.580 164.375 ;
        RECT 77.185 163.315 77.515 163.815 ;
        RECT 77.685 163.485 77.855 163.985 ;
        RECT 78.750 163.700 78.920 164.545 ;
        RECT 79.850 164.385 80.100 164.545 ;
        RECT 79.090 164.115 79.340 164.375 ;
        RECT 80.270 164.115 80.460 164.885 ;
        RECT 79.090 163.865 80.460 164.115 ;
        RECT 80.630 165.055 81.880 165.225 ;
        RECT 80.630 164.295 80.800 165.055 ;
        RECT 81.550 164.935 81.880 165.055 ;
        RECT 80.970 164.475 81.150 164.885 ;
        RECT 82.050 164.715 82.220 165.475 ;
        RECT 82.420 165.385 83.080 165.865 ;
        RECT 83.260 165.270 83.580 165.600 ;
        RECT 82.410 164.945 83.070 165.215 ;
        RECT 82.410 164.885 82.740 164.945 ;
        RECT 82.890 164.715 83.220 164.775 ;
        RECT 81.320 164.545 83.220 164.715 ;
        RECT 80.630 163.985 81.150 164.295 ;
        RECT 81.320 164.035 81.490 164.545 ;
        RECT 83.390 164.375 83.580 165.270 ;
        RECT 81.660 164.205 83.580 164.375 ;
        RECT 83.260 164.185 83.580 164.205 ;
        RECT 83.780 164.955 84.030 165.605 ;
        RECT 84.210 165.405 84.495 165.865 ;
        RECT 84.675 165.155 84.930 165.685 ;
        RECT 85.585 165.385 85.755 165.865 ;
        RECT 85.925 165.215 86.255 165.690 ;
        RECT 86.425 165.385 86.595 165.865 ;
        RECT 86.765 165.215 87.095 165.690 ;
        RECT 87.265 165.385 87.435 165.865 ;
        RECT 87.605 165.215 87.935 165.690 ;
        RECT 88.105 165.385 88.275 165.865 ;
        RECT 88.445 165.215 88.775 165.690 ;
        RECT 88.945 165.385 89.115 165.865 ;
        RECT 89.285 165.215 89.615 165.690 ;
        RECT 89.785 165.385 89.955 165.865 ;
        RECT 90.205 165.690 90.375 165.695 ;
        RECT 90.125 165.215 90.455 165.690 ;
        RECT 90.625 165.385 90.795 165.865 ;
        RECT 91.045 165.690 91.215 165.695 ;
        RECT 90.965 165.215 91.295 165.690 ;
        RECT 91.465 165.385 91.635 165.865 ;
        RECT 91.885 165.690 92.135 165.695 ;
        RECT 91.805 165.215 92.135 165.690 ;
        RECT 92.305 165.385 92.475 165.865 ;
        RECT 92.645 165.215 92.975 165.690 ;
        RECT 93.145 165.385 93.315 165.865 ;
        RECT 93.485 165.215 93.815 165.690 ;
        RECT 93.985 165.385 94.155 165.865 ;
        RECT 94.325 165.215 94.655 165.690 ;
        RECT 94.825 165.385 94.995 165.865 ;
        RECT 95.165 165.215 95.495 165.690 ;
        RECT 95.665 165.385 95.835 165.865 ;
        RECT 96.005 165.215 96.335 165.690 ;
        RECT 83.780 164.625 84.580 164.955 ;
        RECT 81.320 163.865 82.530 164.035 ;
        RECT 78.090 163.530 78.920 163.700 ;
        RECT 79.160 163.315 79.540 163.695 ;
        RECT 79.720 163.575 79.890 163.865 ;
        RECT 81.320 163.785 81.490 163.865 ;
        RECT 80.060 163.315 80.390 163.695 ;
        RECT 80.860 163.535 81.490 163.785 ;
        RECT 81.670 163.315 82.090 163.695 ;
        RECT 82.290 163.575 82.530 163.865 ;
        RECT 82.760 163.315 83.090 164.005 ;
        RECT 83.260 163.575 83.430 164.185 ;
        RECT 83.780 164.035 84.030 164.625 ;
        RECT 84.750 164.295 84.930 165.155 ;
        RECT 85.475 165.045 92.135 165.215 ;
        RECT 92.305 165.045 94.655 165.215 ;
        RECT 94.825 165.045 96.335 165.215 ;
        RECT 96.630 165.235 96.915 165.695 ;
        RECT 97.085 165.405 97.355 165.865 ;
        RECT 96.630 165.065 97.585 165.235 ;
        RECT 85.475 164.505 85.750 165.045 ;
        RECT 92.305 164.875 92.480 165.045 ;
        RECT 94.825 164.875 94.995 165.045 ;
        RECT 85.920 164.675 92.480 164.875 ;
        RECT 92.685 164.675 94.995 164.875 ;
        RECT 95.165 164.675 96.340 164.875 ;
        RECT 92.305 164.505 92.480 164.675 ;
        RECT 94.825 164.505 94.995 164.675 ;
        RECT 85.475 164.335 92.135 164.505 ;
        RECT 92.305 164.335 94.655 164.505 ;
        RECT 94.825 164.335 96.335 164.505 ;
        RECT 96.515 164.335 97.205 164.895 ;
        RECT 84.675 164.165 84.930 164.295 ;
        RECT 83.700 163.525 84.030 164.035 ;
        RECT 84.210 163.315 84.495 164.115 ;
        RECT 84.675 163.995 85.015 164.165 ;
        RECT 84.675 163.625 84.930 163.995 ;
        RECT 85.585 163.315 85.755 164.115 ;
        RECT 85.925 163.485 86.255 164.335 ;
        RECT 86.425 163.315 86.595 164.115 ;
        RECT 86.765 163.485 87.095 164.335 ;
        RECT 87.265 163.315 87.435 164.115 ;
        RECT 87.605 163.485 87.935 164.335 ;
        RECT 88.105 163.315 88.275 164.115 ;
        RECT 88.445 163.485 88.775 164.335 ;
        RECT 88.945 163.315 89.115 164.115 ;
        RECT 89.285 163.485 89.615 164.335 ;
        RECT 89.785 163.315 89.955 164.115 ;
        RECT 90.125 163.485 90.455 164.335 ;
        RECT 90.625 163.315 90.795 164.115 ;
        RECT 90.965 163.485 91.295 164.335 ;
        RECT 91.465 163.315 91.635 164.115 ;
        RECT 91.805 163.485 92.135 164.335 ;
        RECT 92.305 163.315 92.475 164.115 ;
        RECT 92.645 163.485 92.975 164.335 ;
        RECT 93.145 163.315 93.315 164.115 ;
        RECT 93.485 163.485 93.815 164.335 ;
        RECT 93.985 163.315 94.155 164.115 ;
        RECT 94.325 163.485 94.655 164.335 ;
        RECT 94.825 163.315 94.995 164.165 ;
        RECT 95.165 163.485 95.495 164.335 ;
        RECT 95.665 163.315 95.835 164.165 ;
        RECT 96.005 163.485 96.335 164.335 ;
        RECT 97.375 164.165 97.585 165.065 ;
        RECT 96.630 163.945 97.585 164.165 ;
        RECT 97.755 164.895 98.155 165.695 ;
        RECT 98.345 165.235 98.625 165.695 ;
        RECT 99.145 165.405 99.470 165.865 ;
        RECT 98.345 165.065 99.470 165.235 ;
        RECT 99.640 165.125 100.025 165.695 ;
        RECT 100.195 165.140 100.485 165.865 ;
        RECT 99.020 164.955 99.470 165.065 ;
        RECT 97.755 164.335 98.850 164.895 ;
        RECT 99.020 164.625 99.575 164.955 ;
        RECT 96.630 163.485 96.915 163.945 ;
        RECT 97.085 163.315 97.355 163.775 ;
        RECT 97.755 163.485 98.155 164.335 ;
        RECT 99.020 164.165 99.470 164.625 ;
        RECT 99.745 164.455 100.025 165.125 ;
        RECT 100.930 165.055 101.175 165.660 ;
        RECT 101.395 165.330 101.905 165.865 ;
        RECT 100.655 164.885 101.885 165.055 ;
        RECT 98.345 163.945 99.470 164.165 ;
        RECT 98.345 163.485 98.625 163.945 ;
        RECT 99.145 163.315 99.470 163.775 ;
        RECT 99.640 163.485 100.025 164.455 ;
        RECT 100.195 163.315 100.485 164.480 ;
        RECT 100.655 164.075 100.995 164.885 ;
        RECT 101.165 164.320 101.915 164.510 ;
        RECT 100.655 163.665 101.170 164.075 ;
        RECT 101.405 163.315 101.575 164.075 ;
        RECT 101.745 163.655 101.915 164.320 ;
        RECT 102.085 164.335 102.275 165.695 ;
        RECT 102.445 165.185 102.720 165.695 ;
        RECT 102.910 165.330 103.440 165.695 ;
        RECT 103.865 165.465 104.195 165.865 ;
        RECT 103.265 165.295 103.440 165.330 ;
        RECT 102.445 165.015 102.725 165.185 ;
        RECT 102.445 164.535 102.720 165.015 ;
        RECT 102.925 164.335 103.095 165.135 ;
        RECT 102.085 164.165 103.095 164.335 ;
        RECT 103.265 165.125 104.195 165.295 ;
        RECT 104.365 165.125 104.620 165.695 ;
        RECT 103.265 163.995 103.435 165.125 ;
        RECT 104.025 164.955 104.195 165.125 ;
        RECT 102.310 163.825 103.435 163.995 ;
        RECT 103.605 164.625 103.800 164.955 ;
        RECT 104.025 164.625 104.280 164.955 ;
        RECT 103.605 163.655 103.775 164.625 ;
        RECT 104.450 164.455 104.620 165.125 ;
        RECT 104.910 165.235 105.195 165.695 ;
        RECT 105.365 165.405 105.635 165.865 ;
        RECT 104.910 165.065 105.865 165.235 ;
        RECT 101.745 163.485 103.775 163.655 ;
        RECT 103.945 163.315 104.115 164.455 ;
        RECT 104.285 163.485 104.620 164.455 ;
        RECT 104.795 164.335 105.485 164.895 ;
        RECT 105.655 164.165 105.865 165.065 ;
        RECT 104.910 163.945 105.865 164.165 ;
        RECT 106.035 164.895 106.435 165.695 ;
        RECT 106.625 165.235 106.905 165.695 ;
        RECT 107.425 165.405 107.750 165.865 ;
        RECT 106.625 165.065 107.750 165.235 ;
        RECT 107.920 165.125 108.305 165.695 ;
        RECT 107.300 164.955 107.750 165.065 ;
        RECT 106.035 164.335 107.130 164.895 ;
        RECT 107.300 164.625 107.855 164.955 ;
        RECT 104.910 163.485 105.195 163.945 ;
        RECT 105.365 163.315 105.635 163.775 ;
        RECT 106.035 163.485 106.435 164.335 ;
        RECT 107.300 164.165 107.750 164.625 ;
        RECT 108.025 164.455 108.305 165.125 ;
        RECT 106.625 163.945 107.750 164.165 ;
        RECT 106.625 163.485 106.905 163.945 ;
        RECT 107.425 163.315 107.750 163.775 ;
        RECT 107.920 163.485 108.305 164.455 ;
        RECT 108.475 165.190 108.735 165.695 ;
        RECT 108.915 165.485 109.245 165.865 ;
        RECT 109.425 165.315 109.595 165.695 ;
        RECT 108.475 164.390 108.645 165.190 ;
        RECT 108.930 165.145 109.595 165.315 ;
        RECT 108.930 164.890 109.100 165.145 ;
        RECT 110.315 165.095 111.985 165.865 ;
        RECT 112.155 165.115 113.365 165.865 ;
        RECT 108.815 164.560 109.100 164.890 ;
        RECT 109.335 164.595 109.665 164.965 ;
        RECT 108.930 164.415 109.100 164.560 ;
        RECT 108.475 163.485 108.745 164.390 ;
        RECT 108.930 164.245 109.595 164.415 ;
        RECT 108.915 163.315 109.245 164.075 ;
        RECT 109.425 163.485 109.595 164.245 ;
        RECT 110.315 164.405 111.065 164.925 ;
        RECT 111.235 164.575 111.985 165.095 ;
        RECT 112.155 164.405 112.675 164.945 ;
        RECT 112.845 164.575 113.365 165.115 ;
        RECT 110.315 163.315 111.985 164.405 ;
        RECT 112.155 163.315 113.365 164.405 ;
        RECT 11.330 163.145 113.450 163.315 ;
        RECT 11.415 162.055 12.625 163.145 ;
        RECT 11.415 161.345 11.935 161.885 ;
        RECT 12.105 161.515 12.625 162.055 ;
        RECT 12.855 162.005 13.065 163.145 ;
        RECT 13.235 161.995 13.565 162.975 ;
        RECT 13.735 162.005 13.965 163.145 ;
        RECT 14.175 162.310 14.560 163.145 ;
        RECT 14.730 162.140 14.990 162.945 ;
        RECT 15.160 162.310 15.420 163.145 ;
        RECT 15.590 162.140 15.845 162.945 ;
        RECT 16.020 162.310 16.280 163.145 ;
        RECT 16.450 162.140 16.705 162.945 ;
        RECT 16.880 162.310 17.225 163.145 ;
        RECT 11.415 160.595 12.625 161.345 ;
        RECT 12.855 160.595 13.065 161.415 ;
        RECT 13.235 161.395 13.485 161.995 ;
        RECT 14.175 161.970 17.205 162.140 ;
        RECT 13.655 161.585 13.985 161.835 ;
        RECT 13.235 160.765 13.565 161.395 ;
        RECT 13.735 160.595 13.965 161.415 ;
        RECT 14.175 161.405 14.475 161.970 ;
        RECT 14.650 161.575 16.865 161.800 ;
        RECT 17.035 161.405 17.205 161.970 ;
        RECT 14.175 161.235 17.205 161.405 ;
        RECT 17.400 162.005 17.735 162.975 ;
        RECT 17.905 162.005 18.075 163.145 ;
        RECT 18.245 162.805 20.275 162.975 ;
        RECT 17.400 161.335 17.570 162.005 ;
        RECT 18.245 161.835 18.415 162.805 ;
        RECT 17.740 161.505 17.995 161.835 ;
        RECT 18.220 161.505 18.415 161.835 ;
        RECT 18.585 162.465 19.710 162.635 ;
        RECT 17.825 161.335 17.995 161.505 ;
        RECT 18.585 161.335 18.755 162.465 ;
        RECT 14.695 160.595 14.995 161.065 ;
        RECT 15.165 160.790 15.420 161.235 ;
        RECT 15.590 160.595 15.850 161.065 ;
        RECT 16.020 160.790 16.280 161.235 ;
        RECT 16.450 160.595 16.745 161.065 ;
        RECT 17.400 160.765 17.655 161.335 ;
        RECT 17.825 161.165 18.755 161.335 ;
        RECT 18.925 162.125 19.935 162.295 ;
        RECT 18.925 161.325 19.095 162.125 ;
        RECT 18.580 161.130 18.755 161.165 ;
        RECT 17.825 160.595 18.155 160.995 ;
        RECT 18.580 160.765 19.110 161.130 ;
        RECT 19.300 161.105 19.575 161.925 ;
        RECT 19.295 160.935 19.575 161.105 ;
        RECT 19.300 160.765 19.575 160.935 ;
        RECT 19.745 160.765 19.935 162.125 ;
        RECT 20.105 162.140 20.275 162.805 ;
        RECT 20.445 162.385 20.615 163.145 ;
        RECT 20.850 162.385 21.365 162.795 ;
        RECT 20.105 161.950 20.855 162.140 ;
        RECT 21.025 161.575 21.365 162.385 ;
        RECT 20.135 161.405 21.365 161.575 ;
        RECT 22.460 162.005 22.795 162.975 ;
        RECT 22.965 162.005 23.135 163.145 ;
        RECT 23.305 162.805 25.335 162.975 ;
        RECT 20.115 160.595 20.625 161.130 ;
        RECT 20.845 160.800 21.090 161.405 ;
        RECT 22.460 161.335 22.630 162.005 ;
        RECT 23.305 161.835 23.475 162.805 ;
        RECT 22.800 161.505 23.055 161.835 ;
        RECT 23.280 161.505 23.475 161.835 ;
        RECT 23.645 162.465 24.770 162.635 ;
        RECT 22.885 161.335 23.055 161.505 ;
        RECT 23.645 161.335 23.815 162.465 ;
        RECT 22.460 160.765 22.715 161.335 ;
        RECT 22.885 161.165 23.815 161.335 ;
        RECT 23.985 162.125 24.995 162.295 ;
        RECT 23.985 161.325 24.155 162.125 ;
        RECT 24.360 161.785 24.635 161.925 ;
        RECT 24.355 161.615 24.635 161.785 ;
        RECT 23.640 161.130 23.815 161.165 ;
        RECT 22.885 160.595 23.215 160.995 ;
        RECT 23.640 160.765 24.170 161.130 ;
        RECT 24.360 160.765 24.635 161.615 ;
        RECT 24.805 160.765 24.995 162.125 ;
        RECT 25.165 162.140 25.335 162.805 ;
        RECT 25.505 162.385 25.675 163.145 ;
        RECT 25.910 162.385 26.425 162.795 ;
        RECT 25.165 161.950 25.915 162.140 ;
        RECT 26.085 161.575 26.425 162.385 ;
        RECT 26.600 162.475 26.855 162.975 ;
        RECT 27.025 162.645 27.355 163.145 ;
        RECT 26.600 162.305 27.350 162.475 ;
        RECT 25.195 161.405 26.425 161.575 ;
        RECT 26.600 161.485 26.950 162.135 ;
        RECT 25.175 160.595 25.685 161.130 ;
        RECT 25.905 160.800 26.150 161.405 ;
        RECT 27.120 161.315 27.350 162.305 ;
        RECT 26.600 161.145 27.350 161.315 ;
        RECT 26.600 160.855 26.855 161.145 ;
        RECT 27.025 160.595 27.355 160.975 ;
        RECT 27.525 160.855 27.695 162.975 ;
        RECT 27.865 162.175 28.190 162.960 ;
        RECT 28.360 162.685 28.610 163.145 ;
        RECT 28.780 162.645 29.030 162.975 ;
        RECT 29.245 162.645 29.925 162.975 ;
        RECT 28.780 162.515 28.950 162.645 ;
        RECT 28.555 162.345 28.950 162.515 ;
        RECT 27.925 161.125 28.385 162.175 ;
        RECT 28.555 160.985 28.725 162.345 ;
        RECT 29.120 162.085 29.585 162.475 ;
        RECT 28.895 161.275 29.245 161.895 ;
        RECT 29.415 161.495 29.585 162.085 ;
        RECT 29.755 161.865 29.925 162.645 ;
        RECT 30.095 162.545 30.265 162.885 ;
        RECT 30.500 162.715 30.830 163.145 ;
        RECT 31.000 162.545 31.170 162.885 ;
        RECT 31.465 162.685 31.835 163.145 ;
        RECT 30.095 162.375 31.170 162.545 ;
        RECT 32.005 162.515 32.175 162.975 ;
        RECT 32.410 162.635 33.280 162.975 ;
        RECT 33.450 162.685 33.700 163.145 ;
        RECT 31.615 162.345 32.175 162.515 ;
        RECT 31.615 162.205 31.785 162.345 ;
        RECT 30.285 162.035 31.785 162.205 ;
        RECT 32.480 162.175 32.940 162.465 ;
        RECT 29.755 161.695 31.445 161.865 ;
        RECT 29.415 161.275 29.770 161.495 ;
        RECT 29.940 160.985 30.110 161.695 ;
        RECT 30.315 161.275 31.105 161.525 ;
        RECT 31.275 161.515 31.445 161.695 ;
        RECT 31.615 161.345 31.785 162.035 ;
        RECT 28.055 160.595 28.385 160.955 ;
        RECT 28.555 160.815 29.050 160.985 ;
        RECT 29.255 160.815 30.110 160.985 ;
        RECT 30.985 160.595 31.315 161.055 ;
        RECT 31.525 160.955 31.785 161.345 ;
        RECT 31.975 162.165 32.940 162.175 ;
        RECT 33.110 162.255 33.280 162.635 ;
        RECT 33.870 162.595 34.040 162.885 ;
        RECT 34.220 162.765 34.550 163.145 ;
        RECT 33.870 162.425 34.670 162.595 ;
        RECT 31.975 162.005 32.650 162.165 ;
        RECT 33.110 162.085 34.330 162.255 ;
        RECT 31.975 161.215 32.185 162.005 ;
        RECT 33.110 161.995 33.280 162.085 ;
        RECT 32.355 161.215 32.705 161.835 ;
        RECT 32.875 161.825 33.280 161.995 ;
        RECT 32.875 161.045 33.045 161.825 ;
        RECT 33.215 161.375 33.435 161.655 ;
        RECT 33.615 161.545 34.155 161.915 ;
        RECT 34.500 161.835 34.670 162.425 ;
        RECT 34.890 162.005 35.195 163.145 ;
        RECT 35.365 161.955 35.620 162.835 ;
        RECT 35.795 161.980 36.085 163.145 ;
        RECT 36.255 162.385 36.770 162.795 ;
        RECT 37.005 162.385 37.175 163.145 ;
        RECT 37.345 162.805 39.375 162.975 ;
        RECT 34.500 161.805 35.240 161.835 ;
        RECT 33.215 161.205 33.745 161.375 ;
        RECT 31.525 160.785 31.875 160.955 ;
        RECT 32.095 160.765 33.045 161.045 ;
        RECT 33.215 160.595 33.405 161.035 ;
        RECT 33.575 160.975 33.745 161.205 ;
        RECT 33.915 161.145 34.155 161.545 ;
        RECT 34.325 161.505 35.240 161.805 ;
        RECT 34.325 161.330 34.650 161.505 ;
        RECT 34.325 160.975 34.645 161.330 ;
        RECT 35.410 161.305 35.620 161.955 ;
        RECT 36.255 161.575 36.595 162.385 ;
        RECT 37.345 162.140 37.515 162.805 ;
        RECT 37.910 162.465 39.035 162.635 ;
        RECT 36.765 161.950 37.515 162.140 ;
        RECT 37.685 162.125 38.695 162.295 ;
        RECT 36.255 161.405 37.485 161.575 ;
        RECT 33.575 160.805 34.645 160.975 ;
        RECT 34.890 160.595 35.195 161.055 ;
        RECT 35.365 160.775 35.620 161.305 ;
        RECT 35.795 160.595 36.085 161.320 ;
        RECT 36.530 160.800 36.775 161.405 ;
        RECT 36.995 160.595 37.505 161.130 ;
        RECT 37.685 160.765 37.875 162.125 ;
        RECT 38.045 161.785 38.320 161.925 ;
        RECT 38.045 161.615 38.325 161.785 ;
        RECT 38.045 160.765 38.320 161.615 ;
        RECT 38.525 161.325 38.695 162.125 ;
        RECT 38.865 161.335 39.035 162.465 ;
        RECT 39.205 161.835 39.375 162.805 ;
        RECT 39.545 162.005 39.715 163.145 ;
        RECT 39.885 162.005 40.220 162.975 ;
        RECT 39.205 161.505 39.400 161.835 ;
        RECT 39.625 161.505 39.880 161.835 ;
        RECT 39.625 161.335 39.795 161.505 ;
        RECT 40.050 161.335 40.220 162.005 ;
        RECT 38.865 161.165 39.795 161.335 ;
        RECT 38.865 161.130 39.040 161.165 ;
        RECT 38.510 160.765 39.040 161.130 ;
        RECT 39.465 160.595 39.795 160.995 ;
        RECT 39.965 160.765 40.220 161.335 ;
        RECT 40.400 161.955 40.655 162.835 ;
        RECT 40.825 162.005 41.130 163.145 ;
        RECT 41.470 162.765 41.800 163.145 ;
        RECT 41.980 162.595 42.150 162.885 ;
        RECT 42.320 162.685 42.570 163.145 ;
        RECT 41.350 162.425 42.150 162.595 ;
        RECT 42.740 162.635 43.610 162.975 ;
        RECT 40.400 161.305 40.610 161.955 ;
        RECT 41.350 161.835 41.520 162.425 ;
        RECT 42.740 162.255 42.910 162.635 ;
        RECT 43.845 162.515 44.015 162.975 ;
        RECT 44.185 162.685 44.555 163.145 ;
        RECT 44.850 162.545 45.020 162.885 ;
        RECT 45.190 162.715 45.520 163.145 ;
        RECT 45.755 162.545 45.925 162.885 ;
        RECT 41.690 162.085 42.910 162.255 ;
        RECT 43.080 162.175 43.540 162.465 ;
        RECT 43.845 162.345 44.405 162.515 ;
        RECT 44.850 162.375 45.925 162.545 ;
        RECT 46.095 162.645 46.775 162.975 ;
        RECT 46.990 162.645 47.240 162.975 ;
        RECT 47.410 162.685 47.660 163.145 ;
        RECT 44.235 162.205 44.405 162.345 ;
        RECT 43.080 162.165 44.045 162.175 ;
        RECT 42.740 161.995 42.910 162.085 ;
        RECT 43.370 162.005 44.045 162.165 ;
        RECT 40.780 161.805 41.520 161.835 ;
        RECT 40.780 161.505 41.695 161.805 ;
        RECT 41.370 161.330 41.695 161.505 ;
        RECT 40.400 160.775 40.655 161.305 ;
        RECT 40.825 160.595 41.130 161.055 ;
        RECT 41.375 160.975 41.695 161.330 ;
        RECT 41.865 161.545 42.405 161.915 ;
        RECT 42.740 161.825 43.145 161.995 ;
        RECT 41.865 161.145 42.105 161.545 ;
        RECT 42.585 161.375 42.805 161.655 ;
        RECT 42.275 161.205 42.805 161.375 ;
        RECT 42.275 160.975 42.445 161.205 ;
        RECT 42.975 161.045 43.145 161.825 ;
        RECT 43.315 161.215 43.665 161.835 ;
        RECT 43.835 161.215 44.045 162.005 ;
        RECT 44.235 162.035 45.735 162.205 ;
        RECT 44.235 161.345 44.405 162.035 ;
        RECT 46.095 161.865 46.265 162.645 ;
        RECT 47.070 162.515 47.240 162.645 ;
        RECT 44.575 161.695 46.265 161.865 ;
        RECT 46.435 162.085 46.900 162.475 ;
        RECT 47.070 162.345 47.465 162.515 ;
        RECT 44.575 161.515 44.745 161.695 ;
        RECT 41.375 160.805 42.445 160.975 ;
        RECT 42.615 160.595 42.805 161.035 ;
        RECT 42.975 160.765 43.925 161.045 ;
        RECT 44.235 160.955 44.495 161.345 ;
        RECT 44.915 161.275 45.705 161.525 ;
        RECT 44.145 160.785 44.495 160.955 ;
        RECT 44.705 160.595 45.035 161.055 ;
        RECT 45.910 160.985 46.080 161.695 ;
        RECT 46.435 161.495 46.605 162.085 ;
        RECT 46.250 161.275 46.605 161.495 ;
        RECT 46.775 161.275 47.125 161.895 ;
        RECT 47.295 160.985 47.465 162.345 ;
        RECT 47.830 162.175 48.155 162.960 ;
        RECT 47.635 161.125 48.095 162.175 ;
        RECT 45.910 160.815 46.765 160.985 ;
        RECT 46.970 160.815 47.465 160.985 ;
        RECT 47.635 160.595 47.965 160.955 ;
        RECT 48.325 160.855 48.495 162.975 ;
        RECT 48.665 162.645 48.995 163.145 ;
        RECT 49.165 162.475 49.420 162.975 ;
        RECT 48.670 162.305 49.420 162.475 ;
        RECT 48.670 161.315 48.900 162.305 ;
        RECT 49.070 161.485 49.420 162.135 ;
        RECT 49.595 162.070 49.865 162.975 ;
        RECT 50.035 162.385 50.365 163.145 ;
        RECT 50.545 162.215 50.715 162.975 ;
        RECT 50.980 162.710 56.325 163.145 ;
        RECT 48.670 161.145 49.420 161.315 ;
        RECT 48.665 160.595 48.995 160.975 ;
        RECT 49.165 160.855 49.420 161.145 ;
        RECT 49.595 161.270 49.765 162.070 ;
        RECT 50.050 162.045 50.715 162.215 ;
        RECT 50.050 161.900 50.220 162.045 ;
        RECT 49.935 161.570 50.220 161.900 ;
        RECT 50.050 161.315 50.220 161.570 ;
        RECT 50.455 161.495 50.785 161.865 ;
        RECT 52.570 161.460 52.920 162.710 ;
        RECT 56.535 162.005 56.765 163.145 ;
        RECT 56.935 161.995 57.265 162.975 ;
        RECT 57.435 162.005 57.645 163.145 ;
        RECT 57.880 161.995 58.140 163.145 ;
        RECT 58.315 162.070 58.570 162.975 ;
        RECT 58.740 162.385 59.070 163.145 ;
        RECT 59.285 162.215 59.455 162.975 ;
        RECT 49.595 160.765 49.855 161.270 ;
        RECT 50.050 161.145 50.715 161.315 ;
        RECT 50.035 160.595 50.365 160.975 ;
        RECT 50.545 160.765 50.715 161.145 ;
        RECT 54.400 161.140 54.740 161.970 ;
        RECT 56.515 161.585 56.845 161.835 ;
        RECT 50.980 160.595 56.325 161.140 ;
        RECT 56.535 160.595 56.765 161.415 ;
        RECT 57.015 161.395 57.265 161.995 ;
        RECT 56.935 160.765 57.265 161.395 ;
        RECT 57.435 160.595 57.645 161.415 ;
        RECT 57.880 160.595 58.140 161.435 ;
        RECT 58.315 161.340 58.485 162.070 ;
        RECT 58.740 162.045 59.455 162.215 ;
        RECT 58.740 161.835 58.910 162.045 ;
        RECT 59.720 161.995 59.980 163.145 ;
        RECT 60.155 162.070 60.410 162.975 ;
        RECT 60.580 162.385 60.910 163.145 ;
        RECT 61.125 162.215 61.295 162.975 ;
        RECT 58.655 161.505 58.910 161.835 ;
        RECT 58.315 160.765 58.570 161.340 ;
        RECT 58.740 161.315 58.910 161.505 ;
        RECT 59.190 161.495 59.545 161.865 ;
        RECT 58.740 161.145 59.455 161.315 ;
        RECT 58.740 160.595 59.070 160.975 ;
        RECT 59.285 160.765 59.455 161.145 ;
        RECT 59.720 160.595 59.980 161.435 ;
        RECT 60.155 161.340 60.325 162.070 ;
        RECT 60.580 162.045 61.295 162.215 ;
        RECT 60.580 161.835 60.750 162.045 ;
        RECT 61.555 161.980 61.845 163.145 ;
        RECT 62.105 162.215 62.275 162.975 ;
        RECT 62.490 162.385 62.820 163.145 ;
        RECT 62.105 162.045 62.820 162.215 ;
        RECT 62.990 162.070 63.245 162.975 ;
        RECT 60.495 161.505 60.750 161.835 ;
        RECT 60.155 160.765 60.410 161.340 ;
        RECT 60.580 161.315 60.750 161.505 ;
        RECT 61.030 161.495 61.385 161.865 ;
        RECT 62.015 161.495 62.370 161.865 ;
        RECT 62.650 161.835 62.820 162.045 ;
        RECT 62.650 161.505 62.905 161.835 ;
        RECT 60.580 161.145 61.295 161.315 ;
        RECT 60.580 160.595 60.910 160.975 ;
        RECT 61.125 160.765 61.295 161.145 ;
        RECT 61.555 160.595 61.845 161.320 ;
        RECT 62.650 161.315 62.820 161.505 ;
        RECT 63.075 161.340 63.245 162.070 ;
        RECT 63.420 161.995 63.680 163.145 ;
        RECT 63.945 162.215 64.115 162.975 ;
        RECT 64.330 162.385 64.660 163.145 ;
        RECT 63.945 162.045 64.660 162.215 ;
        RECT 64.830 162.070 65.085 162.975 ;
        RECT 63.855 161.495 64.210 161.865 ;
        RECT 64.490 161.835 64.660 162.045 ;
        RECT 64.490 161.505 64.745 161.835 ;
        RECT 62.105 161.145 62.820 161.315 ;
        RECT 62.105 160.765 62.275 161.145 ;
        RECT 62.490 160.595 62.820 160.975 ;
        RECT 62.990 160.765 63.245 161.340 ;
        RECT 63.420 160.595 63.680 161.435 ;
        RECT 64.490 161.315 64.660 161.505 ;
        RECT 64.915 161.340 65.085 162.070 ;
        RECT 65.260 161.995 65.520 163.145 ;
        RECT 66.155 162.055 69.665 163.145 ;
        RECT 69.925 162.215 70.095 162.975 ;
        RECT 70.275 162.385 70.605 163.145 ;
        RECT 66.155 161.535 67.845 162.055 ;
        RECT 69.925 162.045 70.590 162.215 ;
        RECT 70.775 162.070 71.045 162.975 ;
        RECT 70.420 161.900 70.590 162.045 ;
        RECT 63.945 161.145 64.660 161.315 ;
        RECT 63.945 160.765 64.115 161.145 ;
        RECT 64.330 160.595 64.660 160.975 ;
        RECT 64.830 160.765 65.085 161.340 ;
        RECT 65.260 160.595 65.520 161.435 ;
        RECT 68.015 161.365 69.665 161.885 ;
        RECT 69.855 161.495 70.185 161.865 ;
        RECT 70.420 161.570 70.705 161.900 ;
        RECT 66.155 160.595 69.665 161.365 ;
        RECT 70.420 161.315 70.590 161.570 ;
        RECT 69.925 161.145 70.590 161.315 ;
        RECT 70.875 161.270 71.045 162.070 ;
        RECT 69.925 160.765 70.095 161.145 ;
        RECT 70.275 160.595 70.605 160.975 ;
        RECT 70.785 160.765 71.045 161.270 ;
        RECT 71.220 162.005 71.555 162.975 ;
        RECT 71.725 162.005 71.895 163.145 ;
        RECT 72.065 162.805 74.095 162.975 ;
        RECT 71.220 161.335 71.390 162.005 ;
        RECT 72.065 161.835 72.235 162.805 ;
        RECT 71.560 161.505 71.815 161.835 ;
        RECT 72.040 161.505 72.235 161.835 ;
        RECT 72.405 162.465 73.530 162.635 ;
        RECT 71.645 161.335 71.815 161.505 ;
        RECT 72.405 161.335 72.575 162.465 ;
        RECT 71.220 160.765 71.475 161.335 ;
        RECT 71.645 161.165 72.575 161.335 ;
        RECT 72.745 162.125 73.755 162.295 ;
        RECT 72.745 161.325 72.915 162.125 ;
        RECT 72.400 161.130 72.575 161.165 ;
        RECT 71.645 160.595 71.975 160.995 ;
        RECT 72.400 160.765 72.930 161.130 ;
        RECT 73.120 161.105 73.395 161.925 ;
        RECT 73.115 160.935 73.395 161.105 ;
        RECT 73.120 160.765 73.395 160.935 ;
        RECT 73.565 160.765 73.755 162.125 ;
        RECT 73.925 162.140 74.095 162.805 ;
        RECT 74.265 162.385 74.435 163.145 ;
        RECT 74.670 162.385 75.185 162.795 ;
        RECT 73.925 161.950 74.675 162.140 ;
        RECT 74.845 161.575 75.185 162.385 ;
        RECT 75.415 162.005 75.625 163.145 ;
        RECT 73.955 161.405 75.185 161.575 ;
        RECT 75.795 161.995 76.125 162.975 ;
        RECT 76.295 162.005 76.525 163.145 ;
        RECT 76.795 162.005 77.005 163.145 ;
        RECT 77.175 161.995 77.505 162.975 ;
        RECT 77.675 162.005 77.905 163.145 ;
        RECT 79.035 162.385 79.550 162.795 ;
        RECT 79.785 162.385 79.955 163.145 ;
        RECT 80.125 162.805 82.155 162.975 ;
        RECT 73.935 160.595 74.445 161.130 ;
        RECT 74.665 160.800 74.910 161.405 ;
        RECT 75.415 160.595 75.625 161.415 ;
        RECT 75.795 161.395 76.045 161.995 ;
        RECT 76.215 161.585 76.545 161.835 ;
        RECT 75.795 160.765 76.125 161.395 ;
        RECT 76.295 160.595 76.525 161.415 ;
        RECT 76.795 160.595 77.005 161.415 ;
        RECT 77.175 161.395 77.425 161.995 ;
        RECT 77.595 161.585 77.925 161.835 ;
        RECT 79.035 161.575 79.375 162.385 ;
        RECT 80.125 162.140 80.295 162.805 ;
        RECT 80.690 162.465 81.815 162.635 ;
        RECT 79.545 161.950 80.295 162.140 ;
        RECT 80.465 162.125 81.475 162.295 ;
        RECT 77.175 160.765 77.505 161.395 ;
        RECT 77.675 160.595 77.905 161.415 ;
        RECT 79.035 161.405 80.265 161.575 ;
        RECT 79.310 160.800 79.555 161.405 ;
        RECT 79.775 160.595 80.285 161.130 ;
        RECT 80.465 160.765 80.655 162.125 ;
        RECT 80.825 161.105 81.100 161.925 ;
        RECT 81.305 161.325 81.475 162.125 ;
        RECT 81.645 161.335 81.815 162.465 ;
        RECT 81.985 161.835 82.155 162.805 ;
        RECT 82.325 162.005 82.495 163.145 ;
        RECT 82.665 162.005 83.000 162.975 ;
        RECT 81.985 161.505 82.180 161.835 ;
        RECT 82.405 161.505 82.660 161.835 ;
        RECT 82.405 161.335 82.575 161.505 ;
        RECT 82.830 161.335 83.000 162.005 ;
        RECT 83.175 162.385 83.690 162.795 ;
        RECT 83.925 162.385 84.095 163.145 ;
        RECT 84.265 162.805 86.295 162.975 ;
        RECT 83.175 161.575 83.515 162.385 ;
        RECT 84.265 162.140 84.435 162.805 ;
        RECT 84.830 162.465 85.955 162.635 ;
        RECT 83.685 161.950 84.435 162.140 ;
        RECT 84.605 162.125 85.615 162.295 ;
        RECT 83.175 161.405 84.405 161.575 ;
        RECT 81.645 161.165 82.575 161.335 ;
        RECT 81.645 161.130 81.820 161.165 ;
        RECT 80.825 160.935 81.105 161.105 ;
        RECT 80.825 160.765 81.100 160.935 ;
        RECT 81.290 160.765 81.820 161.130 ;
        RECT 82.245 160.595 82.575 160.995 ;
        RECT 82.745 160.765 83.000 161.335 ;
        RECT 83.450 160.800 83.695 161.405 ;
        RECT 83.915 160.595 84.425 161.130 ;
        RECT 84.605 160.765 84.795 162.125 ;
        RECT 84.965 161.445 85.240 161.925 ;
        RECT 84.965 161.275 85.245 161.445 ;
        RECT 85.445 161.325 85.615 162.125 ;
        RECT 85.785 161.335 85.955 162.465 ;
        RECT 86.125 161.835 86.295 162.805 ;
        RECT 86.465 162.005 86.635 163.145 ;
        RECT 86.805 162.005 87.140 162.975 ;
        RECT 86.125 161.505 86.320 161.835 ;
        RECT 86.545 161.505 86.800 161.835 ;
        RECT 86.545 161.335 86.715 161.505 ;
        RECT 86.970 161.335 87.140 162.005 ;
        RECT 87.315 161.980 87.605 163.145 ;
        RECT 87.775 162.005 88.160 162.975 ;
        RECT 88.330 162.685 88.655 163.145 ;
        RECT 89.175 162.515 89.455 162.975 ;
        RECT 88.330 162.295 89.455 162.515 ;
        RECT 84.965 160.765 85.240 161.275 ;
        RECT 85.785 161.165 86.715 161.335 ;
        RECT 85.785 161.130 85.960 161.165 ;
        RECT 85.430 160.765 85.960 161.130 ;
        RECT 86.385 160.595 86.715 160.995 ;
        RECT 86.885 160.765 87.140 161.335 ;
        RECT 87.775 161.335 88.055 162.005 ;
        RECT 88.330 161.835 88.780 162.295 ;
        RECT 89.645 162.125 90.045 162.975 ;
        RECT 90.445 162.685 90.715 163.145 ;
        RECT 90.885 162.515 91.170 162.975 ;
        RECT 88.225 161.505 88.780 161.835 ;
        RECT 88.950 161.565 90.045 162.125 ;
        RECT 88.330 161.395 88.780 161.505 ;
        RECT 87.315 160.595 87.605 161.320 ;
        RECT 87.775 160.765 88.160 161.335 ;
        RECT 88.330 161.225 89.455 161.395 ;
        RECT 88.330 160.595 88.655 161.055 ;
        RECT 89.175 160.765 89.455 161.225 ;
        RECT 89.645 160.765 90.045 161.565 ;
        RECT 90.215 162.295 91.170 162.515 ;
        RECT 90.215 161.395 90.425 162.295 ;
        RECT 90.595 161.565 91.285 162.125 ;
        RECT 91.455 162.070 91.725 162.975 ;
        RECT 91.895 162.385 92.225 163.145 ;
        RECT 92.405 162.215 92.575 162.975 ;
        RECT 90.215 161.225 91.170 161.395 ;
        RECT 90.445 160.595 90.715 161.055 ;
        RECT 90.885 160.765 91.170 161.225 ;
        RECT 91.455 161.270 91.625 162.070 ;
        RECT 91.910 162.045 92.575 162.215 ;
        RECT 92.835 162.385 93.350 162.795 ;
        RECT 93.585 162.385 93.755 163.145 ;
        RECT 93.925 162.805 95.955 162.975 ;
        RECT 91.910 161.900 92.080 162.045 ;
        RECT 91.795 161.570 92.080 161.900 ;
        RECT 91.910 161.315 92.080 161.570 ;
        RECT 92.315 161.495 92.645 161.865 ;
        RECT 92.835 161.575 93.175 162.385 ;
        RECT 93.925 162.140 94.095 162.805 ;
        RECT 94.490 162.465 95.615 162.635 ;
        RECT 93.345 161.950 94.095 162.140 ;
        RECT 94.265 162.125 95.275 162.295 ;
        RECT 92.835 161.405 94.065 161.575 ;
        RECT 91.455 160.765 91.715 161.270 ;
        RECT 91.910 161.145 92.575 161.315 ;
        RECT 91.895 160.595 92.225 160.975 ;
        RECT 92.405 160.765 92.575 161.145 ;
        RECT 93.110 160.800 93.355 161.405 ;
        RECT 93.575 160.595 94.085 161.130 ;
        RECT 94.265 160.765 94.455 162.125 ;
        RECT 94.625 161.785 94.900 161.925 ;
        RECT 94.625 161.615 94.905 161.785 ;
        RECT 94.625 160.765 94.900 161.615 ;
        RECT 95.105 161.325 95.275 162.125 ;
        RECT 95.445 161.335 95.615 162.465 ;
        RECT 95.785 161.835 95.955 162.805 ;
        RECT 96.125 162.005 96.295 163.145 ;
        RECT 96.465 162.005 96.800 162.975 ;
        RECT 95.785 161.505 95.980 161.835 ;
        RECT 96.205 161.505 96.460 161.835 ;
        RECT 96.205 161.335 96.375 161.505 ;
        RECT 96.630 161.335 96.800 162.005 ;
        RECT 95.445 161.165 96.375 161.335 ;
        RECT 95.445 161.130 95.620 161.165 ;
        RECT 95.090 160.765 95.620 161.130 ;
        RECT 96.045 160.595 96.375 160.995 ;
        RECT 96.545 160.765 96.800 161.335 ;
        RECT 97.435 162.005 97.820 162.975 ;
        RECT 97.990 162.685 98.315 163.145 ;
        RECT 98.835 162.515 99.115 162.975 ;
        RECT 97.990 162.295 99.115 162.515 ;
        RECT 97.435 161.335 97.715 162.005 ;
        RECT 97.990 161.835 98.440 162.295 ;
        RECT 99.305 162.125 99.705 162.975 ;
        RECT 100.105 162.685 100.375 163.145 ;
        RECT 100.545 162.515 100.830 162.975 ;
        RECT 97.885 161.505 98.440 161.835 ;
        RECT 98.610 161.565 99.705 162.125 ;
        RECT 97.990 161.395 98.440 161.505 ;
        RECT 97.435 160.765 97.820 161.335 ;
        RECT 97.990 161.225 99.115 161.395 ;
        RECT 97.990 160.595 98.315 161.055 ;
        RECT 98.835 160.765 99.115 161.225 ;
        RECT 99.305 160.765 99.705 161.565 ;
        RECT 99.875 162.295 100.830 162.515 ;
        RECT 101.115 162.385 101.630 162.795 ;
        RECT 101.865 162.385 102.035 163.145 ;
        RECT 102.205 162.805 104.235 162.975 ;
        RECT 99.875 161.395 100.085 162.295 ;
        RECT 100.255 161.565 100.945 162.125 ;
        RECT 101.115 161.575 101.455 162.385 ;
        RECT 102.205 162.140 102.375 162.805 ;
        RECT 102.770 162.465 103.895 162.635 ;
        RECT 101.625 161.950 102.375 162.140 ;
        RECT 102.545 162.125 103.555 162.295 ;
        RECT 101.115 161.405 102.345 161.575 ;
        RECT 99.875 161.225 100.830 161.395 ;
        RECT 100.105 160.595 100.375 161.055 ;
        RECT 100.545 160.765 100.830 161.225 ;
        RECT 101.390 160.800 101.635 161.405 ;
        RECT 101.855 160.595 102.365 161.130 ;
        RECT 102.545 160.765 102.735 162.125 ;
        RECT 102.905 161.785 103.180 161.925 ;
        RECT 102.905 161.615 103.185 161.785 ;
        RECT 102.905 160.765 103.180 161.615 ;
        RECT 103.385 161.325 103.555 162.125 ;
        RECT 103.725 161.335 103.895 162.465 ;
        RECT 104.065 161.835 104.235 162.805 ;
        RECT 104.405 162.005 104.575 163.145 ;
        RECT 104.745 162.005 105.080 162.975 ;
        RECT 105.370 162.515 105.655 162.975 ;
        RECT 105.825 162.685 106.095 163.145 ;
        RECT 105.370 162.295 106.325 162.515 ;
        RECT 104.065 161.505 104.260 161.835 ;
        RECT 104.485 161.505 104.740 161.835 ;
        RECT 104.485 161.335 104.655 161.505 ;
        RECT 104.910 161.335 105.080 162.005 ;
        RECT 105.255 161.565 105.945 162.125 ;
        RECT 106.115 161.395 106.325 162.295 ;
        RECT 103.725 161.165 104.655 161.335 ;
        RECT 103.725 161.130 103.900 161.165 ;
        RECT 103.370 160.765 103.900 161.130 ;
        RECT 104.325 160.595 104.655 160.995 ;
        RECT 104.825 160.765 105.080 161.335 ;
        RECT 105.370 161.225 106.325 161.395 ;
        RECT 106.495 162.125 106.895 162.975 ;
        RECT 107.085 162.515 107.365 162.975 ;
        RECT 107.885 162.685 108.210 163.145 ;
        RECT 107.085 162.295 108.210 162.515 ;
        RECT 106.495 161.565 107.590 162.125 ;
        RECT 107.760 161.835 108.210 162.295 ;
        RECT 108.380 162.005 108.765 162.975 ;
        RECT 105.370 160.765 105.655 161.225 ;
        RECT 105.825 160.595 106.095 161.055 ;
        RECT 106.495 160.765 106.895 161.565 ;
        RECT 107.760 161.505 108.315 161.835 ;
        RECT 107.760 161.395 108.210 161.505 ;
        RECT 107.085 161.225 108.210 161.395 ;
        RECT 108.485 161.335 108.765 162.005 ;
        RECT 108.945 162.165 109.275 162.975 ;
        RECT 109.445 162.345 109.685 163.145 ;
        RECT 108.945 161.995 109.660 162.165 ;
        RECT 108.940 161.585 109.320 161.825 ;
        RECT 109.490 161.755 109.660 161.995 ;
        RECT 109.865 162.125 110.035 162.975 ;
        RECT 110.205 162.345 110.535 163.145 ;
        RECT 110.705 162.125 110.875 162.975 ;
        RECT 109.865 161.955 110.875 162.125 ;
        RECT 111.045 161.995 111.375 163.145 ;
        RECT 112.155 162.055 113.365 163.145 ;
        RECT 109.490 161.585 109.990 161.755 ;
        RECT 109.490 161.415 109.660 161.585 ;
        RECT 110.380 161.445 110.875 161.955 ;
        RECT 112.155 161.515 112.675 162.055 ;
        RECT 110.375 161.415 110.875 161.445 ;
        RECT 107.085 160.765 107.365 161.225 ;
        RECT 107.885 160.595 108.210 161.055 ;
        RECT 108.380 160.765 108.765 161.335 ;
        RECT 109.025 161.245 109.660 161.415 ;
        RECT 109.865 161.245 110.875 161.415 ;
        RECT 109.025 160.765 109.195 161.245 ;
        RECT 109.375 160.595 109.615 161.075 ;
        RECT 109.865 160.765 110.035 161.245 ;
        RECT 110.205 160.595 110.535 161.075 ;
        RECT 110.705 160.765 110.875 161.245 ;
        RECT 111.045 160.595 111.375 161.395 ;
        RECT 112.845 161.345 113.365 161.885 ;
        RECT 112.155 160.595 113.365 161.345 ;
        RECT 11.330 160.425 113.450 160.595 ;
        RECT 11.415 159.675 12.625 160.425 ;
        RECT 13.345 159.875 13.515 160.165 ;
        RECT 13.685 160.045 14.015 160.425 ;
        RECT 13.345 159.705 14.010 159.875 ;
        RECT 11.415 159.135 11.935 159.675 ;
        RECT 12.105 158.965 12.625 159.505 ;
        RECT 11.415 157.875 12.625 158.965 ;
        RECT 13.260 158.885 13.610 159.535 ;
        RECT 13.780 158.715 14.010 159.705 ;
        RECT 13.345 158.545 14.010 158.715 ;
        RECT 13.345 158.045 13.515 158.545 ;
        RECT 13.685 157.875 14.015 158.375 ;
        RECT 14.185 158.045 14.410 160.165 ;
        RECT 14.625 160.045 14.955 160.425 ;
        RECT 15.125 159.875 15.295 160.205 ;
        RECT 15.595 160.045 16.610 160.245 ;
        RECT 14.600 159.685 15.295 159.875 ;
        RECT 14.600 158.715 14.770 159.685 ;
        RECT 14.940 158.885 15.350 159.505 ;
        RECT 15.520 158.935 15.740 159.805 ;
        RECT 15.920 159.495 16.270 159.865 ;
        RECT 16.440 159.315 16.610 160.045 ;
        RECT 16.780 159.985 17.190 160.425 ;
        RECT 17.480 159.785 17.730 160.215 ;
        RECT 17.930 159.965 18.250 160.425 ;
        RECT 18.810 160.035 19.660 160.205 ;
        RECT 16.780 159.445 17.190 159.775 ;
        RECT 17.480 159.445 17.900 159.785 ;
        RECT 16.190 159.275 16.610 159.315 ;
        RECT 16.190 159.105 17.540 159.275 ;
        RECT 14.600 158.545 15.295 158.715 ;
        RECT 15.520 158.555 16.020 158.935 ;
        RECT 14.625 157.875 14.955 158.375 ;
        RECT 15.125 158.045 15.295 158.545 ;
        RECT 16.190 158.260 16.360 159.105 ;
        RECT 17.290 158.945 17.540 159.105 ;
        RECT 16.530 158.675 16.780 158.935 ;
        RECT 17.710 158.675 17.900 159.445 ;
        RECT 16.530 158.425 17.900 158.675 ;
        RECT 18.070 159.615 19.320 159.785 ;
        RECT 18.070 158.855 18.240 159.615 ;
        RECT 18.990 159.495 19.320 159.615 ;
        RECT 18.410 159.035 18.590 159.445 ;
        RECT 19.490 159.275 19.660 160.035 ;
        RECT 19.860 159.945 20.520 160.425 ;
        RECT 20.700 159.830 21.020 160.160 ;
        RECT 19.850 159.505 20.510 159.775 ;
        RECT 19.850 159.445 20.180 159.505 ;
        RECT 20.330 159.275 20.660 159.335 ;
        RECT 18.760 159.105 20.660 159.275 ;
        RECT 18.070 158.545 18.590 158.855 ;
        RECT 18.760 158.595 18.930 159.105 ;
        RECT 20.830 158.935 21.020 159.830 ;
        RECT 19.100 158.765 21.020 158.935 ;
        RECT 20.700 158.745 21.020 158.765 ;
        RECT 21.220 159.515 21.470 160.165 ;
        RECT 21.650 159.965 21.935 160.425 ;
        RECT 22.115 159.715 22.370 160.245 ;
        RECT 21.220 159.185 22.020 159.515 ;
        RECT 18.760 158.425 19.970 158.595 ;
        RECT 15.530 158.090 16.360 158.260 ;
        RECT 16.600 157.875 16.980 158.255 ;
        RECT 17.160 158.135 17.330 158.425 ;
        RECT 18.760 158.345 18.930 158.425 ;
        RECT 17.500 157.875 17.830 158.255 ;
        RECT 18.300 158.095 18.930 158.345 ;
        RECT 19.110 157.875 19.530 158.255 ;
        RECT 19.730 158.135 19.970 158.425 ;
        RECT 20.200 157.875 20.530 158.565 ;
        RECT 20.700 158.135 20.870 158.745 ;
        RECT 21.220 158.595 21.470 159.185 ;
        RECT 22.190 158.855 22.370 159.715 ;
        RECT 22.915 159.700 23.205 160.425 ;
        RECT 23.465 159.875 23.635 160.255 ;
        RECT 23.815 160.045 24.145 160.425 ;
        RECT 23.465 159.705 24.130 159.875 ;
        RECT 24.325 159.750 24.585 160.255 ;
        RECT 23.395 159.155 23.725 159.525 ;
        RECT 23.960 159.450 24.130 159.705 ;
        RECT 23.960 159.120 24.245 159.450 ;
        RECT 21.140 158.085 21.470 158.595 ;
        RECT 21.650 157.875 21.935 158.675 ;
        RECT 22.115 158.385 22.370 158.855 ;
        RECT 22.115 158.215 22.455 158.385 ;
        RECT 22.115 158.185 22.370 158.215 ;
        RECT 22.915 157.875 23.205 159.040 ;
        RECT 23.960 158.975 24.130 159.120 ;
        RECT 23.465 158.805 24.130 158.975 ;
        RECT 24.415 158.950 24.585 159.750 ;
        RECT 23.465 158.045 23.635 158.805 ;
        RECT 23.815 157.875 24.145 158.635 ;
        RECT 24.315 158.045 24.585 158.950 ;
        RECT 24.755 159.685 25.140 160.255 ;
        RECT 25.310 159.965 25.635 160.425 ;
        RECT 26.155 159.795 26.435 160.255 ;
        RECT 24.755 159.015 25.035 159.685 ;
        RECT 25.310 159.625 26.435 159.795 ;
        RECT 25.310 159.515 25.760 159.625 ;
        RECT 25.205 159.185 25.760 159.515 ;
        RECT 26.625 159.455 27.025 160.255 ;
        RECT 27.425 159.965 27.695 160.425 ;
        RECT 27.865 159.795 28.150 160.255 ;
        RECT 24.755 158.045 25.140 159.015 ;
        RECT 25.310 158.725 25.760 159.185 ;
        RECT 25.930 158.895 27.025 159.455 ;
        RECT 25.310 158.505 26.435 158.725 ;
        RECT 25.310 157.875 25.635 158.335 ;
        RECT 26.155 158.045 26.435 158.505 ;
        RECT 26.625 158.045 27.025 158.895 ;
        RECT 27.195 159.625 28.150 159.795 ;
        RECT 28.640 159.645 29.140 160.255 ;
        RECT 27.195 158.725 27.405 159.625 ;
        RECT 27.575 158.895 28.265 159.455 ;
        RECT 28.435 159.185 28.785 159.435 ;
        RECT 28.970 159.015 29.140 159.645 ;
        RECT 29.770 159.775 30.100 160.255 ;
        RECT 30.270 159.965 30.495 160.425 ;
        RECT 30.665 159.775 30.995 160.255 ;
        RECT 29.770 159.605 30.995 159.775 ;
        RECT 31.185 159.625 31.435 160.425 ;
        RECT 31.605 159.625 31.945 160.255 ;
        RECT 29.310 159.235 29.640 159.435 ;
        RECT 29.810 159.235 30.140 159.435 ;
        RECT 30.310 159.235 30.730 159.435 ;
        RECT 30.905 159.265 31.600 159.435 ;
        RECT 30.905 159.015 31.075 159.265 ;
        RECT 31.770 159.015 31.945 159.625 ;
        RECT 32.155 159.605 32.385 160.425 ;
        RECT 32.555 159.625 32.885 160.255 ;
        RECT 32.135 159.185 32.465 159.435 ;
        RECT 32.635 159.025 32.885 159.625 ;
        RECT 33.055 159.605 33.265 160.425 ;
        RECT 33.610 159.795 33.895 160.255 ;
        RECT 34.065 159.965 34.335 160.425 ;
        RECT 33.610 159.625 34.565 159.795 ;
        RECT 28.640 158.845 31.075 159.015 ;
        RECT 27.195 158.505 28.150 158.725 ;
        RECT 27.425 157.875 27.695 158.335 ;
        RECT 27.865 158.045 28.150 158.505 ;
        RECT 28.640 158.045 28.970 158.845 ;
        RECT 29.140 157.875 29.470 158.675 ;
        RECT 29.770 158.045 30.100 158.845 ;
        RECT 30.745 157.875 30.995 158.675 ;
        RECT 31.265 157.875 31.435 159.015 ;
        RECT 31.605 158.045 31.945 159.015 ;
        RECT 32.155 157.875 32.385 159.015 ;
        RECT 32.555 158.045 32.885 159.025 ;
        RECT 33.055 157.875 33.265 159.015 ;
        RECT 33.495 158.895 34.185 159.455 ;
        RECT 34.355 158.725 34.565 159.625 ;
        RECT 33.610 158.505 34.565 158.725 ;
        RECT 34.735 159.455 35.135 160.255 ;
        RECT 35.325 159.795 35.605 160.255 ;
        RECT 36.125 159.965 36.450 160.425 ;
        RECT 35.325 159.625 36.450 159.795 ;
        RECT 36.620 159.685 37.005 160.255 ;
        RECT 36.000 159.515 36.450 159.625 ;
        RECT 34.735 158.895 35.830 159.455 ;
        RECT 36.000 159.185 36.555 159.515 ;
        RECT 33.610 158.045 33.895 158.505 ;
        RECT 34.065 157.875 34.335 158.335 ;
        RECT 34.735 158.045 35.135 158.895 ;
        RECT 36.000 158.725 36.450 159.185 ;
        RECT 36.725 159.015 37.005 159.685 ;
        RECT 37.290 159.795 37.575 160.255 ;
        RECT 37.745 159.965 38.015 160.425 ;
        RECT 37.290 159.625 38.245 159.795 ;
        RECT 35.325 158.505 36.450 158.725 ;
        RECT 35.325 158.045 35.605 158.505 ;
        RECT 36.125 157.875 36.450 158.335 ;
        RECT 36.620 158.045 37.005 159.015 ;
        RECT 37.175 158.895 37.865 159.455 ;
        RECT 38.035 158.725 38.245 159.625 ;
        RECT 37.290 158.505 38.245 158.725 ;
        RECT 38.415 159.455 38.815 160.255 ;
        RECT 39.005 159.795 39.285 160.255 ;
        RECT 39.805 159.965 40.130 160.425 ;
        RECT 39.005 159.625 40.130 159.795 ;
        RECT 40.300 159.685 40.685 160.255 ;
        RECT 39.680 159.515 40.130 159.625 ;
        RECT 38.415 158.895 39.510 159.455 ;
        RECT 39.680 159.185 40.235 159.515 ;
        RECT 37.290 158.045 37.575 158.505 ;
        RECT 37.745 157.875 38.015 158.335 ;
        RECT 38.415 158.045 38.815 158.895 ;
        RECT 39.680 158.725 40.130 159.185 ;
        RECT 40.405 159.015 40.685 159.685 ;
        RECT 39.005 158.505 40.130 158.725 ;
        RECT 39.005 158.045 39.285 158.505 ;
        RECT 39.805 157.875 40.130 158.335 ;
        RECT 40.300 158.045 40.685 159.015 ;
        RECT 40.860 159.685 41.115 160.255 ;
        RECT 41.285 160.025 41.615 160.425 ;
        RECT 42.040 159.890 42.570 160.255 ;
        RECT 42.040 159.855 42.215 159.890 ;
        RECT 41.285 159.685 42.215 159.855 ;
        RECT 42.760 159.745 43.035 160.255 ;
        RECT 40.860 159.015 41.030 159.685 ;
        RECT 41.285 159.515 41.455 159.685 ;
        RECT 41.200 159.185 41.455 159.515 ;
        RECT 41.680 159.185 41.875 159.515 ;
        RECT 40.860 158.045 41.195 159.015 ;
        RECT 41.365 157.875 41.535 159.015 ;
        RECT 41.705 158.215 41.875 159.185 ;
        RECT 42.045 158.555 42.215 159.685 ;
        RECT 42.385 158.895 42.555 159.695 ;
        RECT 42.755 159.575 43.035 159.745 ;
        RECT 42.760 159.095 43.035 159.575 ;
        RECT 43.205 158.895 43.395 160.255 ;
        RECT 43.575 159.890 44.085 160.425 ;
        RECT 44.305 159.615 44.550 160.220 ;
        RECT 45.460 159.660 45.915 160.425 ;
        RECT 46.190 160.045 47.490 160.255 ;
        RECT 47.745 160.065 48.075 160.425 ;
        RECT 47.320 159.895 47.490 160.045 ;
        RECT 48.245 159.925 48.505 160.255 ;
        RECT 43.595 159.445 44.825 159.615 ;
        RECT 42.385 158.725 43.395 158.895 ;
        RECT 43.565 158.880 44.315 159.070 ;
        RECT 42.045 158.385 43.170 158.555 ;
        RECT 43.565 158.215 43.735 158.880 ;
        RECT 44.485 158.635 44.825 159.445 ;
        RECT 46.390 159.435 46.610 159.835 ;
        RECT 45.455 159.235 45.945 159.435 ;
        RECT 46.135 159.225 46.610 159.435 ;
        RECT 46.855 159.435 47.065 159.835 ;
        RECT 47.320 159.770 48.075 159.895 ;
        RECT 47.320 159.725 48.165 159.770 ;
        RECT 47.895 159.605 48.165 159.725 ;
        RECT 46.855 159.225 47.185 159.435 ;
        RECT 47.355 159.165 47.765 159.470 ;
        RECT 41.705 158.045 43.735 158.215 ;
        RECT 43.905 157.875 44.075 158.635 ;
        RECT 44.310 158.225 44.825 158.635 ;
        RECT 45.460 158.995 46.635 159.055 ;
        RECT 47.995 159.030 48.165 159.605 ;
        RECT 47.965 158.995 48.165 159.030 ;
        RECT 45.460 158.885 48.165 158.995 ;
        RECT 45.460 158.265 45.715 158.885 ;
        RECT 46.305 158.825 48.105 158.885 ;
        RECT 46.305 158.795 46.635 158.825 ;
        RECT 48.335 158.725 48.505 159.925 ;
        RECT 48.675 159.700 48.965 160.425 ;
        RECT 50.095 159.605 50.325 160.425 ;
        RECT 50.495 159.625 50.825 160.255 ;
        RECT 50.075 159.185 50.405 159.435 ;
        RECT 45.965 158.625 46.150 158.715 ;
        RECT 46.740 158.625 47.575 158.635 ;
        RECT 45.965 158.425 47.575 158.625 ;
        RECT 45.965 158.385 46.195 158.425 ;
        RECT 45.460 158.045 45.795 158.265 ;
        RECT 46.800 157.875 47.155 158.255 ;
        RECT 47.325 158.045 47.575 158.425 ;
        RECT 47.825 157.875 48.075 158.655 ;
        RECT 48.245 158.045 48.505 158.725 ;
        RECT 48.675 157.875 48.965 159.040 ;
        RECT 50.575 159.025 50.825 159.625 ;
        RECT 50.995 159.605 51.205 160.425 ;
        RECT 51.435 159.625 51.775 160.255 ;
        RECT 51.945 159.625 52.195 160.425 ;
        RECT 52.385 159.775 52.715 160.255 ;
        RECT 52.885 159.965 53.110 160.425 ;
        RECT 53.280 159.775 53.610 160.255 ;
        RECT 50.095 157.875 50.325 159.015 ;
        RECT 50.495 158.045 50.825 159.025 ;
        RECT 51.435 159.065 51.610 159.625 ;
        RECT 52.385 159.605 53.610 159.775 ;
        RECT 54.240 159.645 54.740 160.255 ;
        RECT 55.490 159.715 55.745 160.245 ;
        RECT 55.925 159.965 56.210 160.425 ;
        RECT 51.780 159.265 52.475 159.435 ;
        RECT 51.435 159.015 51.665 159.065 ;
        RECT 52.305 159.015 52.475 159.265 ;
        RECT 52.650 159.235 53.070 159.435 ;
        RECT 53.240 159.235 53.570 159.435 ;
        RECT 53.740 159.235 54.070 159.435 ;
        RECT 54.240 159.015 54.410 159.645 ;
        RECT 54.595 159.185 54.945 159.435 ;
        RECT 55.490 159.065 55.670 159.715 ;
        RECT 56.390 159.515 56.640 160.165 ;
        RECT 55.840 159.185 56.640 159.515 ;
        RECT 50.995 157.875 51.205 159.015 ;
        RECT 51.435 158.045 51.775 159.015 ;
        RECT 51.945 157.875 52.115 159.015 ;
        RECT 52.305 158.845 54.740 159.015 ;
        RECT 55.405 158.895 55.670 159.065 ;
        RECT 52.385 157.875 52.635 158.675 ;
        RECT 53.280 158.045 53.610 158.845 ;
        RECT 53.910 157.875 54.240 158.675 ;
        RECT 54.410 158.045 54.740 158.845 ;
        RECT 55.490 158.855 55.670 158.895 ;
        RECT 55.490 158.185 55.745 158.855 ;
        RECT 55.925 157.875 56.210 158.675 ;
        RECT 56.390 158.595 56.640 159.185 ;
        RECT 56.840 159.830 57.160 160.160 ;
        RECT 57.340 159.945 58.000 160.425 ;
        RECT 58.200 160.035 59.050 160.205 ;
        RECT 56.840 158.935 57.030 159.830 ;
        RECT 57.350 159.505 58.010 159.775 ;
        RECT 57.680 159.445 58.010 159.505 ;
        RECT 57.200 159.275 57.530 159.335 ;
        RECT 58.200 159.275 58.370 160.035 ;
        RECT 59.610 159.965 59.930 160.425 ;
        RECT 60.130 159.785 60.380 160.215 ;
        RECT 60.670 159.985 61.080 160.425 ;
        RECT 61.250 160.045 62.265 160.245 ;
        RECT 58.540 159.615 59.790 159.785 ;
        RECT 58.540 159.495 58.870 159.615 ;
        RECT 57.200 159.105 59.100 159.275 ;
        RECT 56.840 158.765 58.760 158.935 ;
        RECT 56.840 158.745 57.160 158.765 ;
        RECT 56.390 158.085 56.720 158.595 ;
        RECT 56.990 158.135 57.160 158.745 ;
        RECT 58.930 158.595 59.100 159.105 ;
        RECT 59.270 159.035 59.450 159.445 ;
        RECT 59.620 158.855 59.790 159.615 ;
        RECT 57.330 157.875 57.660 158.565 ;
        RECT 57.890 158.425 59.100 158.595 ;
        RECT 59.270 158.545 59.790 158.855 ;
        RECT 59.960 159.445 60.380 159.785 ;
        RECT 60.670 159.445 61.080 159.775 ;
        RECT 59.960 158.675 60.150 159.445 ;
        RECT 61.250 159.315 61.420 160.045 ;
        RECT 62.565 159.875 62.735 160.205 ;
        RECT 62.905 160.045 63.235 160.425 ;
        RECT 61.590 159.495 61.940 159.865 ;
        RECT 61.250 159.275 61.670 159.315 ;
        RECT 60.320 159.105 61.670 159.275 ;
        RECT 60.320 158.945 60.570 159.105 ;
        RECT 61.080 158.675 61.330 158.935 ;
        RECT 59.960 158.425 61.330 158.675 ;
        RECT 57.890 158.135 58.130 158.425 ;
        RECT 58.930 158.345 59.100 158.425 ;
        RECT 58.330 157.875 58.750 158.255 ;
        RECT 58.930 158.095 59.560 158.345 ;
        RECT 60.030 157.875 60.360 158.255 ;
        RECT 60.530 158.135 60.700 158.425 ;
        RECT 61.500 158.260 61.670 159.105 ;
        RECT 62.120 158.935 62.340 159.805 ;
        RECT 62.565 159.685 63.260 159.875 ;
        RECT 61.840 158.555 62.340 158.935 ;
        RECT 62.510 158.885 62.920 159.505 ;
        RECT 63.090 158.715 63.260 159.685 ;
        RECT 62.565 158.545 63.260 158.715 ;
        RECT 60.880 157.875 61.260 158.255 ;
        RECT 61.500 158.090 62.330 158.260 ;
        RECT 62.565 158.045 62.735 158.545 ;
        RECT 62.905 157.875 63.235 158.375 ;
        RECT 63.450 158.045 63.675 160.165 ;
        RECT 63.845 160.045 64.175 160.425 ;
        RECT 64.345 159.875 64.515 160.165 ;
        RECT 63.850 159.705 64.515 159.875 ;
        RECT 63.850 158.715 64.080 159.705 ;
        RECT 64.775 159.675 65.985 160.425 ;
        RECT 64.250 158.885 64.600 159.535 ;
        RECT 64.775 158.965 65.295 159.505 ;
        RECT 65.465 159.135 65.985 159.675 ;
        RECT 66.430 159.615 66.675 160.220 ;
        RECT 66.895 159.890 67.405 160.425 ;
        RECT 66.155 159.445 67.385 159.615 ;
        RECT 63.850 158.545 64.515 158.715 ;
        RECT 63.845 157.875 64.175 158.375 ;
        RECT 64.345 158.045 64.515 158.545 ;
        RECT 64.775 157.875 65.985 158.965 ;
        RECT 66.155 158.635 66.495 159.445 ;
        RECT 66.665 158.880 67.415 159.070 ;
        RECT 66.155 158.225 66.670 158.635 ;
        RECT 66.905 157.875 67.075 158.635 ;
        RECT 67.245 158.215 67.415 158.880 ;
        RECT 67.585 158.895 67.775 160.255 ;
        RECT 67.945 159.745 68.220 160.255 ;
        RECT 68.410 159.890 68.940 160.255 ;
        RECT 69.365 160.025 69.695 160.425 ;
        RECT 68.765 159.855 68.940 159.890 ;
        RECT 67.945 159.575 68.225 159.745 ;
        RECT 67.945 159.095 68.220 159.575 ;
        RECT 68.425 158.895 68.595 159.695 ;
        RECT 67.585 158.725 68.595 158.895 ;
        RECT 68.765 159.685 69.695 159.855 ;
        RECT 69.865 159.685 70.120 160.255 ;
        RECT 68.765 158.555 68.935 159.685 ;
        RECT 69.525 159.515 69.695 159.685 ;
        RECT 67.810 158.385 68.935 158.555 ;
        RECT 69.105 159.185 69.300 159.515 ;
        RECT 69.525 159.185 69.780 159.515 ;
        RECT 69.105 158.215 69.275 159.185 ;
        RECT 69.950 159.015 70.120 159.685 ;
        RECT 70.570 159.615 70.815 160.220 ;
        RECT 71.035 159.890 71.545 160.425 ;
        RECT 67.245 158.045 69.275 158.215 ;
        RECT 69.445 157.875 69.615 159.015 ;
        RECT 69.785 158.045 70.120 159.015 ;
        RECT 70.295 159.445 71.525 159.615 ;
        RECT 70.295 158.635 70.635 159.445 ;
        RECT 70.805 158.880 71.555 159.070 ;
        RECT 70.295 158.225 70.810 158.635 ;
        RECT 71.045 157.875 71.215 158.635 ;
        RECT 71.385 158.215 71.555 158.880 ;
        RECT 71.725 158.895 71.915 160.255 ;
        RECT 72.085 159.745 72.360 160.255 ;
        RECT 72.550 159.890 73.080 160.255 ;
        RECT 73.505 160.025 73.835 160.425 ;
        RECT 72.905 159.855 73.080 159.890 ;
        RECT 72.085 159.575 72.365 159.745 ;
        RECT 72.085 159.095 72.360 159.575 ;
        RECT 72.565 158.895 72.735 159.695 ;
        RECT 71.725 158.725 72.735 158.895 ;
        RECT 72.905 159.685 73.835 159.855 ;
        RECT 74.005 159.685 74.260 160.255 ;
        RECT 74.435 159.700 74.725 160.425 ;
        RECT 75.445 159.875 75.615 160.255 ;
        RECT 75.795 160.045 76.125 160.425 ;
        RECT 75.445 159.705 76.110 159.875 ;
        RECT 76.305 159.750 76.565 160.255 ;
        RECT 72.905 158.555 73.075 159.685 ;
        RECT 73.665 159.515 73.835 159.685 ;
        RECT 71.950 158.385 73.075 158.555 ;
        RECT 73.245 159.185 73.440 159.515 ;
        RECT 73.665 159.185 73.920 159.515 ;
        RECT 73.245 158.215 73.415 159.185 ;
        RECT 74.090 159.015 74.260 159.685 ;
        RECT 75.375 159.155 75.705 159.525 ;
        RECT 75.940 159.450 76.110 159.705 ;
        RECT 75.940 159.120 76.225 159.450 ;
        RECT 71.385 158.045 73.415 158.215 ;
        RECT 73.585 157.875 73.755 159.015 ;
        RECT 73.925 158.045 74.260 159.015 ;
        RECT 74.435 157.875 74.725 159.040 ;
        RECT 75.940 158.975 76.110 159.120 ;
        RECT 75.445 158.805 76.110 158.975 ;
        RECT 76.395 158.950 76.565 159.750 ;
        RECT 75.445 158.045 75.615 158.805 ;
        RECT 75.795 157.875 76.125 158.635 ;
        RECT 76.295 158.045 76.565 158.950 ;
        RECT 77.570 159.715 77.825 160.245 ;
        RECT 78.005 159.965 78.290 160.425 ;
        RECT 77.570 158.855 77.750 159.715 ;
        RECT 78.470 159.515 78.720 160.165 ;
        RECT 77.920 159.185 78.720 159.515 ;
        RECT 77.570 158.725 77.825 158.855 ;
        RECT 77.485 158.555 77.825 158.725 ;
        RECT 77.570 158.185 77.825 158.555 ;
        RECT 78.005 157.875 78.290 158.675 ;
        RECT 78.470 158.595 78.720 159.185 ;
        RECT 78.920 159.830 79.240 160.160 ;
        RECT 79.420 159.945 80.080 160.425 ;
        RECT 80.280 160.035 81.130 160.205 ;
        RECT 78.920 158.935 79.110 159.830 ;
        RECT 79.430 159.505 80.090 159.775 ;
        RECT 79.760 159.445 80.090 159.505 ;
        RECT 79.280 159.275 79.610 159.335 ;
        RECT 80.280 159.275 80.450 160.035 ;
        RECT 81.690 159.965 82.010 160.425 ;
        RECT 82.210 159.785 82.460 160.215 ;
        RECT 82.750 159.985 83.160 160.425 ;
        RECT 83.330 160.045 84.345 160.245 ;
        RECT 80.620 159.615 81.870 159.785 ;
        RECT 80.620 159.495 80.950 159.615 ;
        RECT 79.280 159.105 81.180 159.275 ;
        RECT 78.920 158.765 80.840 158.935 ;
        RECT 78.920 158.745 79.240 158.765 ;
        RECT 78.470 158.085 78.800 158.595 ;
        RECT 79.070 158.135 79.240 158.745 ;
        RECT 81.010 158.595 81.180 159.105 ;
        RECT 81.350 159.035 81.530 159.445 ;
        RECT 81.700 158.855 81.870 159.615 ;
        RECT 79.410 157.875 79.740 158.565 ;
        RECT 79.970 158.425 81.180 158.595 ;
        RECT 81.350 158.545 81.870 158.855 ;
        RECT 82.040 159.445 82.460 159.785 ;
        RECT 82.750 159.445 83.160 159.775 ;
        RECT 82.040 158.675 82.230 159.445 ;
        RECT 83.330 159.315 83.500 160.045 ;
        RECT 84.645 159.875 84.815 160.205 ;
        RECT 84.985 160.045 85.315 160.425 ;
        RECT 83.670 159.495 84.020 159.865 ;
        RECT 83.330 159.275 83.750 159.315 ;
        RECT 82.400 159.105 83.750 159.275 ;
        RECT 82.400 158.945 82.650 159.105 ;
        RECT 83.160 158.675 83.410 158.935 ;
        RECT 82.040 158.425 83.410 158.675 ;
        RECT 79.970 158.135 80.210 158.425 ;
        RECT 81.010 158.345 81.180 158.425 ;
        RECT 80.410 157.875 80.830 158.255 ;
        RECT 81.010 158.095 81.640 158.345 ;
        RECT 82.110 157.875 82.440 158.255 ;
        RECT 82.610 158.135 82.780 158.425 ;
        RECT 83.580 158.260 83.750 159.105 ;
        RECT 84.200 158.935 84.420 159.805 ;
        RECT 84.645 159.685 85.340 159.875 ;
        RECT 83.920 158.555 84.420 158.935 ;
        RECT 84.590 158.885 85.000 159.505 ;
        RECT 85.170 158.715 85.340 159.685 ;
        RECT 84.645 158.545 85.340 158.715 ;
        RECT 82.960 157.875 83.340 158.255 ;
        RECT 83.580 158.090 84.410 158.260 ;
        RECT 84.645 158.045 84.815 158.545 ;
        RECT 84.985 157.875 85.315 158.375 ;
        RECT 85.530 158.045 85.755 160.165 ;
        RECT 85.925 160.045 86.255 160.425 ;
        RECT 86.425 159.875 86.595 160.165 ;
        RECT 85.930 159.705 86.595 159.875 ;
        RECT 85.930 158.715 86.160 159.705 ;
        RECT 87.835 159.605 88.045 160.425 ;
        RECT 88.215 159.625 88.545 160.255 ;
        RECT 86.330 158.885 86.680 159.535 ;
        RECT 88.215 159.025 88.465 159.625 ;
        RECT 88.715 159.605 88.945 160.425 ;
        RECT 89.155 159.655 90.825 160.425 ;
        RECT 88.635 159.185 88.965 159.435 ;
        RECT 85.930 158.545 86.595 158.715 ;
        RECT 85.925 157.875 86.255 158.375 ;
        RECT 86.425 158.045 86.595 158.545 ;
        RECT 87.835 157.875 88.045 159.015 ;
        RECT 88.215 158.045 88.545 159.025 ;
        RECT 88.715 157.875 88.945 159.015 ;
        RECT 89.155 158.965 89.905 159.485 ;
        RECT 90.075 159.135 90.825 159.655 ;
        RECT 91.200 159.645 91.700 160.255 ;
        RECT 90.995 159.185 91.345 159.435 ;
        RECT 91.530 159.015 91.700 159.645 ;
        RECT 92.330 159.775 92.660 160.255 ;
        RECT 92.830 159.965 93.055 160.425 ;
        RECT 93.225 159.775 93.555 160.255 ;
        RECT 92.330 159.605 93.555 159.775 ;
        RECT 93.745 159.625 93.995 160.425 ;
        RECT 94.165 159.625 94.505 160.255 ;
        RECT 91.870 159.235 92.200 159.435 ;
        RECT 92.370 159.235 92.700 159.435 ;
        RECT 92.870 159.235 93.290 159.435 ;
        RECT 93.465 159.265 94.160 159.435 ;
        RECT 93.465 159.015 93.635 159.265 ;
        RECT 94.330 159.015 94.505 159.625 ;
        RECT 89.155 157.875 90.825 158.965 ;
        RECT 91.200 158.845 93.635 159.015 ;
        RECT 91.200 158.045 91.530 158.845 ;
        RECT 91.700 157.875 92.030 158.675 ;
        RECT 92.330 158.045 92.660 158.845 ;
        RECT 93.305 157.875 93.555 158.675 ;
        RECT 93.825 157.875 93.995 159.015 ;
        RECT 94.165 158.045 94.505 159.015 ;
        RECT 94.675 159.625 95.015 160.255 ;
        RECT 95.185 159.625 95.435 160.425 ;
        RECT 95.625 159.775 95.955 160.255 ;
        RECT 96.125 159.965 96.350 160.425 ;
        RECT 96.520 159.775 96.850 160.255 ;
        RECT 94.675 159.015 94.850 159.625 ;
        RECT 95.625 159.605 96.850 159.775 ;
        RECT 97.480 159.645 97.980 160.255 ;
        RECT 98.355 159.655 100.025 160.425 ;
        RECT 100.195 159.700 100.485 160.425 ;
        RECT 100.655 159.655 103.245 160.425 ;
        RECT 95.020 159.265 95.715 159.435 ;
        RECT 95.545 159.015 95.715 159.265 ;
        RECT 95.890 159.235 96.310 159.435 ;
        RECT 96.480 159.235 96.810 159.435 ;
        RECT 96.980 159.235 97.310 159.435 ;
        RECT 97.480 159.015 97.650 159.645 ;
        RECT 97.835 159.185 98.185 159.435 ;
        RECT 94.675 158.045 95.015 159.015 ;
        RECT 95.185 157.875 95.355 159.015 ;
        RECT 95.545 158.845 97.980 159.015 ;
        RECT 95.625 157.875 95.875 158.675 ;
        RECT 96.520 158.045 96.850 158.845 ;
        RECT 97.150 157.875 97.480 158.675 ;
        RECT 97.650 158.045 97.980 158.845 ;
        RECT 98.355 158.965 99.105 159.485 ;
        RECT 99.275 159.135 100.025 159.655 ;
        RECT 98.355 157.875 100.025 158.965 ;
        RECT 100.195 157.875 100.485 159.040 ;
        RECT 100.655 158.965 101.865 159.485 ;
        RECT 102.035 159.135 103.245 159.655 ;
        RECT 103.505 159.775 103.675 160.255 ;
        RECT 103.855 159.945 104.095 160.425 ;
        RECT 104.345 159.775 104.515 160.255 ;
        RECT 104.685 159.945 105.015 160.425 ;
        RECT 105.185 159.775 105.355 160.255 ;
        RECT 103.505 159.605 104.140 159.775 ;
        RECT 104.345 159.605 105.355 159.775 ;
        RECT 105.525 159.625 105.855 160.425 ;
        RECT 106.640 159.880 111.985 160.425 ;
        RECT 103.970 159.435 104.140 159.605 ;
        RECT 103.420 159.195 103.800 159.435 ;
        RECT 103.970 159.265 104.470 159.435 ;
        RECT 103.970 159.025 104.140 159.265 ;
        RECT 104.860 159.065 105.355 159.605 ;
        RECT 100.655 157.875 103.245 158.965 ;
        RECT 103.425 158.855 104.140 159.025 ;
        RECT 104.345 158.895 105.355 159.065 ;
        RECT 103.425 158.045 103.755 158.855 ;
        RECT 103.925 157.875 104.165 158.675 ;
        RECT 104.345 158.045 104.515 158.895 ;
        RECT 104.685 157.875 105.015 158.675 ;
        RECT 105.185 158.045 105.355 158.895 ;
        RECT 105.525 157.875 105.855 159.025 ;
        RECT 108.230 158.310 108.580 159.560 ;
        RECT 110.060 159.050 110.400 159.880 ;
        RECT 112.155 159.675 113.365 160.425 ;
        RECT 112.155 158.965 112.675 159.505 ;
        RECT 112.845 159.135 113.365 159.675 ;
        RECT 106.640 157.875 111.985 158.310 ;
        RECT 112.155 157.875 113.365 158.965 ;
        RECT 11.330 157.705 113.450 157.875 ;
        RECT 11.415 156.615 12.625 157.705 ;
        RECT 11.415 155.905 11.935 156.445 ;
        RECT 12.105 156.075 12.625 156.615 ;
        RECT 12.795 156.615 14.465 157.705 ;
        RECT 14.635 156.630 14.905 157.535 ;
        RECT 15.075 156.945 15.405 157.705 ;
        RECT 15.585 156.775 15.755 157.535 ;
        RECT 12.795 156.095 13.545 156.615 ;
        RECT 13.715 155.925 14.465 156.445 ;
        RECT 11.415 155.155 12.625 155.905 ;
        RECT 12.795 155.155 14.465 155.925 ;
        RECT 14.635 155.830 14.805 156.630 ;
        RECT 15.090 156.605 15.755 156.775 ;
        RECT 15.090 156.460 15.260 156.605 ;
        RECT 14.975 156.130 15.260 156.460 ;
        RECT 16.020 156.565 16.355 157.535 ;
        RECT 16.525 156.565 16.695 157.705 ;
        RECT 16.865 157.365 18.895 157.535 ;
        RECT 15.090 155.875 15.260 156.130 ;
        RECT 15.495 156.055 15.825 156.425 ;
        RECT 16.020 155.895 16.190 156.565 ;
        RECT 16.865 156.395 17.035 157.365 ;
        RECT 16.360 156.065 16.615 156.395 ;
        RECT 16.840 156.065 17.035 156.395 ;
        RECT 17.205 157.025 18.330 157.195 ;
        RECT 16.445 155.895 16.615 156.065 ;
        RECT 17.205 155.895 17.375 157.025 ;
        RECT 14.635 155.325 14.895 155.830 ;
        RECT 15.090 155.705 15.755 155.875 ;
        RECT 15.075 155.155 15.405 155.535 ;
        RECT 15.585 155.325 15.755 155.705 ;
        RECT 16.020 155.325 16.275 155.895 ;
        RECT 16.445 155.725 17.375 155.895 ;
        RECT 17.545 156.685 18.555 156.855 ;
        RECT 17.545 155.885 17.715 156.685 ;
        RECT 17.200 155.690 17.375 155.725 ;
        RECT 16.445 155.155 16.775 155.555 ;
        RECT 17.200 155.325 17.730 155.690 ;
        RECT 17.920 155.665 18.195 156.485 ;
        RECT 17.915 155.495 18.195 155.665 ;
        RECT 17.920 155.325 18.195 155.495 ;
        RECT 18.365 155.325 18.555 156.685 ;
        RECT 18.725 156.700 18.895 157.365 ;
        RECT 19.065 156.945 19.235 157.705 ;
        RECT 19.470 156.945 19.985 157.355 ;
        RECT 20.245 156.960 20.515 157.705 ;
        RECT 21.145 157.700 27.420 157.705 ;
        RECT 18.725 156.510 19.475 156.700 ;
        RECT 19.645 156.135 19.985 156.945 ;
        RECT 20.685 156.790 20.975 157.530 ;
        RECT 21.145 156.975 21.400 157.700 ;
        RECT 21.585 156.805 21.845 157.530 ;
        RECT 22.015 156.975 22.260 157.700 ;
        RECT 22.445 156.805 22.705 157.530 ;
        RECT 22.875 156.975 23.120 157.700 ;
        RECT 23.305 156.805 23.565 157.530 ;
        RECT 23.735 156.975 23.980 157.700 ;
        RECT 24.150 156.805 24.410 157.530 ;
        RECT 24.580 156.975 24.840 157.700 ;
        RECT 25.010 156.805 25.270 157.530 ;
        RECT 25.440 156.975 25.700 157.700 ;
        RECT 25.870 156.805 26.130 157.530 ;
        RECT 26.300 156.975 26.560 157.700 ;
        RECT 26.730 156.805 26.990 157.530 ;
        RECT 27.160 156.905 27.420 157.700 ;
        RECT 21.585 156.790 26.990 156.805 ;
        RECT 18.755 155.965 19.985 156.135 ;
        RECT 20.245 156.565 26.990 156.790 ;
        RECT 20.245 155.975 21.410 156.565 ;
        RECT 27.590 156.395 27.840 157.530 ;
        RECT 28.020 156.895 28.280 157.705 ;
        RECT 28.455 156.395 28.700 157.535 ;
        RECT 28.880 156.895 29.175 157.705 ;
        RECT 29.355 156.565 29.625 157.535 ;
        RECT 29.835 156.905 30.115 157.705 ;
        RECT 30.285 157.195 31.940 157.485 ;
        RECT 32.230 157.075 32.515 157.535 ;
        RECT 32.685 157.245 32.955 157.705 ;
        RECT 30.350 156.855 31.940 157.025 ;
        RECT 32.230 156.855 33.185 157.075 ;
        RECT 30.350 156.735 30.520 156.855 ;
        RECT 29.795 156.565 30.520 156.735 ;
        RECT 21.580 156.145 28.700 156.395 ;
        RECT 18.735 155.155 19.245 155.690 ;
        RECT 19.465 155.360 19.710 155.965 ;
        RECT 20.245 155.805 26.990 155.975 ;
        RECT 20.245 155.155 20.545 155.635 ;
        RECT 20.715 155.350 20.975 155.805 ;
        RECT 21.145 155.155 21.405 155.635 ;
        RECT 21.585 155.350 21.845 155.805 ;
        RECT 22.015 155.155 22.265 155.635 ;
        RECT 22.445 155.350 22.705 155.805 ;
        RECT 22.875 155.155 23.125 155.635 ;
        RECT 23.305 155.350 23.565 155.805 ;
        RECT 23.735 155.155 23.980 155.635 ;
        RECT 24.150 155.350 24.425 155.805 ;
        RECT 24.595 155.155 24.840 155.635 ;
        RECT 25.010 155.350 25.270 155.805 ;
        RECT 25.440 155.155 25.700 155.635 ;
        RECT 25.870 155.350 26.130 155.805 ;
        RECT 26.300 155.155 26.560 155.635 ;
        RECT 26.730 155.350 26.990 155.805 ;
        RECT 27.160 155.155 27.420 155.715 ;
        RECT 27.590 155.335 27.840 156.145 ;
        RECT 28.020 155.155 28.280 155.680 ;
        RECT 28.450 155.335 28.700 156.145 ;
        RECT 28.870 155.835 29.185 156.395 ;
        RECT 29.355 155.830 29.525 156.565 ;
        RECT 29.795 156.395 29.965 156.565 ;
        RECT 29.695 156.065 29.965 156.395 ;
        RECT 30.135 156.065 30.540 156.395 ;
        RECT 30.710 156.065 31.420 156.685 ;
        RECT 31.620 156.565 31.940 156.855 ;
        RECT 29.795 155.895 29.965 156.065 ;
        RECT 28.880 155.155 29.185 155.665 ;
        RECT 29.355 155.485 29.625 155.830 ;
        RECT 29.795 155.725 31.405 155.895 ;
        RECT 31.590 155.825 31.940 156.395 ;
        RECT 32.115 156.125 32.805 156.685 ;
        RECT 32.975 155.955 33.185 156.855 ;
        RECT 29.815 155.155 30.195 155.555 ;
        RECT 30.365 155.375 30.535 155.725 ;
        RECT 30.705 155.155 31.035 155.555 ;
        RECT 31.235 155.375 31.405 155.725 ;
        RECT 32.230 155.785 33.185 155.955 ;
        RECT 33.355 156.685 33.755 157.535 ;
        RECT 33.945 157.075 34.225 157.535 ;
        RECT 34.745 157.245 35.070 157.705 ;
        RECT 33.945 156.855 35.070 157.075 ;
        RECT 33.355 156.125 34.450 156.685 ;
        RECT 34.620 156.395 35.070 156.855 ;
        RECT 35.240 156.565 35.625 157.535 ;
        RECT 31.605 155.155 31.935 155.655 ;
        RECT 32.230 155.325 32.515 155.785 ;
        RECT 32.685 155.155 32.955 155.615 ;
        RECT 33.355 155.325 33.755 156.125 ;
        RECT 34.620 156.065 35.175 156.395 ;
        RECT 34.620 155.955 35.070 156.065 ;
        RECT 33.945 155.785 35.070 155.955 ;
        RECT 35.345 155.895 35.625 156.565 ;
        RECT 35.795 156.540 36.085 157.705 ;
        RECT 36.255 156.565 36.525 157.535 ;
        RECT 36.735 156.905 37.015 157.705 ;
        RECT 37.185 157.195 38.840 157.485 ;
        RECT 37.250 156.855 38.840 157.025 ;
        RECT 37.250 156.735 37.420 156.855 ;
        RECT 36.695 156.565 37.420 156.735 ;
        RECT 33.945 155.325 34.225 155.785 ;
        RECT 34.745 155.155 35.070 155.615 ;
        RECT 35.240 155.325 35.625 155.895 ;
        RECT 35.795 155.155 36.085 155.880 ;
        RECT 36.255 155.830 36.425 156.565 ;
        RECT 36.695 156.395 36.865 156.565 ;
        RECT 37.610 156.515 38.325 156.685 ;
        RECT 38.520 156.565 38.840 156.855 ;
        RECT 39.015 156.565 39.355 157.535 ;
        RECT 39.525 156.565 39.695 157.705 ;
        RECT 39.965 156.905 40.215 157.705 ;
        RECT 40.860 156.735 41.190 157.535 ;
        RECT 41.490 156.905 41.820 157.705 ;
        RECT 41.990 156.735 42.320 157.535 ;
        RECT 39.885 156.565 42.320 156.735 ;
        RECT 43.705 156.775 43.875 157.535 ;
        RECT 44.055 156.945 44.385 157.705 ;
        RECT 43.705 156.605 44.370 156.775 ;
        RECT 44.555 156.630 44.825 157.535 ;
        RECT 39.015 156.515 39.245 156.565 ;
        RECT 36.595 156.065 36.865 156.395 ;
        RECT 37.035 156.065 37.440 156.395 ;
        RECT 37.610 156.065 38.320 156.515 ;
        RECT 36.695 155.895 36.865 156.065 ;
        RECT 36.255 155.485 36.525 155.830 ;
        RECT 36.695 155.725 38.305 155.895 ;
        RECT 38.490 155.825 38.840 156.395 ;
        RECT 39.015 155.955 39.190 156.515 ;
        RECT 39.885 156.315 40.055 156.565 ;
        RECT 39.360 156.145 40.055 156.315 ;
        RECT 40.230 156.145 40.650 156.345 ;
        RECT 40.820 156.145 41.150 156.345 ;
        RECT 41.320 156.145 41.650 156.345 ;
        RECT 36.715 155.155 37.095 155.555 ;
        RECT 37.265 155.375 37.435 155.725 ;
        RECT 37.605 155.155 37.935 155.555 ;
        RECT 38.135 155.375 38.305 155.725 ;
        RECT 38.505 155.155 38.835 155.655 ;
        RECT 39.015 155.325 39.355 155.955 ;
        RECT 39.525 155.155 39.775 155.955 ;
        RECT 39.965 155.805 41.190 155.975 ;
        RECT 39.965 155.325 40.295 155.805 ;
        RECT 40.465 155.155 40.690 155.615 ;
        RECT 40.860 155.325 41.190 155.805 ;
        RECT 41.820 155.935 41.990 156.565 ;
        RECT 44.200 156.460 44.370 156.605 ;
        RECT 42.175 156.145 42.525 156.395 ;
        RECT 43.635 156.055 43.965 156.425 ;
        RECT 44.200 156.130 44.485 156.460 ;
        RECT 41.820 155.325 42.320 155.935 ;
        RECT 44.200 155.875 44.370 156.130 ;
        RECT 43.705 155.705 44.370 155.875 ;
        RECT 44.655 155.830 44.825 156.630 ;
        RECT 43.705 155.325 43.875 155.705 ;
        RECT 44.055 155.155 44.385 155.535 ;
        RECT 44.565 155.325 44.825 155.830 ;
        RECT 44.995 156.565 45.380 157.535 ;
        RECT 45.550 157.245 45.875 157.705 ;
        RECT 46.395 157.075 46.675 157.535 ;
        RECT 45.550 156.855 46.675 157.075 ;
        RECT 44.995 155.895 45.275 156.565 ;
        RECT 45.550 156.395 46.000 156.855 ;
        RECT 46.865 156.685 47.265 157.535 ;
        RECT 47.665 157.245 47.935 157.705 ;
        RECT 48.105 157.075 48.390 157.535 ;
        RECT 45.445 156.065 46.000 156.395 ;
        RECT 46.170 156.125 47.265 156.685 ;
        RECT 45.550 155.955 46.000 156.065 ;
        RECT 44.995 155.325 45.380 155.895 ;
        RECT 45.550 155.785 46.675 155.955 ;
        RECT 45.550 155.155 45.875 155.615 ;
        RECT 46.395 155.325 46.675 155.785 ;
        RECT 46.865 155.325 47.265 156.125 ;
        RECT 47.435 156.855 48.390 157.075 ;
        RECT 47.435 155.955 47.645 156.855 ;
        RECT 47.815 156.125 48.505 156.685 ;
        RECT 48.675 156.615 49.885 157.705 ;
        RECT 50.430 156.725 50.685 157.395 ;
        RECT 50.865 156.905 51.150 157.705 ;
        RECT 51.330 156.985 51.660 157.495 ;
        RECT 50.430 156.685 50.610 156.725 ;
        RECT 48.675 156.075 49.195 156.615 ;
        RECT 50.345 156.515 50.610 156.685 ;
        RECT 47.435 155.785 48.390 155.955 ;
        RECT 49.365 155.905 49.885 156.445 ;
        RECT 47.665 155.155 47.935 155.615 ;
        RECT 48.105 155.325 48.390 155.785 ;
        RECT 48.675 155.155 49.885 155.905 ;
        RECT 50.430 155.865 50.610 156.515 ;
        RECT 51.330 156.395 51.580 156.985 ;
        RECT 51.930 156.835 52.100 157.445 ;
        RECT 52.270 157.015 52.600 157.705 ;
        RECT 52.830 157.155 53.070 157.445 ;
        RECT 53.270 157.325 53.690 157.705 ;
        RECT 53.870 157.235 54.500 157.485 ;
        RECT 54.970 157.325 55.300 157.705 ;
        RECT 53.870 157.155 54.040 157.235 ;
        RECT 55.470 157.155 55.640 157.445 ;
        RECT 55.820 157.325 56.200 157.705 ;
        RECT 56.440 157.320 57.270 157.490 ;
        RECT 52.830 156.985 54.040 157.155 ;
        RECT 50.780 156.065 51.580 156.395 ;
        RECT 50.430 155.335 50.685 155.865 ;
        RECT 50.865 155.155 51.150 155.615 ;
        RECT 51.330 155.415 51.580 156.065 ;
        RECT 51.780 156.815 52.100 156.835 ;
        RECT 51.780 156.645 53.700 156.815 ;
        RECT 51.780 155.750 51.970 156.645 ;
        RECT 53.870 156.475 54.040 156.985 ;
        RECT 54.210 156.725 54.730 157.035 ;
        RECT 52.140 156.305 54.040 156.475 ;
        RECT 52.140 156.245 52.470 156.305 ;
        RECT 52.620 156.075 52.950 156.135 ;
        RECT 52.290 155.805 52.950 156.075 ;
        RECT 51.780 155.420 52.100 155.750 ;
        RECT 52.280 155.155 52.940 155.635 ;
        RECT 53.140 155.545 53.310 156.305 ;
        RECT 54.210 156.135 54.390 156.545 ;
        RECT 53.480 155.965 53.810 156.085 ;
        RECT 54.560 155.965 54.730 156.725 ;
        RECT 53.480 155.795 54.730 155.965 ;
        RECT 54.900 156.905 56.270 157.155 ;
        RECT 54.900 156.135 55.090 156.905 ;
        RECT 56.020 156.645 56.270 156.905 ;
        RECT 55.260 156.475 55.510 156.635 ;
        RECT 56.440 156.475 56.610 157.320 ;
        RECT 57.505 157.035 57.675 157.535 ;
        RECT 57.845 157.205 58.175 157.705 ;
        RECT 56.780 156.645 57.280 157.025 ;
        RECT 57.505 156.865 58.200 157.035 ;
        RECT 55.260 156.305 56.610 156.475 ;
        RECT 56.190 156.265 56.610 156.305 ;
        RECT 54.900 155.795 55.320 156.135 ;
        RECT 55.610 155.805 56.020 156.135 ;
        RECT 53.140 155.375 53.990 155.545 ;
        RECT 54.550 155.155 54.870 155.615 ;
        RECT 55.070 155.365 55.320 155.795 ;
        RECT 55.610 155.155 56.020 155.595 ;
        RECT 56.190 155.535 56.360 156.265 ;
        RECT 56.530 155.715 56.880 156.085 ;
        RECT 57.060 155.775 57.280 156.645 ;
        RECT 57.450 156.075 57.860 156.695 ;
        RECT 58.030 155.895 58.200 156.865 ;
        RECT 57.505 155.705 58.200 155.895 ;
        RECT 56.190 155.335 57.205 155.535 ;
        RECT 57.505 155.375 57.675 155.705 ;
        RECT 57.845 155.155 58.175 155.535 ;
        RECT 58.390 155.415 58.615 157.535 ;
        RECT 58.785 157.205 59.115 157.705 ;
        RECT 59.285 157.035 59.455 157.535 ;
        RECT 58.790 156.865 59.455 157.035 ;
        RECT 58.790 155.875 59.020 156.865 ;
        RECT 60.265 156.775 60.435 157.535 ;
        RECT 60.615 156.945 60.945 157.705 ;
        RECT 59.190 156.045 59.540 156.695 ;
        RECT 60.265 156.605 60.930 156.775 ;
        RECT 61.115 156.630 61.385 157.535 ;
        RECT 60.760 156.460 60.930 156.605 ;
        RECT 60.195 156.055 60.525 156.425 ;
        RECT 60.760 156.130 61.045 156.460 ;
        RECT 60.760 155.875 60.930 156.130 ;
        RECT 58.790 155.705 59.455 155.875 ;
        RECT 58.785 155.155 59.115 155.535 ;
        RECT 59.285 155.415 59.455 155.705 ;
        RECT 60.265 155.705 60.930 155.875 ;
        RECT 61.215 155.830 61.385 156.630 ;
        RECT 61.555 156.540 61.845 157.705 ;
        RECT 62.015 156.615 63.685 157.705 ;
        RECT 62.015 156.095 62.765 156.615 ;
        RECT 63.860 156.555 64.120 157.705 ;
        RECT 64.295 156.630 64.550 157.535 ;
        RECT 64.720 156.945 65.050 157.705 ;
        RECT 65.265 156.775 65.435 157.535 ;
        RECT 62.935 155.925 63.685 156.445 ;
        RECT 60.265 155.325 60.435 155.705 ;
        RECT 60.615 155.155 60.945 155.535 ;
        RECT 61.125 155.325 61.385 155.830 ;
        RECT 61.555 155.155 61.845 155.880 ;
        RECT 62.015 155.155 63.685 155.925 ;
        RECT 63.860 155.155 64.120 155.995 ;
        RECT 64.295 155.900 64.465 156.630 ;
        RECT 64.720 156.605 65.435 156.775 ;
        RECT 65.900 156.735 66.230 157.535 ;
        RECT 66.400 156.905 66.730 157.705 ;
        RECT 67.030 156.735 67.360 157.535 ;
        RECT 68.005 156.905 68.255 157.705 ;
        RECT 64.720 156.395 64.890 156.605 ;
        RECT 65.900 156.565 68.335 156.735 ;
        RECT 68.525 156.565 68.695 157.705 ;
        RECT 68.865 156.565 69.205 157.535 ;
        RECT 69.750 156.725 70.005 157.395 ;
        RECT 70.185 156.905 70.470 157.705 ;
        RECT 70.650 156.985 70.980 157.495 ;
        RECT 69.750 156.685 69.930 156.725 ;
        RECT 64.635 156.065 64.890 156.395 ;
        RECT 64.295 155.325 64.550 155.900 ;
        RECT 64.720 155.875 64.890 156.065 ;
        RECT 65.170 156.055 65.525 156.425 ;
        RECT 65.695 156.145 66.045 156.395 ;
        RECT 66.230 155.935 66.400 156.565 ;
        RECT 66.570 156.145 66.900 156.345 ;
        RECT 67.070 156.145 67.400 156.345 ;
        RECT 67.570 156.145 67.990 156.345 ;
        RECT 68.165 156.315 68.335 156.565 ;
        RECT 68.165 156.145 68.860 156.315 ;
        RECT 64.720 155.705 65.435 155.875 ;
        RECT 64.720 155.155 65.050 155.535 ;
        RECT 65.265 155.325 65.435 155.705 ;
        RECT 65.900 155.325 66.400 155.935 ;
        RECT 67.030 155.805 68.255 155.975 ;
        RECT 69.030 155.955 69.205 156.565 ;
        RECT 69.665 156.515 69.930 156.685 ;
        RECT 67.030 155.325 67.360 155.805 ;
        RECT 67.530 155.155 67.755 155.615 ;
        RECT 67.925 155.325 68.255 155.805 ;
        RECT 68.445 155.155 68.695 155.955 ;
        RECT 68.865 155.325 69.205 155.955 ;
        RECT 69.750 155.865 69.930 156.515 ;
        RECT 70.650 156.395 70.900 156.985 ;
        RECT 71.250 156.835 71.420 157.445 ;
        RECT 71.590 157.015 71.920 157.705 ;
        RECT 72.150 157.155 72.390 157.445 ;
        RECT 72.590 157.325 73.010 157.705 ;
        RECT 73.190 157.235 73.820 157.485 ;
        RECT 74.290 157.325 74.620 157.705 ;
        RECT 73.190 157.155 73.360 157.235 ;
        RECT 74.790 157.155 74.960 157.445 ;
        RECT 75.140 157.325 75.520 157.705 ;
        RECT 75.760 157.320 76.590 157.490 ;
        RECT 72.150 156.985 73.360 157.155 ;
        RECT 70.100 156.065 70.900 156.395 ;
        RECT 69.750 155.335 70.005 155.865 ;
        RECT 70.185 155.155 70.470 155.615 ;
        RECT 70.650 155.415 70.900 156.065 ;
        RECT 71.100 156.815 71.420 156.835 ;
        RECT 71.100 156.645 73.020 156.815 ;
        RECT 71.100 155.750 71.290 156.645 ;
        RECT 73.190 156.475 73.360 156.985 ;
        RECT 73.530 156.725 74.050 157.035 ;
        RECT 71.460 156.305 73.360 156.475 ;
        RECT 71.460 156.245 71.790 156.305 ;
        RECT 71.940 156.075 72.270 156.135 ;
        RECT 71.610 155.805 72.270 156.075 ;
        RECT 71.100 155.420 71.420 155.750 ;
        RECT 71.600 155.155 72.260 155.635 ;
        RECT 72.460 155.545 72.630 156.305 ;
        RECT 73.530 156.135 73.710 156.545 ;
        RECT 72.800 155.965 73.130 156.085 ;
        RECT 73.880 155.965 74.050 156.725 ;
        RECT 72.800 155.795 74.050 155.965 ;
        RECT 74.220 156.905 75.590 157.155 ;
        RECT 74.220 156.135 74.410 156.905 ;
        RECT 75.340 156.645 75.590 156.905 ;
        RECT 74.580 156.475 74.830 156.635 ;
        RECT 75.760 156.475 75.930 157.320 ;
        RECT 76.825 157.035 76.995 157.535 ;
        RECT 77.165 157.205 77.495 157.705 ;
        RECT 76.100 156.645 76.600 157.025 ;
        RECT 76.825 156.865 77.520 157.035 ;
        RECT 74.580 156.305 75.930 156.475 ;
        RECT 75.510 156.265 75.930 156.305 ;
        RECT 74.220 155.795 74.640 156.135 ;
        RECT 74.930 155.805 75.340 156.135 ;
        RECT 72.460 155.375 73.310 155.545 ;
        RECT 73.870 155.155 74.190 155.615 ;
        RECT 74.390 155.365 74.640 155.795 ;
        RECT 74.930 155.155 75.340 155.595 ;
        RECT 75.510 155.535 75.680 156.265 ;
        RECT 75.850 155.715 76.200 156.085 ;
        RECT 76.380 155.775 76.600 156.645 ;
        RECT 76.770 156.075 77.180 156.695 ;
        RECT 77.350 155.895 77.520 156.865 ;
        RECT 76.825 155.705 77.520 155.895 ;
        RECT 75.510 155.335 76.525 155.535 ;
        RECT 76.825 155.375 76.995 155.705 ;
        RECT 77.165 155.155 77.495 155.535 ;
        RECT 77.710 155.415 77.935 157.535 ;
        RECT 78.105 157.205 78.435 157.705 ;
        RECT 78.605 157.035 78.775 157.535 ;
        RECT 78.110 156.865 78.775 157.035 ;
        RECT 78.110 155.875 78.340 156.865 ;
        RECT 78.510 156.045 78.860 156.695 ;
        RECT 79.535 156.565 79.765 157.705 ;
        RECT 79.935 156.555 80.265 157.535 ;
        RECT 80.435 156.565 80.645 157.705 ;
        RECT 80.875 156.945 81.390 157.355 ;
        RECT 81.625 156.945 81.795 157.705 ;
        RECT 81.965 157.365 83.995 157.535 ;
        RECT 79.515 156.145 79.845 156.395 ;
        RECT 78.110 155.705 78.775 155.875 ;
        RECT 78.105 155.155 78.435 155.535 ;
        RECT 78.605 155.415 78.775 155.705 ;
        RECT 79.535 155.155 79.765 155.975 ;
        RECT 80.015 155.955 80.265 156.555 ;
        RECT 80.875 156.135 81.215 156.945 ;
        RECT 81.965 156.700 82.135 157.365 ;
        RECT 82.530 157.025 83.655 157.195 ;
        RECT 81.385 156.510 82.135 156.700 ;
        RECT 82.305 156.685 83.315 156.855 ;
        RECT 79.935 155.325 80.265 155.955 ;
        RECT 80.435 155.155 80.645 155.975 ;
        RECT 80.875 155.965 82.105 156.135 ;
        RECT 81.150 155.360 81.395 155.965 ;
        RECT 81.615 155.155 82.125 155.690 ;
        RECT 82.305 155.325 82.495 156.685 ;
        RECT 82.665 155.665 82.940 156.485 ;
        RECT 83.145 155.885 83.315 156.685 ;
        RECT 83.485 155.895 83.655 157.025 ;
        RECT 83.825 156.395 83.995 157.365 ;
        RECT 84.165 156.565 84.335 157.705 ;
        RECT 84.505 156.565 84.840 157.535 ;
        RECT 83.825 156.065 84.020 156.395 ;
        RECT 84.245 156.065 84.500 156.395 ;
        RECT 84.245 155.895 84.415 156.065 ;
        RECT 84.670 155.895 84.840 156.565 ;
        RECT 83.485 155.725 84.415 155.895 ;
        RECT 83.485 155.690 83.660 155.725 ;
        RECT 82.665 155.495 82.945 155.665 ;
        RECT 82.665 155.325 82.940 155.495 ;
        RECT 83.130 155.325 83.660 155.690 ;
        RECT 84.085 155.155 84.415 155.555 ;
        RECT 84.585 155.325 84.840 155.895 ;
        RECT 85.015 156.630 85.285 157.535 ;
        RECT 85.455 156.945 85.785 157.705 ;
        RECT 85.965 156.775 86.135 157.535 ;
        RECT 85.015 155.830 85.185 156.630 ;
        RECT 85.470 156.605 86.135 156.775 ;
        RECT 85.470 156.460 85.640 156.605 ;
        RECT 87.315 156.540 87.605 157.705 ;
        RECT 88.235 156.615 90.825 157.705 ;
        RECT 91.200 156.735 91.530 157.535 ;
        RECT 91.700 156.905 92.030 157.705 ;
        RECT 92.330 156.735 92.660 157.535 ;
        RECT 93.305 156.905 93.555 157.705 ;
        RECT 85.355 156.130 85.640 156.460 ;
        RECT 85.470 155.875 85.640 156.130 ;
        RECT 85.875 156.055 86.205 156.425 ;
        RECT 88.235 156.095 89.445 156.615 ;
        RECT 91.200 156.565 93.635 156.735 ;
        RECT 93.825 156.565 93.995 157.705 ;
        RECT 94.165 156.565 94.505 157.535 ;
        RECT 89.615 155.925 90.825 156.445 ;
        RECT 90.995 156.145 91.345 156.395 ;
        RECT 91.530 155.935 91.700 156.565 ;
        RECT 91.870 156.145 92.200 156.345 ;
        RECT 92.370 156.145 92.700 156.345 ;
        RECT 92.870 156.145 93.290 156.345 ;
        RECT 93.465 156.315 93.635 156.565 ;
        RECT 93.465 156.145 94.160 156.315 ;
        RECT 85.015 155.325 85.275 155.830 ;
        RECT 85.470 155.705 86.135 155.875 ;
        RECT 85.455 155.155 85.785 155.535 ;
        RECT 85.965 155.325 86.135 155.705 ;
        RECT 87.315 155.155 87.605 155.880 ;
        RECT 88.235 155.155 90.825 155.925 ;
        RECT 91.200 155.325 91.700 155.935 ;
        RECT 92.330 155.805 93.555 155.975 ;
        RECT 94.330 155.955 94.505 156.565 ;
        RECT 94.675 156.615 96.345 157.705 ;
        RECT 94.675 156.095 95.425 156.615 ;
        RECT 96.515 156.565 96.855 157.535 ;
        RECT 97.025 156.565 97.195 157.705 ;
        RECT 97.465 156.905 97.715 157.705 ;
        RECT 98.360 156.735 98.690 157.535 ;
        RECT 98.990 156.905 99.320 157.705 ;
        RECT 99.490 156.735 99.820 157.535 ;
        RECT 97.385 156.565 99.820 156.735 ;
        RECT 100.195 156.565 100.535 157.535 ;
        RECT 100.705 156.565 100.875 157.705 ;
        RECT 101.145 156.905 101.395 157.705 ;
        RECT 102.040 156.735 102.370 157.535 ;
        RECT 102.670 156.905 103.000 157.705 ;
        RECT 103.170 156.735 103.500 157.535 ;
        RECT 101.065 156.565 103.500 156.735 ;
        RECT 104.375 156.565 104.605 157.705 ;
        RECT 92.330 155.325 92.660 155.805 ;
        RECT 92.830 155.155 93.055 155.615 ;
        RECT 93.225 155.325 93.555 155.805 ;
        RECT 93.745 155.155 93.995 155.955 ;
        RECT 94.165 155.325 94.505 155.955 ;
        RECT 95.595 155.925 96.345 156.445 ;
        RECT 94.675 155.155 96.345 155.925 ;
        RECT 96.515 155.955 96.690 156.565 ;
        RECT 97.385 156.315 97.555 156.565 ;
        RECT 96.860 156.145 97.555 156.315 ;
        RECT 97.730 156.145 98.150 156.345 ;
        RECT 98.320 156.145 98.650 156.345 ;
        RECT 98.820 156.145 99.150 156.345 ;
        RECT 96.515 155.325 96.855 155.955 ;
        RECT 97.025 155.155 97.275 155.955 ;
        RECT 97.465 155.805 98.690 155.975 ;
        RECT 97.465 155.325 97.795 155.805 ;
        RECT 97.965 155.155 98.190 155.615 ;
        RECT 98.360 155.325 98.690 155.805 ;
        RECT 99.320 155.935 99.490 156.565 ;
        RECT 99.675 156.145 100.025 156.395 ;
        RECT 100.195 155.955 100.370 156.565 ;
        RECT 101.065 156.315 101.235 156.565 ;
        RECT 100.540 156.145 101.235 156.315 ;
        RECT 101.410 156.145 101.830 156.345 ;
        RECT 102.000 156.145 102.330 156.345 ;
        RECT 102.500 156.145 102.830 156.345 ;
        RECT 99.320 155.325 99.820 155.935 ;
        RECT 100.195 155.325 100.535 155.955 ;
        RECT 100.705 155.155 100.955 155.955 ;
        RECT 101.145 155.805 102.370 155.975 ;
        RECT 101.145 155.325 101.475 155.805 ;
        RECT 101.645 155.155 101.870 155.615 ;
        RECT 102.040 155.325 102.370 155.805 ;
        RECT 103.000 155.935 103.170 156.565 ;
        RECT 104.775 156.555 105.105 157.535 ;
        RECT 105.275 156.565 105.485 157.705 ;
        RECT 105.755 156.565 105.985 157.705 ;
        RECT 106.155 156.555 106.485 157.535 ;
        RECT 106.655 156.565 106.865 157.705 ;
        RECT 107.645 156.775 107.815 157.535 ;
        RECT 107.995 156.945 108.325 157.705 ;
        RECT 107.645 156.605 108.310 156.775 ;
        RECT 108.495 156.630 108.765 157.535 ;
        RECT 103.355 156.145 103.705 156.395 ;
        RECT 104.355 156.145 104.685 156.395 ;
        RECT 103.000 155.325 103.500 155.935 ;
        RECT 104.375 155.155 104.605 155.975 ;
        RECT 104.855 155.955 105.105 156.555 ;
        RECT 105.735 156.145 106.065 156.395 ;
        RECT 104.775 155.325 105.105 155.955 ;
        RECT 105.275 155.155 105.485 155.975 ;
        RECT 105.755 155.155 105.985 155.975 ;
        RECT 106.235 155.955 106.485 156.555 ;
        RECT 108.140 156.460 108.310 156.605 ;
        RECT 107.575 156.055 107.905 156.425 ;
        RECT 108.140 156.130 108.425 156.460 ;
        RECT 106.155 155.325 106.485 155.955 ;
        RECT 106.655 155.155 106.865 155.975 ;
        RECT 108.140 155.875 108.310 156.130 ;
        RECT 107.645 155.705 108.310 155.875 ;
        RECT 108.595 155.830 108.765 156.630 ;
        RECT 109.395 156.615 111.985 157.705 ;
        RECT 112.155 156.615 113.365 157.705 ;
        RECT 109.395 156.095 110.605 156.615 ;
        RECT 110.775 155.925 111.985 156.445 ;
        RECT 112.155 156.075 112.675 156.615 ;
        RECT 107.645 155.325 107.815 155.705 ;
        RECT 107.995 155.155 108.325 155.535 ;
        RECT 108.505 155.325 108.765 155.830 ;
        RECT 109.395 155.155 111.985 155.925 ;
        RECT 112.845 155.905 113.365 156.445 ;
        RECT 112.155 155.155 113.365 155.905 ;
        RECT 11.330 154.985 113.450 155.155 ;
        RECT 11.415 154.235 12.625 154.985 ;
        RECT 12.795 154.235 14.005 154.985 ;
        RECT 11.415 153.695 11.935 154.235 ;
        RECT 12.105 153.525 12.625 154.065 ;
        RECT 11.415 152.435 12.625 153.525 ;
        RECT 12.795 153.525 13.315 154.065 ;
        RECT 13.485 153.695 14.005 154.235 ;
        RECT 14.215 154.165 14.445 154.985 ;
        RECT 14.615 154.185 14.945 154.815 ;
        RECT 14.195 153.745 14.525 153.995 ;
        RECT 14.695 153.585 14.945 154.185 ;
        RECT 15.115 154.165 15.325 154.985 ;
        RECT 15.555 154.310 15.815 154.815 ;
        RECT 15.995 154.605 16.325 154.985 ;
        RECT 16.505 154.435 16.675 154.815 ;
        RECT 12.795 152.435 14.005 153.525 ;
        RECT 14.215 152.435 14.445 153.575 ;
        RECT 14.615 152.605 14.945 153.585 ;
        RECT 15.115 152.435 15.325 153.575 ;
        RECT 15.555 153.510 15.725 154.310 ;
        RECT 16.010 154.265 16.675 154.435 ;
        RECT 16.010 154.010 16.180 154.265 ;
        RECT 16.940 154.245 17.195 154.815 ;
        RECT 17.365 154.585 17.695 154.985 ;
        RECT 18.120 154.450 18.650 154.815 ;
        RECT 18.120 154.415 18.295 154.450 ;
        RECT 17.365 154.245 18.295 154.415 ;
        RECT 15.895 153.680 16.180 154.010 ;
        RECT 16.415 153.715 16.745 154.085 ;
        RECT 16.010 153.535 16.180 153.680 ;
        RECT 16.940 153.575 17.110 154.245 ;
        RECT 17.365 154.075 17.535 154.245 ;
        RECT 17.280 153.745 17.535 154.075 ;
        RECT 17.760 153.745 17.955 154.075 ;
        RECT 15.555 152.605 15.825 153.510 ;
        RECT 16.010 153.365 16.675 153.535 ;
        RECT 15.995 152.435 16.325 153.195 ;
        RECT 16.505 152.605 16.675 153.365 ;
        RECT 16.940 152.605 17.275 153.575 ;
        RECT 17.445 152.435 17.615 153.575 ;
        RECT 17.785 152.775 17.955 153.745 ;
        RECT 18.125 153.115 18.295 154.245 ;
        RECT 18.465 153.455 18.635 154.255 ;
        RECT 18.840 153.965 19.115 154.815 ;
        RECT 18.835 153.795 19.115 153.965 ;
        RECT 18.840 153.655 19.115 153.795 ;
        RECT 19.285 153.455 19.475 154.815 ;
        RECT 19.655 154.450 20.165 154.985 ;
        RECT 20.385 154.175 20.630 154.780 ;
        RECT 21.075 154.215 22.745 154.985 ;
        RECT 22.915 154.260 23.205 154.985 ;
        RECT 19.675 154.005 20.905 154.175 ;
        RECT 18.465 153.285 19.475 153.455 ;
        RECT 19.645 153.440 20.395 153.630 ;
        RECT 18.125 152.945 19.250 153.115 ;
        RECT 19.645 152.775 19.815 153.440 ;
        RECT 20.565 153.195 20.905 154.005 ;
        RECT 17.785 152.605 19.815 152.775 ;
        RECT 19.985 152.435 20.155 153.195 ;
        RECT 20.390 152.785 20.905 153.195 ;
        RECT 21.075 153.525 21.825 154.045 ;
        RECT 21.995 153.695 22.745 154.215 ;
        RECT 23.435 154.165 23.645 154.985 ;
        RECT 23.815 154.185 24.145 154.815 ;
        RECT 21.075 152.435 22.745 153.525 ;
        RECT 22.915 152.435 23.205 153.600 ;
        RECT 23.815 153.585 24.065 154.185 ;
        RECT 24.315 154.165 24.545 154.985 ;
        RECT 24.755 154.185 25.095 154.815 ;
        RECT 25.265 154.185 25.515 154.985 ;
        RECT 25.705 154.335 26.035 154.815 ;
        RECT 26.205 154.525 26.430 154.985 ;
        RECT 26.600 154.335 26.930 154.815 ;
        RECT 24.235 153.745 24.565 153.995 ;
        RECT 23.435 152.435 23.645 153.575 ;
        RECT 23.815 152.605 24.145 153.585 ;
        RECT 24.755 153.575 24.930 154.185 ;
        RECT 25.705 154.165 26.930 154.335 ;
        RECT 27.560 154.205 28.060 154.815 ;
        RECT 28.640 154.205 29.140 154.815 ;
        RECT 25.100 153.825 25.795 153.995 ;
        RECT 25.625 153.575 25.795 153.825 ;
        RECT 25.970 153.795 26.390 153.995 ;
        RECT 26.560 153.795 26.890 153.995 ;
        RECT 27.060 153.795 27.390 153.995 ;
        RECT 27.560 153.575 27.730 154.205 ;
        RECT 27.915 153.745 28.265 153.995 ;
        RECT 28.435 153.745 28.785 153.995 ;
        RECT 28.970 153.575 29.140 154.205 ;
        RECT 29.770 154.335 30.100 154.815 ;
        RECT 30.270 154.525 30.495 154.985 ;
        RECT 30.665 154.335 30.995 154.815 ;
        RECT 29.770 154.165 30.995 154.335 ;
        RECT 31.185 154.185 31.435 154.985 ;
        RECT 31.605 154.185 31.945 154.815 ;
        RECT 29.310 153.795 29.640 153.995 ;
        RECT 29.810 153.795 30.140 153.995 ;
        RECT 30.310 153.795 30.730 153.995 ;
        RECT 30.905 153.825 31.600 153.995 ;
        RECT 30.905 153.575 31.075 153.825 ;
        RECT 31.770 153.575 31.945 154.185 ;
        RECT 32.155 154.165 32.385 154.985 ;
        RECT 32.555 154.185 32.885 154.815 ;
        RECT 32.135 153.745 32.465 153.995 ;
        RECT 32.635 153.585 32.885 154.185 ;
        RECT 33.055 154.165 33.265 154.985 ;
        RECT 33.700 154.205 34.200 154.815 ;
        RECT 33.495 153.745 33.845 153.995 ;
        RECT 24.315 152.435 24.545 153.575 ;
        RECT 24.755 152.605 25.095 153.575 ;
        RECT 25.265 152.435 25.435 153.575 ;
        RECT 25.625 153.405 28.060 153.575 ;
        RECT 25.705 152.435 25.955 153.235 ;
        RECT 26.600 152.605 26.930 153.405 ;
        RECT 27.230 152.435 27.560 153.235 ;
        RECT 27.730 152.605 28.060 153.405 ;
        RECT 28.640 153.405 31.075 153.575 ;
        RECT 28.640 152.605 28.970 153.405 ;
        RECT 29.140 152.435 29.470 153.235 ;
        RECT 29.770 152.605 30.100 153.405 ;
        RECT 30.745 152.435 30.995 153.235 ;
        RECT 31.265 152.435 31.435 153.575 ;
        RECT 31.605 152.605 31.945 153.575 ;
        RECT 32.155 152.435 32.385 153.575 ;
        RECT 32.555 152.605 32.885 153.585 ;
        RECT 34.030 153.575 34.200 154.205 ;
        RECT 34.830 154.335 35.160 154.815 ;
        RECT 35.330 154.525 35.555 154.985 ;
        RECT 35.725 154.335 36.055 154.815 ;
        RECT 34.830 154.165 36.055 154.335 ;
        RECT 36.245 154.185 36.495 154.985 ;
        RECT 36.665 154.185 37.005 154.815 ;
        RECT 37.380 154.205 37.880 154.815 ;
        RECT 34.370 153.795 34.700 153.995 ;
        RECT 34.870 153.795 35.200 153.995 ;
        RECT 35.370 153.795 35.790 153.995 ;
        RECT 35.965 153.825 36.660 153.995 ;
        RECT 35.965 153.575 36.135 153.825 ;
        RECT 36.830 153.575 37.005 154.185 ;
        RECT 37.175 153.745 37.525 153.995 ;
        RECT 37.710 153.575 37.880 154.205 ;
        RECT 38.510 154.335 38.840 154.815 ;
        RECT 39.010 154.525 39.235 154.985 ;
        RECT 39.405 154.335 39.735 154.815 ;
        RECT 38.510 154.165 39.735 154.335 ;
        RECT 39.925 154.185 40.175 154.985 ;
        RECT 40.345 154.185 40.685 154.815 ;
        RECT 38.050 153.795 38.380 153.995 ;
        RECT 38.550 153.795 38.880 153.995 ;
        RECT 39.050 153.795 39.470 153.995 ;
        RECT 39.645 153.825 40.340 153.995 ;
        RECT 39.645 153.575 39.815 153.825 ;
        RECT 40.510 153.575 40.685 154.185 ;
        RECT 33.055 152.435 33.265 153.575 ;
        RECT 33.700 153.405 36.135 153.575 ;
        RECT 33.700 152.605 34.030 153.405 ;
        RECT 34.200 152.435 34.530 153.235 ;
        RECT 34.830 152.605 35.160 153.405 ;
        RECT 35.805 152.435 36.055 153.235 ;
        RECT 36.325 152.435 36.495 153.575 ;
        RECT 36.665 152.605 37.005 153.575 ;
        RECT 37.380 153.405 39.815 153.575 ;
        RECT 37.380 152.605 37.710 153.405 ;
        RECT 37.880 152.435 38.210 153.235 ;
        RECT 38.510 152.605 38.840 153.405 ;
        RECT 39.485 152.435 39.735 153.235 ;
        RECT 40.005 152.435 40.175 153.575 ;
        RECT 40.345 152.605 40.685 153.575 ;
        RECT 40.855 154.185 41.195 154.815 ;
        RECT 41.365 154.185 41.615 154.985 ;
        RECT 41.805 154.335 42.135 154.815 ;
        RECT 42.305 154.525 42.530 154.985 ;
        RECT 42.700 154.335 43.030 154.815 ;
        RECT 40.855 153.575 41.030 154.185 ;
        RECT 41.805 154.165 43.030 154.335 ;
        RECT 43.660 154.205 44.160 154.815 ;
        RECT 44.650 154.355 44.935 154.815 ;
        RECT 45.105 154.525 45.375 154.985 ;
        RECT 41.200 153.825 41.895 153.995 ;
        RECT 41.725 153.575 41.895 153.825 ;
        RECT 42.070 153.795 42.490 153.995 ;
        RECT 42.660 153.795 42.990 153.995 ;
        RECT 43.160 153.795 43.490 153.995 ;
        RECT 43.660 153.575 43.830 154.205 ;
        RECT 44.650 154.185 45.605 154.355 ;
        RECT 44.015 153.745 44.365 153.995 ;
        RECT 40.855 152.605 41.195 153.575 ;
        RECT 41.365 152.435 41.535 153.575 ;
        RECT 41.725 153.405 44.160 153.575 ;
        RECT 44.535 153.455 45.225 154.015 ;
        RECT 41.805 152.435 42.055 153.235 ;
        RECT 42.700 152.605 43.030 153.405 ;
        RECT 43.330 152.435 43.660 153.235 ;
        RECT 43.830 152.605 44.160 153.405 ;
        RECT 45.395 153.285 45.605 154.185 ;
        RECT 44.650 153.065 45.605 153.285 ;
        RECT 45.775 154.015 46.175 154.815 ;
        RECT 46.365 154.355 46.645 154.815 ;
        RECT 47.165 154.525 47.490 154.985 ;
        RECT 46.365 154.185 47.490 154.355 ;
        RECT 47.660 154.245 48.045 154.815 ;
        RECT 48.675 154.260 48.965 154.985 ;
        RECT 47.040 154.075 47.490 154.185 ;
        RECT 45.775 153.455 46.870 154.015 ;
        RECT 47.040 153.745 47.595 154.075 ;
        RECT 44.650 152.605 44.935 153.065 ;
        RECT 45.105 152.435 45.375 152.895 ;
        RECT 45.775 152.605 46.175 153.455 ;
        RECT 47.040 153.285 47.490 153.745 ;
        RECT 47.765 153.575 48.045 154.245 ;
        RECT 49.140 154.245 49.395 154.815 ;
        RECT 49.565 154.585 49.895 154.985 ;
        RECT 50.320 154.450 50.850 154.815 ;
        RECT 50.320 154.415 50.495 154.450 ;
        RECT 49.565 154.245 50.495 154.415 ;
        RECT 51.040 154.305 51.315 154.815 ;
        RECT 46.365 153.065 47.490 153.285 ;
        RECT 46.365 152.605 46.645 153.065 ;
        RECT 47.165 152.435 47.490 152.895 ;
        RECT 47.660 152.605 48.045 153.575 ;
        RECT 48.675 152.435 48.965 153.600 ;
        RECT 49.140 153.575 49.310 154.245 ;
        RECT 49.565 154.075 49.735 154.245 ;
        RECT 49.480 153.745 49.735 154.075 ;
        RECT 49.960 153.745 50.155 154.075 ;
        RECT 49.140 152.605 49.475 153.575 ;
        RECT 49.645 152.435 49.815 153.575 ;
        RECT 49.985 152.775 50.155 153.745 ;
        RECT 50.325 153.115 50.495 154.245 ;
        RECT 50.665 153.455 50.835 154.255 ;
        RECT 51.035 154.135 51.315 154.305 ;
        RECT 51.040 153.655 51.315 154.135 ;
        RECT 51.485 153.455 51.675 154.815 ;
        RECT 51.855 154.450 52.365 154.985 ;
        RECT 52.585 154.175 52.830 154.780 ;
        RECT 53.365 154.505 53.665 154.985 ;
        RECT 53.835 154.335 54.095 154.790 ;
        RECT 54.265 154.505 54.525 154.985 ;
        RECT 54.705 154.335 54.965 154.790 ;
        RECT 55.135 154.505 55.385 154.985 ;
        RECT 55.565 154.335 55.825 154.790 ;
        RECT 55.995 154.505 56.245 154.985 ;
        RECT 56.425 154.335 56.685 154.790 ;
        RECT 56.855 154.505 57.100 154.985 ;
        RECT 57.270 154.335 57.545 154.790 ;
        RECT 57.715 154.505 57.960 154.985 ;
        RECT 58.130 154.335 58.390 154.790 ;
        RECT 58.560 154.505 58.820 154.985 ;
        RECT 58.990 154.335 59.250 154.790 ;
        RECT 59.420 154.505 59.680 154.985 ;
        RECT 59.850 154.335 60.110 154.790 ;
        RECT 60.280 154.425 60.540 154.985 ;
        RECT 51.875 154.005 53.105 154.175 ;
        RECT 50.665 153.285 51.675 153.455 ;
        RECT 51.845 153.440 52.595 153.630 ;
        RECT 50.325 152.945 51.450 153.115 ;
        RECT 51.845 152.775 52.015 153.440 ;
        RECT 52.765 153.195 53.105 154.005 ;
        RECT 53.365 154.165 60.110 154.335 ;
        RECT 53.365 153.575 54.530 154.165 ;
        RECT 60.710 153.995 60.960 154.805 ;
        RECT 61.140 154.460 61.400 154.985 ;
        RECT 61.570 153.995 61.820 154.805 ;
        RECT 62.000 154.475 62.305 154.985 ;
        RECT 54.700 153.745 61.820 153.995 ;
        RECT 61.990 153.745 62.305 154.305 ;
        RECT 62.475 154.235 63.685 154.985 ;
        RECT 53.365 153.350 60.110 153.575 ;
        RECT 49.985 152.605 52.015 152.775 ;
        RECT 52.185 152.435 52.355 153.195 ;
        RECT 52.590 152.785 53.105 153.195 ;
        RECT 53.365 152.435 53.635 153.180 ;
        RECT 53.805 152.610 54.095 153.350 ;
        RECT 54.705 153.335 60.110 153.350 ;
        RECT 54.265 152.440 54.520 153.165 ;
        RECT 54.705 152.610 54.965 153.335 ;
        RECT 55.135 152.440 55.380 153.165 ;
        RECT 55.565 152.610 55.825 153.335 ;
        RECT 55.995 152.440 56.240 153.165 ;
        RECT 56.425 152.610 56.685 153.335 ;
        RECT 56.855 152.440 57.100 153.165 ;
        RECT 57.270 152.610 57.530 153.335 ;
        RECT 57.700 152.440 57.960 153.165 ;
        RECT 58.130 152.610 58.390 153.335 ;
        RECT 58.560 152.440 58.820 153.165 ;
        RECT 58.990 152.610 59.250 153.335 ;
        RECT 59.420 152.440 59.680 153.165 ;
        RECT 59.850 152.610 60.110 153.335 ;
        RECT 60.280 152.440 60.540 153.235 ;
        RECT 60.710 152.610 60.960 153.745 ;
        RECT 54.265 152.435 60.540 152.440 ;
        RECT 61.140 152.435 61.400 153.245 ;
        RECT 61.575 152.605 61.820 153.745 ;
        RECT 62.475 153.525 62.995 154.065 ;
        RECT 63.165 153.695 63.685 154.235 ;
        RECT 63.855 154.185 64.195 154.815 ;
        RECT 64.365 154.185 64.615 154.985 ;
        RECT 64.805 154.335 65.135 154.815 ;
        RECT 65.305 154.525 65.530 154.985 ;
        RECT 65.700 154.335 66.030 154.815 ;
        RECT 63.855 153.575 64.030 154.185 ;
        RECT 64.805 154.165 66.030 154.335 ;
        RECT 66.660 154.205 67.160 154.815 ;
        RECT 67.740 154.205 68.240 154.815 ;
        RECT 64.200 153.825 64.895 153.995 ;
        RECT 64.725 153.575 64.895 153.825 ;
        RECT 65.070 153.795 65.490 153.995 ;
        RECT 65.660 153.795 65.990 153.995 ;
        RECT 66.160 153.795 66.490 153.995 ;
        RECT 66.660 153.575 66.830 154.205 ;
        RECT 67.015 153.745 67.365 153.995 ;
        RECT 67.535 153.745 67.885 153.995 ;
        RECT 68.070 153.575 68.240 154.205 ;
        RECT 68.870 154.335 69.200 154.815 ;
        RECT 69.370 154.525 69.595 154.985 ;
        RECT 69.765 154.335 70.095 154.815 ;
        RECT 68.870 154.165 70.095 154.335 ;
        RECT 70.285 154.185 70.535 154.985 ;
        RECT 70.705 154.185 71.045 154.815 ;
        RECT 71.215 154.215 72.885 154.985 ;
        RECT 68.410 153.795 68.740 153.995 ;
        RECT 68.910 153.795 69.240 153.995 ;
        RECT 69.410 153.965 69.830 153.995 ;
        RECT 69.410 153.795 69.835 153.965 ;
        RECT 70.005 153.825 70.700 153.995 ;
        RECT 70.005 153.575 70.175 153.825 ;
        RECT 70.870 153.575 71.045 154.185 ;
        RECT 62.000 152.435 62.295 153.245 ;
        RECT 62.475 152.435 63.685 153.525 ;
        RECT 63.855 152.605 64.195 153.575 ;
        RECT 64.365 152.435 64.535 153.575 ;
        RECT 64.725 153.405 67.160 153.575 ;
        RECT 64.805 152.435 65.055 153.235 ;
        RECT 65.700 152.605 66.030 153.405 ;
        RECT 66.330 152.435 66.660 153.235 ;
        RECT 66.830 152.605 67.160 153.405 ;
        RECT 67.740 153.405 70.175 153.575 ;
        RECT 67.740 152.605 68.070 153.405 ;
        RECT 68.240 152.435 68.570 153.235 ;
        RECT 68.870 152.605 69.200 153.405 ;
        RECT 69.845 152.435 70.095 153.235 ;
        RECT 70.365 152.435 70.535 153.575 ;
        RECT 70.705 152.605 71.045 153.575 ;
        RECT 71.215 153.525 71.965 154.045 ;
        RECT 72.135 153.695 72.885 154.215 ;
        RECT 73.115 154.165 73.325 154.985 ;
        RECT 73.495 154.185 73.825 154.815 ;
        RECT 73.495 153.585 73.745 154.185 ;
        RECT 73.995 154.165 74.225 154.985 ;
        RECT 74.435 154.260 74.725 154.985 ;
        RECT 75.815 154.215 79.325 154.985 ;
        RECT 79.500 154.440 84.845 154.985 ;
        RECT 73.915 153.745 74.245 153.995 ;
        RECT 71.215 152.435 72.885 153.525 ;
        RECT 73.115 152.435 73.325 153.575 ;
        RECT 73.495 152.605 73.825 153.585 ;
        RECT 73.995 152.435 74.225 153.575 ;
        RECT 74.435 152.435 74.725 153.600 ;
        RECT 75.815 153.525 77.505 154.045 ;
        RECT 77.675 153.695 79.325 154.215 ;
        RECT 75.815 152.435 79.325 153.525 ;
        RECT 81.090 152.870 81.440 154.120 ;
        RECT 82.920 153.610 83.260 154.440 ;
        RECT 85.015 154.185 85.355 154.815 ;
        RECT 85.525 154.185 85.775 154.985 ;
        RECT 85.965 154.335 86.295 154.815 ;
        RECT 86.465 154.525 86.690 154.985 ;
        RECT 86.860 154.335 87.190 154.815 ;
        RECT 85.015 153.575 85.190 154.185 ;
        RECT 85.965 154.165 87.190 154.335 ;
        RECT 87.820 154.205 88.320 154.815 ;
        RECT 88.695 154.235 89.905 154.985 ;
        RECT 85.360 153.825 86.055 153.995 ;
        RECT 85.885 153.575 86.055 153.825 ;
        RECT 86.230 153.795 86.650 153.995 ;
        RECT 86.820 153.795 87.150 153.995 ;
        RECT 87.320 153.795 87.650 153.995 ;
        RECT 87.820 153.575 87.990 154.205 ;
        RECT 88.175 153.745 88.525 153.995 ;
        RECT 79.500 152.435 84.845 152.870 ;
        RECT 85.015 152.605 85.355 153.575 ;
        RECT 85.525 152.435 85.695 153.575 ;
        RECT 85.885 153.405 88.320 153.575 ;
        RECT 85.965 152.435 86.215 153.235 ;
        RECT 86.860 152.605 87.190 153.405 ;
        RECT 87.490 152.435 87.820 153.235 ;
        RECT 87.990 152.605 88.320 153.405 ;
        RECT 88.695 153.525 89.215 154.065 ;
        RECT 89.385 153.695 89.905 154.235 ;
        RECT 90.075 154.310 90.345 154.655 ;
        RECT 90.535 154.585 90.915 154.985 ;
        RECT 91.085 154.415 91.255 154.765 ;
        RECT 91.425 154.585 91.755 154.985 ;
        RECT 91.955 154.415 92.125 154.765 ;
        RECT 92.325 154.485 92.655 154.985 ;
        RECT 90.075 153.575 90.245 154.310 ;
        RECT 90.515 154.245 92.125 154.415 ;
        RECT 90.515 154.075 90.685 154.245 ;
        RECT 90.415 153.745 90.685 154.075 ;
        RECT 90.855 153.745 91.260 154.075 ;
        RECT 90.515 153.575 90.685 153.745 ;
        RECT 88.695 152.435 89.905 153.525 ;
        RECT 90.075 152.605 90.345 153.575 ;
        RECT 90.515 153.405 91.240 153.575 ;
        RECT 91.430 153.455 92.140 154.075 ;
        RECT 92.310 153.745 92.660 154.315 ;
        RECT 93.040 154.205 93.540 154.815 ;
        RECT 92.835 153.745 93.185 153.995 ;
        RECT 93.370 153.575 93.540 154.205 ;
        RECT 94.170 154.335 94.500 154.815 ;
        RECT 94.670 154.525 94.895 154.985 ;
        RECT 95.065 154.335 95.395 154.815 ;
        RECT 94.170 154.165 95.395 154.335 ;
        RECT 95.585 154.185 95.835 154.985 ;
        RECT 96.005 154.185 96.345 154.815 ;
        RECT 96.630 154.355 96.915 154.815 ;
        RECT 97.085 154.525 97.355 154.985 ;
        RECT 96.630 154.185 97.585 154.355 ;
        RECT 93.710 153.795 94.040 153.995 ;
        RECT 94.210 153.795 94.540 153.995 ;
        RECT 94.710 153.795 95.130 153.995 ;
        RECT 95.305 153.825 96.000 153.995 ;
        RECT 95.305 153.575 95.475 153.825 ;
        RECT 96.170 153.575 96.345 154.185 ;
        RECT 91.070 153.285 91.240 153.405 ;
        RECT 92.340 153.285 92.660 153.575 ;
        RECT 90.555 152.435 90.835 153.235 ;
        RECT 91.070 153.115 92.660 153.285 ;
        RECT 93.040 153.405 95.475 153.575 ;
        RECT 91.005 152.655 92.660 152.945 ;
        RECT 93.040 152.605 93.370 153.405 ;
        RECT 93.540 152.435 93.870 153.235 ;
        RECT 94.170 152.605 94.500 153.405 ;
        RECT 95.145 152.435 95.395 153.235 ;
        RECT 95.665 152.435 95.835 153.575 ;
        RECT 96.005 152.605 96.345 153.575 ;
        RECT 96.515 153.455 97.205 154.015 ;
        RECT 97.375 153.285 97.585 154.185 ;
        RECT 96.630 153.065 97.585 153.285 ;
        RECT 97.755 154.015 98.155 154.815 ;
        RECT 98.345 154.355 98.625 154.815 ;
        RECT 99.145 154.525 99.470 154.985 ;
        RECT 98.345 154.185 99.470 154.355 ;
        RECT 99.640 154.245 100.025 154.815 ;
        RECT 100.195 154.260 100.485 154.985 ;
        RECT 99.020 154.075 99.470 154.185 ;
        RECT 97.755 153.455 98.850 154.015 ;
        RECT 99.020 153.745 99.575 154.075 ;
        RECT 96.630 152.605 96.915 153.065 ;
        RECT 97.085 152.435 97.355 152.895 ;
        RECT 97.755 152.605 98.155 153.455 ;
        RECT 99.020 153.285 99.470 153.745 ;
        RECT 99.745 153.575 100.025 154.245 ;
        RECT 100.655 154.215 102.325 154.985 ;
        RECT 98.345 153.065 99.470 153.285 ;
        RECT 98.345 152.605 98.625 153.065 ;
        RECT 99.145 152.435 99.470 152.895 ;
        RECT 99.640 152.605 100.025 153.575 ;
        RECT 100.195 152.435 100.485 153.600 ;
        RECT 100.655 153.525 101.405 154.045 ;
        RECT 101.575 153.695 102.325 154.215 ;
        RECT 102.500 154.275 102.755 154.805 ;
        RECT 102.925 154.525 103.230 154.985 ;
        RECT 103.475 154.605 104.545 154.775 ;
        RECT 102.500 153.625 102.710 154.275 ;
        RECT 103.475 154.250 103.795 154.605 ;
        RECT 103.470 154.075 103.795 154.250 ;
        RECT 102.880 153.775 103.795 154.075 ;
        RECT 103.965 154.035 104.205 154.435 ;
        RECT 104.375 154.375 104.545 154.605 ;
        RECT 104.715 154.545 104.905 154.985 ;
        RECT 105.075 154.535 106.025 154.815 ;
        RECT 106.245 154.625 106.595 154.795 ;
        RECT 104.375 154.205 104.905 154.375 ;
        RECT 102.880 153.745 103.620 153.775 ;
        RECT 100.655 152.435 102.325 153.525 ;
        RECT 102.500 152.745 102.755 153.625 ;
        RECT 102.925 152.435 103.230 153.575 ;
        RECT 103.450 153.155 103.620 153.745 ;
        RECT 103.965 153.665 104.505 154.035 ;
        RECT 104.685 153.925 104.905 154.205 ;
        RECT 105.075 153.755 105.245 154.535 ;
        RECT 104.840 153.585 105.245 153.755 ;
        RECT 105.415 153.745 105.765 154.365 ;
        RECT 104.840 153.495 105.010 153.585 ;
        RECT 105.935 153.575 106.145 154.365 ;
        RECT 103.790 153.325 105.010 153.495 ;
        RECT 105.470 153.415 106.145 153.575 ;
        RECT 103.450 152.985 104.250 153.155 ;
        RECT 103.570 152.435 103.900 152.815 ;
        RECT 104.080 152.695 104.250 152.985 ;
        RECT 104.840 152.945 105.010 153.325 ;
        RECT 105.180 153.405 106.145 153.415 ;
        RECT 106.335 154.235 106.595 154.625 ;
        RECT 106.805 154.525 107.135 154.985 ;
        RECT 108.010 154.595 108.865 154.765 ;
        RECT 109.070 154.595 109.565 154.765 ;
        RECT 109.735 154.625 110.065 154.985 ;
        RECT 106.335 153.545 106.505 154.235 ;
        RECT 106.675 153.885 106.845 154.065 ;
        RECT 107.015 154.055 107.805 154.305 ;
        RECT 108.010 153.885 108.180 154.595 ;
        RECT 108.350 154.085 108.705 154.305 ;
        RECT 106.675 153.715 108.365 153.885 ;
        RECT 105.180 153.115 105.640 153.405 ;
        RECT 106.335 153.375 107.835 153.545 ;
        RECT 106.335 153.235 106.505 153.375 ;
        RECT 105.945 153.065 106.505 153.235 ;
        RECT 104.420 152.435 104.670 152.895 ;
        RECT 104.840 152.605 105.710 152.945 ;
        RECT 105.945 152.605 106.115 153.065 ;
        RECT 106.950 153.035 108.025 153.205 ;
        RECT 106.285 152.435 106.655 152.895 ;
        RECT 106.950 152.695 107.120 153.035 ;
        RECT 107.290 152.435 107.620 152.865 ;
        RECT 107.855 152.695 108.025 153.035 ;
        RECT 108.195 152.935 108.365 153.715 ;
        RECT 108.535 153.495 108.705 154.085 ;
        RECT 108.875 153.685 109.225 154.305 ;
        RECT 108.535 153.105 109.000 153.495 ;
        RECT 109.395 153.235 109.565 154.595 ;
        RECT 109.735 153.405 110.195 154.455 ;
        RECT 109.170 153.065 109.565 153.235 ;
        RECT 109.170 152.935 109.340 153.065 ;
        RECT 108.195 152.605 108.875 152.935 ;
        RECT 109.090 152.605 109.340 152.935 ;
        RECT 109.510 152.435 109.760 152.895 ;
        RECT 109.930 152.620 110.255 153.405 ;
        RECT 110.425 152.605 110.595 154.725 ;
        RECT 110.765 154.605 111.095 154.985 ;
        RECT 111.265 154.435 111.520 154.725 ;
        RECT 110.770 154.265 111.520 154.435 ;
        RECT 110.770 153.275 111.000 154.265 ;
        RECT 112.155 154.235 113.365 154.985 ;
        RECT 111.170 153.445 111.520 154.095 ;
        RECT 112.155 153.525 112.675 154.065 ;
        RECT 112.845 153.695 113.365 154.235 ;
        RECT 110.770 153.105 111.520 153.275 ;
        RECT 110.765 152.435 111.095 152.935 ;
        RECT 111.265 152.605 111.520 153.105 ;
        RECT 112.155 152.435 113.365 153.525 ;
        RECT 11.330 152.265 113.450 152.435 ;
        RECT 11.415 151.175 12.625 152.265 ;
        RECT 12.885 151.595 13.055 152.095 ;
        RECT 13.225 151.765 13.555 152.265 ;
        RECT 12.885 151.425 13.550 151.595 ;
        RECT 11.415 150.465 11.935 151.005 ;
        RECT 12.105 150.635 12.625 151.175 ;
        RECT 12.800 150.605 13.150 151.255 ;
        RECT 11.415 149.715 12.625 150.465 ;
        RECT 13.320 150.435 13.550 151.425 ;
        RECT 12.885 150.265 13.550 150.435 ;
        RECT 12.885 149.975 13.055 150.265 ;
        RECT 13.225 149.715 13.555 150.095 ;
        RECT 13.725 149.975 13.950 152.095 ;
        RECT 14.165 151.765 14.495 152.265 ;
        RECT 14.665 151.595 14.835 152.095 ;
        RECT 15.070 151.880 15.900 152.050 ;
        RECT 16.140 151.885 16.520 152.265 ;
        RECT 14.140 151.425 14.835 151.595 ;
        RECT 14.140 150.455 14.310 151.425 ;
        RECT 14.480 150.635 14.890 151.255 ;
        RECT 15.060 151.205 15.560 151.585 ;
        RECT 14.140 150.265 14.835 150.455 ;
        RECT 15.060 150.335 15.280 151.205 ;
        RECT 15.730 151.035 15.900 151.880 ;
        RECT 16.700 151.715 16.870 152.005 ;
        RECT 17.040 151.885 17.370 152.265 ;
        RECT 17.840 151.795 18.470 152.045 ;
        RECT 18.650 151.885 19.070 152.265 ;
        RECT 18.300 151.715 18.470 151.795 ;
        RECT 19.270 151.715 19.510 152.005 ;
        RECT 16.070 151.465 17.440 151.715 ;
        RECT 16.070 151.205 16.320 151.465 ;
        RECT 16.830 151.035 17.080 151.195 ;
        RECT 15.730 150.865 17.080 151.035 ;
        RECT 15.730 150.825 16.150 150.865 ;
        RECT 15.460 150.275 15.810 150.645 ;
        RECT 14.165 149.715 14.495 150.095 ;
        RECT 14.665 149.935 14.835 150.265 ;
        RECT 15.980 150.095 16.150 150.825 ;
        RECT 17.250 150.695 17.440 151.465 ;
        RECT 16.320 150.365 16.730 150.695 ;
        RECT 17.020 150.355 17.440 150.695 ;
        RECT 17.610 151.285 18.130 151.595 ;
        RECT 18.300 151.545 19.510 151.715 ;
        RECT 19.740 151.575 20.070 152.265 ;
        RECT 17.610 150.525 17.780 151.285 ;
        RECT 17.950 150.695 18.130 151.105 ;
        RECT 18.300 151.035 18.470 151.545 ;
        RECT 20.240 151.395 20.410 152.005 ;
        RECT 20.680 151.545 21.010 152.055 ;
        RECT 20.240 151.375 20.560 151.395 ;
        RECT 18.640 151.205 20.560 151.375 ;
        RECT 18.300 150.865 20.200 151.035 ;
        RECT 18.530 150.525 18.860 150.645 ;
        RECT 17.610 150.355 18.860 150.525 ;
        RECT 15.135 149.895 16.150 150.095 ;
        RECT 16.320 149.715 16.730 150.155 ;
        RECT 17.020 149.925 17.270 150.355 ;
        RECT 17.470 149.715 17.790 150.175 ;
        RECT 19.030 150.105 19.200 150.865 ;
        RECT 19.870 150.805 20.200 150.865 ;
        RECT 19.390 150.635 19.720 150.695 ;
        RECT 19.390 150.365 20.050 150.635 ;
        RECT 20.370 150.310 20.560 151.205 ;
        RECT 18.350 149.935 19.200 150.105 ;
        RECT 19.400 149.715 20.060 150.195 ;
        RECT 20.240 149.980 20.560 150.310 ;
        RECT 20.760 150.955 21.010 151.545 ;
        RECT 21.190 151.465 21.475 152.265 ;
        RECT 21.655 151.925 21.910 151.955 ;
        RECT 21.655 151.755 21.995 151.925 ;
        RECT 21.655 151.285 21.910 151.755 ;
        RECT 20.760 150.625 21.560 150.955 ;
        RECT 20.760 149.975 21.010 150.625 ;
        RECT 21.730 150.425 21.910 151.285 ;
        RECT 21.190 149.715 21.475 150.175 ;
        RECT 21.655 149.895 21.910 150.425 ;
        RECT 22.920 151.075 23.175 151.955 ;
        RECT 23.345 151.125 23.650 152.265 ;
        RECT 23.990 151.885 24.320 152.265 ;
        RECT 24.500 151.715 24.670 152.005 ;
        RECT 24.840 151.805 25.090 152.265 ;
        RECT 23.870 151.545 24.670 151.715 ;
        RECT 25.260 151.755 26.130 152.095 ;
        RECT 22.920 150.425 23.130 151.075 ;
        RECT 23.870 150.955 24.040 151.545 ;
        RECT 25.260 151.375 25.430 151.755 ;
        RECT 26.365 151.635 26.535 152.095 ;
        RECT 26.705 151.805 27.075 152.265 ;
        RECT 27.370 151.665 27.540 152.005 ;
        RECT 27.710 151.835 28.040 152.265 ;
        RECT 28.275 151.665 28.445 152.005 ;
        RECT 24.210 151.205 25.430 151.375 ;
        RECT 25.600 151.295 26.060 151.585 ;
        RECT 26.365 151.465 26.925 151.635 ;
        RECT 27.370 151.495 28.445 151.665 ;
        RECT 28.615 151.765 29.295 152.095 ;
        RECT 29.510 151.765 29.760 152.095 ;
        RECT 29.930 151.805 30.180 152.265 ;
        RECT 26.755 151.325 26.925 151.465 ;
        RECT 25.600 151.285 26.565 151.295 ;
        RECT 25.260 151.115 25.430 151.205 ;
        RECT 25.890 151.125 26.565 151.285 ;
        RECT 23.300 150.925 24.040 150.955 ;
        RECT 23.300 150.625 24.215 150.925 ;
        RECT 23.890 150.450 24.215 150.625 ;
        RECT 22.920 149.895 23.175 150.425 ;
        RECT 23.345 149.715 23.650 150.175 ;
        RECT 23.895 150.095 24.215 150.450 ;
        RECT 24.385 150.665 24.925 151.035 ;
        RECT 25.260 150.945 25.665 151.115 ;
        RECT 24.385 150.265 24.625 150.665 ;
        RECT 25.105 150.495 25.325 150.775 ;
        RECT 24.795 150.325 25.325 150.495 ;
        RECT 24.795 150.095 24.965 150.325 ;
        RECT 25.495 150.165 25.665 150.945 ;
        RECT 25.835 150.335 26.185 150.955 ;
        RECT 26.355 150.335 26.565 151.125 ;
        RECT 26.755 151.155 28.255 151.325 ;
        RECT 26.755 150.465 26.925 151.155 ;
        RECT 28.615 150.985 28.785 151.765 ;
        RECT 29.590 151.635 29.760 151.765 ;
        RECT 27.095 150.815 28.785 150.985 ;
        RECT 28.955 151.205 29.420 151.595 ;
        RECT 29.590 151.465 29.985 151.635 ;
        RECT 27.095 150.635 27.265 150.815 ;
        RECT 23.895 149.925 24.965 150.095 ;
        RECT 25.135 149.715 25.325 150.155 ;
        RECT 25.495 149.885 26.445 150.165 ;
        RECT 26.755 150.075 27.015 150.465 ;
        RECT 27.435 150.395 28.225 150.645 ;
        RECT 26.665 149.905 27.015 150.075 ;
        RECT 27.225 149.715 27.555 150.175 ;
        RECT 28.430 150.105 28.600 150.815 ;
        RECT 28.955 150.615 29.125 151.205 ;
        RECT 28.770 150.395 29.125 150.615 ;
        RECT 29.295 150.395 29.645 151.015 ;
        RECT 29.815 150.105 29.985 151.465 ;
        RECT 30.350 151.295 30.675 152.080 ;
        RECT 30.155 150.245 30.615 151.295 ;
        RECT 28.430 149.935 29.285 150.105 ;
        RECT 29.490 149.935 29.985 150.105 ;
        RECT 30.155 149.715 30.485 150.075 ;
        RECT 30.845 149.975 31.015 152.095 ;
        RECT 31.185 151.765 31.515 152.265 ;
        RECT 31.685 151.595 31.940 152.095 ;
        RECT 31.190 151.425 31.940 151.595 ;
        RECT 31.190 150.435 31.420 151.425 ;
        RECT 32.320 151.295 32.650 152.095 ;
        RECT 32.820 151.465 33.150 152.265 ;
        RECT 33.450 151.295 33.780 152.095 ;
        RECT 34.425 151.465 34.675 152.265 ;
        RECT 31.590 150.605 31.940 151.255 ;
        RECT 32.320 151.125 34.755 151.295 ;
        RECT 34.945 151.125 35.115 152.265 ;
        RECT 35.285 151.125 35.625 152.095 ;
        RECT 32.115 150.705 32.465 150.955 ;
        RECT 32.650 150.495 32.820 151.125 ;
        RECT 32.990 150.705 33.320 150.905 ;
        RECT 33.490 150.705 33.820 150.905 ;
        RECT 33.990 150.705 34.410 150.905 ;
        RECT 34.585 150.875 34.755 151.125 ;
        RECT 34.585 150.705 35.280 150.875 ;
        RECT 31.190 150.265 31.940 150.435 ;
        RECT 31.185 149.715 31.515 150.095 ;
        RECT 31.685 149.975 31.940 150.265 ;
        RECT 32.320 149.885 32.820 150.495 ;
        RECT 33.450 150.365 34.675 150.535 ;
        RECT 35.450 150.515 35.625 151.125 ;
        RECT 35.795 151.100 36.085 152.265 ;
        RECT 36.315 151.125 36.525 152.265 ;
        RECT 36.695 151.115 37.025 152.095 ;
        RECT 37.195 151.125 37.425 152.265 ;
        RECT 37.640 151.125 37.975 152.095 ;
        RECT 38.145 151.125 38.315 152.265 ;
        RECT 38.485 151.925 40.515 152.095 ;
        RECT 33.450 149.885 33.780 150.365 ;
        RECT 33.950 149.715 34.175 150.175 ;
        RECT 34.345 149.885 34.675 150.365 ;
        RECT 34.865 149.715 35.115 150.515 ;
        RECT 35.285 149.885 35.625 150.515 ;
        RECT 35.795 149.715 36.085 150.440 ;
        RECT 36.315 149.715 36.525 150.535 ;
        RECT 36.695 150.515 36.945 151.115 ;
        RECT 37.115 150.705 37.445 150.955 ;
        RECT 36.695 149.885 37.025 150.515 ;
        RECT 37.195 149.715 37.425 150.535 ;
        RECT 37.640 150.455 37.810 151.125 ;
        RECT 38.485 150.955 38.655 151.925 ;
        RECT 37.980 150.625 38.235 150.955 ;
        RECT 38.460 150.625 38.655 150.955 ;
        RECT 38.825 151.585 39.950 151.755 ;
        RECT 38.065 150.455 38.235 150.625 ;
        RECT 38.825 150.455 38.995 151.585 ;
        RECT 37.640 149.885 37.895 150.455 ;
        RECT 38.065 150.285 38.995 150.455 ;
        RECT 39.165 151.245 40.175 151.415 ;
        RECT 39.165 150.445 39.335 151.245 ;
        RECT 39.540 150.565 39.815 151.045 ;
        RECT 39.535 150.395 39.815 150.565 ;
        RECT 38.820 150.250 38.995 150.285 ;
        RECT 38.065 149.715 38.395 150.115 ;
        RECT 38.820 149.885 39.350 150.250 ;
        RECT 39.540 149.885 39.815 150.395 ;
        RECT 39.985 149.885 40.175 151.245 ;
        RECT 40.345 151.260 40.515 151.925 ;
        RECT 40.685 151.505 40.855 152.265 ;
        RECT 41.090 151.505 41.605 151.915 ;
        RECT 40.345 151.070 41.095 151.260 ;
        RECT 41.265 150.695 41.605 151.505 ;
        RECT 40.375 150.525 41.605 150.695 ;
        RECT 42.235 151.175 44.825 152.265 ;
        RECT 42.235 150.655 43.445 151.175 ;
        RECT 45.000 151.075 45.255 151.955 ;
        RECT 45.425 151.125 45.730 152.265 ;
        RECT 46.070 151.885 46.400 152.265 ;
        RECT 46.580 151.715 46.750 152.005 ;
        RECT 46.920 151.805 47.170 152.265 ;
        RECT 45.950 151.545 46.750 151.715 ;
        RECT 47.340 151.755 48.210 152.095 ;
        RECT 40.355 149.715 40.865 150.250 ;
        RECT 41.085 149.920 41.330 150.525 ;
        RECT 43.615 150.485 44.825 151.005 ;
        RECT 42.235 149.715 44.825 150.485 ;
        RECT 45.000 150.425 45.210 151.075 ;
        RECT 45.950 150.955 46.120 151.545 ;
        RECT 47.340 151.375 47.510 151.755 ;
        RECT 48.445 151.635 48.615 152.095 ;
        RECT 48.785 151.805 49.155 152.265 ;
        RECT 49.450 151.665 49.620 152.005 ;
        RECT 49.790 151.835 50.120 152.265 ;
        RECT 50.355 151.665 50.525 152.005 ;
        RECT 46.290 151.205 47.510 151.375 ;
        RECT 47.680 151.295 48.140 151.585 ;
        RECT 48.445 151.465 49.005 151.635 ;
        RECT 49.450 151.495 50.525 151.665 ;
        RECT 50.695 151.765 51.375 152.095 ;
        RECT 51.590 151.765 51.840 152.095 ;
        RECT 52.010 151.805 52.260 152.265 ;
        RECT 48.835 151.325 49.005 151.465 ;
        RECT 47.680 151.285 48.645 151.295 ;
        RECT 47.340 151.115 47.510 151.205 ;
        RECT 47.970 151.125 48.645 151.285 ;
        RECT 45.380 150.925 46.120 150.955 ;
        RECT 45.380 150.625 46.295 150.925 ;
        RECT 45.970 150.450 46.295 150.625 ;
        RECT 45.000 149.895 45.255 150.425 ;
        RECT 45.425 149.715 45.730 150.175 ;
        RECT 45.975 150.095 46.295 150.450 ;
        RECT 46.465 150.665 47.005 151.035 ;
        RECT 47.340 150.945 47.745 151.115 ;
        RECT 46.465 150.265 46.705 150.665 ;
        RECT 47.185 150.495 47.405 150.775 ;
        RECT 46.875 150.325 47.405 150.495 ;
        RECT 46.875 150.095 47.045 150.325 ;
        RECT 47.575 150.165 47.745 150.945 ;
        RECT 47.915 150.335 48.265 150.955 ;
        RECT 48.435 150.335 48.645 151.125 ;
        RECT 48.835 151.155 50.335 151.325 ;
        RECT 48.835 150.465 49.005 151.155 ;
        RECT 50.695 150.985 50.865 151.765 ;
        RECT 51.670 151.635 51.840 151.765 ;
        RECT 49.175 150.815 50.865 150.985 ;
        RECT 51.035 151.205 51.500 151.595 ;
        RECT 51.670 151.465 52.065 151.635 ;
        RECT 49.175 150.635 49.345 150.815 ;
        RECT 45.975 149.925 47.045 150.095 ;
        RECT 47.215 149.715 47.405 150.155 ;
        RECT 47.575 149.885 48.525 150.165 ;
        RECT 48.835 150.075 49.095 150.465 ;
        RECT 49.515 150.395 50.305 150.645 ;
        RECT 48.745 149.905 49.095 150.075 ;
        RECT 49.305 149.715 49.635 150.175 ;
        RECT 50.510 150.105 50.680 150.815 ;
        RECT 51.035 150.615 51.205 151.205 ;
        RECT 50.850 150.395 51.205 150.615 ;
        RECT 51.375 150.395 51.725 151.015 ;
        RECT 51.895 150.105 52.065 151.465 ;
        RECT 52.430 151.295 52.755 152.080 ;
        RECT 52.235 150.245 52.695 151.295 ;
        RECT 50.510 149.935 51.365 150.105 ;
        RECT 51.570 149.935 52.065 150.105 ;
        RECT 52.235 149.715 52.565 150.075 ;
        RECT 52.925 149.975 53.095 152.095 ;
        RECT 53.265 151.765 53.595 152.265 ;
        RECT 53.765 151.595 54.020 152.095 ;
        RECT 53.270 151.425 54.020 151.595 ;
        RECT 53.270 150.435 53.500 151.425 ;
        RECT 53.670 150.605 54.020 151.255 ;
        RECT 54.195 151.175 55.865 152.265 ;
        RECT 56.035 151.505 56.550 151.915 ;
        RECT 56.785 151.505 56.955 152.265 ;
        RECT 57.125 151.925 59.155 152.095 ;
        RECT 54.195 150.655 54.945 151.175 ;
        RECT 55.115 150.485 55.865 151.005 ;
        RECT 56.035 150.695 56.375 151.505 ;
        RECT 57.125 151.260 57.295 151.925 ;
        RECT 57.690 151.585 58.815 151.755 ;
        RECT 56.545 151.070 57.295 151.260 ;
        RECT 57.465 151.245 58.475 151.415 ;
        RECT 56.035 150.525 57.265 150.695 ;
        RECT 53.270 150.265 54.020 150.435 ;
        RECT 53.265 149.715 53.595 150.095 ;
        RECT 53.765 149.975 54.020 150.265 ;
        RECT 54.195 149.715 55.865 150.485 ;
        RECT 56.310 149.920 56.555 150.525 ;
        RECT 56.775 149.715 57.285 150.250 ;
        RECT 57.465 149.885 57.655 151.245 ;
        RECT 57.825 150.225 58.100 151.045 ;
        RECT 58.305 150.445 58.475 151.245 ;
        RECT 58.645 150.455 58.815 151.585 ;
        RECT 58.985 150.955 59.155 151.925 ;
        RECT 59.325 151.125 59.495 152.265 ;
        RECT 59.665 151.125 60.000 152.095 ;
        RECT 58.985 150.625 59.180 150.955 ;
        RECT 59.405 150.625 59.660 150.955 ;
        RECT 59.405 150.455 59.575 150.625 ;
        RECT 59.830 150.455 60.000 151.125 ;
        RECT 60.175 151.175 61.385 152.265 ;
        RECT 60.175 150.635 60.695 151.175 ;
        RECT 61.555 151.100 61.845 152.265 ;
        RECT 62.070 151.395 62.355 152.265 ;
        RECT 62.525 151.635 62.785 152.095 ;
        RECT 62.960 151.805 63.215 152.265 ;
        RECT 63.385 151.635 63.645 152.095 ;
        RECT 62.525 151.465 63.645 151.635 ;
        RECT 63.815 151.465 64.125 152.265 ;
        RECT 62.525 151.215 62.785 151.465 ;
        RECT 64.295 151.295 64.605 152.095 ;
        RECT 62.030 151.045 62.785 151.215 ;
        RECT 63.575 151.125 64.605 151.295 ;
        RECT 60.865 150.465 61.385 151.005 ;
        RECT 58.645 150.285 59.575 150.455 ;
        RECT 58.645 150.250 58.820 150.285 ;
        RECT 57.825 150.055 58.105 150.225 ;
        RECT 57.825 149.885 58.100 150.055 ;
        RECT 58.290 149.885 58.820 150.250 ;
        RECT 59.245 149.715 59.575 150.115 ;
        RECT 59.745 149.885 60.000 150.455 ;
        RECT 60.175 149.715 61.385 150.465 ;
        RECT 62.030 150.535 62.435 151.045 ;
        RECT 63.575 150.875 63.745 151.125 ;
        RECT 62.605 150.705 63.745 150.875 ;
        RECT 61.555 149.715 61.845 150.440 ;
        RECT 62.030 150.365 63.680 150.535 ;
        RECT 63.915 150.385 64.265 150.955 ;
        RECT 62.075 149.715 62.355 150.195 ;
        RECT 62.525 149.975 62.785 150.365 ;
        RECT 62.960 149.715 63.215 150.195 ;
        RECT 63.385 149.975 63.680 150.365 ;
        RECT 64.435 150.215 64.605 151.125 ;
        RECT 64.780 151.115 65.040 152.265 ;
        RECT 65.215 151.190 65.470 152.095 ;
        RECT 65.640 151.505 65.970 152.265 ;
        RECT 66.185 151.335 66.355 152.095 ;
        RECT 63.860 149.715 64.135 150.195 ;
        RECT 64.305 149.885 64.605 150.215 ;
        RECT 64.780 149.715 65.040 150.555 ;
        RECT 65.215 150.460 65.385 151.190 ;
        RECT 65.640 151.165 66.355 151.335 ;
        RECT 65.640 150.955 65.810 151.165 ;
        RECT 66.620 151.115 66.880 152.265 ;
        RECT 67.055 151.190 67.310 152.095 ;
        RECT 67.480 151.505 67.810 152.265 ;
        RECT 68.025 151.335 68.195 152.095 ;
        RECT 65.555 150.625 65.810 150.955 ;
        RECT 65.215 149.885 65.470 150.460 ;
        RECT 65.640 150.435 65.810 150.625 ;
        RECT 66.090 150.615 66.445 150.985 ;
        RECT 65.640 150.265 66.355 150.435 ;
        RECT 65.640 149.715 65.970 150.095 ;
        RECT 66.185 149.885 66.355 150.265 ;
        RECT 66.620 149.715 66.880 150.555 ;
        RECT 67.055 150.460 67.225 151.190 ;
        RECT 67.480 151.165 68.195 151.335 ;
        RECT 67.480 150.955 67.650 151.165 ;
        RECT 68.455 151.125 68.795 152.095 ;
        RECT 68.965 151.125 69.135 152.265 ;
        RECT 69.405 151.465 69.655 152.265 ;
        RECT 70.300 151.295 70.630 152.095 ;
        RECT 70.930 151.465 71.260 152.265 ;
        RECT 71.430 151.295 71.760 152.095 ;
        RECT 69.325 151.125 71.760 151.295 ;
        RECT 72.225 151.335 72.395 152.095 ;
        RECT 72.610 151.505 72.940 152.265 ;
        RECT 72.225 151.165 72.940 151.335 ;
        RECT 73.110 151.190 73.365 152.095 ;
        RECT 67.395 150.625 67.650 150.955 ;
        RECT 67.055 149.885 67.310 150.460 ;
        RECT 67.480 150.435 67.650 150.625 ;
        RECT 67.930 150.615 68.285 150.985 ;
        RECT 68.455 150.515 68.630 151.125 ;
        RECT 69.325 150.875 69.495 151.125 ;
        RECT 68.800 150.705 69.495 150.875 ;
        RECT 69.670 150.705 70.090 150.905 ;
        RECT 70.260 150.705 70.590 150.905 ;
        RECT 70.760 150.705 71.090 150.905 ;
        RECT 67.480 150.265 68.195 150.435 ;
        RECT 67.480 149.715 67.810 150.095 ;
        RECT 68.025 149.885 68.195 150.265 ;
        RECT 68.455 149.885 68.795 150.515 ;
        RECT 68.965 149.715 69.215 150.515 ;
        RECT 69.405 150.365 70.630 150.535 ;
        RECT 69.405 149.885 69.735 150.365 ;
        RECT 69.905 149.715 70.130 150.175 ;
        RECT 70.300 149.885 70.630 150.365 ;
        RECT 71.260 150.495 71.430 151.125 ;
        RECT 71.615 150.705 71.965 150.955 ;
        RECT 72.135 150.615 72.490 150.985 ;
        RECT 72.770 150.955 72.940 151.165 ;
        RECT 72.770 150.625 73.025 150.955 ;
        RECT 71.260 149.885 71.760 150.495 ;
        RECT 72.770 150.435 72.940 150.625 ;
        RECT 73.195 150.460 73.365 151.190 ;
        RECT 73.540 151.115 73.800 152.265 ;
        RECT 73.975 151.175 77.485 152.265 ;
        RECT 77.660 151.830 83.005 152.265 ;
        RECT 73.975 150.655 75.665 151.175 ;
        RECT 72.225 150.265 72.940 150.435 ;
        RECT 72.225 149.885 72.395 150.265 ;
        RECT 72.610 149.715 72.940 150.095 ;
        RECT 73.110 149.885 73.365 150.460 ;
        RECT 73.540 149.715 73.800 150.555 ;
        RECT 75.835 150.485 77.485 151.005 ;
        RECT 79.250 150.580 79.600 151.830 ;
        RECT 83.235 151.125 83.445 152.265 ;
        RECT 83.615 151.115 83.945 152.095 ;
        RECT 84.115 151.125 84.345 152.265 ;
        RECT 85.565 151.335 85.735 152.095 ;
        RECT 85.915 151.505 86.245 152.265 ;
        RECT 85.565 151.165 86.230 151.335 ;
        RECT 86.415 151.190 86.685 152.095 ;
        RECT 73.975 149.715 77.485 150.485 ;
        RECT 81.080 150.260 81.420 151.090 ;
        RECT 77.660 149.715 83.005 150.260 ;
        RECT 83.235 149.715 83.445 150.535 ;
        RECT 83.615 150.515 83.865 151.115 ;
        RECT 86.060 151.020 86.230 151.165 ;
        RECT 84.035 150.705 84.365 150.955 ;
        RECT 85.495 150.615 85.825 150.985 ;
        RECT 86.060 150.690 86.345 151.020 ;
        RECT 83.615 149.885 83.945 150.515 ;
        RECT 84.115 149.715 84.345 150.535 ;
        RECT 86.060 150.435 86.230 150.690 ;
        RECT 85.565 150.265 86.230 150.435 ;
        RECT 86.515 150.390 86.685 151.190 ;
        RECT 87.315 151.100 87.605 152.265 ;
        RECT 88.235 151.175 91.745 152.265 ;
        RECT 91.920 151.755 93.575 152.045 ;
        RECT 91.920 151.415 93.510 151.585 ;
        RECT 93.745 151.465 94.025 152.265 ;
        RECT 88.235 150.655 89.925 151.175 ;
        RECT 91.920 151.125 92.240 151.415 ;
        RECT 93.340 151.295 93.510 151.415 ;
        RECT 92.435 151.075 93.150 151.245 ;
        RECT 93.340 151.125 94.065 151.295 ;
        RECT 94.235 151.125 94.505 152.095 ;
        RECT 94.880 151.295 95.210 152.095 ;
        RECT 95.380 151.465 95.710 152.265 ;
        RECT 96.010 151.295 96.340 152.095 ;
        RECT 96.985 151.465 97.235 152.265 ;
        RECT 94.880 151.125 97.315 151.295 ;
        RECT 97.505 151.125 97.675 152.265 ;
        RECT 97.845 151.125 98.185 152.095 ;
        RECT 90.095 150.485 91.745 151.005 ;
        RECT 85.565 149.885 85.735 150.265 ;
        RECT 85.915 149.715 86.245 150.095 ;
        RECT 86.425 149.885 86.685 150.390 ;
        RECT 87.315 149.715 87.605 150.440 ;
        RECT 88.235 149.715 91.745 150.485 ;
        RECT 91.920 150.385 92.270 150.955 ;
        RECT 92.440 150.625 93.150 151.075 ;
        RECT 93.895 150.955 94.065 151.125 ;
        RECT 93.320 150.625 93.725 150.955 ;
        RECT 93.895 150.625 94.165 150.955 ;
        RECT 93.895 150.455 94.065 150.625 ;
        RECT 92.455 150.285 94.065 150.455 ;
        RECT 94.335 150.390 94.505 151.125 ;
        RECT 94.675 150.705 95.025 150.955 ;
        RECT 95.210 150.495 95.380 151.125 ;
        RECT 95.550 150.705 95.880 150.905 ;
        RECT 96.050 150.705 96.380 150.905 ;
        RECT 96.550 150.705 96.970 150.905 ;
        RECT 97.145 150.875 97.315 151.125 ;
        RECT 97.145 150.705 97.840 150.875 ;
        RECT 91.925 149.715 92.255 150.215 ;
        RECT 92.455 149.935 92.625 150.285 ;
        RECT 92.825 149.715 93.155 150.115 ;
        RECT 93.325 149.935 93.495 150.285 ;
        RECT 93.665 149.715 94.045 150.115 ;
        RECT 94.235 150.045 94.505 150.390 ;
        RECT 94.880 149.885 95.380 150.495 ;
        RECT 96.010 150.365 97.235 150.535 ;
        RECT 98.010 150.515 98.185 151.125 ;
        RECT 98.355 151.505 98.870 151.915 ;
        RECT 99.105 151.505 99.275 152.265 ;
        RECT 99.445 151.925 101.475 152.095 ;
        RECT 98.355 150.695 98.695 151.505 ;
        RECT 99.445 151.260 99.615 151.925 ;
        RECT 100.010 151.585 101.135 151.755 ;
        RECT 98.865 151.070 99.615 151.260 ;
        RECT 99.785 151.245 100.795 151.415 ;
        RECT 98.355 150.525 99.585 150.695 ;
        RECT 96.010 149.885 96.340 150.365 ;
        RECT 96.510 149.715 96.735 150.175 ;
        RECT 96.905 149.885 97.235 150.365 ;
        RECT 97.425 149.715 97.675 150.515 ;
        RECT 97.845 149.885 98.185 150.515 ;
        RECT 98.630 149.920 98.875 150.525 ;
        RECT 99.095 149.715 99.605 150.250 ;
        RECT 99.785 149.885 99.975 151.245 ;
        RECT 100.145 150.905 100.420 151.045 ;
        RECT 100.145 150.735 100.425 150.905 ;
        RECT 100.145 149.885 100.420 150.735 ;
        RECT 100.625 150.445 100.795 151.245 ;
        RECT 100.965 150.455 101.135 151.585 ;
        RECT 101.305 150.955 101.475 151.925 ;
        RECT 101.645 151.125 101.815 152.265 ;
        RECT 101.985 151.125 102.320 152.095 ;
        RECT 101.305 150.625 101.500 150.955 ;
        RECT 101.725 150.625 101.980 150.955 ;
        RECT 101.725 150.455 101.895 150.625 ;
        RECT 102.150 150.455 102.320 151.125 ;
        RECT 102.870 151.285 103.125 151.955 ;
        RECT 103.305 151.465 103.590 152.265 ;
        RECT 103.770 151.545 104.100 152.055 ;
        RECT 102.870 150.565 103.050 151.285 ;
        RECT 103.770 150.955 104.020 151.545 ;
        RECT 104.370 151.395 104.540 152.005 ;
        RECT 104.710 151.575 105.040 152.265 ;
        RECT 105.270 151.715 105.510 152.005 ;
        RECT 105.710 151.885 106.130 152.265 ;
        RECT 106.310 151.795 106.940 152.045 ;
        RECT 107.410 151.885 107.740 152.265 ;
        RECT 106.310 151.715 106.480 151.795 ;
        RECT 107.910 151.715 108.080 152.005 ;
        RECT 108.260 151.885 108.640 152.265 ;
        RECT 108.880 151.880 109.710 152.050 ;
        RECT 105.270 151.545 106.480 151.715 ;
        RECT 103.220 150.625 104.020 150.955 ;
        RECT 100.965 150.285 101.895 150.455 ;
        RECT 100.965 150.250 101.140 150.285 ;
        RECT 100.610 149.885 101.140 150.250 ;
        RECT 101.565 149.715 101.895 150.115 ;
        RECT 102.065 149.885 102.320 150.455 ;
        RECT 102.785 150.425 103.050 150.565 ;
        RECT 102.785 150.395 103.125 150.425 ;
        RECT 102.870 149.895 103.125 150.395 ;
        RECT 103.305 149.715 103.590 150.175 ;
        RECT 103.770 149.975 104.020 150.625 ;
        RECT 104.220 151.375 104.540 151.395 ;
        RECT 104.220 151.205 106.140 151.375 ;
        RECT 104.220 150.310 104.410 151.205 ;
        RECT 106.310 151.035 106.480 151.545 ;
        RECT 106.650 151.285 107.170 151.595 ;
        RECT 104.580 150.865 106.480 151.035 ;
        RECT 104.580 150.805 104.910 150.865 ;
        RECT 105.060 150.635 105.390 150.695 ;
        RECT 104.730 150.365 105.390 150.635 ;
        RECT 104.220 149.980 104.540 150.310 ;
        RECT 104.720 149.715 105.380 150.195 ;
        RECT 105.580 150.105 105.750 150.865 ;
        RECT 106.650 150.695 106.830 151.105 ;
        RECT 105.920 150.525 106.250 150.645 ;
        RECT 107.000 150.525 107.170 151.285 ;
        RECT 105.920 150.355 107.170 150.525 ;
        RECT 107.340 151.465 108.710 151.715 ;
        RECT 107.340 150.695 107.530 151.465 ;
        RECT 108.460 151.205 108.710 151.465 ;
        RECT 107.700 151.035 107.950 151.195 ;
        RECT 108.880 151.035 109.050 151.880 ;
        RECT 109.945 151.595 110.115 152.095 ;
        RECT 110.285 151.765 110.615 152.265 ;
        RECT 109.220 151.205 109.720 151.585 ;
        RECT 109.945 151.425 110.640 151.595 ;
        RECT 107.700 150.865 109.050 151.035 ;
        RECT 108.630 150.825 109.050 150.865 ;
        RECT 107.340 150.355 107.760 150.695 ;
        RECT 108.050 150.365 108.460 150.695 ;
        RECT 105.580 149.935 106.430 150.105 ;
        RECT 106.990 149.715 107.310 150.175 ;
        RECT 107.510 149.925 107.760 150.355 ;
        RECT 108.050 149.715 108.460 150.155 ;
        RECT 108.630 150.095 108.800 150.825 ;
        RECT 108.970 150.275 109.320 150.645 ;
        RECT 109.500 150.335 109.720 151.205 ;
        RECT 109.890 150.635 110.300 151.255 ;
        RECT 110.470 150.455 110.640 151.425 ;
        RECT 109.945 150.265 110.640 150.455 ;
        RECT 108.630 149.895 109.645 150.095 ;
        RECT 109.945 149.935 110.115 150.265 ;
        RECT 110.285 149.715 110.615 150.095 ;
        RECT 110.830 149.975 111.055 152.095 ;
        RECT 111.225 151.765 111.555 152.265 ;
        RECT 111.725 151.595 111.895 152.095 ;
        RECT 111.230 151.425 111.895 151.595 ;
        RECT 111.230 150.435 111.460 151.425 ;
        RECT 111.630 150.605 111.980 151.255 ;
        RECT 112.155 151.175 113.365 152.265 ;
        RECT 112.155 150.635 112.675 151.175 ;
        RECT 112.845 150.465 113.365 151.005 ;
        RECT 111.230 150.265 111.895 150.435 ;
        RECT 111.225 149.715 111.555 150.095 ;
        RECT 111.725 149.975 111.895 150.265 ;
        RECT 112.155 149.715 113.365 150.465 ;
        RECT 11.330 149.545 113.450 149.715 ;
        RECT 11.415 148.795 12.625 149.545 ;
        RECT 13.345 148.995 13.515 149.285 ;
        RECT 13.685 149.165 14.015 149.545 ;
        RECT 13.345 148.825 14.010 148.995 ;
        RECT 11.415 148.255 11.935 148.795 ;
        RECT 12.105 148.085 12.625 148.625 ;
        RECT 11.415 146.995 12.625 148.085 ;
        RECT 13.260 148.005 13.610 148.655 ;
        RECT 13.780 147.835 14.010 148.825 ;
        RECT 13.345 147.665 14.010 147.835 ;
        RECT 13.345 147.165 13.515 147.665 ;
        RECT 13.685 146.995 14.015 147.495 ;
        RECT 14.185 147.165 14.410 149.285 ;
        RECT 14.625 149.165 14.955 149.545 ;
        RECT 15.125 148.995 15.295 149.325 ;
        RECT 15.595 149.165 16.610 149.365 ;
        RECT 14.600 148.805 15.295 148.995 ;
        RECT 14.600 147.835 14.770 148.805 ;
        RECT 14.940 148.005 15.350 148.625 ;
        RECT 15.520 148.055 15.740 148.925 ;
        RECT 15.920 148.615 16.270 148.985 ;
        RECT 16.440 148.435 16.610 149.165 ;
        RECT 16.780 149.105 17.190 149.545 ;
        RECT 17.480 148.905 17.730 149.335 ;
        RECT 17.930 149.085 18.250 149.545 ;
        RECT 18.810 149.155 19.660 149.325 ;
        RECT 16.780 148.565 17.190 148.895 ;
        RECT 17.480 148.565 17.900 148.905 ;
        RECT 16.190 148.395 16.610 148.435 ;
        RECT 16.190 148.225 17.540 148.395 ;
        RECT 14.600 147.665 15.295 147.835 ;
        RECT 15.520 147.675 16.020 148.055 ;
        RECT 14.625 146.995 14.955 147.495 ;
        RECT 15.125 147.165 15.295 147.665 ;
        RECT 16.190 147.380 16.360 148.225 ;
        RECT 17.290 148.065 17.540 148.225 ;
        RECT 16.530 147.795 16.780 148.055 ;
        RECT 17.710 147.795 17.900 148.565 ;
        RECT 16.530 147.545 17.900 147.795 ;
        RECT 18.070 148.735 19.320 148.905 ;
        RECT 18.070 147.975 18.240 148.735 ;
        RECT 18.990 148.615 19.320 148.735 ;
        RECT 18.410 148.155 18.590 148.565 ;
        RECT 19.490 148.395 19.660 149.155 ;
        RECT 19.860 149.065 20.520 149.545 ;
        RECT 20.700 148.950 21.020 149.280 ;
        RECT 19.850 148.625 20.510 148.895 ;
        RECT 19.850 148.565 20.180 148.625 ;
        RECT 20.330 148.395 20.660 148.455 ;
        RECT 18.760 148.225 20.660 148.395 ;
        RECT 18.070 147.665 18.590 147.975 ;
        RECT 18.760 147.715 18.930 148.225 ;
        RECT 20.830 148.055 21.020 148.950 ;
        RECT 19.100 147.885 21.020 148.055 ;
        RECT 20.700 147.865 21.020 147.885 ;
        RECT 21.220 148.635 21.470 149.285 ;
        RECT 21.650 149.085 21.935 149.545 ;
        RECT 22.115 149.205 22.370 149.365 ;
        RECT 22.115 149.035 22.455 149.205 ;
        RECT 22.115 148.835 22.370 149.035 ;
        RECT 21.220 148.305 22.020 148.635 ;
        RECT 18.760 147.545 19.970 147.715 ;
        RECT 15.530 147.210 16.360 147.380 ;
        RECT 16.600 146.995 16.980 147.375 ;
        RECT 17.160 147.255 17.330 147.545 ;
        RECT 18.760 147.465 18.930 147.545 ;
        RECT 17.500 146.995 17.830 147.375 ;
        RECT 18.300 147.215 18.930 147.465 ;
        RECT 19.110 146.995 19.530 147.375 ;
        RECT 19.730 147.255 19.970 147.545 ;
        RECT 20.200 146.995 20.530 147.685 ;
        RECT 20.700 147.255 20.870 147.865 ;
        RECT 21.220 147.715 21.470 148.305 ;
        RECT 22.190 147.975 22.370 148.835 ;
        RECT 22.915 148.820 23.205 149.545 ;
        RECT 24.295 148.870 24.565 149.215 ;
        RECT 24.755 149.145 25.135 149.545 ;
        RECT 25.305 148.975 25.475 149.325 ;
        RECT 25.645 149.145 25.975 149.545 ;
        RECT 26.175 148.975 26.345 149.325 ;
        RECT 26.545 149.045 26.875 149.545 ;
        RECT 21.140 147.205 21.470 147.715 ;
        RECT 21.650 146.995 21.935 147.795 ;
        RECT 22.115 147.305 22.370 147.975 ;
        RECT 22.915 146.995 23.205 148.160 ;
        RECT 24.295 148.135 24.465 148.870 ;
        RECT 24.735 148.805 26.345 148.975 ;
        RECT 24.735 148.635 24.905 148.805 ;
        RECT 24.635 148.305 24.905 148.635 ;
        RECT 25.075 148.305 25.480 148.635 ;
        RECT 24.735 148.135 24.905 148.305 ;
        RECT 25.650 148.185 26.360 148.635 ;
        RECT 26.530 148.305 26.880 148.875 ;
        RECT 27.330 148.735 27.575 149.340 ;
        RECT 27.795 149.010 28.305 149.545 ;
        RECT 27.055 148.565 28.285 148.735 ;
        RECT 24.295 147.165 24.565 148.135 ;
        RECT 24.735 147.965 25.460 148.135 ;
        RECT 25.650 148.015 26.365 148.185 ;
        RECT 25.290 147.845 25.460 147.965 ;
        RECT 26.560 147.845 26.880 148.135 ;
        RECT 24.775 146.995 25.055 147.795 ;
        RECT 25.290 147.675 26.880 147.845 ;
        RECT 27.055 147.755 27.395 148.565 ;
        RECT 27.565 148.000 28.315 148.190 ;
        RECT 25.225 147.215 26.880 147.505 ;
        RECT 27.055 147.345 27.570 147.755 ;
        RECT 27.805 146.995 27.975 147.755 ;
        RECT 28.145 147.335 28.315 148.000 ;
        RECT 28.485 148.015 28.675 149.375 ;
        RECT 28.845 149.205 29.120 149.375 ;
        RECT 28.845 149.035 29.125 149.205 ;
        RECT 28.845 148.215 29.120 149.035 ;
        RECT 29.310 149.010 29.840 149.375 ;
        RECT 30.265 149.145 30.595 149.545 ;
        RECT 29.665 148.975 29.840 149.010 ;
        RECT 29.325 148.015 29.495 148.815 ;
        RECT 28.485 147.845 29.495 148.015 ;
        RECT 29.665 148.805 30.595 148.975 ;
        RECT 30.765 148.805 31.020 149.375 ;
        RECT 31.200 148.995 31.455 149.285 ;
        RECT 31.625 149.165 31.955 149.545 ;
        RECT 31.200 148.825 31.950 148.995 ;
        RECT 29.665 147.675 29.835 148.805 ;
        RECT 30.425 148.635 30.595 148.805 ;
        RECT 28.710 147.505 29.835 147.675 ;
        RECT 30.005 148.305 30.200 148.635 ;
        RECT 30.425 148.305 30.680 148.635 ;
        RECT 30.005 147.335 30.175 148.305 ;
        RECT 30.850 148.135 31.020 148.805 ;
        RECT 28.145 147.165 30.175 147.335 ;
        RECT 30.345 146.995 30.515 148.135 ;
        RECT 30.685 147.165 31.020 148.135 ;
        RECT 31.200 148.005 31.550 148.655 ;
        RECT 31.720 147.835 31.950 148.825 ;
        RECT 31.200 147.665 31.950 147.835 ;
        RECT 31.200 147.165 31.455 147.665 ;
        RECT 31.625 146.995 31.955 147.495 ;
        RECT 32.125 147.165 32.295 149.285 ;
        RECT 32.655 149.185 32.985 149.545 ;
        RECT 33.155 149.155 33.650 149.325 ;
        RECT 33.855 149.155 34.710 149.325 ;
        RECT 32.525 147.965 32.985 149.015 ;
        RECT 32.465 147.180 32.790 147.965 ;
        RECT 33.155 147.795 33.325 149.155 ;
        RECT 33.495 148.245 33.845 148.865 ;
        RECT 34.015 148.645 34.370 148.865 ;
        RECT 34.015 148.055 34.185 148.645 ;
        RECT 34.540 148.445 34.710 149.155 ;
        RECT 35.585 149.085 35.915 149.545 ;
        RECT 36.125 149.185 36.475 149.355 ;
        RECT 34.915 148.615 35.705 148.865 ;
        RECT 36.125 148.795 36.385 149.185 ;
        RECT 36.695 149.095 37.645 149.375 ;
        RECT 37.815 149.105 38.005 149.545 ;
        RECT 38.175 149.165 39.245 149.335 ;
        RECT 35.875 148.445 36.045 148.625 ;
        RECT 33.155 147.625 33.550 147.795 ;
        RECT 33.720 147.665 34.185 148.055 ;
        RECT 34.355 148.275 36.045 148.445 ;
        RECT 33.380 147.495 33.550 147.625 ;
        RECT 34.355 147.495 34.525 148.275 ;
        RECT 36.215 148.105 36.385 148.795 ;
        RECT 34.885 147.935 36.385 148.105 ;
        RECT 36.575 148.135 36.785 148.925 ;
        RECT 36.955 148.305 37.305 148.925 ;
        RECT 37.475 148.315 37.645 149.095 ;
        RECT 38.175 148.935 38.345 149.165 ;
        RECT 37.815 148.765 38.345 148.935 ;
        RECT 37.815 148.485 38.035 148.765 ;
        RECT 38.515 148.595 38.755 148.995 ;
        RECT 37.475 148.145 37.880 148.315 ;
        RECT 38.215 148.225 38.755 148.595 ;
        RECT 38.925 148.810 39.245 149.165 ;
        RECT 39.490 149.085 39.795 149.545 ;
        RECT 39.965 148.835 40.220 149.365 ;
        RECT 38.925 148.635 39.250 148.810 ;
        RECT 38.925 148.335 39.840 148.635 ;
        RECT 39.100 148.305 39.840 148.335 ;
        RECT 36.575 147.975 37.250 148.135 ;
        RECT 37.710 148.055 37.880 148.145 ;
        RECT 36.575 147.965 37.540 147.975 ;
        RECT 36.215 147.795 36.385 147.935 ;
        RECT 32.960 146.995 33.210 147.455 ;
        RECT 33.380 147.165 33.630 147.495 ;
        RECT 33.845 147.165 34.525 147.495 ;
        RECT 34.695 147.595 35.770 147.765 ;
        RECT 36.215 147.625 36.775 147.795 ;
        RECT 37.080 147.675 37.540 147.965 ;
        RECT 37.710 147.885 38.930 148.055 ;
        RECT 34.695 147.255 34.865 147.595 ;
        RECT 35.100 146.995 35.430 147.425 ;
        RECT 35.600 147.255 35.770 147.595 ;
        RECT 36.065 146.995 36.435 147.455 ;
        RECT 36.605 147.165 36.775 147.625 ;
        RECT 37.710 147.505 37.880 147.885 ;
        RECT 39.100 147.715 39.270 148.305 ;
        RECT 40.010 148.185 40.220 148.835 ;
        RECT 41.060 148.765 41.560 149.375 ;
        RECT 40.855 148.305 41.205 148.555 ;
        RECT 37.010 147.165 37.880 147.505 ;
        RECT 38.470 147.545 39.270 147.715 ;
        RECT 38.050 146.995 38.300 147.455 ;
        RECT 38.470 147.255 38.640 147.545 ;
        RECT 38.820 146.995 39.150 147.375 ;
        RECT 39.490 146.995 39.795 148.135 ;
        RECT 39.965 147.305 40.220 148.185 ;
        RECT 41.390 148.135 41.560 148.765 ;
        RECT 42.190 148.895 42.520 149.375 ;
        RECT 42.690 149.085 42.915 149.545 ;
        RECT 43.085 148.895 43.415 149.375 ;
        RECT 42.190 148.725 43.415 148.895 ;
        RECT 43.605 148.745 43.855 149.545 ;
        RECT 44.025 148.745 44.365 149.375 ;
        RECT 44.535 148.775 47.125 149.545 ;
        RECT 41.730 148.355 42.060 148.555 ;
        RECT 42.230 148.355 42.560 148.555 ;
        RECT 42.730 148.355 43.150 148.555 ;
        RECT 43.325 148.385 44.020 148.555 ;
        RECT 43.325 148.135 43.495 148.385 ;
        RECT 44.190 148.135 44.365 148.745 ;
        RECT 41.060 147.965 43.495 148.135 ;
        RECT 41.060 147.165 41.390 147.965 ;
        RECT 41.560 146.995 41.890 147.795 ;
        RECT 42.190 147.165 42.520 147.965 ;
        RECT 43.165 146.995 43.415 147.795 ;
        RECT 43.685 146.995 43.855 148.135 ;
        RECT 44.025 147.165 44.365 148.135 ;
        RECT 44.535 148.085 45.745 148.605 ;
        RECT 45.915 148.255 47.125 148.775 ;
        RECT 47.335 148.725 47.565 149.545 ;
        RECT 47.735 148.745 48.065 149.375 ;
        RECT 47.315 148.305 47.645 148.555 ;
        RECT 47.815 148.145 48.065 148.745 ;
        RECT 48.235 148.725 48.445 149.545 ;
        RECT 48.675 148.820 48.965 149.545 ;
        RECT 49.135 148.795 50.345 149.545 ;
        RECT 50.605 148.995 50.775 149.375 ;
        RECT 50.955 149.165 51.285 149.545 ;
        RECT 50.605 148.825 51.270 148.995 ;
        RECT 51.465 148.870 51.725 149.375 ;
        RECT 44.535 146.995 47.125 148.085 ;
        RECT 47.335 146.995 47.565 148.135 ;
        RECT 47.735 147.165 48.065 148.145 ;
        RECT 48.235 146.995 48.445 148.135 ;
        RECT 48.675 146.995 48.965 148.160 ;
        RECT 49.135 148.085 49.655 148.625 ;
        RECT 49.825 148.255 50.345 148.795 ;
        RECT 50.535 148.275 50.865 148.645 ;
        RECT 51.100 148.570 51.270 148.825 ;
        RECT 51.100 148.240 51.385 148.570 ;
        RECT 51.100 148.095 51.270 148.240 ;
        RECT 49.135 146.995 50.345 148.085 ;
        RECT 50.605 147.925 51.270 148.095 ;
        RECT 51.555 148.070 51.725 148.870 ;
        RECT 50.605 147.165 50.775 147.925 ;
        RECT 50.955 146.995 51.285 147.755 ;
        RECT 51.455 147.165 51.725 148.070 ;
        RECT 51.895 148.745 52.235 149.375 ;
        RECT 52.405 148.745 52.655 149.545 ;
        RECT 52.845 148.895 53.175 149.375 ;
        RECT 53.345 149.085 53.570 149.545 ;
        RECT 53.740 148.895 54.070 149.375 ;
        RECT 51.895 148.695 52.125 148.745 ;
        RECT 52.845 148.725 54.070 148.895 ;
        RECT 54.700 148.765 55.200 149.375 ;
        RECT 56.870 148.835 57.125 149.365 ;
        RECT 57.305 149.085 57.590 149.545 ;
        RECT 51.895 148.135 52.070 148.695 ;
        RECT 52.240 148.385 52.935 148.555 ;
        RECT 52.765 148.135 52.935 148.385 ;
        RECT 53.110 148.355 53.530 148.555 ;
        RECT 53.700 148.355 54.030 148.555 ;
        RECT 54.200 148.355 54.530 148.555 ;
        RECT 54.700 148.135 54.870 148.765 ;
        RECT 55.055 148.305 55.405 148.555 ;
        RECT 56.870 148.185 57.050 148.835 ;
        RECT 57.770 148.635 58.020 149.285 ;
        RECT 57.220 148.305 58.020 148.635 ;
        RECT 51.895 147.165 52.235 148.135 ;
        RECT 52.405 146.995 52.575 148.135 ;
        RECT 52.765 147.965 55.200 148.135 ;
        RECT 56.785 148.015 57.050 148.185 ;
        RECT 52.845 146.995 53.095 147.795 ;
        RECT 53.740 147.165 54.070 147.965 ;
        RECT 54.370 146.995 54.700 147.795 ;
        RECT 54.870 147.165 55.200 147.965 ;
        RECT 56.870 147.975 57.050 148.015 ;
        RECT 56.870 147.305 57.125 147.975 ;
        RECT 57.305 146.995 57.590 147.795 ;
        RECT 57.770 147.715 58.020 148.305 ;
        RECT 58.220 148.950 58.540 149.280 ;
        RECT 58.720 149.065 59.380 149.545 ;
        RECT 59.580 149.155 60.430 149.325 ;
        RECT 58.220 148.055 58.410 148.950 ;
        RECT 58.730 148.625 59.390 148.895 ;
        RECT 59.060 148.565 59.390 148.625 ;
        RECT 58.580 148.395 58.910 148.455 ;
        RECT 59.580 148.395 59.750 149.155 ;
        RECT 60.990 149.085 61.310 149.545 ;
        RECT 61.510 148.905 61.760 149.335 ;
        RECT 62.050 149.105 62.460 149.545 ;
        RECT 62.630 149.165 63.645 149.365 ;
        RECT 59.920 148.735 61.170 148.905 ;
        RECT 59.920 148.615 60.250 148.735 ;
        RECT 58.580 148.225 60.480 148.395 ;
        RECT 58.220 147.885 60.140 148.055 ;
        RECT 58.220 147.865 58.540 147.885 ;
        RECT 57.770 147.205 58.100 147.715 ;
        RECT 58.370 147.255 58.540 147.865 ;
        RECT 60.310 147.715 60.480 148.225 ;
        RECT 60.650 148.155 60.830 148.565 ;
        RECT 61.000 147.975 61.170 148.735 ;
        RECT 58.710 146.995 59.040 147.685 ;
        RECT 59.270 147.545 60.480 147.715 ;
        RECT 60.650 147.665 61.170 147.975 ;
        RECT 61.340 148.565 61.760 148.905 ;
        RECT 62.050 148.565 62.460 148.895 ;
        RECT 61.340 147.795 61.530 148.565 ;
        RECT 62.630 148.435 62.800 149.165 ;
        RECT 63.945 148.995 64.115 149.325 ;
        RECT 64.285 149.165 64.615 149.545 ;
        RECT 62.970 148.615 63.320 148.985 ;
        RECT 62.630 148.395 63.050 148.435 ;
        RECT 61.700 148.225 63.050 148.395 ;
        RECT 61.700 148.065 61.950 148.225 ;
        RECT 62.460 147.795 62.710 148.055 ;
        RECT 61.340 147.545 62.710 147.795 ;
        RECT 59.270 147.255 59.510 147.545 ;
        RECT 60.310 147.465 60.480 147.545 ;
        RECT 59.710 146.995 60.130 147.375 ;
        RECT 60.310 147.215 60.940 147.465 ;
        RECT 61.410 146.995 61.740 147.375 ;
        RECT 61.910 147.255 62.080 147.545 ;
        RECT 62.880 147.380 63.050 148.225 ;
        RECT 63.500 148.055 63.720 148.925 ;
        RECT 63.945 148.805 64.640 148.995 ;
        RECT 63.220 147.675 63.720 148.055 ;
        RECT 63.890 148.005 64.300 148.625 ;
        RECT 64.470 147.835 64.640 148.805 ;
        RECT 63.945 147.665 64.640 147.835 ;
        RECT 62.260 146.995 62.640 147.375 ;
        RECT 62.880 147.210 63.710 147.380 ;
        RECT 63.945 147.165 64.115 147.665 ;
        RECT 64.285 146.995 64.615 147.495 ;
        RECT 64.830 147.165 65.055 149.285 ;
        RECT 65.225 149.165 65.555 149.545 ;
        RECT 65.725 148.995 65.895 149.285 ;
        RECT 65.230 148.825 65.895 148.995 ;
        RECT 66.165 149.015 66.495 149.375 ;
        RECT 66.665 149.185 66.995 149.545 ;
        RECT 67.195 149.015 67.525 149.375 ;
        RECT 65.230 147.835 65.460 148.825 ;
        RECT 66.165 148.805 67.525 149.015 ;
        RECT 68.035 148.785 68.745 149.375 ;
        RECT 65.630 148.005 65.980 148.655 ;
        RECT 66.155 148.305 66.465 148.635 ;
        RECT 66.675 148.305 67.050 148.635 ;
        RECT 67.370 148.305 67.865 148.635 ;
        RECT 65.230 147.665 65.895 147.835 ;
        RECT 65.225 146.995 65.555 147.495 ;
        RECT 65.725 147.165 65.895 147.665 ;
        RECT 66.165 146.995 66.495 148.055 ;
        RECT 66.675 147.380 66.845 148.305 ;
        RECT 67.015 147.815 67.345 148.035 ;
        RECT 67.540 148.015 67.865 148.305 ;
        RECT 68.040 148.015 68.370 148.555 ;
        RECT 68.540 147.815 68.745 148.785 ;
        RECT 67.015 147.585 68.745 147.815 ;
        RECT 67.015 147.185 67.345 147.585 ;
        RECT 67.515 146.995 67.845 147.355 ;
        RECT 68.045 147.165 68.745 147.585 ;
        RECT 68.915 149.045 69.215 149.375 ;
        RECT 69.385 149.065 69.660 149.545 ;
        RECT 68.915 148.135 69.085 149.045 ;
        RECT 69.840 148.895 70.135 149.285 ;
        RECT 70.305 149.065 70.560 149.545 ;
        RECT 70.735 148.895 70.995 149.285 ;
        RECT 71.165 149.065 71.445 149.545 ;
        RECT 69.255 148.305 69.605 148.875 ;
        RECT 69.840 148.725 71.490 148.895 ;
        RECT 71.675 148.775 74.265 149.545 ;
        RECT 74.435 148.820 74.725 149.545 ;
        RECT 74.895 148.795 76.105 149.545 ;
        RECT 69.775 148.385 70.915 148.555 ;
        RECT 69.775 148.135 69.945 148.385 ;
        RECT 71.085 148.215 71.490 148.725 ;
        RECT 68.915 147.965 69.945 148.135 ;
        RECT 70.735 148.045 71.490 148.215 ;
        RECT 71.675 148.085 72.885 148.605 ;
        RECT 73.055 148.255 74.265 148.775 ;
        RECT 68.915 147.165 69.225 147.965 ;
        RECT 70.735 147.795 70.995 148.045 ;
        RECT 69.395 146.995 69.705 147.795 ;
        RECT 69.875 147.625 70.995 147.795 ;
        RECT 69.875 147.165 70.135 147.625 ;
        RECT 70.305 146.995 70.560 147.455 ;
        RECT 70.735 147.165 70.995 147.625 ;
        RECT 71.165 146.995 71.450 147.865 ;
        RECT 71.675 146.995 74.265 148.085 ;
        RECT 74.435 146.995 74.725 148.160 ;
        RECT 74.895 148.085 75.415 148.625 ;
        RECT 75.585 148.255 76.105 148.795 ;
        RECT 76.550 148.735 76.795 149.340 ;
        RECT 77.015 149.010 77.525 149.545 ;
        RECT 76.275 148.565 77.505 148.735 ;
        RECT 74.895 146.995 76.105 148.085 ;
        RECT 76.275 147.755 76.615 148.565 ;
        RECT 76.785 148.000 77.535 148.190 ;
        RECT 76.275 147.345 76.790 147.755 ;
        RECT 77.025 146.995 77.195 147.755 ;
        RECT 77.365 147.335 77.535 148.000 ;
        RECT 77.705 148.015 77.895 149.375 ;
        RECT 78.065 148.525 78.340 149.375 ;
        RECT 78.530 149.010 79.060 149.375 ;
        RECT 79.485 149.145 79.815 149.545 ;
        RECT 78.885 148.975 79.060 149.010 ;
        RECT 78.065 148.355 78.345 148.525 ;
        RECT 78.065 148.215 78.340 148.355 ;
        RECT 78.545 148.015 78.715 148.815 ;
        RECT 77.705 147.845 78.715 148.015 ;
        RECT 78.885 148.805 79.815 148.975 ;
        RECT 79.985 148.805 80.240 149.375 ;
        RECT 78.885 147.675 79.055 148.805 ;
        RECT 79.645 148.635 79.815 148.805 ;
        RECT 77.930 147.505 79.055 147.675 ;
        RECT 79.225 148.305 79.420 148.635 ;
        RECT 79.645 148.305 79.900 148.635 ;
        RECT 79.225 147.335 79.395 148.305 ;
        RECT 80.070 148.135 80.240 148.805 ;
        RECT 77.365 147.165 79.395 147.335 ;
        RECT 79.565 146.995 79.735 148.135 ;
        RECT 79.905 147.165 80.240 148.135 ;
        RECT 80.420 148.835 80.675 149.365 ;
        RECT 80.845 149.085 81.150 149.545 ;
        RECT 81.395 149.165 82.465 149.335 ;
        RECT 80.420 148.185 80.630 148.835 ;
        RECT 81.395 148.810 81.715 149.165 ;
        RECT 81.390 148.635 81.715 148.810 ;
        RECT 80.800 148.335 81.715 148.635 ;
        RECT 81.885 148.595 82.125 148.995 ;
        RECT 82.295 148.935 82.465 149.165 ;
        RECT 82.635 149.105 82.825 149.545 ;
        RECT 82.995 149.095 83.945 149.375 ;
        RECT 84.165 149.185 84.515 149.355 ;
        RECT 82.295 148.765 82.825 148.935 ;
        RECT 80.800 148.305 81.540 148.335 ;
        RECT 80.420 147.305 80.675 148.185 ;
        RECT 80.845 146.995 81.150 148.135 ;
        RECT 81.370 147.715 81.540 148.305 ;
        RECT 81.885 148.225 82.425 148.595 ;
        RECT 82.605 148.485 82.825 148.765 ;
        RECT 82.995 148.315 83.165 149.095 ;
        RECT 82.760 148.145 83.165 148.315 ;
        RECT 83.335 148.305 83.685 148.925 ;
        RECT 82.760 148.055 82.930 148.145 ;
        RECT 83.855 148.135 84.065 148.925 ;
        RECT 81.710 147.885 82.930 148.055 ;
        RECT 83.390 147.975 84.065 148.135 ;
        RECT 81.370 147.545 82.170 147.715 ;
        RECT 81.490 146.995 81.820 147.375 ;
        RECT 82.000 147.255 82.170 147.545 ;
        RECT 82.760 147.505 82.930 147.885 ;
        RECT 83.100 147.965 84.065 147.975 ;
        RECT 84.255 148.795 84.515 149.185 ;
        RECT 84.725 149.085 85.055 149.545 ;
        RECT 85.930 149.155 86.785 149.325 ;
        RECT 86.990 149.155 87.485 149.325 ;
        RECT 87.655 149.185 87.985 149.545 ;
        RECT 84.255 148.105 84.425 148.795 ;
        RECT 84.595 148.445 84.765 148.625 ;
        RECT 84.935 148.615 85.725 148.865 ;
        RECT 85.930 148.445 86.100 149.155 ;
        RECT 86.270 148.645 86.625 148.865 ;
        RECT 84.595 148.275 86.285 148.445 ;
        RECT 83.100 147.675 83.560 147.965 ;
        RECT 84.255 147.935 85.755 148.105 ;
        RECT 84.255 147.795 84.425 147.935 ;
        RECT 83.865 147.625 84.425 147.795 ;
        RECT 82.340 146.995 82.590 147.455 ;
        RECT 82.760 147.165 83.630 147.505 ;
        RECT 83.865 147.165 84.035 147.625 ;
        RECT 84.870 147.595 85.945 147.765 ;
        RECT 84.205 146.995 84.575 147.455 ;
        RECT 84.870 147.255 85.040 147.595 ;
        RECT 85.210 146.995 85.540 147.425 ;
        RECT 85.775 147.255 85.945 147.595 ;
        RECT 86.115 147.495 86.285 148.275 ;
        RECT 86.455 148.055 86.625 148.645 ;
        RECT 86.795 148.245 87.145 148.865 ;
        RECT 86.455 147.665 86.920 148.055 ;
        RECT 87.315 147.795 87.485 149.155 ;
        RECT 87.655 147.965 88.115 149.015 ;
        RECT 87.090 147.625 87.485 147.795 ;
        RECT 87.090 147.495 87.260 147.625 ;
        RECT 86.115 147.165 86.795 147.495 ;
        RECT 87.010 147.165 87.260 147.495 ;
        RECT 87.430 146.995 87.680 147.455 ;
        RECT 87.850 147.180 88.175 147.965 ;
        RECT 88.345 147.165 88.515 149.285 ;
        RECT 88.685 149.165 89.015 149.545 ;
        RECT 89.185 148.995 89.440 149.285 ;
        RECT 88.690 148.825 89.440 148.995 ;
        RECT 89.730 148.915 90.015 149.375 ;
        RECT 90.185 149.085 90.455 149.545 ;
        RECT 88.690 147.835 88.920 148.825 ;
        RECT 89.730 148.745 90.685 148.915 ;
        RECT 89.090 148.005 89.440 148.655 ;
        RECT 89.615 148.015 90.305 148.575 ;
        RECT 90.475 147.845 90.685 148.745 ;
        RECT 88.690 147.665 89.440 147.835 ;
        RECT 88.685 146.995 89.015 147.495 ;
        RECT 89.185 147.165 89.440 147.665 ;
        RECT 89.730 147.625 90.685 147.845 ;
        RECT 90.855 148.575 91.255 149.375 ;
        RECT 91.445 148.915 91.725 149.375 ;
        RECT 92.245 149.085 92.570 149.545 ;
        RECT 91.445 148.745 92.570 148.915 ;
        RECT 92.740 148.805 93.125 149.375 ;
        RECT 92.120 148.635 92.570 148.745 ;
        RECT 90.855 148.015 91.950 148.575 ;
        RECT 92.120 148.305 92.675 148.635 ;
        RECT 89.730 147.165 90.015 147.625 ;
        RECT 90.185 146.995 90.455 147.455 ;
        RECT 90.855 147.165 91.255 148.015 ;
        RECT 92.120 147.845 92.570 148.305 ;
        RECT 92.845 148.135 93.125 148.805 ;
        RECT 91.445 147.625 92.570 147.845 ;
        RECT 91.445 147.165 91.725 147.625 ;
        RECT 92.245 146.995 92.570 147.455 ;
        RECT 92.740 147.165 93.125 148.135 ;
        RECT 93.755 148.745 94.095 149.375 ;
        RECT 94.265 148.745 94.515 149.545 ;
        RECT 94.705 148.895 95.035 149.375 ;
        RECT 95.205 149.085 95.430 149.545 ;
        RECT 95.600 148.895 95.930 149.375 ;
        RECT 93.755 148.695 93.985 148.745 ;
        RECT 94.705 148.725 95.930 148.895 ;
        RECT 96.560 148.765 97.060 149.375 ;
        RECT 97.445 149.045 97.775 149.545 ;
        RECT 97.975 148.975 98.145 149.325 ;
        RECT 98.345 149.145 98.675 149.545 ;
        RECT 98.845 148.975 99.015 149.325 ;
        RECT 99.185 149.145 99.565 149.545 ;
        RECT 93.755 148.135 93.930 148.695 ;
        RECT 94.100 148.385 94.795 148.555 ;
        RECT 94.625 148.135 94.795 148.385 ;
        RECT 94.970 148.355 95.390 148.555 ;
        RECT 95.560 148.355 95.890 148.555 ;
        RECT 96.060 148.355 96.390 148.555 ;
        RECT 96.560 148.135 96.730 148.765 ;
        RECT 96.915 148.305 97.265 148.555 ;
        RECT 97.440 148.305 97.790 148.875 ;
        RECT 97.975 148.805 99.585 148.975 ;
        RECT 99.755 148.870 100.025 149.215 ;
        RECT 99.415 148.635 99.585 148.805 ;
        RECT 97.960 148.185 98.670 148.635 ;
        RECT 98.840 148.305 99.245 148.635 ;
        RECT 99.415 148.305 99.685 148.635 ;
        RECT 93.755 147.165 94.095 148.135 ;
        RECT 94.265 146.995 94.435 148.135 ;
        RECT 94.625 147.965 97.060 148.135 ;
        RECT 94.705 146.995 94.955 147.795 ;
        RECT 95.600 147.165 95.930 147.965 ;
        RECT 96.230 146.995 96.560 147.795 ;
        RECT 96.730 147.165 97.060 147.965 ;
        RECT 97.440 147.845 97.760 148.135 ;
        RECT 97.955 148.015 98.670 148.185 ;
        RECT 99.415 148.135 99.585 148.305 ;
        RECT 99.855 148.135 100.025 148.870 ;
        RECT 100.195 148.820 100.485 149.545 ;
        RECT 100.655 148.775 102.325 149.545 ;
        RECT 98.860 147.965 99.585 148.135 ;
        RECT 98.860 147.845 99.030 147.965 ;
        RECT 97.440 147.675 99.030 147.845 ;
        RECT 97.440 147.215 99.095 147.505 ;
        RECT 99.265 146.995 99.545 147.795 ;
        RECT 99.755 147.165 100.025 148.135 ;
        RECT 100.195 146.995 100.485 148.160 ;
        RECT 100.655 148.085 101.405 148.605 ;
        RECT 101.575 148.255 102.325 148.775 ;
        RECT 102.770 148.735 103.015 149.340 ;
        RECT 103.235 149.010 103.745 149.545 ;
        RECT 102.495 148.565 103.725 148.735 ;
        RECT 100.655 146.995 102.325 148.085 ;
        RECT 102.495 147.755 102.835 148.565 ;
        RECT 103.005 148.000 103.755 148.190 ;
        RECT 102.495 147.345 103.010 147.755 ;
        RECT 103.245 146.995 103.415 147.755 ;
        RECT 103.585 147.335 103.755 148.000 ;
        RECT 103.925 148.015 104.115 149.375 ;
        RECT 104.285 148.865 104.560 149.375 ;
        RECT 104.750 149.010 105.280 149.375 ;
        RECT 105.705 149.145 106.035 149.545 ;
        RECT 105.105 148.975 105.280 149.010 ;
        RECT 104.285 148.695 104.565 148.865 ;
        RECT 104.285 148.215 104.560 148.695 ;
        RECT 104.765 148.015 104.935 148.815 ;
        RECT 103.925 147.845 104.935 148.015 ;
        RECT 105.105 148.805 106.035 148.975 ;
        RECT 106.205 148.805 106.460 149.375 ;
        RECT 105.105 147.675 105.275 148.805 ;
        RECT 105.865 148.635 106.035 148.805 ;
        RECT 104.150 147.505 105.275 147.675 ;
        RECT 105.445 148.305 105.640 148.635 ;
        RECT 105.865 148.305 106.120 148.635 ;
        RECT 105.445 147.335 105.615 148.305 ;
        RECT 106.290 148.135 106.460 148.805 ;
        RECT 106.635 148.795 107.845 149.545 ;
        RECT 108.105 148.995 108.275 149.375 ;
        RECT 108.455 149.165 108.785 149.545 ;
        RECT 108.105 148.825 108.770 148.995 ;
        RECT 108.965 148.870 109.225 149.375 ;
        RECT 103.585 147.165 105.615 147.335 ;
        RECT 105.785 146.995 105.955 148.135 ;
        RECT 106.125 147.165 106.460 148.135 ;
        RECT 106.635 148.085 107.155 148.625 ;
        RECT 107.325 148.255 107.845 148.795 ;
        RECT 108.035 148.275 108.365 148.645 ;
        RECT 108.600 148.570 108.770 148.825 ;
        RECT 108.600 148.240 108.885 148.570 ;
        RECT 108.600 148.095 108.770 148.240 ;
        RECT 106.635 146.995 107.845 148.085 ;
        RECT 108.105 147.925 108.770 148.095 ;
        RECT 109.055 148.070 109.225 148.870 ;
        RECT 109.395 148.775 111.985 149.545 ;
        RECT 112.155 148.795 113.365 149.545 ;
        RECT 108.105 147.165 108.275 147.925 ;
        RECT 108.455 146.995 108.785 147.755 ;
        RECT 108.955 147.165 109.225 148.070 ;
        RECT 109.395 148.085 110.605 148.605 ;
        RECT 110.775 148.255 111.985 148.775 ;
        RECT 112.155 148.085 112.675 148.625 ;
        RECT 112.845 148.255 113.365 148.795 ;
        RECT 109.395 146.995 111.985 148.085 ;
        RECT 112.155 146.995 113.365 148.085 ;
        RECT 11.330 146.825 113.450 146.995 ;
        RECT 11.415 145.735 12.625 146.825 ;
        RECT 11.415 145.025 11.935 145.565 ;
        RECT 12.105 145.195 12.625 145.735 ;
        RECT 13.755 145.685 13.985 146.825 ;
        RECT 14.155 145.675 14.485 146.655 ;
        RECT 14.655 145.685 14.865 146.825 ;
        RECT 15.095 145.750 15.365 146.655 ;
        RECT 15.535 146.065 15.865 146.825 ;
        RECT 16.045 145.895 16.215 146.655 ;
        RECT 16.590 146.195 16.875 146.655 ;
        RECT 17.045 146.365 17.315 146.825 ;
        RECT 16.590 145.975 17.545 146.195 ;
        RECT 13.735 145.265 14.065 145.515 ;
        RECT 11.415 144.275 12.625 145.025 ;
        RECT 13.755 144.275 13.985 145.095 ;
        RECT 14.235 145.075 14.485 145.675 ;
        RECT 14.155 144.445 14.485 145.075 ;
        RECT 14.655 144.275 14.865 145.095 ;
        RECT 15.095 144.950 15.265 145.750 ;
        RECT 15.550 145.725 16.215 145.895 ;
        RECT 15.550 145.580 15.720 145.725 ;
        RECT 15.435 145.250 15.720 145.580 ;
        RECT 15.550 144.995 15.720 145.250 ;
        RECT 15.955 145.175 16.285 145.545 ;
        RECT 16.475 145.245 17.165 145.805 ;
        RECT 17.335 145.075 17.545 145.975 ;
        RECT 15.095 144.445 15.355 144.950 ;
        RECT 15.550 144.825 16.215 144.995 ;
        RECT 15.535 144.275 15.865 144.655 ;
        RECT 16.045 144.445 16.215 144.825 ;
        RECT 16.590 144.905 17.545 145.075 ;
        RECT 17.715 145.805 18.115 146.655 ;
        RECT 18.305 146.195 18.585 146.655 ;
        RECT 19.105 146.365 19.430 146.825 ;
        RECT 18.305 145.975 19.430 146.195 ;
        RECT 17.715 145.245 18.810 145.805 ;
        RECT 18.980 145.515 19.430 145.975 ;
        RECT 19.600 145.685 19.985 146.655 ;
        RECT 16.590 144.445 16.875 144.905 ;
        RECT 17.045 144.275 17.315 144.735 ;
        RECT 17.715 144.445 18.115 145.245 ;
        RECT 18.980 145.185 19.535 145.515 ;
        RECT 18.980 145.075 19.430 145.185 ;
        RECT 18.305 144.905 19.430 145.075 ;
        RECT 19.705 145.015 19.985 145.685 ;
        RECT 18.305 144.445 18.585 144.905 ;
        RECT 19.105 144.275 19.430 144.735 ;
        RECT 19.600 144.445 19.985 145.015 ;
        RECT 20.160 145.685 20.495 146.655 ;
        RECT 20.665 145.685 20.835 146.825 ;
        RECT 21.005 146.485 23.035 146.655 ;
        RECT 20.160 145.015 20.330 145.685 ;
        RECT 21.005 145.515 21.175 146.485 ;
        RECT 20.500 145.185 20.755 145.515 ;
        RECT 20.980 145.185 21.175 145.515 ;
        RECT 21.345 146.145 22.470 146.315 ;
        RECT 20.585 145.015 20.755 145.185 ;
        RECT 21.345 145.015 21.515 146.145 ;
        RECT 20.160 144.445 20.415 145.015 ;
        RECT 20.585 144.845 21.515 145.015 ;
        RECT 21.685 145.805 22.695 145.975 ;
        RECT 21.685 145.005 21.855 145.805 ;
        RECT 22.060 145.465 22.335 145.605 ;
        RECT 22.055 145.295 22.335 145.465 ;
        RECT 21.340 144.810 21.515 144.845 ;
        RECT 20.585 144.275 20.915 144.675 ;
        RECT 21.340 144.445 21.870 144.810 ;
        RECT 22.060 144.445 22.335 145.295 ;
        RECT 22.505 144.445 22.695 145.805 ;
        RECT 22.865 145.820 23.035 146.485 ;
        RECT 23.205 146.065 23.375 146.825 ;
        RECT 23.610 146.065 24.125 146.475 ;
        RECT 22.865 145.630 23.615 145.820 ;
        RECT 23.785 145.255 24.125 146.065 ;
        RECT 22.895 145.085 24.125 145.255 ;
        RECT 24.295 145.735 26.885 146.825 ;
        RECT 27.170 146.195 27.455 146.655 ;
        RECT 27.625 146.365 27.895 146.825 ;
        RECT 27.170 145.975 28.125 146.195 ;
        RECT 24.295 145.215 25.505 145.735 ;
        RECT 22.875 144.275 23.385 144.810 ;
        RECT 23.605 144.480 23.850 145.085 ;
        RECT 25.675 145.045 26.885 145.565 ;
        RECT 27.055 145.245 27.745 145.805 ;
        RECT 27.915 145.075 28.125 145.975 ;
        RECT 24.295 144.275 26.885 145.045 ;
        RECT 27.170 144.905 28.125 145.075 ;
        RECT 28.295 145.805 28.695 146.655 ;
        RECT 28.885 146.195 29.165 146.655 ;
        RECT 29.685 146.365 30.010 146.825 ;
        RECT 28.885 145.975 30.010 146.195 ;
        RECT 28.295 145.245 29.390 145.805 ;
        RECT 29.560 145.515 30.010 145.975 ;
        RECT 30.180 145.685 30.565 146.655 ;
        RECT 27.170 144.445 27.455 144.905 ;
        RECT 27.625 144.275 27.895 144.735 ;
        RECT 28.295 144.445 28.695 145.245 ;
        RECT 29.560 145.185 30.115 145.515 ;
        RECT 29.560 145.075 30.010 145.185 ;
        RECT 28.885 144.905 30.010 145.075 ;
        RECT 30.285 145.015 30.565 145.685 ;
        RECT 28.885 144.445 29.165 144.905 ;
        RECT 29.685 144.275 30.010 144.735 ;
        RECT 30.180 144.445 30.565 145.015 ;
        RECT 30.735 145.685 31.120 146.655 ;
        RECT 31.290 146.365 31.615 146.825 ;
        RECT 32.135 146.195 32.415 146.655 ;
        RECT 31.290 145.975 32.415 146.195 ;
        RECT 30.735 145.015 31.015 145.685 ;
        RECT 31.290 145.515 31.740 145.975 ;
        RECT 32.605 145.805 33.005 146.655 ;
        RECT 33.405 146.365 33.675 146.825 ;
        RECT 33.845 146.195 34.130 146.655 ;
        RECT 31.185 145.185 31.740 145.515 ;
        RECT 31.910 145.245 33.005 145.805 ;
        RECT 31.290 145.075 31.740 145.185 ;
        RECT 30.735 144.445 31.120 145.015 ;
        RECT 31.290 144.905 32.415 145.075 ;
        RECT 31.290 144.275 31.615 144.735 ;
        RECT 32.135 144.445 32.415 144.905 ;
        RECT 32.605 144.445 33.005 145.245 ;
        RECT 33.175 145.975 34.130 146.195 ;
        RECT 33.175 145.075 33.385 145.975 ;
        RECT 33.555 145.245 34.245 145.805 ;
        RECT 34.415 145.750 34.685 146.655 ;
        RECT 34.855 146.065 35.185 146.825 ;
        RECT 35.365 145.895 35.535 146.655 ;
        RECT 33.175 144.905 34.130 145.075 ;
        RECT 33.405 144.275 33.675 144.735 ;
        RECT 33.845 144.445 34.130 144.905 ;
        RECT 34.415 144.950 34.585 145.750 ;
        RECT 34.870 145.725 35.535 145.895 ;
        RECT 34.870 145.580 35.040 145.725 ;
        RECT 35.795 145.660 36.085 146.825 ;
        RECT 37.175 145.750 37.445 146.655 ;
        RECT 37.615 146.065 37.945 146.825 ;
        RECT 38.125 145.895 38.295 146.655 ;
        RECT 34.755 145.250 35.040 145.580 ;
        RECT 34.870 144.995 35.040 145.250 ;
        RECT 35.275 145.175 35.605 145.545 ;
        RECT 34.415 144.445 34.675 144.950 ;
        RECT 34.870 144.825 35.535 144.995 ;
        RECT 34.855 144.275 35.185 144.655 ;
        RECT 35.365 144.445 35.535 144.825 ;
        RECT 35.795 144.275 36.085 145.000 ;
        RECT 37.175 144.950 37.345 145.750 ;
        RECT 37.630 145.725 38.295 145.895 ;
        RECT 38.760 145.855 39.090 146.655 ;
        RECT 39.260 146.025 39.590 146.825 ;
        RECT 39.890 145.855 40.220 146.655 ;
        RECT 40.865 146.025 41.115 146.825 ;
        RECT 37.630 145.580 37.800 145.725 ;
        RECT 38.760 145.685 41.195 145.855 ;
        RECT 41.385 145.685 41.555 146.825 ;
        RECT 41.725 145.685 42.065 146.655 ;
        RECT 37.515 145.250 37.800 145.580 ;
        RECT 37.630 144.995 37.800 145.250 ;
        RECT 38.035 145.175 38.365 145.545 ;
        RECT 38.555 145.265 38.905 145.515 ;
        RECT 39.090 145.055 39.260 145.685 ;
        RECT 39.430 145.265 39.760 145.465 ;
        RECT 39.930 145.265 40.260 145.465 ;
        RECT 40.430 145.265 40.850 145.465 ;
        RECT 41.025 145.435 41.195 145.685 ;
        RECT 41.025 145.265 41.720 145.435 ;
        RECT 37.175 144.445 37.435 144.950 ;
        RECT 37.630 144.825 38.295 144.995 ;
        RECT 37.615 144.275 37.945 144.655 ;
        RECT 38.125 144.445 38.295 144.825 ;
        RECT 38.760 144.445 39.260 145.055 ;
        RECT 39.890 144.925 41.115 145.095 ;
        RECT 41.890 145.075 42.065 145.685 ;
        RECT 42.695 145.735 45.285 146.825 ;
        RECT 45.460 146.390 50.805 146.825 ;
        RECT 42.695 145.215 43.905 145.735 ;
        RECT 39.890 144.445 40.220 144.925 ;
        RECT 40.390 144.275 40.615 144.735 ;
        RECT 40.785 144.445 41.115 144.925 ;
        RECT 41.305 144.275 41.555 145.075 ;
        RECT 41.725 144.445 42.065 145.075 ;
        RECT 44.075 145.045 45.285 145.565 ;
        RECT 47.050 145.140 47.400 146.390 ;
        RECT 50.975 145.685 51.315 146.655 ;
        RECT 51.485 145.685 51.655 146.825 ;
        RECT 51.925 146.025 52.175 146.825 ;
        RECT 52.820 145.855 53.150 146.655 ;
        RECT 53.450 146.025 53.780 146.825 ;
        RECT 53.950 145.855 54.280 146.655 ;
        RECT 51.845 145.685 54.280 145.855 ;
        RECT 54.655 145.735 55.865 146.825 ;
        RECT 56.035 146.065 56.550 146.475 ;
        RECT 56.785 146.065 56.955 146.825 ;
        RECT 57.125 146.485 59.155 146.655 ;
        RECT 42.695 144.275 45.285 145.045 ;
        RECT 48.880 144.820 49.220 145.650 ;
        RECT 50.975 145.075 51.150 145.685 ;
        RECT 51.845 145.435 52.015 145.685 ;
        RECT 51.320 145.265 52.015 145.435 ;
        RECT 52.190 145.265 52.610 145.465 ;
        RECT 52.780 145.265 53.110 145.465 ;
        RECT 53.280 145.265 53.610 145.465 ;
        RECT 45.460 144.275 50.805 144.820 ;
        RECT 50.975 144.445 51.315 145.075 ;
        RECT 51.485 144.275 51.735 145.075 ;
        RECT 51.925 144.925 53.150 145.095 ;
        RECT 51.925 144.445 52.255 144.925 ;
        RECT 52.425 144.275 52.650 144.735 ;
        RECT 52.820 144.445 53.150 144.925 ;
        RECT 53.780 145.055 53.950 145.685 ;
        RECT 54.135 145.265 54.485 145.515 ;
        RECT 54.655 145.195 55.175 145.735 ;
        RECT 53.780 144.445 54.280 145.055 ;
        RECT 55.345 145.025 55.865 145.565 ;
        RECT 56.035 145.255 56.375 146.065 ;
        RECT 57.125 145.820 57.295 146.485 ;
        RECT 57.690 146.145 58.815 146.315 ;
        RECT 56.545 145.630 57.295 145.820 ;
        RECT 57.465 145.805 58.475 145.975 ;
        RECT 56.035 145.085 57.265 145.255 ;
        RECT 54.655 144.275 55.865 145.025 ;
        RECT 56.310 144.480 56.555 145.085 ;
        RECT 56.775 144.275 57.285 144.810 ;
        RECT 57.465 144.445 57.655 145.805 ;
        RECT 57.825 145.125 58.100 145.605 ;
        RECT 57.825 144.955 58.105 145.125 ;
        RECT 58.305 145.005 58.475 145.805 ;
        RECT 58.645 145.015 58.815 146.145 ;
        RECT 58.985 145.515 59.155 146.485 ;
        RECT 59.325 145.685 59.495 146.825 ;
        RECT 59.665 145.685 60.000 146.655 ;
        RECT 60.235 145.685 60.445 146.825 ;
        RECT 58.985 145.185 59.180 145.515 ;
        RECT 59.405 145.185 59.660 145.515 ;
        RECT 59.405 145.015 59.575 145.185 ;
        RECT 59.830 145.015 60.000 145.685 ;
        RECT 60.615 145.675 60.945 146.655 ;
        RECT 61.115 145.685 61.345 146.825 ;
        RECT 57.825 144.445 58.100 144.955 ;
        RECT 58.645 144.845 59.575 145.015 ;
        RECT 58.645 144.810 58.820 144.845 ;
        RECT 58.290 144.445 58.820 144.810 ;
        RECT 59.245 144.275 59.575 144.675 ;
        RECT 59.745 144.445 60.000 145.015 ;
        RECT 60.235 144.275 60.445 145.095 ;
        RECT 60.615 145.075 60.865 145.675 ;
        RECT 61.555 145.660 61.845 146.825 ;
        RECT 62.480 145.675 62.740 146.825 ;
        RECT 62.915 145.750 63.170 146.655 ;
        RECT 63.340 146.065 63.670 146.825 ;
        RECT 63.885 145.895 64.055 146.655 ;
        RECT 61.035 145.265 61.365 145.515 ;
        RECT 60.615 144.445 60.945 145.075 ;
        RECT 61.115 144.275 61.345 145.095 ;
        RECT 61.555 144.275 61.845 145.000 ;
        RECT 62.480 144.275 62.740 145.115 ;
        RECT 62.915 145.020 63.085 145.750 ;
        RECT 63.340 145.725 64.055 145.895 ;
        RECT 64.405 145.895 64.575 146.655 ;
        RECT 64.790 146.065 65.120 146.825 ;
        RECT 64.405 145.725 65.120 145.895 ;
        RECT 65.290 145.750 65.545 146.655 ;
        RECT 63.340 145.515 63.510 145.725 ;
        RECT 63.255 145.185 63.510 145.515 ;
        RECT 62.915 144.445 63.170 145.020 ;
        RECT 63.340 144.995 63.510 145.185 ;
        RECT 63.790 145.175 64.145 145.545 ;
        RECT 64.315 145.175 64.670 145.545 ;
        RECT 64.950 145.515 65.120 145.725 ;
        RECT 64.950 145.185 65.205 145.515 ;
        RECT 64.950 144.995 65.120 145.185 ;
        RECT 65.375 145.020 65.545 145.750 ;
        RECT 65.720 145.675 65.980 146.825 ;
        RECT 66.245 145.895 66.415 146.655 ;
        RECT 66.630 146.065 66.960 146.825 ;
        RECT 66.245 145.725 66.960 145.895 ;
        RECT 67.130 145.750 67.385 146.655 ;
        RECT 66.155 145.175 66.510 145.545 ;
        RECT 66.790 145.515 66.960 145.725 ;
        RECT 66.790 145.185 67.045 145.515 ;
        RECT 63.340 144.825 64.055 144.995 ;
        RECT 63.340 144.275 63.670 144.655 ;
        RECT 63.885 144.445 64.055 144.825 ;
        RECT 64.405 144.825 65.120 144.995 ;
        RECT 64.405 144.445 64.575 144.825 ;
        RECT 64.790 144.275 65.120 144.655 ;
        RECT 65.290 144.445 65.545 145.020 ;
        RECT 65.720 144.275 65.980 145.115 ;
        RECT 66.790 144.995 66.960 145.185 ;
        RECT 67.215 145.020 67.385 145.750 ;
        RECT 67.560 145.675 67.820 146.825 ;
        RECT 68.915 145.735 72.425 146.825 ;
        RECT 68.915 145.215 70.605 145.735 ;
        RECT 72.655 145.685 72.865 146.825 ;
        RECT 73.035 145.675 73.365 146.655 ;
        RECT 73.535 145.685 73.765 146.825 ;
        RECT 74.350 145.845 74.605 146.515 ;
        RECT 74.785 146.025 75.070 146.825 ;
        RECT 75.250 146.105 75.580 146.615 ;
        RECT 66.245 144.825 66.960 144.995 ;
        RECT 66.245 144.445 66.415 144.825 ;
        RECT 66.630 144.275 66.960 144.655 ;
        RECT 67.130 144.445 67.385 145.020 ;
        RECT 67.560 144.275 67.820 145.115 ;
        RECT 70.775 145.045 72.425 145.565 ;
        RECT 68.915 144.275 72.425 145.045 ;
        RECT 72.655 144.275 72.865 145.095 ;
        RECT 73.035 145.075 73.285 145.675 ;
        RECT 73.455 145.265 73.785 145.515 ;
        RECT 74.350 145.465 74.530 145.845 ;
        RECT 75.250 145.515 75.500 146.105 ;
        RECT 75.850 145.955 76.020 146.565 ;
        RECT 76.190 146.135 76.520 146.825 ;
        RECT 76.750 146.275 76.990 146.565 ;
        RECT 77.190 146.445 77.610 146.825 ;
        RECT 77.790 146.355 78.420 146.605 ;
        RECT 78.890 146.445 79.220 146.825 ;
        RECT 77.790 146.275 77.960 146.355 ;
        RECT 79.390 146.275 79.560 146.565 ;
        RECT 79.740 146.445 80.120 146.825 ;
        RECT 80.360 146.440 81.190 146.610 ;
        RECT 76.750 146.105 77.960 146.275 ;
        RECT 74.265 145.295 74.530 145.465 ;
        RECT 73.035 144.445 73.365 145.075 ;
        RECT 73.535 144.275 73.765 145.095 ;
        RECT 74.350 144.985 74.530 145.295 ;
        RECT 74.700 145.185 75.500 145.515 ;
        RECT 74.350 144.455 74.605 144.985 ;
        RECT 74.785 144.275 75.070 144.735 ;
        RECT 75.250 144.535 75.500 145.185 ;
        RECT 75.700 145.935 76.020 145.955 ;
        RECT 75.700 145.765 77.620 145.935 ;
        RECT 75.700 144.870 75.890 145.765 ;
        RECT 77.790 145.595 77.960 146.105 ;
        RECT 78.130 145.845 78.650 146.155 ;
        RECT 76.060 145.425 77.960 145.595 ;
        RECT 76.060 145.365 76.390 145.425 ;
        RECT 76.540 145.195 76.870 145.255 ;
        RECT 76.210 144.925 76.870 145.195 ;
        RECT 75.700 144.540 76.020 144.870 ;
        RECT 76.200 144.275 76.860 144.755 ;
        RECT 77.060 144.665 77.230 145.425 ;
        RECT 78.130 145.255 78.310 145.665 ;
        RECT 77.400 145.085 77.730 145.205 ;
        RECT 78.480 145.085 78.650 145.845 ;
        RECT 77.400 144.915 78.650 145.085 ;
        RECT 78.820 146.025 80.190 146.275 ;
        RECT 78.820 145.255 79.010 146.025 ;
        RECT 79.940 145.765 80.190 146.025 ;
        RECT 79.180 145.595 79.430 145.755 ;
        RECT 80.360 145.595 80.530 146.440 ;
        RECT 81.425 146.155 81.595 146.655 ;
        RECT 81.765 146.325 82.095 146.825 ;
        RECT 80.700 145.765 81.200 146.145 ;
        RECT 81.425 145.985 82.120 146.155 ;
        RECT 79.180 145.425 80.530 145.595 ;
        RECT 80.110 145.385 80.530 145.425 ;
        RECT 78.820 144.915 79.240 145.255 ;
        RECT 79.530 144.925 79.940 145.255 ;
        RECT 77.060 144.495 77.910 144.665 ;
        RECT 78.470 144.275 78.790 144.735 ;
        RECT 78.990 144.485 79.240 144.915 ;
        RECT 79.530 144.275 79.940 144.715 ;
        RECT 80.110 144.655 80.280 145.385 ;
        RECT 80.450 144.835 80.800 145.205 ;
        RECT 80.980 144.895 81.200 145.765 ;
        RECT 81.370 145.195 81.780 145.815 ;
        RECT 81.950 145.015 82.120 145.985 ;
        RECT 81.425 144.825 82.120 145.015 ;
        RECT 80.110 144.455 81.125 144.655 ;
        RECT 81.425 144.495 81.595 144.825 ;
        RECT 81.765 144.275 82.095 144.655 ;
        RECT 82.310 144.535 82.535 146.655 ;
        RECT 82.705 146.325 83.035 146.825 ;
        RECT 83.205 146.155 83.375 146.655 ;
        RECT 82.710 145.985 83.375 146.155 ;
        RECT 82.710 144.995 82.940 145.985 ;
        RECT 83.110 145.165 83.460 145.815 ;
        RECT 83.635 145.735 87.145 146.825 ;
        RECT 83.635 145.215 85.325 145.735 ;
        RECT 87.315 145.660 87.605 146.825 ;
        RECT 87.775 145.735 91.285 146.825 ;
        RECT 85.495 145.045 87.145 145.565 ;
        RECT 87.775 145.215 89.465 145.735 ;
        RECT 91.455 145.685 91.725 146.655 ;
        RECT 91.935 146.025 92.215 146.825 ;
        RECT 92.385 146.315 94.040 146.605 ;
        RECT 92.450 145.975 94.040 146.145 ;
        RECT 92.450 145.855 92.620 145.975 ;
        RECT 91.895 145.685 92.620 145.855 ;
        RECT 89.635 145.045 91.285 145.565 ;
        RECT 82.710 144.825 83.375 144.995 ;
        RECT 82.705 144.275 83.035 144.655 ;
        RECT 83.205 144.535 83.375 144.825 ;
        RECT 83.635 144.275 87.145 145.045 ;
        RECT 87.315 144.275 87.605 145.000 ;
        RECT 87.775 144.275 91.285 145.045 ;
        RECT 91.455 144.950 91.625 145.685 ;
        RECT 91.895 145.515 92.065 145.685 ;
        RECT 92.810 145.635 93.525 145.805 ;
        RECT 93.720 145.685 94.040 145.975 ;
        RECT 94.215 145.735 96.805 146.825 ;
        RECT 97.180 145.855 97.510 146.655 ;
        RECT 97.680 146.025 98.010 146.825 ;
        RECT 98.310 145.855 98.640 146.655 ;
        RECT 99.285 146.025 99.535 146.825 ;
        RECT 91.795 145.185 92.065 145.515 ;
        RECT 92.235 145.185 92.640 145.515 ;
        RECT 92.810 145.185 93.520 145.635 ;
        RECT 91.895 145.015 92.065 145.185 ;
        RECT 91.455 144.605 91.725 144.950 ;
        RECT 91.895 144.845 93.505 145.015 ;
        RECT 93.690 144.945 94.040 145.515 ;
        RECT 94.215 145.215 95.425 145.735 ;
        RECT 97.180 145.685 99.615 145.855 ;
        RECT 99.805 145.685 99.975 146.825 ;
        RECT 100.145 145.685 100.485 146.655 ;
        RECT 95.595 145.045 96.805 145.565 ;
        RECT 96.975 145.265 97.325 145.515 ;
        RECT 97.510 145.055 97.680 145.685 ;
        RECT 97.850 145.265 98.180 145.465 ;
        RECT 98.350 145.265 98.680 145.465 ;
        RECT 98.850 145.265 99.270 145.465 ;
        RECT 99.445 145.435 99.615 145.685 ;
        RECT 99.445 145.265 100.140 145.435 ;
        RECT 91.915 144.275 92.295 144.675 ;
        RECT 92.465 144.495 92.635 144.845 ;
        RECT 92.805 144.275 93.135 144.675 ;
        RECT 93.335 144.495 93.505 144.845 ;
        RECT 93.705 144.275 94.035 144.775 ;
        RECT 94.215 144.275 96.805 145.045 ;
        RECT 97.180 144.445 97.680 145.055 ;
        RECT 98.310 144.925 99.535 145.095 ;
        RECT 100.310 145.075 100.485 145.685 ;
        RECT 100.655 145.735 102.325 146.825 ;
        RECT 102.495 146.065 103.010 146.475 ;
        RECT 103.245 146.065 103.415 146.825 ;
        RECT 103.585 146.485 105.615 146.655 ;
        RECT 100.655 145.215 101.405 145.735 ;
        RECT 98.310 144.445 98.640 144.925 ;
        RECT 98.810 144.275 99.035 144.735 ;
        RECT 99.205 144.445 99.535 144.925 ;
        RECT 99.725 144.275 99.975 145.075 ;
        RECT 100.145 144.445 100.485 145.075 ;
        RECT 101.575 145.045 102.325 145.565 ;
        RECT 102.495 145.255 102.835 146.065 ;
        RECT 103.585 145.820 103.755 146.485 ;
        RECT 104.150 146.145 105.275 146.315 ;
        RECT 103.005 145.630 103.755 145.820 ;
        RECT 103.925 145.805 104.935 145.975 ;
        RECT 102.495 145.085 103.725 145.255 ;
        RECT 100.655 144.275 102.325 145.045 ;
        RECT 102.770 144.480 103.015 145.085 ;
        RECT 103.235 144.275 103.745 144.810 ;
        RECT 103.925 144.445 104.115 145.805 ;
        RECT 104.285 145.465 104.560 145.605 ;
        RECT 104.285 145.295 104.565 145.465 ;
        RECT 104.285 144.445 104.560 145.295 ;
        RECT 104.765 145.005 104.935 145.805 ;
        RECT 105.105 145.015 105.275 146.145 ;
        RECT 105.445 145.515 105.615 146.485 ;
        RECT 105.785 145.685 105.955 146.825 ;
        RECT 106.125 145.685 106.460 146.655 ;
        RECT 106.695 145.685 106.905 146.825 ;
        RECT 105.445 145.185 105.640 145.515 ;
        RECT 105.865 145.185 106.120 145.515 ;
        RECT 105.865 145.015 106.035 145.185 ;
        RECT 106.290 145.015 106.460 145.685 ;
        RECT 107.075 145.675 107.405 146.655 ;
        RECT 107.575 145.685 107.805 146.825 ;
        RECT 108.105 145.895 108.275 146.655 ;
        RECT 108.455 146.065 108.785 146.825 ;
        RECT 108.105 145.725 108.770 145.895 ;
        RECT 108.955 145.750 109.225 146.655 ;
        RECT 105.105 144.845 106.035 145.015 ;
        RECT 105.105 144.810 105.280 144.845 ;
        RECT 104.750 144.445 105.280 144.810 ;
        RECT 105.705 144.275 106.035 144.675 ;
        RECT 106.205 144.445 106.460 145.015 ;
        RECT 106.695 144.275 106.905 145.095 ;
        RECT 107.075 145.075 107.325 145.675 ;
        RECT 108.600 145.580 108.770 145.725 ;
        RECT 107.495 145.265 107.825 145.515 ;
        RECT 108.035 145.175 108.365 145.545 ;
        RECT 108.600 145.250 108.885 145.580 ;
        RECT 107.075 144.445 107.405 145.075 ;
        RECT 107.575 144.275 107.805 145.095 ;
        RECT 108.600 144.995 108.770 145.250 ;
        RECT 108.105 144.825 108.770 144.995 ;
        RECT 109.055 144.950 109.225 145.750 ;
        RECT 109.395 145.735 111.985 146.825 ;
        RECT 112.155 145.735 113.365 146.825 ;
        RECT 109.395 145.215 110.605 145.735 ;
        RECT 110.775 145.045 111.985 145.565 ;
        RECT 112.155 145.195 112.675 145.735 ;
        RECT 108.105 144.445 108.275 144.825 ;
        RECT 108.455 144.275 108.785 144.655 ;
        RECT 108.965 144.445 109.225 144.950 ;
        RECT 109.395 144.275 111.985 145.045 ;
        RECT 112.845 145.025 113.365 145.565 ;
        RECT 112.155 144.275 113.365 145.025 ;
        RECT 11.330 144.105 113.450 144.275 ;
        RECT 11.415 143.355 12.625 144.105 ;
        RECT 11.415 142.815 11.935 143.355 ;
        RECT 13.715 143.335 17.225 144.105 ;
        RECT 17.400 143.560 22.745 144.105 ;
        RECT 12.105 142.645 12.625 143.185 ;
        RECT 11.415 141.555 12.625 142.645 ;
        RECT 13.715 142.645 15.405 143.165 ;
        RECT 15.575 142.815 17.225 143.335 ;
        RECT 13.715 141.555 17.225 142.645 ;
        RECT 18.990 141.990 19.340 143.240 ;
        RECT 20.820 142.730 21.160 143.560 ;
        RECT 22.915 143.380 23.205 144.105 ;
        RECT 23.840 143.560 29.185 144.105 ;
        RECT 17.400 141.555 22.745 141.990 ;
        RECT 22.915 141.555 23.205 142.720 ;
        RECT 25.430 141.990 25.780 143.240 ;
        RECT 27.260 142.730 27.600 143.560 ;
        RECT 29.355 143.430 29.625 143.775 ;
        RECT 29.815 143.705 30.195 144.105 ;
        RECT 30.365 143.535 30.535 143.885 ;
        RECT 30.705 143.705 31.035 144.105 ;
        RECT 31.235 143.535 31.405 143.885 ;
        RECT 31.605 143.605 31.935 144.105 ;
        RECT 32.580 143.560 37.925 144.105 ;
        RECT 38.100 143.560 43.445 144.105 ;
        RECT 29.355 142.695 29.525 143.430 ;
        RECT 29.795 143.365 31.405 143.535 ;
        RECT 29.795 143.195 29.965 143.365 ;
        RECT 29.695 142.865 29.965 143.195 ;
        RECT 30.135 142.865 30.540 143.195 ;
        RECT 29.795 142.695 29.965 142.865 ;
        RECT 23.840 141.555 29.185 141.990 ;
        RECT 29.355 141.725 29.625 142.695 ;
        RECT 29.795 142.525 30.520 142.695 ;
        RECT 30.710 142.575 31.420 143.195 ;
        RECT 31.590 142.865 31.940 143.435 ;
        RECT 30.350 142.405 30.520 142.525 ;
        RECT 31.620 142.405 31.940 142.695 ;
        RECT 29.835 141.555 30.115 142.355 ;
        RECT 30.350 142.235 31.940 142.405 ;
        RECT 30.285 141.775 31.940 142.065 ;
        RECT 34.170 141.990 34.520 143.240 ;
        RECT 36.000 142.730 36.340 143.560 ;
        RECT 39.690 141.990 40.040 143.240 ;
        RECT 41.520 142.730 41.860 143.560 ;
        RECT 43.615 143.305 43.955 143.935 ;
        RECT 44.125 143.305 44.375 144.105 ;
        RECT 44.565 143.455 44.895 143.935 ;
        RECT 45.065 143.645 45.290 144.105 ;
        RECT 45.460 143.455 45.790 143.935 ;
        RECT 43.615 142.695 43.790 143.305 ;
        RECT 44.565 143.285 45.790 143.455 ;
        RECT 46.420 143.325 46.920 143.935 ;
        RECT 47.295 143.355 48.505 144.105 ;
        RECT 48.675 143.380 48.965 144.105 ;
        RECT 49.135 143.355 50.345 144.105 ;
        RECT 43.960 142.945 44.655 143.115 ;
        RECT 44.485 142.695 44.655 142.945 ;
        RECT 44.830 142.915 45.250 143.115 ;
        RECT 45.420 142.915 45.750 143.115 ;
        RECT 45.920 142.915 46.250 143.115 ;
        RECT 46.420 142.695 46.590 143.325 ;
        RECT 46.775 142.865 47.125 143.115 ;
        RECT 32.580 141.555 37.925 141.990 ;
        RECT 38.100 141.555 43.445 141.990 ;
        RECT 43.615 141.725 43.955 142.695 ;
        RECT 44.125 141.555 44.295 142.695 ;
        RECT 44.485 142.525 46.920 142.695 ;
        RECT 44.565 141.555 44.815 142.355 ;
        RECT 45.460 141.725 45.790 142.525 ;
        RECT 46.090 141.555 46.420 142.355 ;
        RECT 46.590 141.725 46.920 142.525 ;
        RECT 47.295 142.645 47.815 143.185 ;
        RECT 47.985 142.815 48.505 143.355 ;
        RECT 47.295 141.555 48.505 142.645 ;
        RECT 48.675 141.555 48.965 142.720 ;
        RECT 49.135 142.645 49.655 143.185 ;
        RECT 49.825 142.815 50.345 143.355 ;
        RECT 50.790 143.295 51.035 143.900 ;
        RECT 51.255 143.570 51.765 144.105 ;
        RECT 50.515 143.125 51.745 143.295 ;
        RECT 49.135 141.555 50.345 142.645 ;
        RECT 50.515 142.315 50.855 143.125 ;
        RECT 51.025 142.560 51.775 142.750 ;
        RECT 50.515 141.905 51.030 142.315 ;
        RECT 51.265 141.555 51.435 142.315 ;
        RECT 51.605 141.895 51.775 142.560 ;
        RECT 51.945 142.575 52.135 143.935 ;
        RECT 52.305 143.085 52.580 143.935 ;
        RECT 52.770 143.570 53.300 143.935 ;
        RECT 53.725 143.705 54.055 144.105 ;
        RECT 53.125 143.535 53.300 143.570 ;
        RECT 52.305 142.915 52.585 143.085 ;
        RECT 52.305 142.775 52.580 142.915 ;
        RECT 52.785 142.575 52.955 143.375 ;
        RECT 51.945 142.405 52.955 142.575 ;
        RECT 53.125 143.365 54.055 143.535 ;
        RECT 54.225 143.365 54.480 143.935 ;
        RECT 55.205 143.555 55.375 143.935 ;
        RECT 55.555 143.725 55.885 144.105 ;
        RECT 55.205 143.385 55.870 143.555 ;
        RECT 56.065 143.430 56.325 143.935 ;
        RECT 53.125 142.235 53.295 143.365 ;
        RECT 53.885 143.195 54.055 143.365 ;
        RECT 52.170 142.065 53.295 142.235 ;
        RECT 53.465 142.865 53.660 143.195 ;
        RECT 53.885 142.865 54.140 143.195 ;
        RECT 53.465 141.895 53.635 142.865 ;
        RECT 54.310 142.695 54.480 143.365 ;
        RECT 55.135 142.835 55.465 143.205 ;
        RECT 55.700 143.130 55.870 143.385 ;
        RECT 51.605 141.725 53.635 141.895 ;
        RECT 53.805 141.555 53.975 142.695 ;
        RECT 54.145 141.725 54.480 142.695 ;
        RECT 55.700 142.800 55.985 143.130 ;
        RECT 55.700 142.655 55.870 142.800 ;
        RECT 55.205 142.485 55.870 142.655 ;
        RECT 56.155 142.630 56.325 143.430 ;
        RECT 56.495 143.355 57.705 144.105 ;
        RECT 55.205 141.725 55.375 142.485 ;
        RECT 55.555 141.555 55.885 142.315 ;
        RECT 56.055 141.725 56.325 142.630 ;
        RECT 56.495 142.645 57.015 143.185 ;
        RECT 57.185 142.815 57.705 143.355 ;
        RECT 57.875 143.335 61.385 144.105 ;
        RECT 61.645 143.555 61.815 143.935 ;
        RECT 61.995 143.725 62.325 144.105 ;
        RECT 61.645 143.385 62.310 143.555 ;
        RECT 62.505 143.430 62.765 143.935 ;
        RECT 57.875 142.645 59.565 143.165 ;
        RECT 59.735 142.815 61.385 143.335 ;
        RECT 61.575 142.835 61.905 143.205 ;
        RECT 62.140 143.130 62.310 143.385 ;
        RECT 62.140 142.800 62.425 143.130 ;
        RECT 62.140 142.655 62.310 142.800 ;
        RECT 56.495 141.555 57.705 142.645 ;
        RECT 57.875 141.555 61.385 142.645 ;
        RECT 61.645 142.485 62.310 142.655 ;
        RECT 62.595 142.630 62.765 143.430 ;
        RECT 63.855 143.335 67.365 144.105 ;
        RECT 61.645 141.725 61.815 142.485 ;
        RECT 61.995 141.555 62.325 142.315 ;
        RECT 62.495 141.725 62.765 142.630 ;
        RECT 63.855 142.645 65.545 143.165 ;
        RECT 65.715 142.815 67.365 143.335 ;
        RECT 67.535 143.430 67.805 143.775 ;
        RECT 67.995 143.705 68.375 144.105 ;
        RECT 68.545 143.535 68.715 143.885 ;
        RECT 68.885 143.705 69.215 144.105 ;
        RECT 69.415 143.535 69.585 143.885 ;
        RECT 69.785 143.605 70.115 144.105 ;
        RECT 67.535 142.695 67.705 143.430 ;
        RECT 67.975 143.365 69.585 143.535 ;
        RECT 67.975 143.195 68.145 143.365 ;
        RECT 67.875 142.865 68.145 143.195 ;
        RECT 68.315 142.865 68.720 143.195 ;
        RECT 67.975 142.695 68.145 142.865 ;
        RECT 63.855 141.555 67.365 142.645 ;
        RECT 67.535 141.725 67.805 142.695 ;
        RECT 67.975 142.525 68.700 142.695 ;
        RECT 68.890 142.575 69.600 143.195 ;
        RECT 69.770 142.865 70.120 143.435 ;
        RECT 70.295 143.305 70.635 143.935 ;
        RECT 70.805 143.305 71.055 144.105 ;
        RECT 71.245 143.455 71.575 143.935 ;
        RECT 71.745 143.645 71.970 144.105 ;
        RECT 72.140 143.455 72.470 143.935 ;
        RECT 70.295 143.255 70.525 143.305 ;
        RECT 71.245 143.285 72.470 143.455 ;
        RECT 73.100 143.325 73.600 143.935 ;
        RECT 74.435 143.380 74.725 144.105 ;
        RECT 70.295 142.695 70.470 143.255 ;
        RECT 70.640 142.945 71.335 143.115 ;
        RECT 71.165 142.695 71.335 142.945 ;
        RECT 71.510 142.915 71.930 143.115 ;
        RECT 72.100 142.915 72.430 143.115 ;
        RECT 72.600 142.915 72.930 143.115 ;
        RECT 73.100 142.695 73.270 143.325 ;
        RECT 75.630 143.295 75.875 143.900 ;
        RECT 76.095 143.570 76.605 144.105 ;
        RECT 75.355 143.125 76.585 143.295 ;
        RECT 73.455 142.865 73.805 143.115 ;
        RECT 68.530 142.405 68.700 142.525 ;
        RECT 69.800 142.405 70.120 142.695 ;
        RECT 68.015 141.555 68.295 142.355 ;
        RECT 68.530 142.235 70.120 142.405 ;
        RECT 68.465 141.775 70.120 142.065 ;
        RECT 70.295 141.725 70.635 142.695 ;
        RECT 70.805 141.555 70.975 142.695 ;
        RECT 71.165 142.525 73.600 142.695 ;
        RECT 71.245 141.555 71.495 142.355 ;
        RECT 72.140 141.725 72.470 142.525 ;
        RECT 72.770 141.555 73.100 142.355 ;
        RECT 73.270 141.725 73.600 142.525 ;
        RECT 74.435 141.555 74.725 142.720 ;
        RECT 75.355 142.315 75.695 143.125 ;
        RECT 75.865 142.560 76.615 142.750 ;
        RECT 75.355 141.905 75.870 142.315 ;
        RECT 76.105 141.555 76.275 142.315 ;
        RECT 76.445 141.895 76.615 142.560 ;
        RECT 76.785 142.575 76.975 143.935 ;
        RECT 77.145 143.085 77.420 143.935 ;
        RECT 77.610 143.570 78.140 143.935 ;
        RECT 78.565 143.705 78.895 144.105 ;
        RECT 77.965 143.535 78.140 143.570 ;
        RECT 77.145 142.915 77.425 143.085 ;
        RECT 77.145 142.775 77.420 142.915 ;
        RECT 77.625 142.575 77.795 143.375 ;
        RECT 76.785 142.405 77.795 142.575 ;
        RECT 77.965 143.365 78.895 143.535 ;
        RECT 79.065 143.365 79.320 143.935 ;
        RECT 79.585 143.555 79.755 143.935 ;
        RECT 79.935 143.725 80.265 144.105 ;
        RECT 79.585 143.385 80.250 143.555 ;
        RECT 80.445 143.430 80.705 143.935 ;
        RECT 77.965 142.235 78.135 143.365 ;
        RECT 78.725 143.195 78.895 143.365 ;
        RECT 77.010 142.065 78.135 142.235 ;
        RECT 78.305 142.865 78.500 143.195 ;
        RECT 78.725 142.865 78.980 143.195 ;
        RECT 78.305 141.895 78.475 142.865 ;
        RECT 79.150 142.695 79.320 143.365 ;
        RECT 79.515 142.835 79.845 143.205 ;
        RECT 80.080 143.130 80.250 143.385 ;
        RECT 76.445 141.725 78.475 141.895 ;
        RECT 78.645 141.555 78.815 142.695 ;
        RECT 78.985 141.725 79.320 142.695 ;
        RECT 80.080 142.800 80.365 143.130 ;
        RECT 80.080 142.655 80.250 142.800 ;
        RECT 79.585 142.485 80.250 142.655 ;
        RECT 80.535 142.630 80.705 143.430 ;
        RECT 81.335 143.335 84.845 144.105 ;
        RECT 79.585 141.725 79.755 142.485 ;
        RECT 79.935 141.555 80.265 142.315 ;
        RECT 80.435 141.725 80.705 142.630 ;
        RECT 81.335 142.645 83.025 143.165 ;
        RECT 83.195 142.815 84.845 143.335 ;
        RECT 85.015 143.430 85.285 143.775 ;
        RECT 85.475 143.705 85.855 144.105 ;
        RECT 86.025 143.535 86.195 143.885 ;
        RECT 86.365 143.705 86.695 144.105 ;
        RECT 86.895 143.535 87.065 143.885 ;
        RECT 87.265 143.605 87.595 144.105 ;
        RECT 85.015 142.695 85.185 143.430 ;
        RECT 85.455 143.365 87.065 143.535 ;
        RECT 85.455 143.195 85.625 143.365 ;
        RECT 85.355 142.865 85.625 143.195 ;
        RECT 85.795 142.865 86.200 143.195 ;
        RECT 85.455 142.695 85.625 142.865 ;
        RECT 86.370 142.745 87.080 143.195 ;
        RECT 87.250 142.865 87.600 143.435 ;
        RECT 87.775 143.305 88.115 143.935 ;
        RECT 88.285 143.305 88.535 144.105 ;
        RECT 88.725 143.455 89.055 143.935 ;
        RECT 89.225 143.645 89.450 144.105 ;
        RECT 89.620 143.455 89.950 143.935 ;
        RECT 87.775 143.255 88.005 143.305 ;
        RECT 88.725 143.285 89.950 143.455 ;
        RECT 90.580 143.325 91.080 143.935 ;
        RECT 91.915 143.335 93.585 144.105 ;
        RECT 81.335 141.555 84.845 142.645 ;
        RECT 85.015 141.725 85.285 142.695 ;
        RECT 85.455 142.525 86.180 142.695 ;
        RECT 86.370 142.575 87.085 142.745 ;
        RECT 87.775 142.695 87.950 143.255 ;
        RECT 88.120 142.945 88.815 143.115 ;
        RECT 88.645 142.695 88.815 142.945 ;
        RECT 88.990 142.915 89.410 143.115 ;
        RECT 89.580 142.915 89.910 143.115 ;
        RECT 90.080 142.915 90.410 143.115 ;
        RECT 90.580 142.695 90.750 143.325 ;
        RECT 90.935 142.865 91.285 143.115 ;
        RECT 86.010 142.405 86.180 142.525 ;
        RECT 87.280 142.405 87.600 142.695 ;
        RECT 85.495 141.555 85.775 142.355 ;
        RECT 86.010 142.235 87.600 142.405 ;
        RECT 85.945 141.775 87.600 142.065 ;
        RECT 87.775 141.725 88.115 142.695 ;
        RECT 88.285 141.555 88.455 142.695 ;
        RECT 88.645 142.525 91.080 142.695 ;
        RECT 88.725 141.555 88.975 142.355 ;
        RECT 89.620 141.725 89.950 142.525 ;
        RECT 90.250 141.555 90.580 142.355 ;
        RECT 90.750 141.725 91.080 142.525 ;
        RECT 91.915 142.645 92.665 143.165 ;
        RECT 92.835 142.815 93.585 143.335 ;
        RECT 93.755 143.305 94.095 143.935 ;
        RECT 94.265 143.305 94.515 144.105 ;
        RECT 94.705 143.455 95.035 143.935 ;
        RECT 95.205 143.645 95.430 144.105 ;
        RECT 95.600 143.455 95.930 143.935 ;
        RECT 93.755 142.695 93.930 143.305 ;
        RECT 94.705 143.285 95.930 143.455 ;
        RECT 96.560 143.325 97.060 143.935 ;
        RECT 97.435 143.430 97.705 143.775 ;
        RECT 97.895 143.705 98.275 144.105 ;
        RECT 98.445 143.535 98.615 143.885 ;
        RECT 98.785 143.705 99.115 144.105 ;
        RECT 99.315 143.535 99.485 143.885 ;
        RECT 99.685 143.605 100.015 144.105 ;
        RECT 94.100 142.945 94.795 143.115 ;
        RECT 94.625 142.695 94.795 142.945 ;
        RECT 94.970 142.915 95.390 143.115 ;
        RECT 95.560 142.915 95.890 143.115 ;
        RECT 96.060 142.915 96.390 143.115 ;
        RECT 96.560 142.695 96.730 143.325 ;
        RECT 96.915 142.865 97.265 143.115 ;
        RECT 97.435 142.695 97.605 143.430 ;
        RECT 97.875 143.365 99.485 143.535 ;
        RECT 97.875 143.195 98.045 143.365 ;
        RECT 97.775 142.865 98.045 143.195 ;
        RECT 98.215 142.865 98.620 143.195 ;
        RECT 97.875 142.695 98.045 142.865 ;
        RECT 98.790 142.745 99.500 143.195 ;
        RECT 99.670 142.865 100.020 143.435 ;
        RECT 100.195 143.380 100.485 144.105 ;
        RECT 101.155 143.285 101.385 144.105 ;
        RECT 101.555 143.305 101.885 143.935 ;
        RECT 101.135 142.865 101.465 143.115 ;
        RECT 91.915 141.555 93.585 142.645 ;
        RECT 93.755 141.725 94.095 142.695 ;
        RECT 94.265 141.555 94.435 142.695 ;
        RECT 94.625 142.525 97.060 142.695 ;
        RECT 94.705 141.555 94.955 142.355 ;
        RECT 95.600 141.725 95.930 142.525 ;
        RECT 96.230 141.555 96.560 142.355 ;
        RECT 96.730 141.725 97.060 142.525 ;
        RECT 97.435 141.725 97.705 142.695 ;
        RECT 97.875 142.525 98.600 142.695 ;
        RECT 98.790 142.575 99.505 142.745 ;
        RECT 98.430 142.405 98.600 142.525 ;
        RECT 99.700 142.405 100.020 142.695 ;
        RECT 97.915 141.555 98.195 142.355 ;
        RECT 98.430 142.235 100.020 142.405 ;
        RECT 98.365 141.775 100.020 142.065 ;
        RECT 100.195 141.555 100.485 142.720 ;
        RECT 101.635 142.705 101.885 143.305 ;
        RECT 102.055 143.285 102.265 144.105 ;
        RECT 102.870 143.425 103.125 143.925 ;
        RECT 103.305 143.645 103.590 144.105 ;
        RECT 102.785 143.395 103.125 143.425 ;
        RECT 102.785 143.255 103.050 143.395 ;
        RECT 101.155 141.555 101.385 142.695 ;
        RECT 101.555 141.725 101.885 142.705 ;
        RECT 102.055 141.555 102.265 142.695 ;
        RECT 102.870 142.535 103.050 143.255 ;
        RECT 103.770 143.195 104.020 143.845 ;
        RECT 103.220 142.865 104.020 143.195 ;
        RECT 102.870 141.865 103.125 142.535 ;
        RECT 103.305 141.555 103.590 142.355 ;
        RECT 103.770 142.275 104.020 142.865 ;
        RECT 104.220 143.510 104.540 143.840 ;
        RECT 104.720 143.625 105.380 144.105 ;
        RECT 105.580 143.715 106.430 143.885 ;
        RECT 104.220 142.615 104.410 143.510 ;
        RECT 104.730 143.185 105.390 143.455 ;
        RECT 105.060 143.125 105.390 143.185 ;
        RECT 104.580 142.955 104.910 143.015 ;
        RECT 105.580 142.955 105.750 143.715 ;
        RECT 106.990 143.645 107.310 144.105 ;
        RECT 107.510 143.465 107.760 143.895 ;
        RECT 108.050 143.665 108.460 144.105 ;
        RECT 108.630 143.725 109.645 143.925 ;
        RECT 105.920 143.295 107.170 143.465 ;
        RECT 105.920 143.175 106.250 143.295 ;
        RECT 104.580 142.785 106.480 142.955 ;
        RECT 104.220 142.445 106.140 142.615 ;
        RECT 104.220 142.425 104.540 142.445 ;
        RECT 103.770 141.765 104.100 142.275 ;
        RECT 104.370 141.815 104.540 142.425 ;
        RECT 106.310 142.275 106.480 142.785 ;
        RECT 106.650 142.715 106.830 143.125 ;
        RECT 107.000 142.535 107.170 143.295 ;
        RECT 104.710 141.555 105.040 142.245 ;
        RECT 105.270 142.105 106.480 142.275 ;
        RECT 106.650 142.225 107.170 142.535 ;
        RECT 107.340 143.125 107.760 143.465 ;
        RECT 108.050 143.125 108.460 143.455 ;
        RECT 107.340 142.355 107.530 143.125 ;
        RECT 108.630 142.995 108.800 143.725 ;
        RECT 109.945 143.555 110.115 143.885 ;
        RECT 110.285 143.725 110.615 144.105 ;
        RECT 108.970 143.175 109.320 143.545 ;
        RECT 108.630 142.955 109.050 142.995 ;
        RECT 107.700 142.785 109.050 142.955 ;
        RECT 107.700 142.625 107.950 142.785 ;
        RECT 108.460 142.355 108.710 142.615 ;
        RECT 107.340 142.105 108.710 142.355 ;
        RECT 105.270 141.815 105.510 142.105 ;
        RECT 106.310 142.025 106.480 142.105 ;
        RECT 105.710 141.555 106.130 141.935 ;
        RECT 106.310 141.775 106.940 142.025 ;
        RECT 107.410 141.555 107.740 141.935 ;
        RECT 107.910 141.815 108.080 142.105 ;
        RECT 108.880 141.940 109.050 142.785 ;
        RECT 109.500 142.615 109.720 143.485 ;
        RECT 109.945 143.365 110.640 143.555 ;
        RECT 109.220 142.235 109.720 142.615 ;
        RECT 109.890 142.565 110.300 143.185 ;
        RECT 110.470 142.395 110.640 143.365 ;
        RECT 109.945 142.225 110.640 142.395 ;
        RECT 108.260 141.555 108.640 141.935 ;
        RECT 108.880 141.770 109.710 141.940 ;
        RECT 109.945 141.725 110.115 142.225 ;
        RECT 110.285 141.555 110.615 142.055 ;
        RECT 110.830 141.725 111.055 143.845 ;
        RECT 111.225 143.725 111.555 144.105 ;
        RECT 111.725 143.555 111.895 143.845 ;
        RECT 111.230 143.385 111.895 143.555 ;
        RECT 111.230 142.395 111.460 143.385 ;
        RECT 112.155 143.355 113.365 144.105 ;
        RECT 111.630 142.565 111.980 143.215 ;
        RECT 112.155 142.645 112.675 143.185 ;
        RECT 112.845 142.815 113.365 143.355 ;
        RECT 111.230 142.225 111.895 142.395 ;
        RECT 111.225 141.555 111.555 142.055 ;
        RECT 111.725 141.725 111.895 142.225 ;
        RECT 112.155 141.555 113.365 142.645 ;
        RECT 11.330 141.385 113.450 141.555 ;
        RECT 11.415 140.295 12.625 141.385 ;
        RECT 11.415 139.585 11.935 140.125 ;
        RECT 12.105 139.755 12.625 140.295 ;
        RECT 13.255 140.295 16.765 141.385 ;
        RECT 13.255 139.775 14.945 140.295 ;
        RECT 16.995 140.245 17.205 141.385 ;
        RECT 17.375 140.235 17.705 141.215 ;
        RECT 17.875 140.245 18.105 141.385 ;
        RECT 19.240 140.245 19.575 141.215 ;
        RECT 19.745 140.245 19.915 141.385 ;
        RECT 20.085 141.045 22.115 141.215 ;
        RECT 15.115 139.605 16.765 140.125 ;
        RECT 11.415 138.835 12.625 139.585 ;
        RECT 13.255 138.835 16.765 139.605 ;
        RECT 16.995 138.835 17.205 139.655 ;
        RECT 17.375 139.635 17.625 140.235 ;
        RECT 17.795 139.825 18.125 140.075 ;
        RECT 17.375 139.005 17.705 139.635 ;
        RECT 17.875 138.835 18.105 139.655 ;
        RECT 19.240 139.575 19.410 140.245 ;
        RECT 20.085 140.075 20.255 141.045 ;
        RECT 19.580 139.745 19.835 140.075 ;
        RECT 20.060 139.745 20.255 140.075 ;
        RECT 20.425 140.705 21.550 140.875 ;
        RECT 19.665 139.575 19.835 139.745 ;
        RECT 20.425 139.575 20.595 140.705 ;
        RECT 19.240 139.005 19.495 139.575 ;
        RECT 19.665 139.405 20.595 139.575 ;
        RECT 20.765 140.365 21.775 140.535 ;
        RECT 20.765 139.565 20.935 140.365 ;
        RECT 21.140 140.025 21.415 140.165 ;
        RECT 21.135 139.855 21.415 140.025 ;
        RECT 20.420 139.370 20.595 139.405 ;
        RECT 19.665 138.835 19.995 139.235 ;
        RECT 20.420 139.005 20.950 139.370 ;
        RECT 21.140 139.005 21.415 139.855 ;
        RECT 21.585 139.005 21.775 140.365 ;
        RECT 21.945 140.380 22.115 141.045 ;
        RECT 22.285 140.625 22.455 141.385 ;
        RECT 22.690 140.625 23.205 141.035 ;
        RECT 21.945 140.190 22.695 140.380 ;
        RECT 22.865 139.815 23.205 140.625 ;
        RECT 24.335 140.245 24.565 141.385 ;
        RECT 24.735 140.235 25.065 141.215 ;
        RECT 25.235 140.245 25.445 141.385 ;
        RECT 26.135 140.665 26.595 141.215 ;
        RECT 26.785 140.665 27.115 141.385 ;
        RECT 24.315 139.825 24.645 140.075 ;
        RECT 21.975 139.645 23.205 139.815 ;
        RECT 21.955 138.835 22.465 139.370 ;
        RECT 22.685 139.040 22.930 139.645 ;
        RECT 24.335 138.835 24.565 139.655 ;
        RECT 24.815 139.635 25.065 140.235 ;
        RECT 24.735 139.005 25.065 139.635 ;
        RECT 25.235 138.835 25.445 139.655 ;
        RECT 26.135 139.295 26.385 140.665 ;
        RECT 27.315 140.495 27.615 141.045 ;
        RECT 27.785 140.715 28.065 141.385 ;
        RECT 28.635 140.715 28.915 141.385 ;
        RECT 26.675 140.325 27.615 140.495 ;
        RECT 29.085 140.495 29.385 141.045 ;
        RECT 29.585 140.665 29.915 141.385 ;
        RECT 30.105 140.665 30.565 141.215 ;
        RECT 26.675 140.075 26.845 140.325 ;
        RECT 27.985 140.075 28.250 140.435 ;
        RECT 26.555 139.745 26.845 140.075 ;
        RECT 27.015 139.825 27.355 140.075 ;
        RECT 27.575 139.825 28.250 140.075 ;
        RECT 28.450 140.075 28.715 140.435 ;
        RECT 29.085 140.325 30.025 140.495 ;
        RECT 29.855 140.075 30.025 140.325 ;
        RECT 28.450 139.825 29.125 140.075 ;
        RECT 29.345 139.825 29.685 140.075 ;
        RECT 26.675 139.655 26.845 139.745 ;
        RECT 29.855 139.745 30.145 140.075 ;
        RECT 29.855 139.655 30.025 139.745 ;
        RECT 26.675 139.465 28.065 139.655 ;
        RECT 26.135 139.005 26.695 139.295 ;
        RECT 26.865 138.835 27.115 139.295 ;
        RECT 27.735 139.105 28.065 139.465 ;
        RECT 28.635 139.465 30.025 139.655 ;
        RECT 28.635 139.105 28.965 139.465 ;
        RECT 30.315 139.295 30.565 140.665 ;
        RECT 30.735 140.295 31.945 141.385 ;
        RECT 32.115 140.295 35.625 141.385 ;
        RECT 30.735 139.755 31.255 140.295 ;
        RECT 31.425 139.585 31.945 140.125 ;
        RECT 32.115 139.775 33.805 140.295 ;
        RECT 35.795 140.220 36.085 141.385 ;
        RECT 36.715 140.295 38.385 141.385 ;
        RECT 38.560 140.875 40.215 141.165 ;
        RECT 38.560 140.535 40.150 140.705 ;
        RECT 40.385 140.585 40.665 141.385 ;
        RECT 33.975 139.605 35.625 140.125 ;
        RECT 36.715 139.775 37.465 140.295 ;
        RECT 38.560 140.245 38.880 140.535 ;
        RECT 39.980 140.415 40.150 140.535 ;
        RECT 37.635 139.605 38.385 140.125 ;
        RECT 29.585 138.835 29.835 139.295 ;
        RECT 30.005 139.005 30.565 139.295 ;
        RECT 30.735 138.835 31.945 139.585 ;
        RECT 32.115 138.835 35.625 139.605 ;
        RECT 35.795 138.835 36.085 139.560 ;
        RECT 36.715 138.835 38.385 139.605 ;
        RECT 38.560 139.505 38.910 140.075 ;
        RECT 39.080 139.745 39.790 140.365 ;
        RECT 39.980 140.245 40.705 140.415 ;
        RECT 40.875 140.245 41.145 141.215 ;
        RECT 41.320 140.875 42.975 141.165 ;
        RECT 41.320 140.535 42.910 140.705 ;
        RECT 43.145 140.585 43.425 141.385 ;
        RECT 41.320 140.245 41.640 140.535 ;
        RECT 42.740 140.415 42.910 140.535 ;
        RECT 40.535 140.075 40.705 140.245 ;
        RECT 39.960 139.745 40.365 140.075 ;
        RECT 40.535 139.745 40.805 140.075 ;
        RECT 40.535 139.575 40.705 139.745 ;
        RECT 39.095 139.405 40.705 139.575 ;
        RECT 40.975 139.510 41.145 140.245 ;
        RECT 38.565 138.835 38.895 139.335 ;
        RECT 39.095 139.055 39.265 139.405 ;
        RECT 39.465 138.835 39.795 139.235 ;
        RECT 39.965 139.055 40.135 139.405 ;
        RECT 40.305 138.835 40.685 139.235 ;
        RECT 40.875 139.165 41.145 139.510 ;
        RECT 41.320 139.505 41.670 140.075 ;
        RECT 41.840 139.745 42.550 140.365 ;
        RECT 42.740 140.245 43.465 140.415 ;
        RECT 43.635 140.245 43.905 141.215 ;
        RECT 43.295 140.075 43.465 140.245 ;
        RECT 42.720 139.745 43.125 140.075 ;
        RECT 43.295 139.745 43.565 140.075 ;
        RECT 43.295 139.575 43.465 139.745 ;
        RECT 41.855 139.405 43.465 139.575 ;
        RECT 43.735 139.510 43.905 140.245 ;
        RECT 44.075 140.295 45.285 141.385 ;
        RECT 44.075 139.755 44.595 140.295 ;
        RECT 45.455 140.245 45.795 141.215 ;
        RECT 45.965 140.245 46.135 141.385 ;
        RECT 46.405 140.585 46.655 141.385 ;
        RECT 47.300 140.415 47.630 141.215 ;
        RECT 47.930 140.585 48.260 141.385 ;
        RECT 48.430 140.415 48.760 141.215 ;
        RECT 46.325 140.245 48.760 140.415 ;
        RECT 49.510 140.405 49.765 141.075 ;
        RECT 49.945 140.585 50.230 141.385 ;
        RECT 50.410 140.665 50.740 141.175 ;
        RECT 44.765 139.585 45.285 140.125 ;
        RECT 41.325 138.835 41.655 139.335 ;
        RECT 41.855 139.055 42.025 139.405 ;
        RECT 42.225 138.835 42.555 139.235 ;
        RECT 42.725 139.055 42.895 139.405 ;
        RECT 43.065 138.835 43.445 139.235 ;
        RECT 43.635 139.165 43.905 139.510 ;
        RECT 44.075 138.835 45.285 139.585 ;
        RECT 45.455 139.685 45.630 140.245 ;
        RECT 46.325 139.995 46.495 140.245 ;
        RECT 45.800 139.825 46.495 139.995 ;
        RECT 46.670 139.825 47.090 140.025 ;
        RECT 47.260 139.825 47.590 140.025 ;
        RECT 47.760 139.825 48.090 140.025 ;
        RECT 45.455 139.635 45.685 139.685 ;
        RECT 45.455 139.005 45.795 139.635 ;
        RECT 45.965 138.835 46.215 139.635 ;
        RECT 46.405 139.485 47.630 139.655 ;
        RECT 46.405 139.005 46.735 139.485 ;
        RECT 46.905 138.835 47.130 139.295 ;
        RECT 47.300 139.005 47.630 139.485 ;
        RECT 48.260 139.615 48.430 140.245 ;
        RECT 48.615 139.825 48.965 140.075 ;
        RECT 48.260 139.005 48.760 139.615 ;
        RECT 49.510 139.545 49.690 140.405 ;
        RECT 50.410 140.075 50.660 140.665 ;
        RECT 51.010 140.515 51.180 141.125 ;
        RECT 51.350 140.695 51.680 141.385 ;
        RECT 51.910 140.835 52.150 141.125 ;
        RECT 52.350 141.005 52.770 141.385 ;
        RECT 52.950 140.915 53.580 141.165 ;
        RECT 54.050 141.005 54.380 141.385 ;
        RECT 52.950 140.835 53.120 140.915 ;
        RECT 54.550 140.835 54.720 141.125 ;
        RECT 54.900 141.005 55.280 141.385 ;
        RECT 55.520 141.000 56.350 141.170 ;
        RECT 51.910 140.665 53.120 140.835 ;
        RECT 49.860 139.745 50.660 140.075 ;
        RECT 49.510 139.345 49.765 139.545 ;
        RECT 49.425 139.175 49.765 139.345 ;
        RECT 49.510 139.015 49.765 139.175 ;
        RECT 49.945 138.835 50.230 139.295 ;
        RECT 50.410 139.095 50.660 139.745 ;
        RECT 50.860 140.495 51.180 140.515 ;
        RECT 50.860 140.325 52.780 140.495 ;
        RECT 50.860 139.430 51.050 140.325 ;
        RECT 52.950 140.155 53.120 140.665 ;
        RECT 53.290 140.405 53.810 140.715 ;
        RECT 51.220 139.985 53.120 140.155 ;
        RECT 51.220 139.925 51.550 139.985 ;
        RECT 51.700 139.755 52.030 139.815 ;
        RECT 51.370 139.485 52.030 139.755 ;
        RECT 50.860 139.100 51.180 139.430 ;
        RECT 51.360 138.835 52.020 139.315 ;
        RECT 52.220 139.225 52.390 139.985 ;
        RECT 53.290 139.815 53.470 140.225 ;
        RECT 52.560 139.645 52.890 139.765 ;
        RECT 53.640 139.645 53.810 140.405 ;
        RECT 52.560 139.475 53.810 139.645 ;
        RECT 53.980 140.585 55.350 140.835 ;
        RECT 53.980 139.815 54.170 140.585 ;
        RECT 55.100 140.325 55.350 140.585 ;
        RECT 54.340 140.155 54.590 140.315 ;
        RECT 55.520 140.155 55.690 141.000 ;
        RECT 56.585 140.715 56.755 141.215 ;
        RECT 56.925 140.885 57.255 141.385 ;
        RECT 55.860 140.325 56.360 140.705 ;
        RECT 56.585 140.545 57.280 140.715 ;
        RECT 54.340 139.985 55.690 140.155 ;
        RECT 55.270 139.945 55.690 139.985 ;
        RECT 53.980 139.475 54.400 139.815 ;
        RECT 54.690 139.485 55.100 139.815 ;
        RECT 52.220 139.055 53.070 139.225 ;
        RECT 53.630 138.835 53.950 139.295 ;
        RECT 54.150 139.045 54.400 139.475 ;
        RECT 54.690 138.835 55.100 139.275 ;
        RECT 55.270 139.215 55.440 139.945 ;
        RECT 55.610 139.395 55.960 139.765 ;
        RECT 56.140 139.455 56.360 140.325 ;
        RECT 56.530 139.755 56.940 140.375 ;
        RECT 57.110 139.575 57.280 140.545 ;
        RECT 56.585 139.385 57.280 139.575 ;
        RECT 55.270 139.015 56.285 139.215 ;
        RECT 56.585 139.055 56.755 139.385 ;
        RECT 56.925 138.835 57.255 139.215 ;
        RECT 57.470 139.095 57.695 141.215 ;
        RECT 57.865 140.885 58.195 141.385 ;
        RECT 58.365 140.715 58.535 141.215 ;
        RECT 57.870 140.545 58.535 140.715 ;
        RECT 57.870 139.555 58.100 140.545 ;
        RECT 58.270 139.725 58.620 140.375 ;
        RECT 58.795 140.295 61.385 141.385 ;
        RECT 58.795 139.775 60.005 140.295 ;
        RECT 61.555 140.220 61.845 141.385 ;
        RECT 62.015 140.295 63.685 141.385 ;
        RECT 63.860 140.950 69.205 141.385 ;
        RECT 60.175 139.605 61.385 140.125 ;
        RECT 62.015 139.775 62.765 140.295 ;
        RECT 62.935 139.605 63.685 140.125 ;
        RECT 65.450 139.700 65.800 140.950 ;
        RECT 69.375 140.245 69.715 141.215 ;
        RECT 69.885 140.245 70.055 141.385 ;
        RECT 70.325 140.585 70.575 141.385 ;
        RECT 71.220 140.415 71.550 141.215 ;
        RECT 71.850 140.585 72.180 141.385 ;
        RECT 72.350 140.415 72.680 141.215 ;
        RECT 70.245 140.245 72.680 140.415 ;
        RECT 73.055 140.295 74.725 141.385 ;
        RECT 74.895 140.625 75.410 141.035 ;
        RECT 75.645 140.625 75.815 141.385 ;
        RECT 75.985 141.045 78.015 141.215 ;
        RECT 57.870 139.385 58.535 139.555 ;
        RECT 57.865 138.835 58.195 139.215 ;
        RECT 58.365 139.095 58.535 139.385 ;
        RECT 58.795 138.835 61.385 139.605 ;
        RECT 61.555 138.835 61.845 139.560 ;
        RECT 62.015 138.835 63.685 139.605 ;
        RECT 67.280 139.380 67.620 140.210 ;
        RECT 69.375 139.635 69.550 140.245 ;
        RECT 70.245 139.995 70.415 140.245 ;
        RECT 69.720 139.825 70.415 139.995 ;
        RECT 70.590 139.825 71.010 140.025 ;
        RECT 71.180 139.825 71.510 140.025 ;
        RECT 71.680 139.825 72.010 140.025 ;
        RECT 63.860 138.835 69.205 139.380 ;
        RECT 69.375 139.005 69.715 139.635 ;
        RECT 69.885 138.835 70.135 139.635 ;
        RECT 70.325 139.485 71.550 139.655 ;
        RECT 70.325 139.005 70.655 139.485 ;
        RECT 70.825 138.835 71.050 139.295 ;
        RECT 71.220 139.005 71.550 139.485 ;
        RECT 72.180 139.615 72.350 140.245 ;
        RECT 72.535 139.825 72.885 140.075 ;
        RECT 73.055 139.775 73.805 140.295 ;
        RECT 72.180 139.005 72.680 139.615 ;
        RECT 73.975 139.605 74.725 140.125 ;
        RECT 74.895 139.815 75.235 140.625 ;
        RECT 75.985 140.380 76.155 141.045 ;
        RECT 76.550 140.705 77.675 140.875 ;
        RECT 75.405 140.190 76.155 140.380 ;
        RECT 76.325 140.365 77.335 140.535 ;
        RECT 74.895 139.645 76.125 139.815 ;
        RECT 73.055 138.835 74.725 139.605 ;
        RECT 75.170 139.040 75.415 139.645 ;
        RECT 75.635 138.835 76.145 139.370 ;
        RECT 76.325 139.005 76.515 140.365 ;
        RECT 76.685 139.345 76.960 140.165 ;
        RECT 77.165 139.565 77.335 140.365 ;
        RECT 77.505 139.575 77.675 140.705 ;
        RECT 77.845 140.075 78.015 141.045 ;
        RECT 78.185 140.245 78.355 141.385 ;
        RECT 78.525 140.245 78.860 141.215 ;
        RECT 79.585 140.455 79.755 141.215 ;
        RECT 79.935 140.625 80.265 141.385 ;
        RECT 79.585 140.285 80.250 140.455 ;
        RECT 80.435 140.310 80.705 141.215 ;
        RECT 77.845 139.745 78.040 140.075 ;
        RECT 78.265 139.745 78.520 140.075 ;
        RECT 78.265 139.575 78.435 139.745 ;
        RECT 78.690 139.575 78.860 140.245 ;
        RECT 80.080 140.140 80.250 140.285 ;
        RECT 79.515 139.735 79.845 140.105 ;
        RECT 80.080 139.810 80.365 140.140 ;
        RECT 77.505 139.405 78.435 139.575 ;
        RECT 77.505 139.370 77.680 139.405 ;
        RECT 76.685 139.175 76.965 139.345 ;
        RECT 76.685 139.005 76.960 139.175 ;
        RECT 77.150 139.005 77.680 139.370 ;
        RECT 78.105 138.835 78.435 139.235 ;
        RECT 78.605 139.005 78.860 139.575 ;
        RECT 80.080 139.555 80.250 139.810 ;
        RECT 79.585 139.385 80.250 139.555 ;
        RECT 80.535 139.510 80.705 140.310 ;
        RECT 80.965 140.455 81.135 141.215 ;
        RECT 81.315 140.625 81.645 141.385 ;
        RECT 80.965 140.285 81.630 140.455 ;
        RECT 81.815 140.310 82.085 141.215 ;
        RECT 81.460 140.140 81.630 140.285 ;
        RECT 80.895 139.735 81.225 140.105 ;
        RECT 81.460 139.810 81.745 140.140 ;
        RECT 81.460 139.555 81.630 139.810 ;
        RECT 79.585 139.005 79.755 139.385 ;
        RECT 79.935 138.835 80.265 139.215 ;
        RECT 80.445 139.005 80.705 139.510 ;
        RECT 80.965 139.385 81.630 139.555 ;
        RECT 81.915 139.510 82.085 140.310 ;
        RECT 82.255 140.295 83.465 141.385 ;
        RECT 83.635 140.295 87.145 141.385 ;
        RECT 82.255 139.755 82.775 140.295 ;
        RECT 82.945 139.585 83.465 140.125 ;
        RECT 83.635 139.775 85.325 140.295 ;
        RECT 87.315 140.220 87.605 141.385 ;
        RECT 87.780 140.950 93.125 141.385 ;
        RECT 85.495 139.605 87.145 140.125 ;
        RECT 89.370 139.700 89.720 140.950 ;
        RECT 93.295 140.625 93.810 141.035 ;
        RECT 94.045 140.625 94.215 141.385 ;
        RECT 94.385 141.045 96.415 141.215 ;
        RECT 80.965 139.005 81.135 139.385 ;
        RECT 81.315 138.835 81.645 139.215 ;
        RECT 81.825 139.005 82.085 139.510 ;
        RECT 82.255 138.835 83.465 139.585 ;
        RECT 83.635 138.835 87.145 139.605 ;
        RECT 87.315 138.835 87.605 139.560 ;
        RECT 91.200 139.380 91.540 140.210 ;
        RECT 93.295 139.815 93.635 140.625 ;
        RECT 94.385 140.380 94.555 141.045 ;
        RECT 94.950 140.705 96.075 140.875 ;
        RECT 93.805 140.190 94.555 140.380 ;
        RECT 94.725 140.365 95.735 140.535 ;
        RECT 93.295 139.645 94.525 139.815 ;
        RECT 87.780 138.835 93.125 139.380 ;
        RECT 93.570 139.040 93.815 139.645 ;
        RECT 94.035 138.835 94.545 139.370 ;
        RECT 94.725 139.005 94.915 140.365 ;
        RECT 95.085 140.025 95.360 140.165 ;
        RECT 95.085 139.855 95.365 140.025 ;
        RECT 95.085 139.005 95.360 139.855 ;
        RECT 95.565 139.565 95.735 140.365 ;
        RECT 95.905 139.575 96.075 140.705 ;
        RECT 96.245 140.075 96.415 141.045 ;
        RECT 96.585 140.245 96.755 141.385 ;
        RECT 96.925 140.245 97.260 141.215 ;
        RECT 96.245 139.745 96.440 140.075 ;
        RECT 96.665 139.745 96.920 140.075 ;
        RECT 96.665 139.575 96.835 139.745 ;
        RECT 97.090 139.575 97.260 140.245 ;
        RECT 97.895 140.295 100.485 141.385 ;
        RECT 101.030 140.705 101.285 141.075 ;
        RECT 100.945 140.535 101.285 140.705 ;
        RECT 101.465 140.585 101.750 141.385 ;
        RECT 101.930 140.665 102.260 141.175 ;
        RECT 101.030 140.405 101.285 140.535 ;
        RECT 97.895 139.775 99.105 140.295 ;
        RECT 99.275 139.605 100.485 140.125 ;
        RECT 95.905 139.405 96.835 139.575 ;
        RECT 95.905 139.370 96.080 139.405 ;
        RECT 95.550 139.005 96.080 139.370 ;
        RECT 96.505 138.835 96.835 139.235 ;
        RECT 97.005 139.005 97.260 139.575 ;
        RECT 97.895 138.835 100.485 139.605 ;
        RECT 101.030 139.545 101.210 140.405 ;
        RECT 101.930 140.075 102.180 140.665 ;
        RECT 102.530 140.515 102.700 141.125 ;
        RECT 102.870 140.695 103.200 141.385 ;
        RECT 103.430 140.835 103.670 141.125 ;
        RECT 103.870 141.005 104.290 141.385 ;
        RECT 104.470 140.915 105.100 141.165 ;
        RECT 105.570 141.005 105.900 141.385 ;
        RECT 104.470 140.835 104.640 140.915 ;
        RECT 106.070 140.835 106.240 141.125 ;
        RECT 106.420 141.005 106.800 141.385 ;
        RECT 107.040 141.000 107.870 141.170 ;
        RECT 103.430 140.665 104.640 140.835 ;
        RECT 101.380 139.745 102.180 140.075 ;
        RECT 101.030 139.015 101.285 139.545 ;
        RECT 101.465 138.835 101.750 139.295 ;
        RECT 101.930 139.095 102.180 139.745 ;
        RECT 102.380 140.495 102.700 140.515 ;
        RECT 102.380 140.325 104.300 140.495 ;
        RECT 102.380 139.430 102.570 140.325 ;
        RECT 104.470 140.155 104.640 140.665 ;
        RECT 104.810 140.405 105.330 140.715 ;
        RECT 102.740 139.985 104.640 140.155 ;
        RECT 102.740 139.925 103.070 139.985 ;
        RECT 103.220 139.755 103.550 139.815 ;
        RECT 102.890 139.485 103.550 139.755 ;
        RECT 102.380 139.100 102.700 139.430 ;
        RECT 102.880 138.835 103.540 139.315 ;
        RECT 103.740 139.225 103.910 139.985 ;
        RECT 104.810 139.815 104.990 140.225 ;
        RECT 104.080 139.645 104.410 139.765 ;
        RECT 105.160 139.645 105.330 140.405 ;
        RECT 104.080 139.475 105.330 139.645 ;
        RECT 105.500 140.585 106.870 140.835 ;
        RECT 105.500 139.815 105.690 140.585 ;
        RECT 106.620 140.325 106.870 140.585 ;
        RECT 105.860 140.155 106.110 140.315 ;
        RECT 107.040 140.155 107.210 141.000 ;
        RECT 108.105 140.715 108.275 141.215 ;
        RECT 108.445 140.885 108.775 141.385 ;
        RECT 107.380 140.325 107.880 140.705 ;
        RECT 108.105 140.545 108.800 140.715 ;
        RECT 105.860 139.985 107.210 140.155 ;
        RECT 106.790 139.945 107.210 139.985 ;
        RECT 105.500 139.475 105.920 139.815 ;
        RECT 106.210 139.485 106.620 139.815 ;
        RECT 103.740 139.055 104.590 139.225 ;
        RECT 105.150 138.835 105.470 139.295 ;
        RECT 105.670 139.045 105.920 139.475 ;
        RECT 106.210 138.835 106.620 139.275 ;
        RECT 106.790 139.215 106.960 139.945 ;
        RECT 107.130 139.395 107.480 139.765 ;
        RECT 107.660 139.455 107.880 140.325 ;
        RECT 108.050 139.755 108.460 140.375 ;
        RECT 108.630 139.575 108.800 140.545 ;
        RECT 108.105 139.385 108.800 139.575 ;
        RECT 106.790 139.015 107.805 139.215 ;
        RECT 108.105 139.055 108.275 139.385 ;
        RECT 108.445 138.835 108.775 139.215 ;
        RECT 108.990 139.095 109.215 141.215 ;
        RECT 109.385 140.885 109.715 141.385 ;
        RECT 109.885 140.715 110.055 141.215 ;
        RECT 109.390 140.545 110.055 140.715 ;
        RECT 109.390 139.555 109.620 140.545 ;
        RECT 109.790 139.725 110.140 140.375 ;
        RECT 110.315 140.295 111.985 141.385 ;
        RECT 112.155 140.295 113.365 141.385 ;
        RECT 110.315 139.775 111.065 140.295 ;
        RECT 111.235 139.605 111.985 140.125 ;
        RECT 112.155 139.755 112.675 140.295 ;
        RECT 109.390 139.385 110.055 139.555 ;
        RECT 109.385 138.835 109.715 139.215 ;
        RECT 109.885 139.095 110.055 139.385 ;
        RECT 110.315 138.835 111.985 139.605 ;
        RECT 112.845 139.585 113.365 140.125 ;
        RECT 112.155 138.835 113.365 139.585 ;
        RECT 11.330 138.665 113.450 138.835 ;
        RECT 11.415 137.915 12.625 138.665 ;
        RECT 13.630 138.325 13.885 138.485 ;
        RECT 13.545 138.155 13.885 138.325 ;
        RECT 14.065 138.205 14.350 138.665 ;
        RECT 13.630 137.955 13.885 138.155 ;
        RECT 11.415 137.375 11.935 137.915 ;
        RECT 12.105 137.205 12.625 137.745 ;
        RECT 11.415 136.115 12.625 137.205 ;
        RECT 13.630 137.095 13.810 137.955 ;
        RECT 14.530 137.755 14.780 138.405 ;
        RECT 13.980 137.425 14.780 137.755 ;
        RECT 13.630 136.425 13.885 137.095 ;
        RECT 14.065 136.115 14.350 136.915 ;
        RECT 14.530 136.835 14.780 137.425 ;
        RECT 14.980 138.070 15.300 138.400 ;
        RECT 15.480 138.185 16.140 138.665 ;
        RECT 16.340 138.275 17.190 138.445 ;
        RECT 14.980 137.175 15.170 138.070 ;
        RECT 15.490 137.745 16.150 138.015 ;
        RECT 15.820 137.685 16.150 137.745 ;
        RECT 15.340 137.515 15.670 137.575 ;
        RECT 16.340 137.515 16.510 138.275 ;
        RECT 17.750 138.205 18.070 138.665 ;
        RECT 18.270 138.025 18.520 138.455 ;
        RECT 18.810 138.225 19.220 138.665 ;
        RECT 19.390 138.285 20.405 138.485 ;
        RECT 16.680 137.855 17.930 138.025 ;
        RECT 16.680 137.735 17.010 137.855 ;
        RECT 15.340 137.345 17.240 137.515 ;
        RECT 14.980 137.005 16.900 137.175 ;
        RECT 14.980 136.985 15.300 137.005 ;
        RECT 14.530 136.325 14.860 136.835 ;
        RECT 15.130 136.375 15.300 136.985 ;
        RECT 17.070 136.835 17.240 137.345 ;
        RECT 17.410 137.275 17.590 137.685 ;
        RECT 17.760 137.095 17.930 137.855 ;
        RECT 15.470 136.115 15.800 136.805 ;
        RECT 16.030 136.665 17.240 136.835 ;
        RECT 17.410 136.785 17.930 137.095 ;
        RECT 18.100 137.685 18.520 138.025 ;
        RECT 18.810 137.685 19.220 138.015 ;
        RECT 18.100 136.915 18.290 137.685 ;
        RECT 19.390 137.555 19.560 138.285 ;
        RECT 20.705 138.115 20.875 138.445 ;
        RECT 21.045 138.285 21.375 138.665 ;
        RECT 19.730 137.735 20.080 138.105 ;
        RECT 19.390 137.515 19.810 137.555 ;
        RECT 18.460 137.345 19.810 137.515 ;
        RECT 18.460 137.185 18.710 137.345 ;
        RECT 19.220 136.915 19.470 137.175 ;
        RECT 18.100 136.665 19.470 136.915 ;
        RECT 16.030 136.375 16.270 136.665 ;
        RECT 17.070 136.585 17.240 136.665 ;
        RECT 16.470 136.115 16.890 136.495 ;
        RECT 17.070 136.335 17.700 136.585 ;
        RECT 18.170 136.115 18.500 136.495 ;
        RECT 18.670 136.375 18.840 136.665 ;
        RECT 19.640 136.500 19.810 137.345 ;
        RECT 20.260 137.175 20.480 138.045 ;
        RECT 20.705 137.925 21.400 138.115 ;
        RECT 19.980 136.795 20.480 137.175 ;
        RECT 20.650 137.125 21.060 137.745 ;
        RECT 21.230 136.955 21.400 137.925 ;
        RECT 20.705 136.785 21.400 136.955 ;
        RECT 19.020 136.115 19.400 136.495 ;
        RECT 19.640 136.330 20.470 136.500 ;
        RECT 20.705 136.285 20.875 136.785 ;
        RECT 21.045 136.115 21.375 136.615 ;
        RECT 21.590 136.285 21.815 138.405 ;
        RECT 21.985 138.285 22.315 138.665 ;
        RECT 22.485 138.115 22.655 138.405 ;
        RECT 21.990 137.945 22.655 138.115 ;
        RECT 21.990 136.955 22.220 137.945 ;
        RECT 22.915 137.940 23.205 138.665 ;
        RECT 23.750 138.325 24.005 138.485 ;
        RECT 23.665 138.155 24.005 138.325 ;
        RECT 24.185 138.205 24.470 138.665 ;
        RECT 23.750 137.955 24.005 138.155 ;
        RECT 22.390 137.125 22.740 137.775 ;
        RECT 21.990 136.785 22.655 136.955 ;
        RECT 21.985 136.115 22.315 136.615 ;
        RECT 22.485 136.285 22.655 136.785 ;
        RECT 22.915 136.115 23.205 137.280 ;
        RECT 23.750 137.095 23.930 137.955 ;
        RECT 24.650 137.755 24.900 138.405 ;
        RECT 24.100 137.425 24.900 137.755 ;
        RECT 23.750 136.425 24.005 137.095 ;
        RECT 24.185 136.115 24.470 136.915 ;
        RECT 24.650 136.835 24.900 137.425 ;
        RECT 25.100 138.070 25.420 138.400 ;
        RECT 25.600 138.185 26.260 138.665 ;
        RECT 26.460 138.275 27.310 138.445 ;
        RECT 25.100 137.175 25.290 138.070 ;
        RECT 25.610 137.745 26.270 138.015 ;
        RECT 25.940 137.685 26.270 137.745 ;
        RECT 25.460 137.515 25.790 137.575 ;
        RECT 26.460 137.515 26.630 138.275 ;
        RECT 27.870 138.205 28.190 138.665 ;
        RECT 28.390 138.025 28.640 138.455 ;
        RECT 28.930 138.225 29.340 138.665 ;
        RECT 29.510 138.285 30.525 138.485 ;
        RECT 26.800 137.855 28.050 138.025 ;
        RECT 26.800 137.735 27.130 137.855 ;
        RECT 25.460 137.345 27.360 137.515 ;
        RECT 25.100 137.005 27.020 137.175 ;
        RECT 25.100 136.985 25.420 137.005 ;
        RECT 24.650 136.325 24.980 136.835 ;
        RECT 25.250 136.375 25.420 136.985 ;
        RECT 27.190 136.835 27.360 137.345 ;
        RECT 27.530 137.275 27.710 137.685 ;
        RECT 27.880 137.095 28.050 137.855 ;
        RECT 25.590 136.115 25.920 136.805 ;
        RECT 26.150 136.665 27.360 136.835 ;
        RECT 27.530 136.785 28.050 137.095 ;
        RECT 28.220 137.685 28.640 138.025 ;
        RECT 28.930 137.685 29.340 138.015 ;
        RECT 28.220 136.915 28.410 137.685 ;
        RECT 29.510 137.555 29.680 138.285 ;
        RECT 30.825 138.115 30.995 138.445 ;
        RECT 31.165 138.285 31.495 138.665 ;
        RECT 29.850 137.735 30.200 138.105 ;
        RECT 29.510 137.515 29.930 137.555 ;
        RECT 28.580 137.345 29.930 137.515 ;
        RECT 28.580 137.185 28.830 137.345 ;
        RECT 29.340 136.915 29.590 137.175 ;
        RECT 28.220 136.665 29.590 136.915 ;
        RECT 26.150 136.375 26.390 136.665 ;
        RECT 27.190 136.585 27.360 136.665 ;
        RECT 26.590 136.115 27.010 136.495 ;
        RECT 27.190 136.335 27.820 136.585 ;
        RECT 28.290 136.115 28.620 136.495 ;
        RECT 28.790 136.375 28.960 136.665 ;
        RECT 29.760 136.500 29.930 137.345 ;
        RECT 30.380 137.175 30.600 138.045 ;
        RECT 30.825 137.925 31.520 138.115 ;
        RECT 30.100 136.795 30.600 137.175 ;
        RECT 30.770 137.125 31.180 137.745 ;
        RECT 31.350 136.955 31.520 137.925 ;
        RECT 30.825 136.785 31.520 136.955 ;
        RECT 29.140 136.115 29.520 136.495 ;
        RECT 29.760 136.330 30.590 136.500 ;
        RECT 30.825 136.285 30.995 136.785 ;
        RECT 31.165 136.115 31.495 136.615 ;
        RECT 31.710 136.285 31.935 138.405 ;
        RECT 32.105 138.285 32.435 138.665 ;
        RECT 32.605 138.115 32.775 138.405 ;
        RECT 32.110 137.945 32.775 138.115 ;
        RECT 33.035 138.205 33.595 138.495 ;
        RECT 33.765 138.205 34.015 138.665 ;
        RECT 32.110 136.955 32.340 137.945 ;
        RECT 32.510 137.125 32.860 137.775 ;
        RECT 32.110 136.785 32.775 136.955 ;
        RECT 32.105 136.115 32.435 136.615 ;
        RECT 32.605 136.285 32.775 136.785 ;
        RECT 33.035 136.835 33.285 138.205 ;
        RECT 34.635 138.035 34.965 138.395 ;
        RECT 33.575 137.845 34.965 138.035 ;
        RECT 36.255 137.990 36.525 138.335 ;
        RECT 36.715 138.265 37.095 138.665 ;
        RECT 37.265 138.095 37.435 138.445 ;
        RECT 37.605 138.265 37.935 138.665 ;
        RECT 38.135 138.095 38.305 138.445 ;
        RECT 38.505 138.165 38.835 138.665 ;
        RECT 39.480 138.120 44.825 138.665 ;
        RECT 33.575 137.755 33.745 137.845 ;
        RECT 33.455 137.425 33.745 137.755 ;
        RECT 33.915 137.425 34.255 137.675 ;
        RECT 34.475 137.425 35.150 137.675 ;
        RECT 33.575 137.175 33.745 137.425 ;
        RECT 33.575 137.005 34.515 137.175 ;
        RECT 34.885 137.065 35.150 137.425 ;
        RECT 36.255 137.255 36.425 137.990 ;
        RECT 36.695 137.925 38.305 138.095 ;
        RECT 36.695 137.755 36.865 137.925 ;
        RECT 36.595 137.425 36.865 137.755 ;
        RECT 37.035 137.425 37.440 137.755 ;
        RECT 36.695 137.255 36.865 137.425 ;
        RECT 33.035 136.285 33.495 136.835 ;
        RECT 33.685 136.115 34.015 136.835 ;
        RECT 34.215 136.455 34.515 137.005 ;
        RECT 34.685 136.115 34.965 136.785 ;
        RECT 36.255 136.285 36.525 137.255 ;
        RECT 36.695 137.085 37.420 137.255 ;
        RECT 37.610 137.135 38.320 137.755 ;
        RECT 38.490 137.425 38.840 137.995 ;
        RECT 37.250 136.965 37.420 137.085 ;
        RECT 38.520 136.965 38.840 137.255 ;
        RECT 36.735 136.115 37.015 136.915 ;
        RECT 37.250 136.795 38.840 136.965 ;
        RECT 37.185 136.335 38.840 136.625 ;
        RECT 41.070 136.550 41.420 137.800 ;
        RECT 42.900 137.290 43.240 138.120 ;
        RECT 44.995 137.865 45.335 138.495 ;
        RECT 45.505 137.865 45.755 138.665 ;
        RECT 45.945 138.015 46.275 138.495 ;
        RECT 46.445 138.205 46.670 138.665 ;
        RECT 46.840 138.015 47.170 138.495 ;
        RECT 44.995 137.255 45.170 137.865 ;
        RECT 45.945 137.845 47.170 138.015 ;
        RECT 47.800 137.885 48.300 138.495 ;
        RECT 48.675 137.940 48.965 138.665 ;
        RECT 49.595 137.895 51.265 138.665 ;
        RECT 45.340 137.505 46.035 137.675 ;
        RECT 45.865 137.255 46.035 137.505 ;
        RECT 46.210 137.475 46.630 137.675 ;
        RECT 46.800 137.475 47.130 137.675 ;
        RECT 47.300 137.475 47.630 137.675 ;
        RECT 47.800 137.255 47.970 137.885 ;
        RECT 48.155 137.425 48.505 137.675 ;
        RECT 39.480 136.115 44.825 136.550 ;
        RECT 44.995 136.285 45.335 137.255 ;
        RECT 45.505 136.115 45.675 137.255 ;
        RECT 45.865 137.085 48.300 137.255 ;
        RECT 45.945 136.115 46.195 136.915 ;
        RECT 46.840 136.285 47.170 137.085 ;
        RECT 47.470 136.115 47.800 136.915 ;
        RECT 47.970 136.285 48.300 137.085 ;
        RECT 48.675 136.115 48.965 137.280 ;
        RECT 49.595 137.205 50.345 137.725 ;
        RECT 50.515 137.375 51.265 137.895 ;
        RECT 51.475 137.845 51.705 138.665 ;
        RECT 51.875 137.865 52.205 138.495 ;
        RECT 51.455 137.425 51.785 137.675 ;
        RECT 51.955 137.265 52.205 137.865 ;
        RECT 52.375 137.845 52.585 138.665 ;
        RECT 53.090 137.855 53.335 138.460 ;
        RECT 53.555 138.130 54.065 138.665 ;
        RECT 49.595 136.115 51.265 137.205 ;
        RECT 51.475 136.115 51.705 137.255 ;
        RECT 51.875 136.285 52.205 137.265 ;
        RECT 52.815 137.685 54.045 137.855 ;
        RECT 52.375 136.115 52.585 137.255 ;
        RECT 52.815 136.875 53.155 137.685 ;
        RECT 53.325 137.120 54.075 137.310 ;
        RECT 52.815 136.465 53.330 136.875 ;
        RECT 53.565 136.115 53.735 136.875 ;
        RECT 53.905 136.455 54.075 137.120 ;
        RECT 54.245 137.135 54.435 138.495 ;
        RECT 54.605 138.325 54.880 138.495 ;
        RECT 54.605 138.155 54.885 138.325 ;
        RECT 54.605 137.335 54.880 138.155 ;
        RECT 55.070 138.130 55.600 138.495 ;
        RECT 56.025 138.265 56.355 138.665 ;
        RECT 55.425 138.095 55.600 138.130 ;
        RECT 55.085 137.135 55.255 137.935 ;
        RECT 54.245 136.965 55.255 137.135 ;
        RECT 55.425 137.925 56.355 138.095 ;
        RECT 56.525 137.925 56.780 138.495 ;
        RECT 57.965 138.115 58.135 138.495 ;
        RECT 58.315 138.285 58.645 138.665 ;
        RECT 57.965 137.945 58.630 138.115 ;
        RECT 58.825 137.990 59.085 138.495 ;
        RECT 55.425 136.795 55.595 137.925 ;
        RECT 56.185 137.755 56.355 137.925 ;
        RECT 54.470 136.625 55.595 136.795 ;
        RECT 55.765 137.425 55.960 137.755 ;
        RECT 56.185 137.425 56.440 137.755 ;
        RECT 55.765 136.455 55.935 137.425 ;
        RECT 56.610 137.255 56.780 137.925 ;
        RECT 57.895 137.395 58.225 137.765 ;
        RECT 58.460 137.690 58.630 137.945 ;
        RECT 53.905 136.285 55.935 136.455 ;
        RECT 56.105 136.115 56.275 137.255 ;
        RECT 56.445 136.285 56.780 137.255 ;
        RECT 58.460 137.360 58.745 137.690 ;
        RECT 58.460 137.215 58.630 137.360 ;
        RECT 57.965 137.045 58.630 137.215 ;
        RECT 58.915 137.190 59.085 137.990 ;
        RECT 59.255 137.895 62.765 138.665 ;
        RECT 62.940 138.265 63.275 138.665 ;
        RECT 63.445 138.095 63.650 138.495 ;
        RECT 63.860 138.185 64.135 138.665 ;
        RECT 64.345 138.165 64.605 138.495 ;
        RECT 57.965 136.285 58.135 137.045 ;
        RECT 58.315 136.115 58.645 136.875 ;
        RECT 58.815 136.285 59.085 137.190 ;
        RECT 59.255 137.205 60.945 137.725 ;
        RECT 61.115 137.375 62.765 137.895 ;
        RECT 62.965 137.925 63.650 138.095 ;
        RECT 59.255 136.115 62.765 137.205 ;
        RECT 62.965 136.895 63.305 137.925 ;
        RECT 63.475 137.255 63.725 137.755 ;
        RECT 63.905 137.425 64.265 138.005 ;
        RECT 64.435 137.255 64.605 138.165 ;
        RECT 65.235 137.895 67.825 138.665 ;
        RECT 63.475 137.085 64.605 137.255 ;
        RECT 62.965 136.720 63.630 136.895 ;
        RECT 62.940 136.115 63.275 136.540 ;
        RECT 63.445 136.315 63.630 136.720 ;
        RECT 63.835 136.115 64.165 136.895 ;
        RECT 64.335 136.315 64.605 137.085 ;
        RECT 65.235 137.205 66.445 137.725 ;
        RECT 66.615 137.375 67.825 137.895 ;
        RECT 67.995 137.990 68.265 138.335 ;
        RECT 68.455 138.265 68.835 138.665 ;
        RECT 69.005 138.095 69.175 138.445 ;
        RECT 69.345 138.265 69.675 138.665 ;
        RECT 69.875 138.095 70.045 138.445 ;
        RECT 70.245 138.165 70.575 138.665 ;
        RECT 67.995 137.255 68.165 137.990 ;
        RECT 68.435 137.925 70.045 138.095 ;
        RECT 68.435 137.755 68.605 137.925 ;
        RECT 68.335 137.425 68.605 137.755 ;
        RECT 68.775 137.425 69.180 137.755 ;
        RECT 68.435 137.255 68.605 137.425 ;
        RECT 65.235 136.115 67.825 137.205 ;
        RECT 67.995 136.285 68.265 137.255 ;
        RECT 68.435 137.085 69.160 137.255 ;
        RECT 69.350 137.135 70.060 137.755 ;
        RECT 70.230 137.425 70.580 137.995 ;
        RECT 71.215 137.895 72.885 138.665 ;
        RECT 68.990 136.965 69.160 137.085 ;
        RECT 70.260 136.965 70.580 137.255 ;
        RECT 68.475 136.115 68.755 136.915 ;
        RECT 68.990 136.795 70.580 136.965 ;
        RECT 71.215 137.205 71.965 137.725 ;
        RECT 72.135 137.375 72.885 137.895 ;
        RECT 73.115 137.845 73.325 138.665 ;
        RECT 73.495 137.865 73.825 138.495 ;
        RECT 73.495 137.265 73.745 137.865 ;
        RECT 73.995 137.845 74.225 138.665 ;
        RECT 74.435 137.940 74.725 138.665 ;
        RECT 75.270 138.325 75.525 138.485 ;
        RECT 75.185 138.155 75.525 138.325 ;
        RECT 75.705 138.205 75.990 138.665 ;
        RECT 75.270 137.955 75.525 138.155 ;
        RECT 73.915 137.425 74.245 137.675 ;
        RECT 68.925 136.335 70.580 136.625 ;
        RECT 71.215 136.115 72.885 137.205 ;
        RECT 73.115 136.115 73.325 137.255 ;
        RECT 73.495 136.285 73.825 137.265 ;
        RECT 73.995 136.115 74.225 137.255 ;
        RECT 74.435 136.115 74.725 137.280 ;
        RECT 75.270 137.095 75.450 137.955 ;
        RECT 76.170 137.755 76.420 138.405 ;
        RECT 75.620 137.425 76.420 137.755 ;
        RECT 75.270 136.425 75.525 137.095 ;
        RECT 75.705 136.115 75.990 136.915 ;
        RECT 76.170 136.835 76.420 137.425 ;
        RECT 76.620 138.070 76.940 138.400 ;
        RECT 77.120 138.185 77.780 138.665 ;
        RECT 77.980 138.275 78.830 138.445 ;
        RECT 76.620 137.175 76.810 138.070 ;
        RECT 77.130 137.745 77.790 138.015 ;
        RECT 77.460 137.685 77.790 137.745 ;
        RECT 76.980 137.515 77.310 137.575 ;
        RECT 77.980 137.515 78.150 138.275 ;
        RECT 79.390 138.205 79.710 138.665 ;
        RECT 79.910 138.025 80.160 138.455 ;
        RECT 80.450 138.225 80.860 138.665 ;
        RECT 81.030 138.285 82.045 138.485 ;
        RECT 78.320 137.855 79.570 138.025 ;
        RECT 78.320 137.735 78.650 137.855 ;
        RECT 76.980 137.345 78.880 137.515 ;
        RECT 76.620 137.005 78.540 137.175 ;
        RECT 76.620 136.985 76.940 137.005 ;
        RECT 76.170 136.325 76.500 136.835 ;
        RECT 76.770 136.375 76.940 136.985 ;
        RECT 78.710 136.835 78.880 137.345 ;
        RECT 79.050 137.275 79.230 137.685 ;
        RECT 79.400 137.095 79.570 137.855 ;
        RECT 77.110 136.115 77.440 136.805 ;
        RECT 77.670 136.665 78.880 136.835 ;
        RECT 79.050 136.785 79.570 137.095 ;
        RECT 79.740 137.685 80.160 138.025 ;
        RECT 80.450 137.685 80.860 138.015 ;
        RECT 79.740 136.915 79.930 137.685 ;
        RECT 81.030 137.555 81.200 138.285 ;
        RECT 82.345 138.115 82.515 138.445 ;
        RECT 82.685 138.285 83.015 138.665 ;
        RECT 81.370 137.735 81.720 138.105 ;
        RECT 81.030 137.515 81.450 137.555 ;
        RECT 80.100 137.345 81.450 137.515 ;
        RECT 80.100 137.185 80.350 137.345 ;
        RECT 80.860 136.915 81.110 137.175 ;
        RECT 79.740 136.665 81.110 136.915 ;
        RECT 77.670 136.375 77.910 136.665 ;
        RECT 78.710 136.585 78.880 136.665 ;
        RECT 78.110 136.115 78.530 136.495 ;
        RECT 78.710 136.335 79.340 136.585 ;
        RECT 79.810 136.115 80.140 136.495 ;
        RECT 80.310 136.375 80.480 136.665 ;
        RECT 81.280 136.500 81.450 137.345 ;
        RECT 81.900 137.175 82.120 138.045 ;
        RECT 82.345 137.925 83.040 138.115 ;
        RECT 81.620 136.795 82.120 137.175 ;
        RECT 82.290 137.125 82.700 137.745 ;
        RECT 82.870 136.955 83.040 137.925 ;
        RECT 82.345 136.785 83.040 136.955 ;
        RECT 80.660 136.115 81.040 136.495 ;
        RECT 81.280 136.330 82.110 136.500 ;
        RECT 82.345 136.285 82.515 136.785 ;
        RECT 82.685 136.115 83.015 136.615 ;
        RECT 83.230 136.285 83.455 138.405 ;
        RECT 83.625 138.285 83.955 138.665 ;
        RECT 84.125 138.115 84.295 138.405 ;
        RECT 83.630 137.945 84.295 138.115 ;
        RECT 83.630 136.955 83.860 137.945 ;
        RECT 85.290 137.855 85.535 138.460 ;
        RECT 85.755 138.130 86.265 138.665 ;
        RECT 84.030 137.125 84.380 137.775 ;
        RECT 85.015 137.685 86.245 137.855 ;
        RECT 83.630 136.785 84.295 136.955 ;
        RECT 83.625 136.115 83.955 136.615 ;
        RECT 84.125 136.285 84.295 136.785 ;
        RECT 85.015 136.875 85.355 137.685 ;
        RECT 85.525 137.120 86.275 137.310 ;
        RECT 85.015 136.465 85.530 136.875 ;
        RECT 85.765 136.115 85.935 136.875 ;
        RECT 86.105 136.455 86.275 137.120 ;
        RECT 86.445 137.135 86.635 138.495 ;
        RECT 86.805 138.325 87.080 138.495 ;
        RECT 86.805 138.155 87.085 138.325 ;
        RECT 86.805 137.335 87.080 138.155 ;
        RECT 87.270 138.130 87.800 138.495 ;
        RECT 88.225 138.265 88.555 138.665 ;
        RECT 87.625 138.095 87.800 138.130 ;
        RECT 87.285 137.135 87.455 137.935 ;
        RECT 86.445 136.965 87.455 137.135 ;
        RECT 87.625 137.925 88.555 138.095 ;
        RECT 88.725 137.925 88.980 138.495 ;
        RECT 89.530 138.325 89.785 138.485 ;
        RECT 89.445 138.155 89.785 138.325 ;
        RECT 89.965 138.205 90.250 138.665 ;
        RECT 87.625 136.795 87.795 137.925 ;
        RECT 88.385 137.755 88.555 137.925 ;
        RECT 86.670 136.625 87.795 136.795 ;
        RECT 87.965 137.425 88.160 137.755 ;
        RECT 88.385 137.425 88.640 137.755 ;
        RECT 87.965 136.455 88.135 137.425 ;
        RECT 88.810 137.255 88.980 137.925 ;
        RECT 86.105 136.285 88.135 136.455 ;
        RECT 88.305 136.115 88.475 137.255 ;
        RECT 88.645 136.285 88.980 137.255 ;
        RECT 89.530 137.955 89.785 138.155 ;
        RECT 89.530 137.095 89.710 137.955 ;
        RECT 90.430 137.755 90.680 138.405 ;
        RECT 89.880 137.425 90.680 137.755 ;
        RECT 89.530 136.425 89.785 137.095 ;
        RECT 89.965 136.115 90.250 136.915 ;
        RECT 90.430 136.835 90.680 137.425 ;
        RECT 90.880 138.070 91.200 138.400 ;
        RECT 91.380 138.185 92.040 138.665 ;
        RECT 92.240 138.275 93.090 138.445 ;
        RECT 90.880 137.175 91.070 138.070 ;
        RECT 91.390 137.745 92.050 138.015 ;
        RECT 91.720 137.685 92.050 137.745 ;
        RECT 91.240 137.515 91.570 137.575 ;
        RECT 92.240 137.515 92.410 138.275 ;
        RECT 93.650 138.205 93.970 138.665 ;
        RECT 94.170 138.025 94.420 138.455 ;
        RECT 94.710 138.225 95.120 138.665 ;
        RECT 95.290 138.285 96.305 138.485 ;
        RECT 92.580 137.855 93.830 138.025 ;
        RECT 92.580 137.735 92.910 137.855 ;
        RECT 91.240 137.345 93.140 137.515 ;
        RECT 90.880 137.005 92.800 137.175 ;
        RECT 90.880 136.985 91.200 137.005 ;
        RECT 90.430 136.325 90.760 136.835 ;
        RECT 91.030 136.375 91.200 136.985 ;
        RECT 92.970 136.835 93.140 137.345 ;
        RECT 93.310 137.275 93.490 137.685 ;
        RECT 93.660 137.095 93.830 137.855 ;
        RECT 91.370 136.115 91.700 136.805 ;
        RECT 91.930 136.665 93.140 136.835 ;
        RECT 93.310 136.785 93.830 137.095 ;
        RECT 94.000 137.685 94.420 138.025 ;
        RECT 94.710 137.685 95.120 138.015 ;
        RECT 94.000 136.915 94.190 137.685 ;
        RECT 95.290 137.555 95.460 138.285 ;
        RECT 96.605 138.115 96.775 138.445 ;
        RECT 96.945 138.285 97.275 138.665 ;
        RECT 95.630 137.735 95.980 138.105 ;
        RECT 95.290 137.515 95.710 137.555 ;
        RECT 94.360 137.345 95.710 137.515 ;
        RECT 94.360 137.185 94.610 137.345 ;
        RECT 95.120 136.915 95.370 137.175 ;
        RECT 94.000 136.665 95.370 136.915 ;
        RECT 91.930 136.375 92.170 136.665 ;
        RECT 92.970 136.585 93.140 136.665 ;
        RECT 92.370 136.115 92.790 136.495 ;
        RECT 92.970 136.335 93.600 136.585 ;
        RECT 94.070 136.115 94.400 136.495 ;
        RECT 94.570 136.375 94.740 136.665 ;
        RECT 95.540 136.500 95.710 137.345 ;
        RECT 96.160 137.175 96.380 138.045 ;
        RECT 96.605 137.925 97.300 138.115 ;
        RECT 95.880 136.795 96.380 137.175 ;
        RECT 96.550 137.125 96.960 137.745 ;
        RECT 97.130 136.955 97.300 137.925 ;
        RECT 96.605 136.785 97.300 136.955 ;
        RECT 94.920 136.115 95.300 136.495 ;
        RECT 95.540 136.330 96.370 136.500 ;
        RECT 96.605 136.285 96.775 136.785 ;
        RECT 96.945 136.115 97.275 136.615 ;
        RECT 97.490 136.285 97.715 138.405 ;
        RECT 97.885 138.285 98.215 138.665 ;
        RECT 98.385 138.115 98.555 138.405 ;
        RECT 97.890 137.945 98.555 138.115 ;
        RECT 97.890 136.955 98.120 137.945 ;
        RECT 98.815 137.915 100.025 138.665 ;
        RECT 100.195 137.940 100.485 138.665 ;
        RECT 98.290 137.125 98.640 137.775 ;
        RECT 98.815 137.205 99.335 137.745 ;
        RECT 99.505 137.375 100.025 137.915 ;
        RECT 101.390 137.855 101.635 138.460 ;
        RECT 101.855 138.130 102.365 138.665 ;
        RECT 101.115 137.685 102.345 137.855 ;
        RECT 97.890 136.785 98.555 136.955 ;
        RECT 97.885 136.115 98.215 136.615 ;
        RECT 98.385 136.285 98.555 136.785 ;
        RECT 98.815 136.115 100.025 137.205 ;
        RECT 100.195 136.115 100.485 137.280 ;
        RECT 101.115 136.875 101.455 137.685 ;
        RECT 101.625 137.120 102.375 137.310 ;
        RECT 101.115 136.465 101.630 136.875 ;
        RECT 101.865 136.115 102.035 136.875 ;
        RECT 102.205 136.455 102.375 137.120 ;
        RECT 102.545 137.135 102.735 138.495 ;
        RECT 102.905 138.325 103.180 138.495 ;
        RECT 102.905 138.155 103.185 138.325 ;
        RECT 102.905 137.335 103.180 138.155 ;
        RECT 103.370 138.130 103.900 138.495 ;
        RECT 104.325 138.265 104.655 138.665 ;
        RECT 103.725 138.095 103.900 138.130 ;
        RECT 103.385 137.135 103.555 137.935 ;
        RECT 102.545 136.965 103.555 137.135 ;
        RECT 103.725 137.925 104.655 138.095 ;
        RECT 104.825 137.925 105.080 138.495 ;
        RECT 106.265 138.115 106.435 138.495 ;
        RECT 106.615 138.285 106.945 138.665 ;
        RECT 106.265 137.945 106.930 138.115 ;
        RECT 107.125 137.990 107.385 138.495 ;
        RECT 103.725 136.795 103.895 137.925 ;
        RECT 104.485 137.755 104.655 137.925 ;
        RECT 102.770 136.625 103.895 136.795 ;
        RECT 104.065 137.425 104.260 137.755 ;
        RECT 104.485 137.425 104.740 137.755 ;
        RECT 104.065 136.455 104.235 137.425 ;
        RECT 104.910 137.255 105.080 137.925 ;
        RECT 106.195 137.395 106.525 137.765 ;
        RECT 106.760 137.690 106.930 137.945 ;
        RECT 102.205 136.285 104.235 136.455 ;
        RECT 104.405 136.115 104.575 137.255 ;
        RECT 104.745 136.285 105.080 137.255 ;
        RECT 106.760 137.360 107.045 137.690 ;
        RECT 106.760 137.215 106.930 137.360 ;
        RECT 106.265 137.045 106.930 137.215 ;
        RECT 107.215 137.190 107.385 137.990 ;
        RECT 108.475 137.895 111.985 138.665 ;
        RECT 112.155 137.915 113.365 138.665 ;
        RECT 106.265 136.285 106.435 137.045 ;
        RECT 106.615 136.115 106.945 136.875 ;
        RECT 107.115 136.285 107.385 137.190 ;
        RECT 108.475 137.205 110.165 137.725 ;
        RECT 110.335 137.375 111.985 137.895 ;
        RECT 112.155 137.205 112.675 137.745 ;
        RECT 112.845 137.375 113.365 137.915 ;
        RECT 108.475 136.115 111.985 137.205 ;
        RECT 112.155 136.115 113.365 137.205 ;
        RECT 11.330 135.945 113.450 136.115 ;
        RECT 11.415 134.855 12.625 135.945 ;
        RECT 11.415 134.145 11.935 134.685 ;
        RECT 12.105 134.315 12.625 134.855 ;
        RECT 12.795 134.855 16.305 135.945 ;
        RECT 16.475 135.185 16.990 135.595 ;
        RECT 17.225 135.185 17.395 135.945 ;
        RECT 17.565 135.605 19.595 135.775 ;
        RECT 12.795 134.335 14.485 134.855 ;
        RECT 14.655 134.165 16.305 134.685 ;
        RECT 16.475 134.375 16.815 135.185 ;
        RECT 17.565 134.940 17.735 135.605 ;
        RECT 18.130 135.265 19.255 135.435 ;
        RECT 16.985 134.750 17.735 134.940 ;
        RECT 17.905 134.925 18.915 135.095 ;
        RECT 16.475 134.205 17.705 134.375 ;
        RECT 11.415 133.395 12.625 134.145 ;
        RECT 12.795 133.395 16.305 134.165 ;
        RECT 16.750 133.600 16.995 134.205 ;
        RECT 17.215 133.395 17.725 133.930 ;
        RECT 17.905 133.565 18.095 134.925 ;
        RECT 18.265 134.585 18.540 134.725 ;
        RECT 18.265 134.415 18.545 134.585 ;
        RECT 18.265 133.565 18.540 134.415 ;
        RECT 18.745 134.125 18.915 134.925 ;
        RECT 19.085 134.135 19.255 135.265 ;
        RECT 19.425 134.635 19.595 135.605 ;
        RECT 19.765 134.805 19.935 135.945 ;
        RECT 20.105 134.805 20.440 135.775 ;
        RECT 19.425 134.305 19.620 134.635 ;
        RECT 19.845 134.305 20.100 134.635 ;
        RECT 19.845 134.135 20.015 134.305 ;
        RECT 20.270 134.135 20.440 134.805 ;
        RECT 19.085 133.965 20.015 134.135 ;
        RECT 19.085 133.930 19.260 133.965 ;
        RECT 18.730 133.565 19.260 133.930 ;
        RECT 19.685 133.395 20.015 133.795 ;
        RECT 20.185 133.565 20.440 134.135 ;
        RECT 21.075 134.870 21.345 135.775 ;
        RECT 21.515 135.185 21.845 135.945 ;
        RECT 22.025 135.015 22.195 135.775 ;
        RECT 21.075 134.070 21.245 134.870 ;
        RECT 21.530 134.845 22.195 135.015 ;
        RECT 22.455 134.855 25.045 135.945 ;
        RECT 25.305 135.015 25.475 135.775 ;
        RECT 25.655 135.185 25.985 135.945 ;
        RECT 21.530 134.700 21.700 134.845 ;
        RECT 21.415 134.370 21.700 134.700 ;
        RECT 21.530 134.115 21.700 134.370 ;
        RECT 21.935 134.295 22.265 134.665 ;
        RECT 22.455 134.335 23.665 134.855 ;
        RECT 25.305 134.845 25.970 135.015 ;
        RECT 26.155 134.870 26.425 135.775 ;
        RECT 25.800 134.700 25.970 134.845 ;
        RECT 23.835 134.165 25.045 134.685 ;
        RECT 25.235 134.295 25.565 134.665 ;
        RECT 25.800 134.370 26.085 134.700 ;
        RECT 21.075 133.565 21.335 134.070 ;
        RECT 21.530 133.945 22.195 134.115 ;
        RECT 21.515 133.395 21.845 133.775 ;
        RECT 22.025 133.565 22.195 133.945 ;
        RECT 22.455 133.395 25.045 134.165 ;
        RECT 25.800 134.115 25.970 134.370 ;
        RECT 25.305 133.945 25.970 134.115 ;
        RECT 26.255 134.070 26.425 134.870 ;
        RECT 25.305 133.565 25.475 133.945 ;
        RECT 25.655 133.395 25.985 133.775 ;
        RECT 26.165 133.565 26.425 134.070 ;
        RECT 26.600 134.805 26.935 135.775 ;
        RECT 27.105 134.805 27.275 135.945 ;
        RECT 27.445 135.605 29.475 135.775 ;
        RECT 26.600 134.135 26.770 134.805 ;
        RECT 27.445 134.635 27.615 135.605 ;
        RECT 26.940 134.305 27.195 134.635 ;
        RECT 27.420 134.305 27.615 134.635 ;
        RECT 27.785 135.265 28.910 135.435 ;
        RECT 27.025 134.135 27.195 134.305 ;
        RECT 27.785 134.135 27.955 135.265 ;
        RECT 26.600 133.565 26.855 134.135 ;
        RECT 27.025 133.965 27.955 134.135 ;
        RECT 28.125 134.925 29.135 135.095 ;
        RECT 28.125 134.125 28.295 134.925 ;
        RECT 28.500 134.585 28.775 134.725 ;
        RECT 28.495 134.415 28.775 134.585 ;
        RECT 27.780 133.930 27.955 133.965 ;
        RECT 27.025 133.395 27.355 133.795 ;
        RECT 27.780 133.565 28.310 133.930 ;
        RECT 28.500 133.565 28.775 134.415 ;
        RECT 28.945 133.565 29.135 134.925 ;
        RECT 29.305 134.940 29.475 135.605 ;
        RECT 29.645 135.185 29.815 135.945 ;
        RECT 30.050 135.185 30.565 135.595 ;
        RECT 29.305 134.750 30.055 134.940 ;
        RECT 30.225 134.375 30.565 135.185 ;
        RECT 29.335 134.205 30.565 134.375 ;
        RECT 30.735 134.855 33.325 135.945 ;
        RECT 33.695 135.275 33.975 135.945 ;
        RECT 34.145 135.055 34.445 135.605 ;
        RECT 34.645 135.225 34.975 135.945 ;
        RECT 35.165 135.225 35.625 135.775 ;
        RECT 30.735 134.335 31.945 134.855 ;
        RECT 29.315 133.395 29.825 133.930 ;
        RECT 30.045 133.600 30.290 134.205 ;
        RECT 32.115 134.165 33.325 134.685 ;
        RECT 33.510 134.635 33.775 134.995 ;
        RECT 34.145 134.885 35.085 135.055 ;
        RECT 34.915 134.635 35.085 134.885 ;
        RECT 33.510 134.385 34.185 134.635 ;
        RECT 34.405 134.385 34.745 134.635 ;
        RECT 34.915 134.305 35.205 134.635 ;
        RECT 34.915 134.215 35.085 134.305 ;
        RECT 30.735 133.395 33.325 134.165 ;
        RECT 33.695 134.025 35.085 134.215 ;
        RECT 33.695 133.665 34.025 134.025 ;
        RECT 35.375 133.855 35.625 135.225 ;
        RECT 35.795 134.780 36.085 135.945 ;
        RECT 37.175 134.805 37.445 135.775 ;
        RECT 37.655 135.145 37.935 135.945 ;
        RECT 38.105 135.435 39.760 135.725 ;
        RECT 38.170 135.095 39.760 135.265 ;
        RECT 38.170 134.975 38.340 135.095 ;
        RECT 37.615 134.805 38.340 134.975 ;
        RECT 34.645 133.395 34.895 133.855 ;
        RECT 35.065 133.565 35.625 133.855 ;
        RECT 35.795 133.395 36.085 134.120 ;
        RECT 37.175 134.070 37.345 134.805 ;
        RECT 37.615 134.635 37.785 134.805 ;
        RECT 38.530 134.755 39.245 134.925 ;
        RECT 39.440 134.805 39.760 135.095 ;
        RECT 39.935 134.805 40.275 135.775 ;
        RECT 40.445 134.805 40.615 135.945 ;
        RECT 40.885 135.145 41.135 135.945 ;
        RECT 41.780 134.975 42.110 135.775 ;
        RECT 42.410 135.145 42.740 135.945 ;
        RECT 42.910 134.975 43.240 135.775 ;
        RECT 40.805 134.805 43.240 134.975 ;
        RECT 43.615 134.805 43.955 135.775 ;
        RECT 44.125 134.805 44.295 135.945 ;
        RECT 44.565 135.145 44.815 135.945 ;
        RECT 45.460 134.975 45.790 135.775 ;
        RECT 46.090 135.145 46.420 135.945 ;
        RECT 46.590 134.975 46.920 135.775 ;
        RECT 44.485 134.805 46.920 134.975 ;
        RECT 47.295 134.805 47.635 135.775 ;
        RECT 47.805 134.805 47.975 135.945 ;
        RECT 48.245 135.145 48.495 135.945 ;
        RECT 49.140 134.975 49.470 135.775 ;
        RECT 49.770 135.145 50.100 135.945 ;
        RECT 50.270 134.975 50.600 135.775 ;
        RECT 48.165 134.805 50.600 134.975 ;
        RECT 52.270 134.965 52.525 135.635 ;
        RECT 52.705 135.145 52.990 135.945 ;
        RECT 53.170 135.225 53.500 135.735 ;
        RECT 52.270 134.925 52.450 134.965 ;
        RECT 37.515 134.305 37.785 134.635 ;
        RECT 37.955 134.305 38.360 134.635 ;
        RECT 38.530 134.305 39.240 134.755 ;
        RECT 37.615 134.135 37.785 134.305 ;
        RECT 37.175 133.725 37.445 134.070 ;
        RECT 37.615 133.965 39.225 134.135 ;
        RECT 39.410 134.065 39.760 134.635 ;
        RECT 39.935 134.245 40.110 134.805 ;
        RECT 40.805 134.555 40.975 134.805 ;
        RECT 40.280 134.385 40.975 134.555 ;
        RECT 41.150 134.385 41.570 134.585 ;
        RECT 41.740 134.385 42.070 134.585 ;
        RECT 42.240 134.385 42.570 134.585 ;
        RECT 39.935 134.195 40.165 134.245 ;
        RECT 37.635 133.395 38.015 133.795 ;
        RECT 38.185 133.615 38.355 133.965 ;
        RECT 38.525 133.395 38.855 133.795 ;
        RECT 39.055 133.615 39.225 133.965 ;
        RECT 39.425 133.395 39.755 133.895 ;
        RECT 39.935 133.565 40.275 134.195 ;
        RECT 40.445 133.395 40.695 134.195 ;
        RECT 40.885 134.045 42.110 134.215 ;
        RECT 40.885 133.565 41.215 134.045 ;
        RECT 41.385 133.395 41.610 133.855 ;
        RECT 41.780 133.565 42.110 134.045 ;
        RECT 42.740 134.175 42.910 134.805 ;
        RECT 43.095 134.385 43.445 134.635 ;
        RECT 43.615 134.195 43.790 134.805 ;
        RECT 44.485 134.555 44.655 134.805 ;
        RECT 43.960 134.385 44.655 134.555 ;
        RECT 44.830 134.385 45.250 134.585 ;
        RECT 45.420 134.385 45.750 134.585 ;
        RECT 45.920 134.385 46.250 134.585 ;
        RECT 42.740 133.565 43.240 134.175 ;
        RECT 43.615 133.565 43.955 134.195 ;
        RECT 44.125 133.395 44.375 134.195 ;
        RECT 44.565 134.045 45.790 134.215 ;
        RECT 44.565 133.565 44.895 134.045 ;
        RECT 45.065 133.395 45.290 133.855 ;
        RECT 45.460 133.565 45.790 134.045 ;
        RECT 46.420 134.175 46.590 134.805 ;
        RECT 46.775 134.385 47.125 134.635 ;
        RECT 47.295 134.195 47.470 134.805 ;
        RECT 48.165 134.555 48.335 134.805 ;
        RECT 47.640 134.385 48.335 134.555 ;
        RECT 48.510 134.385 48.930 134.585 ;
        RECT 49.100 134.385 49.430 134.585 ;
        RECT 49.600 134.385 49.930 134.585 ;
        RECT 46.420 133.565 46.920 134.175 ;
        RECT 47.295 133.565 47.635 134.195 ;
        RECT 47.805 133.395 48.055 134.195 ;
        RECT 48.245 134.045 49.470 134.215 ;
        RECT 48.245 133.565 48.575 134.045 ;
        RECT 48.745 133.395 48.970 133.855 ;
        RECT 49.140 133.565 49.470 134.045 ;
        RECT 50.100 134.175 50.270 134.805 ;
        RECT 52.185 134.755 52.450 134.925 ;
        RECT 50.455 134.385 50.805 134.635 ;
        RECT 50.100 133.565 50.600 134.175 ;
        RECT 52.270 134.105 52.450 134.755 ;
        RECT 53.170 134.635 53.420 135.225 ;
        RECT 53.770 135.075 53.940 135.685 ;
        RECT 54.110 135.255 54.440 135.945 ;
        RECT 54.670 135.395 54.910 135.685 ;
        RECT 55.110 135.565 55.530 135.945 ;
        RECT 55.710 135.475 56.340 135.725 ;
        RECT 56.810 135.565 57.140 135.945 ;
        RECT 55.710 135.395 55.880 135.475 ;
        RECT 57.310 135.395 57.480 135.685 ;
        RECT 57.660 135.565 58.040 135.945 ;
        RECT 58.280 135.560 59.110 135.730 ;
        RECT 54.670 135.225 55.880 135.395 ;
        RECT 52.620 134.305 53.420 134.635 ;
        RECT 52.270 133.575 52.525 134.105 ;
        RECT 52.705 133.395 52.990 133.855 ;
        RECT 53.170 133.655 53.420 134.305 ;
        RECT 53.620 135.055 53.940 135.075 ;
        RECT 53.620 134.885 55.540 135.055 ;
        RECT 53.620 133.990 53.810 134.885 ;
        RECT 55.710 134.715 55.880 135.225 ;
        RECT 56.050 134.965 56.570 135.275 ;
        RECT 53.980 134.545 55.880 134.715 ;
        RECT 53.980 134.485 54.310 134.545 ;
        RECT 54.460 134.315 54.790 134.375 ;
        RECT 54.130 134.045 54.790 134.315 ;
        RECT 53.620 133.660 53.940 133.990 ;
        RECT 54.120 133.395 54.780 133.875 ;
        RECT 54.980 133.785 55.150 134.545 ;
        RECT 56.050 134.375 56.230 134.785 ;
        RECT 55.320 134.205 55.650 134.325 ;
        RECT 56.400 134.205 56.570 134.965 ;
        RECT 55.320 134.035 56.570 134.205 ;
        RECT 56.740 135.145 58.110 135.395 ;
        RECT 56.740 134.375 56.930 135.145 ;
        RECT 57.860 134.885 58.110 135.145 ;
        RECT 57.100 134.715 57.350 134.875 ;
        RECT 58.280 134.715 58.450 135.560 ;
        RECT 59.345 135.275 59.515 135.775 ;
        RECT 59.685 135.445 60.015 135.945 ;
        RECT 58.620 134.885 59.120 135.265 ;
        RECT 59.345 135.105 60.040 135.275 ;
        RECT 57.100 134.545 58.450 134.715 ;
        RECT 58.030 134.505 58.450 134.545 ;
        RECT 56.740 134.035 57.160 134.375 ;
        RECT 57.450 134.045 57.860 134.375 ;
        RECT 54.980 133.615 55.830 133.785 ;
        RECT 56.390 133.395 56.710 133.855 ;
        RECT 56.910 133.605 57.160 134.035 ;
        RECT 57.450 133.395 57.860 133.835 ;
        RECT 58.030 133.775 58.200 134.505 ;
        RECT 58.370 133.955 58.720 134.325 ;
        RECT 58.900 134.015 59.120 134.885 ;
        RECT 59.290 134.315 59.700 134.935 ;
        RECT 59.870 134.135 60.040 135.105 ;
        RECT 59.345 133.945 60.040 134.135 ;
        RECT 58.030 133.575 59.045 133.775 ;
        RECT 59.345 133.615 59.515 133.945 ;
        RECT 59.685 133.395 60.015 133.775 ;
        RECT 60.230 133.655 60.455 135.775 ;
        RECT 60.625 135.445 60.955 135.945 ;
        RECT 61.125 135.275 61.295 135.775 ;
        RECT 60.630 135.105 61.295 135.275 ;
        RECT 60.630 134.115 60.860 135.105 ;
        RECT 61.030 134.285 61.380 134.935 ;
        RECT 61.555 134.780 61.845 135.945 ;
        RECT 62.015 134.855 63.225 135.945 ;
        RECT 62.015 134.315 62.535 134.855 ;
        RECT 63.395 134.805 63.665 135.775 ;
        RECT 63.875 135.145 64.155 135.945 ;
        RECT 64.325 135.435 65.980 135.725 ;
        RECT 64.390 135.095 65.980 135.265 ;
        RECT 64.390 134.975 64.560 135.095 ;
        RECT 63.835 134.805 64.560 134.975 ;
        RECT 62.705 134.145 63.225 134.685 ;
        RECT 60.630 133.945 61.295 134.115 ;
        RECT 60.625 133.395 60.955 133.775 ;
        RECT 61.125 133.655 61.295 133.945 ;
        RECT 61.555 133.395 61.845 134.120 ;
        RECT 62.015 133.395 63.225 134.145 ;
        RECT 63.395 134.070 63.565 134.805 ;
        RECT 63.835 134.635 64.005 134.805 ;
        RECT 64.750 134.755 65.465 134.925 ;
        RECT 65.660 134.805 65.980 135.095 ;
        RECT 66.155 134.805 66.495 135.775 ;
        RECT 66.665 134.805 66.835 135.945 ;
        RECT 67.105 135.145 67.355 135.945 ;
        RECT 68.000 134.975 68.330 135.775 ;
        RECT 68.630 135.145 68.960 135.945 ;
        RECT 69.130 134.975 69.460 135.775 ;
        RECT 67.025 134.805 69.460 134.975 ;
        RECT 69.835 134.805 70.175 135.775 ;
        RECT 70.345 134.805 70.515 135.945 ;
        RECT 70.785 135.145 71.035 135.945 ;
        RECT 71.680 134.975 72.010 135.775 ;
        RECT 72.310 135.145 72.640 135.945 ;
        RECT 72.810 134.975 73.140 135.775 ;
        RECT 70.705 134.805 73.140 134.975 ;
        RECT 73.515 135.185 74.030 135.595 ;
        RECT 74.265 135.185 74.435 135.945 ;
        RECT 74.605 135.605 76.635 135.775 ;
        RECT 63.735 134.305 64.005 134.635 ;
        RECT 64.175 134.305 64.580 134.635 ;
        RECT 64.750 134.305 65.460 134.755 ;
        RECT 63.835 134.135 64.005 134.305 ;
        RECT 63.395 133.725 63.665 134.070 ;
        RECT 63.835 133.965 65.445 134.135 ;
        RECT 65.630 134.065 65.980 134.635 ;
        RECT 66.155 134.245 66.330 134.805 ;
        RECT 67.025 134.555 67.195 134.805 ;
        RECT 66.500 134.385 67.195 134.555 ;
        RECT 67.370 134.385 67.790 134.585 ;
        RECT 67.960 134.385 68.290 134.585 ;
        RECT 68.460 134.385 68.790 134.585 ;
        RECT 66.155 134.195 66.385 134.245 ;
        RECT 63.855 133.395 64.235 133.795 ;
        RECT 64.405 133.615 64.575 133.965 ;
        RECT 64.745 133.395 65.075 133.795 ;
        RECT 65.275 133.615 65.445 133.965 ;
        RECT 65.645 133.395 65.975 133.895 ;
        RECT 66.155 133.565 66.495 134.195 ;
        RECT 66.665 133.395 66.915 134.195 ;
        RECT 67.105 134.045 68.330 134.215 ;
        RECT 67.105 133.565 67.435 134.045 ;
        RECT 67.605 133.395 67.830 133.855 ;
        RECT 68.000 133.565 68.330 134.045 ;
        RECT 68.960 134.175 69.130 134.805 ;
        RECT 69.315 134.385 69.665 134.635 ;
        RECT 69.835 134.195 70.010 134.805 ;
        RECT 70.705 134.555 70.875 134.805 ;
        RECT 70.180 134.385 70.875 134.555 ;
        RECT 71.050 134.385 71.470 134.585 ;
        RECT 71.640 134.385 71.970 134.585 ;
        RECT 72.140 134.385 72.470 134.585 ;
        RECT 68.960 133.565 69.460 134.175 ;
        RECT 69.835 133.565 70.175 134.195 ;
        RECT 70.345 133.395 70.595 134.195 ;
        RECT 70.785 134.045 72.010 134.215 ;
        RECT 70.785 133.565 71.115 134.045 ;
        RECT 71.285 133.395 71.510 133.855 ;
        RECT 71.680 133.565 72.010 134.045 ;
        RECT 72.640 134.175 72.810 134.805 ;
        RECT 72.995 134.385 73.345 134.635 ;
        RECT 73.515 134.375 73.855 135.185 ;
        RECT 74.605 134.940 74.775 135.605 ;
        RECT 75.170 135.265 76.295 135.435 ;
        RECT 74.025 134.750 74.775 134.940 ;
        RECT 74.945 134.925 75.955 135.095 ;
        RECT 73.515 134.205 74.745 134.375 ;
        RECT 72.640 133.565 73.140 134.175 ;
        RECT 73.790 133.600 74.035 134.205 ;
        RECT 74.255 133.395 74.765 133.930 ;
        RECT 74.945 133.565 75.135 134.925 ;
        RECT 75.305 134.585 75.580 134.725 ;
        RECT 75.305 134.415 75.585 134.585 ;
        RECT 75.305 133.565 75.580 134.415 ;
        RECT 75.785 134.125 75.955 134.925 ;
        RECT 76.125 134.135 76.295 135.265 ;
        RECT 76.465 134.635 76.635 135.605 ;
        RECT 76.805 134.805 76.975 135.945 ;
        RECT 77.145 134.805 77.480 135.775 ;
        RECT 78.030 135.605 78.285 135.635 ;
        RECT 77.945 135.435 78.285 135.605 ;
        RECT 76.465 134.305 76.660 134.635 ;
        RECT 76.885 134.305 77.140 134.635 ;
        RECT 76.885 134.135 77.055 134.305 ;
        RECT 77.310 134.135 77.480 134.805 ;
        RECT 76.125 133.965 77.055 134.135 ;
        RECT 76.125 133.930 76.300 133.965 ;
        RECT 75.770 133.565 76.300 133.930 ;
        RECT 76.725 133.395 77.055 133.795 ;
        RECT 77.225 133.565 77.480 134.135 ;
        RECT 78.030 134.965 78.285 135.435 ;
        RECT 78.465 135.145 78.750 135.945 ;
        RECT 78.930 135.225 79.260 135.735 ;
        RECT 78.030 134.105 78.210 134.965 ;
        RECT 78.930 134.635 79.180 135.225 ;
        RECT 79.530 135.075 79.700 135.685 ;
        RECT 79.870 135.255 80.200 135.945 ;
        RECT 80.430 135.395 80.670 135.685 ;
        RECT 80.870 135.565 81.290 135.945 ;
        RECT 81.470 135.475 82.100 135.725 ;
        RECT 82.570 135.565 82.900 135.945 ;
        RECT 81.470 135.395 81.640 135.475 ;
        RECT 83.070 135.395 83.240 135.685 ;
        RECT 83.420 135.565 83.800 135.945 ;
        RECT 84.040 135.560 84.870 135.730 ;
        RECT 80.430 135.225 81.640 135.395 ;
        RECT 78.380 134.305 79.180 134.635 ;
        RECT 78.030 133.575 78.285 134.105 ;
        RECT 78.465 133.395 78.750 133.855 ;
        RECT 78.930 133.655 79.180 134.305 ;
        RECT 79.380 135.055 79.700 135.075 ;
        RECT 79.380 134.885 81.300 135.055 ;
        RECT 79.380 133.990 79.570 134.885 ;
        RECT 81.470 134.715 81.640 135.225 ;
        RECT 81.810 134.965 82.330 135.275 ;
        RECT 79.740 134.545 81.640 134.715 ;
        RECT 79.740 134.485 80.070 134.545 ;
        RECT 80.220 134.315 80.550 134.375 ;
        RECT 79.890 134.045 80.550 134.315 ;
        RECT 79.380 133.660 79.700 133.990 ;
        RECT 79.880 133.395 80.540 133.875 ;
        RECT 80.740 133.785 80.910 134.545 ;
        RECT 81.810 134.375 81.990 134.785 ;
        RECT 81.080 134.205 81.410 134.325 ;
        RECT 82.160 134.205 82.330 134.965 ;
        RECT 81.080 134.035 82.330 134.205 ;
        RECT 82.500 135.145 83.870 135.395 ;
        RECT 82.500 134.375 82.690 135.145 ;
        RECT 83.620 134.885 83.870 135.145 ;
        RECT 82.860 134.715 83.110 134.875 ;
        RECT 84.040 134.715 84.210 135.560 ;
        RECT 85.105 135.275 85.275 135.775 ;
        RECT 85.445 135.445 85.775 135.945 ;
        RECT 84.380 134.885 84.880 135.265 ;
        RECT 85.105 135.105 85.800 135.275 ;
        RECT 82.860 134.545 84.210 134.715 ;
        RECT 83.790 134.505 84.210 134.545 ;
        RECT 82.500 134.035 82.920 134.375 ;
        RECT 83.210 134.045 83.620 134.375 ;
        RECT 80.740 133.615 81.590 133.785 ;
        RECT 82.150 133.395 82.470 133.855 ;
        RECT 82.670 133.605 82.920 134.035 ;
        RECT 83.210 133.395 83.620 133.835 ;
        RECT 83.790 133.775 83.960 134.505 ;
        RECT 84.130 133.955 84.480 134.325 ;
        RECT 84.660 134.015 84.880 134.885 ;
        RECT 85.050 134.315 85.460 134.935 ;
        RECT 85.630 134.135 85.800 135.105 ;
        RECT 85.105 133.945 85.800 134.135 ;
        RECT 83.790 133.575 84.805 133.775 ;
        RECT 85.105 133.615 85.275 133.945 ;
        RECT 85.445 133.395 85.775 133.775 ;
        RECT 85.990 133.655 86.215 135.775 ;
        RECT 86.385 135.445 86.715 135.945 ;
        RECT 86.885 135.275 87.055 135.775 ;
        RECT 86.390 135.105 87.055 135.275 ;
        RECT 86.390 134.115 86.620 135.105 ;
        RECT 86.790 134.285 87.140 134.935 ;
        RECT 87.315 134.780 87.605 135.945 ;
        RECT 87.835 134.805 88.045 135.945 ;
        RECT 88.215 134.795 88.545 135.775 ;
        RECT 88.715 134.805 88.945 135.945 ;
        RECT 89.155 134.870 89.425 135.775 ;
        RECT 89.595 135.185 89.925 135.945 ;
        RECT 90.105 135.015 90.275 135.775 ;
        RECT 86.390 133.945 87.055 134.115 ;
        RECT 86.385 133.395 86.715 133.775 ;
        RECT 86.885 133.655 87.055 133.945 ;
        RECT 87.315 133.395 87.605 134.120 ;
        RECT 87.835 133.395 88.045 134.215 ;
        RECT 88.215 134.195 88.465 134.795 ;
        RECT 88.635 134.385 88.965 134.635 ;
        RECT 88.215 133.565 88.545 134.195 ;
        RECT 88.715 133.395 88.945 134.215 ;
        RECT 89.155 134.070 89.325 134.870 ;
        RECT 89.610 134.845 90.275 135.015 ;
        RECT 90.995 134.855 92.665 135.945 ;
        RECT 89.610 134.700 89.780 134.845 ;
        RECT 89.495 134.370 89.780 134.700 ;
        RECT 89.610 134.115 89.780 134.370 ;
        RECT 90.015 134.295 90.345 134.665 ;
        RECT 90.995 134.335 91.745 134.855 ;
        RECT 92.895 134.805 93.105 135.945 ;
        RECT 93.275 134.795 93.605 135.775 ;
        RECT 93.775 134.805 94.005 135.945 ;
        RECT 94.215 134.855 95.885 135.945 ;
        RECT 96.055 134.870 96.325 135.775 ;
        RECT 96.495 135.185 96.825 135.945 ;
        RECT 97.005 135.015 97.175 135.775 ;
        RECT 91.915 134.165 92.665 134.685 ;
        RECT 89.155 133.565 89.415 134.070 ;
        RECT 89.610 133.945 90.275 134.115 ;
        RECT 89.595 133.395 89.925 133.775 ;
        RECT 90.105 133.565 90.275 133.945 ;
        RECT 90.995 133.395 92.665 134.165 ;
        RECT 92.895 133.395 93.105 134.215 ;
        RECT 93.275 134.195 93.525 134.795 ;
        RECT 93.695 134.385 94.025 134.635 ;
        RECT 94.215 134.335 94.965 134.855 ;
        RECT 93.275 133.565 93.605 134.195 ;
        RECT 93.775 133.395 94.005 134.215 ;
        RECT 95.135 134.165 95.885 134.685 ;
        RECT 94.215 133.395 95.885 134.165 ;
        RECT 96.055 134.070 96.225 134.870 ;
        RECT 96.510 134.845 97.175 135.015 ;
        RECT 97.435 134.855 100.945 135.945 ;
        RECT 101.120 135.510 106.465 135.945 ;
        RECT 106.640 135.510 111.985 135.945 ;
        RECT 96.510 134.700 96.680 134.845 ;
        RECT 96.395 134.370 96.680 134.700 ;
        RECT 96.510 134.115 96.680 134.370 ;
        RECT 96.915 134.295 97.245 134.665 ;
        RECT 97.435 134.335 99.125 134.855 ;
        RECT 99.295 134.165 100.945 134.685 ;
        RECT 102.710 134.260 103.060 135.510 ;
        RECT 96.055 133.565 96.315 134.070 ;
        RECT 96.510 133.945 97.175 134.115 ;
        RECT 96.495 133.395 96.825 133.775 ;
        RECT 97.005 133.565 97.175 133.945 ;
        RECT 97.435 133.395 100.945 134.165 ;
        RECT 104.540 133.940 104.880 134.770 ;
        RECT 108.230 134.260 108.580 135.510 ;
        RECT 112.155 134.855 113.365 135.945 ;
        RECT 110.060 133.940 110.400 134.770 ;
        RECT 112.155 134.315 112.675 134.855 ;
        RECT 112.845 134.145 113.365 134.685 ;
        RECT 101.120 133.395 106.465 133.940 ;
        RECT 106.640 133.395 111.985 133.940 ;
        RECT 112.155 133.395 113.365 134.145 ;
        RECT 11.330 133.225 113.450 133.395 ;
        RECT 11.415 132.475 12.625 133.225 ;
        RECT 13.170 132.515 13.425 133.045 ;
        RECT 13.605 132.765 13.890 133.225 ;
        RECT 11.415 131.935 11.935 132.475 ;
        RECT 12.105 131.765 12.625 132.305 ;
        RECT 13.170 131.865 13.350 132.515 ;
        RECT 14.070 132.315 14.320 132.965 ;
        RECT 13.520 131.985 14.320 132.315 ;
        RECT 11.415 130.675 12.625 131.765 ;
        RECT 13.085 131.695 13.350 131.865 ;
        RECT 13.170 131.655 13.350 131.695 ;
        RECT 13.170 130.985 13.425 131.655 ;
        RECT 13.605 130.675 13.890 131.475 ;
        RECT 14.070 131.395 14.320 131.985 ;
        RECT 14.520 132.630 14.840 132.960 ;
        RECT 15.020 132.745 15.680 133.225 ;
        RECT 15.880 132.835 16.730 133.005 ;
        RECT 14.520 131.735 14.710 132.630 ;
        RECT 15.030 132.305 15.690 132.575 ;
        RECT 15.360 132.245 15.690 132.305 ;
        RECT 14.880 132.075 15.210 132.135 ;
        RECT 15.880 132.075 16.050 132.835 ;
        RECT 17.290 132.765 17.610 133.225 ;
        RECT 17.810 132.585 18.060 133.015 ;
        RECT 18.350 132.785 18.760 133.225 ;
        RECT 18.930 132.845 19.945 133.045 ;
        RECT 16.220 132.415 17.470 132.585 ;
        RECT 16.220 132.295 16.550 132.415 ;
        RECT 14.880 131.905 16.780 132.075 ;
        RECT 14.520 131.565 16.440 131.735 ;
        RECT 14.520 131.545 14.840 131.565 ;
        RECT 14.070 130.885 14.400 131.395 ;
        RECT 14.670 130.935 14.840 131.545 ;
        RECT 16.610 131.395 16.780 131.905 ;
        RECT 16.950 131.835 17.130 132.245 ;
        RECT 17.300 131.655 17.470 132.415 ;
        RECT 15.010 130.675 15.340 131.365 ;
        RECT 15.570 131.225 16.780 131.395 ;
        RECT 16.950 131.345 17.470 131.655 ;
        RECT 17.640 132.245 18.060 132.585 ;
        RECT 18.350 132.245 18.760 132.575 ;
        RECT 17.640 131.475 17.830 132.245 ;
        RECT 18.930 132.115 19.100 132.845 ;
        RECT 20.245 132.675 20.415 133.005 ;
        RECT 20.585 132.845 20.915 133.225 ;
        RECT 19.270 132.295 19.620 132.665 ;
        RECT 18.930 132.075 19.350 132.115 ;
        RECT 18.000 131.905 19.350 132.075 ;
        RECT 18.000 131.745 18.250 131.905 ;
        RECT 18.760 131.475 19.010 131.735 ;
        RECT 17.640 131.225 19.010 131.475 ;
        RECT 15.570 130.935 15.810 131.225 ;
        RECT 16.610 131.145 16.780 131.225 ;
        RECT 16.010 130.675 16.430 131.055 ;
        RECT 16.610 130.895 17.240 131.145 ;
        RECT 17.710 130.675 18.040 131.055 ;
        RECT 18.210 130.935 18.380 131.225 ;
        RECT 19.180 131.060 19.350 131.905 ;
        RECT 19.800 131.735 20.020 132.605 ;
        RECT 20.245 132.485 20.940 132.675 ;
        RECT 19.520 131.355 20.020 131.735 ;
        RECT 20.190 131.685 20.600 132.305 ;
        RECT 20.770 131.515 20.940 132.485 ;
        RECT 20.245 131.345 20.940 131.515 ;
        RECT 18.560 130.675 18.940 131.055 ;
        RECT 19.180 130.890 20.010 131.060 ;
        RECT 20.245 130.845 20.415 131.345 ;
        RECT 20.585 130.675 20.915 131.175 ;
        RECT 21.130 130.845 21.355 132.965 ;
        RECT 21.525 132.845 21.855 133.225 ;
        RECT 22.025 132.675 22.195 132.965 ;
        RECT 21.530 132.505 22.195 132.675 ;
        RECT 21.530 131.515 21.760 132.505 ;
        RECT 22.915 132.500 23.205 133.225 ;
        RECT 23.415 132.405 23.645 133.225 ;
        RECT 23.815 132.425 24.145 133.055 ;
        RECT 21.930 131.685 22.280 132.335 ;
        RECT 23.395 131.985 23.725 132.235 ;
        RECT 21.530 131.345 22.195 131.515 ;
        RECT 21.525 130.675 21.855 131.175 ;
        RECT 22.025 130.845 22.195 131.345 ;
        RECT 22.915 130.675 23.205 131.840 ;
        RECT 23.895 131.825 24.145 132.425 ;
        RECT 24.315 132.405 24.525 133.225 ;
        RECT 25.675 132.455 29.185 133.225 ;
        RECT 23.415 130.675 23.645 131.815 ;
        RECT 23.815 130.845 24.145 131.825 ;
        RECT 24.315 130.675 24.525 131.815 ;
        RECT 25.675 131.765 27.365 132.285 ;
        RECT 27.535 131.935 29.185 132.455 ;
        RECT 29.360 132.485 29.615 133.055 ;
        RECT 29.785 132.825 30.115 133.225 ;
        RECT 30.540 132.690 31.070 133.055 ;
        RECT 30.540 132.655 30.715 132.690 ;
        RECT 29.785 132.485 30.715 132.655 ;
        RECT 31.260 132.545 31.535 133.055 ;
        RECT 29.360 131.815 29.530 132.485 ;
        RECT 29.785 132.315 29.955 132.485 ;
        RECT 29.700 131.985 29.955 132.315 ;
        RECT 30.180 131.985 30.375 132.315 ;
        RECT 25.675 130.675 29.185 131.765 ;
        RECT 29.360 130.845 29.695 131.815 ;
        RECT 29.865 130.675 30.035 131.815 ;
        RECT 30.205 131.015 30.375 131.985 ;
        RECT 30.545 131.355 30.715 132.485 ;
        RECT 30.885 131.695 31.055 132.495 ;
        RECT 31.255 132.375 31.535 132.545 ;
        RECT 31.260 131.895 31.535 132.375 ;
        RECT 31.705 131.695 31.895 133.055 ;
        RECT 32.075 132.690 32.585 133.225 ;
        RECT 32.805 132.415 33.050 133.020 ;
        RECT 34.155 132.595 34.485 132.955 ;
        RECT 35.105 132.765 35.355 133.225 ;
        RECT 35.525 132.765 36.085 133.055 ;
        RECT 32.095 132.245 33.325 132.415 ;
        RECT 34.155 132.405 35.545 132.595 ;
        RECT 30.885 131.525 31.895 131.695 ;
        RECT 32.065 131.680 32.815 131.870 ;
        RECT 30.545 131.185 31.670 131.355 ;
        RECT 32.065 131.015 32.235 131.680 ;
        RECT 32.985 131.435 33.325 132.245 ;
        RECT 35.375 132.315 35.545 132.405 ;
        RECT 33.970 131.985 34.645 132.235 ;
        RECT 34.865 131.985 35.205 132.235 ;
        RECT 35.375 131.985 35.665 132.315 ;
        RECT 33.970 131.625 34.235 131.985 ;
        RECT 35.375 131.735 35.545 131.985 ;
        RECT 30.205 130.845 32.235 131.015 ;
        RECT 32.405 130.675 32.575 131.435 ;
        RECT 32.810 131.025 33.325 131.435 ;
        RECT 34.605 131.565 35.545 131.735 ;
        RECT 34.155 130.675 34.435 131.345 ;
        RECT 34.605 131.015 34.905 131.565 ;
        RECT 35.835 131.395 36.085 132.765 ;
        RECT 36.455 132.595 36.785 132.955 ;
        RECT 37.405 132.765 37.655 133.225 ;
        RECT 37.825 132.765 38.385 133.055 ;
        RECT 36.455 132.405 37.845 132.595 ;
        RECT 37.675 132.315 37.845 132.405 ;
        RECT 36.270 131.985 36.945 132.235 ;
        RECT 37.165 131.985 37.505 132.235 ;
        RECT 37.675 131.985 37.965 132.315 ;
        RECT 36.270 131.625 36.535 131.985 ;
        RECT 37.675 131.735 37.845 131.985 ;
        RECT 35.105 130.675 35.435 131.395 ;
        RECT 35.625 130.845 36.085 131.395 ;
        RECT 36.905 131.565 37.845 131.735 ;
        RECT 36.455 130.675 36.735 131.345 ;
        RECT 36.905 131.015 37.205 131.565 ;
        RECT 38.135 131.395 38.385 132.765 ;
        RECT 38.555 132.455 40.225 133.225 ;
        RECT 40.405 132.725 40.735 133.225 ;
        RECT 40.935 132.655 41.105 133.005 ;
        RECT 41.305 132.825 41.635 133.225 ;
        RECT 41.805 132.655 41.975 133.005 ;
        RECT 42.145 132.825 42.525 133.225 ;
        RECT 37.405 130.675 37.735 131.395 ;
        RECT 37.925 130.845 38.385 131.395 ;
        RECT 38.555 131.765 39.305 132.285 ;
        RECT 39.475 131.935 40.225 132.455 ;
        RECT 40.400 131.985 40.750 132.555 ;
        RECT 40.935 132.485 42.545 132.655 ;
        RECT 42.715 132.550 42.985 132.895 ;
        RECT 42.375 132.315 42.545 132.485 ;
        RECT 38.555 130.675 40.225 131.765 ;
        RECT 40.400 131.525 40.720 131.815 ;
        RECT 40.920 131.695 41.630 132.315 ;
        RECT 41.800 131.985 42.205 132.315 ;
        RECT 42.375 131.985 42.645 132.315 ;
        RECT 42.375 131.815 42.545 131.985 ;
        RECT 42.815 131.815 42.985 132.550 ;
        RECT 41.820 131.645 42.545 131.815 ;
        RECT 41.820 131.525 41.990 131.645 ;
        RECT 40.400 131.355 41.990 131.525 ;
        RECT 40.400 130.895 42.055 131.185 ;
        RECT 42.225 130.675 42.505 131.475 ;
        RECT 42.715 130.845 42.985 131.815 ;
        RECT 43.155 132.550 43.425 132.895 ;
        RECT 43.615 132.825 43.995 133.225 ;
        RECT 44.165 132.655 44.335 133.005 ;
        RECT 44.505 132.825 44.835 133.225 ;
        RECT 45.035 132.655 45.205 133.005 ;
        RECT 45.405 132.725 45.735 133.225 ;
        RECT 43.155 131.815 43.325 132.550 ;
        RECT 43.595 132.485 45.205 132.655 ;
        RECT 43.595 132.315 43.765 132.485 ;
        RECT 43.495 131.985 43.765 132.315 ;
        RECT 43.935 131.985 44.340 132.315 ;
        RECT 43.595 131.815 43.765 131.985 ;
        RECT 44.510 131.865 45.220 132.315 ;
        RECT 45.390 131.985 45.740 132.555 ;
        RECT 45.915 132.455 48.505 133.225 ;
        RECT 48.675 132.500 48.965 133.225 ;
        RECT 49.135 132.455 50.805 133.225 ;
        RECT 43.155 130.845 43.425 131.815 ;
        RECT 43.595 131.645 44.320 131.815 ;
        RECT 44.510 131.695 45.225 131.865 ;
        RECT 44.150 131.525 44.320 131.645 ;
        RECT 45.420 131.525 45.740 131.815 ;
        RECT 43.635 130.675 43.915 131.475 ;
        RECT 44.150 131.355 45.740 131.525 ;
        RECT 45.915 131.765 47.125 132.285 ;
        RECT 47.295 131.935 48.505 132.455 ;
        RECT 44.085 130.895 45.740 131.185 ;
        RECT 45.915 130.675 48.505 131.765 ;
        RECT 48.675 130.675 48.965 131.840 ;
        RECT 49.135 131.765 49.885 132.285 ;
        RECT 50.055 131.935 50.805 132.455 ;
        RECT 51.015 132.405 51.245 133.225 ;
        RECT 51.415 132.425 51.745 133.055 ;
        RECT 50.995 131.985 51.325 132.235 ;
        RECT 51.495 131.825 51.745 132.425 ;
        RECT 51.915 132.405 52.125 133.225 ;
        RECT 52.630 132.415 52.875 133.020 ;
        RECT 53.095 132.690 53.605 133.225 ;
        RECT 49.135 130.675 50.805 131.765 ;
        RECT 51.015 130.675 51.245 131.815 ;
        RECT 51.415 130.845 51.745 131.825 ;
        RECT 52.355 132.245 53.585 132.415 ;
        RECT 51.915 130.675 52.125 131.815 ;
        RECT 52.355 131.435 52.695 132.245 ;
        RECT 52.865 131.680 53.615 131.870 ;
        RECT 52.355 131.025 52.870 131.435 ;
        RECT 53.105 130.675 53.275 131.435 ;
        RECT 53.445 131.015 53.615 131.680 ;
        RECT 53.785 131.695 53.975 133.055 ;
        RECT 54.145 132.885 54.420 133.055 ;
        RECT 54.145 132.715 54.425 132.885 ;
        RECT 54.145 131.895 54.420 132.715 ;
        RECT 54.610 132.690 55.140 133.055 ;
        RECT 55.565 132.825 55.895 133.225 ;
        RECT 54.965 132.655 55.140 132.690 ;
        RECT 54.625 131.695 54.795 132.495 ;
        RECT 53.785 131.525 54.795 131.695 ;
        RECT 54.965 132.485 55.895 132.655 ;
        RECT 56.065 132.485 56.320 133.055 ;
        RECT 57.505 132.675 57.675 133.055 ;
        RECT 57.855 132.845 58.185 133.225 ;
        RECT 57.505 132.505 58.170 132.675 ;
        RECT 58.365 132.550 58.625 133.055 ;
        RECT 54.965 131.355 55.135 132.485 ;
        RECT 55.725 132.315 55.895 132.485 ;
        RECT 54.010 131.185 55.135 131.355 ;
        RECT 55.305 131.985 55.500 132.315 ;
        RECT 55.725 131.985 55.980 132.315 ;
        RECT 55.305 131.015 55.475 131.985 ;
        RECT 56.150 131.815 56.320 132.485 ;
        RECT 57.435 131.955 57.765 132.325 ;
        RECT 58.000 132.250 58.170 132.505 ;
        RECT 53.445 130.845 55.475 131.015 ;
        RECT 55.645 130.675 55.815 131.815 ;
        RECT 55.985 130.845 56.320 131.815 ;
        RECT 58.000 131.920 58.285 132.250 ;
        RECT 58.000 131.775 58.170 131.920 ;
        RECT 57.505 131.605 58.170 131.775 ;
        RECT 58.455 131.750 58.625 132.550 ;
        RECT 58.795 132.455 61.385 133.225 ;
        RECT 61.560 132.825 61.895 133.225 ;
        RECT 62.065 132.655 62.270 133.055 ;
        RECT 62.480 132.745 62.755 133.225 ;
        RECT 62.965 132.725 63.225 133.055 ;
        RECT 57.505 130.845 57.675 131.605 ;
        RECT 57.855 130.675 58.185 131.435 ;
        RECT 58.355 130.845 58.625 131.750 ;
        RECT 58.795 131.765 60.005 132.285 ;
        RECT 60.175 131.935 61.385 132.455 ;
        RECT 61.585 132.485 62.270 132.655 ;
        RECT 58.795 130.675 61.385 131.765 ;
        RECT 61.585 131.455 61.925 132.485 ;
        RECT 62.095 131.815 62.345 132.315 ;
        RECT 62.525 131.985 62.885 132.565 ;
        RECT 63.055 131.815 63.225 132.725 ;
        RECT 62.095 131.645 63.225 131.815 ;
        RECT 61.585 131.280 62.250 131.455 ;
        RECT 61.560 130.675 61.895 131.100 ;
        RECT 62.065 130.875 62.250 131.280 ;
        RECT 62.455 130.675 62.785 131.455 ;
        RECT 62.955 130.875 63.225 131.645 ;
        RECT 63.395 132.765 63.955 133.055 ;
        RECT 64.125 132.765 64.375 133.225 ;
        RECT 63.395 131.395 63.645 132.765 ;
        RECT 64.995 132.595 65.325 132.955 ;
        RECT 63.935 132.405 65.325 132.595 ;
        RECT 66.155 132.455 67.825 133.225 ;
        RECT 68.005 132.725 68.335 133.225 ;
        RECT 68.535 132.655 68.705 133.005 ;
        RECT 68.905 132.825 69.235 133.225 ;
        RECT 69.405 132.655 69.575 133.005 ;
        RECT 69.745 132.825 70.125 133.225 ;
        RECT 63.935 132.315 64.105 132.405 ;
        RECT 63.815 131.985 64.105 132.315 ;
        RECT 64.275 131.985 64.615 132.235 ;
        RECT 64.835 131.985 65.510 132.235 ;
        RECT 63.935 131.735 64.105 131.985 ;
        RECT 63.935 131.565 64.875 131.735 ;
        RECT 65.245 131.625 65.510 131.985 ;
        RECT 66.155 131.765 66.905 132.285 ;
        RECT 67.075 131.935 67.825 132.455 ;
        RECT 68.000 131.985 68.350 132.555 ;
        RECT 68.535 132.485 70.145 132.655 ;
        RECT 70.315 132.550 70.585 132.895 ;
        RECT 69.975 132.315 70.145 132.485 ;
        RECT 63.395 130.845 63.855 131.395 ;
        RECT 64.045 130.675 64.375 131.395 ;
        RECT 64.575 131.015 64.875 131.565 ;
        RECT 65.045 130.675 65.325 131.345 ;
        RECT 66.155 130.675 67.825 131.765 ;
        RECT 68.000 131.525 68.320 131.815 ;
        RECT 68.520 131.695 69.230 132.315 ;
        RECT 69.400 131.985 69.805 132.315 ;
        RECT 69.975 131.985 70.245 132.315 ;
        RECT 69.975 131.815 70.145 131.985 ;
        RECT 70.415 131.815 70.585 132.550 ;
        RECT 69.420 131.645 70.145 131.815 ;
        RECT 69.420 131.525 69.590 131.645 ;
        RECT 68.000 131.355 69.590 131.525 ;
        RECT 68.000 130.895 69.655 131.185 ;
        RECT 69.825 130.675 70.105 131.475 ;
        RECT 70.315 130.845 70.585 131.815 ;
        RECT 70.755 132.765 71.315 133.055 ;
        RECT 71.485 132.765 71.735 133.225 ;
        RECT 70.755 131.395 71.005 132.765 ;
        RECT 72.355 132.595 72.685 132.955 ;
        RECT 71.295 132.405 72.685 132.595 ;
        RECT 73.055 132.475 74.265 133.225 ;
        RECT 74.435 132.500 74.725 133.225 ;
        RECT 75.270 132.885 75.525 133.045 ;
        RECT 75.185 132.715 75.525 132.885 ;
        RECT 75.705 132.765 75.990 133.225 ;
        RECT 75.270 132.515 75.525 132.715 ;
        RECT 71.295 132.315 71.465 132.405 ;
        RECT 71.175 131.985 71.465 132.315 ;
        RECT 71.635 131.985 71.975 132.235 ;
        RECT 72.195 131.985 72.870 132.235 ;
        RECT 71.295 131.735 71.465 131.985 ;
        RECT 71.295 131.565 72.235 131.735 ;
        RECT 72.605 131.625 72.870 131.985 ;
        RECT 73.055 131.765 73.575 132.305 ;
        RECT 73.745 131.935 74.265 132.475 ;
        RECT 70.755 130.845 71.215 131.395 ;
        RECT 71.405 130.675 71.735 131.395 ;
        RECT 71.935 131.015 72.235 131.565 ;
        RECT 72.405 130.675 72.685 131.345 ;
        RECT 73.055 130.675 74.265 131.765 ;
        RECT 74.435 130.675 74.725 131.840 ;
        RECT 75.270 131.655 75.450 132.515 ;
        RECT 76.170 132.315 76.420 132.965 ;
        RECT 75.620 131.985 76.420 132.315 ;
        RECT 75.270 130.985 75.525 131.655 ;
        RECT 75.705 130.675 75.990 131.475 ;
        RECT 76.170 131.395 76.420 131.985 ;
        RECT 76.620 132.630 76.940 132.960 ;
        RECT 77.120 132.745 77.780 133.225 ;
        RECT 77.980 132.835 78.830 133.005 ;
        RECT 76.620 131.735 76.810 132.630 ;
        RECT 77.130 132.305 77.790 132.575 ;
        RECT 77.460 132.245 77.790 132.305 ;
        RECT 76.980 132.075 77.310 132.135 ;
        RECT 77.980 132.075 78.150 132.835 ;
        RECT 79.390 132.765 79.710 133.225 ;
        RECT 79.910 132.585 80.160 133.015 ;
        RECT 80.450 132.785 80.860 133.225 ;
        RECT 81.030 132.845 82.045 133.045 ;
        RECT 78.320 132.415 79.570 132.585 ;
        RECT 78.320 132.295 78.650 132.415 ;
        RECT 76.980 131.905 78.880 132.075 ;
        RECT 76.620 131.565 78.540 131.735 ;
        RECT 76.620 131.545 76.940 131.565 ;
        RECT 76.170 130.885 76.500 131.395 ;
        RECT 76.770 130.935 76.940 131.545 ;
        RECT 78.710 131.395 78.880 131.905 ;
        RECT 79.050 131.835 79.230 132.245 ;
        RECT 79.400 131.655 79.570 132.415 ;
        RECT 77.110 130.675 77.440 131.365 ;
        RECT 77.670 131.225 78.880 131.395 ;
        RECT 79.050 131.345 79.570 131.655 ;
        RECT 79.740 132.245 80.160 132.585 ;
        RECT 80.450 132.245 80.860 132.575 ;
        RECT 79.740 131.475 79.930 132.245 ;
        RECT 81.030 132.115 81.200 132.845 ;
        RECT 82.345 132.675 82.515 133.005 ;
        RECT 82.685 132.845 83.015 133.225 ;
        RECT 81.370 132.295 81.720 132.665 ;
        RECT 81.030 132.075 81.450 132.115 ;
        RECT 80.100 131.905 81.450 132.075 ;
        RECT 80.100 131.745 80.350 131.905 ;
        RECT 80.860 131.475 81.110 131.735 ;
        RECT 79.740 131.225 81.110 131.475 ;
        RECT 77.670 130.935 77.910 131.225 ;
        RECT 78.710 131.145 78.880 131.225 ;
        RECT 78.110 130.675 78.530 131.055 ;
        RECT 78.710 130.895 79.340 131.145 ;
        RECT 79.810 130.675 80.140 131.055 ;
        RECT 80.310 130.935 80.480 131.225 ;
        RECT 81.280 131.060 81.450 131.905 ;
        RECT 81.900 131.735 82.120 132.605 ;
        RECT 82.345 132.485 83.040 132.675 ;
        RECT 81.620 131.355 82.120 131.735 ;
        RECT 82.290 131.685 82.700 132.305 ;
        RECT 82.870 131.515 83.040 132.485 ;
        RECT 82.345 131.345 83.040 131.515 ;
        RECT 80.660 130.675 81.040 131.055 ;
        RECT 81.280 130.890 82.110 131.060 ;
        RECT 82.345 130.845 82.515 131.345 ;
        RECT 82.685 130.675 83.015 131.175 ;
        RECT 83.230 130.845 83.455 132.965 ;
        RECT 83.625 132.845 83.955 133.225 ;
        RECT 84.125 132.675 84.295 132.965 ;
        RECT 84.560 132.680 89.905 133.225 ;
        RECT 83.630 132.505 84.295 132.675 ;
        RECT 83.630 131.515 83.860 132.505 ;
        RECT 84.030 131.685 84.380 132.335 ;
        RECT 83.630 131.345 84.295 131.515 ;
        RECT 83.625 130.675 83.955 131.175 ;
        RECT 84.125 130.845 84.295 131.345 ;
        RECT 86.150 131.110 86.500 132.360 ;
        RECT 87.980 131.850 88.320 132.680 ;
        RECT 90.275 132.595 90.605 132.955 ;
        RECT 91.225 132.765 91.475 133.225 ;
        RECT 91.645 132.765 92.205 133.055 ;
        RECT 90.275 132.405 91.665 132.595 ;
        RECT 91.495 132.315 91.665 132.405 ;
        RECT 90.090 131.985 90.765 132.235 ;
        RECT 90.985 131.985 91.325 132.235 ;
        RECT 91.495 131.985 91.785 132.315 ;
        RECT 90.090 131.625 90.355 131.985 ;
        RECT 91.495 131.735 91.665 131.985 ;
        RECT 90.725 131.565 91.665 131.735 ;
        RECT 84.560 130.675 89.905 131.110 ;
        RECT 90.275 130.675 90.555 131.345 ;
        RECT 90.725 131.015 91.025 131.565 ;
        RECT 91.955 131.395 92.205 132.765 ;
        RECT 91.225 130.675 91.555 131.395 ;
        RECT 91.745 130.845 92.205 131.395 ;
        RECT 93.295 132.765 93.855 133.055 ;
        RECT 94.025 132.765 94.275 133.225 ;
        RECT 93.295 131.395 93.545 132.765 ;
        RECT 94.895 132.595 95.225 132.955 ;
        RECT 93.835 132.405 95.225 132.595 ;
        RECT 95.795 132.595 96.125 132.955 ;
        RECT 96.745 132.765 96.995 133.225 ;
        RECT 97.165 132.765 97.725 133.055 ;
        RECT 95.795 132.405 97.185 132.595 ;
        RECT 93.835 132.315 94.005 132.405 ;
        RECT 93.715 131.985 94.005 132.315 ;
        RECT 97.015 132.315 97.185 132.405 ;
        RECT 94.175 131.985 94.515 132.235 ;
        RECT 94.735 131.985 95.410 132.235 ;
        RECT 93.835 131.735 94.005 131.985 ;
        RECT 93.835 131.565 94.775 131.735 ;
        RECT 95.145 131.625 95.410 131.985 ;
        RECT 95.610 131.985 96.285 132.235 ;
        RECT 96.505 131.985 96.845 132.235 ;
        RECT 97.015 131.985 97.305 132.315 ;
        RECT 95.610 131.625 95.875 131.985 ;
        RECT 97.015 131.735 97.185 131.985 ;
        RECT 93.295 130.845 93.755 131.395 ;
        RECT 93.945 130.675 94.275 131.395 ;
        RECT 94.475 131.015 94.775 131.565 ;
        RECT 96.245 131.565 97.185 131.735 ;
        RECT 94.945 130.675 95.225 131.345 ;
        RECT 95.795 130.675 96.075 131.345 ;
        RECT 96.245 131.015 96.545 131.565 ;
        RECT 97.475 131.395 97.725 132.765 ;
        RECT 96.745 130.675 97.075 131.395 ;
        RECT 97.265 130.845 97.725 131.395 ;
        RECT 97.895 132.765 98.455 133.055 ;
        RECT 98.625 132.765 98.875 133.225 ;
        RECT 97.895 131.395 98.145 132.765 ;
        RECT 99.495 132.595 99.825 132.955 ;
        RECT 98.435 132.405 99.825 132.595 ;
        RECT 100.195 132.500 100.485 133.225 ;
        RECT 101.115 132.455 104.625 133.225 ;
        RECT 98.435 132.315 98.605 132.405 ;
        RECT 98.315 131.985 98.605 132.315 ;
        RECT 98.775 131.985 99.115 132.235 ;
        RECT 99.335 131.985 100.010 132.235 ;
        RECT 98.435 131.735 98.605 131.985 ;
        RECT 98.435 131.565 99.375 131.735 ;
        RECT 99.745 131.625 100.010 131.985 ;
        RECT 97.895 130.845 98.355 131.395 ;
        RECT 98.545 130.675 98.875 131.395 ;
        RECT 99.075 131.015 99.375 131.565 ;
        RECT 99.545 130.675 99.825 131.345 ;
        RECT 100.195 130.675 100.485 131.840 ;
        RECT 101.115 131.765 102.805 132.285 ;
        RECT 102.975 131.935 104.625 132.455 ;
        RECT 104.835 132.405 105.065 133.225 ;
        RECT 105.235 132.425 105.565 133.055 ;
        RECT 104.815 131.985 105.145 132.235 ;
        RECT 105.315 131.825 105.565 132.425 ;
        RECT 105.735 132.405 105.945 133.225 ;
        RECT 107.185 132.675 107.355 133.055 ;
        RECT 107.535 132.845 107.865 133.225 ;
        RECT 107.185 132.505 107.850 132.675 ;
        RECT 108.045 132.550 108.305 133.055 ;
        RECT 107.115 131.955 107.445 132.325 ;
        RECT 107.680 132.250 107.850 132.505 ;
        RECT 101.115 130.675 104.625 131.765 ;
        RECT 104.835 130.675 105.065 131.815 ;
        RECT 105.235 130.845 105.565 131.825 ;
        RECT 107.680 131.920 107.965 132.250 ;
        RECT 105.735 130.675 105.945 131.815 ;
        RECT 107.680 131.775 107.850 131.920 ;
        RECT 107.185 131.605 107.850 131.775 ;
        RECT 108.135 131.750 108.305 132.550 ;
        RECT 108.475 132.455 111.985 133.225 ;
        RECT 112.155 132.475 113.365 133.225 ;
        RECT 107.185 130.845 107.355 131.605 ;
        RECT 107.535 130.675 107.865 131.435 ;
        RECT 108.035 130.845 108.305 131.750 ;
        RECT 108.475 131.765 110.165 132.285 ;
        RECT 110.335 131.935 111.985 132.455 ;
        RECT 112.155 131.765 112.675 132.305 ;
        RECT 112.845 131.935 113.365 132.475 ;
        RECT 108.475 130.675 111.985 131.765 ;
        RECT 112.155 130.675 113.365 131.765 ;
        RECT 11.330 130.505 113.450 130.675 ;
        RECT 11.415 129.415 12.625 130.505 ;
        RECT 11.415 128.705 11.935 129.245 ;
        RECT 12.105 128.875 12.625 129.415 ;
        RECT 12.795 129.415 16.305 130.505 ;
        RECT 12.795 128.895 14.485 129.415 ;
        RECT 16.535 129.365 16.745 130.505 ;
        RECT 16.915 129.355 17.245 130.335 ;
        RECT 17.415 129.365 17.645 130.505 ;
        RECT 17.855 129.415 19.065 130.505 ;
        RECT 19.325 129.575 19.495 130.335 ;
        RECT 19.675 129.745 20.005 130.505 ;
        RECT 14.655 128.725 16.305 129.245 ;
        RECT 11.415 127.955 12.625 128.705 ;
        RECT 12.795 127.955 16.305 128.725 ;
        RECT 16.535 127.955 16.745 128.775 ;
        RECT 16.915 128.755 17.165 129.355 ;
        RECT 17.335 128.945 17.665 129.195 ;
        RECT 17.855 128.875 18.375 129.415 ;
        RECT 19.325 129.405 19.990 129.575 ;
        RECT 20.175 129.430 20.445 130.335 ;
        RECT 19.820 129.260 19.990 129.405 ;
        RECT 16.915 128.125 17.245 128.755 ;
        RECT 17.415 127.955 17.645 128.775 ;
        RECT 18.545 128.705 19.065 129.245 ;
        RECT 19.255 128.855 19.585 129.225 ;
        RECT 19.820 128.930 20.105 129.260 ;
        RECT 17.855 127.955 19.065 128.705 ;
        RECT 19.820 128.675 19.990 128.930 ;
        RECT 19.325 128.505 19.990 128.675 ;
        RECT 20.275 128.630 20.445 129.430 ;
        RECT 21.625 129.575 21.795 130.335 ;
        RECT 21.975 129.745 22.305 130.505 ;
        RECT 21.625 129.405 22.290 129.575 ;
        RECT 22.475 129.430 22.745 130.335 ;
        RECT 23.115 129.835 23.395 130.505 ;
        RECT 23.565 129.615 23.865 130.165 ;
        RECT 24.065 129.785 24.395 130.505 ;
        RECT 24.585 129.785 25.045 130.335 ;
        RECT 22.120 129.260 22.290 129.405 ;
        RECT 21.555 128.855 21.885 129.225 ;
        RECT 22.120 128.930 22.405 129.260 ;
        RECT 22.120 128.675 22.290 128.930 ;
        RECT 19.325 128.125 19.495 128.505 ;
        RECT 19.675 127.955 20.005 128.335 ;
        RECT 20.185 128.125 20.445 128.630 ;
        RECT 21.625 128.505 22.290 128.675 ;
        RECT 22.575 128.630 22.745 129.430 ;
        RECT 22.930 129.195 23.195 129.555 ;
        RECT 23.565 129.445 24.505 129.615 ;
        RECT 24.335 129.195 24.505 129.445 ;
        RECT 22.930 128.945 23.605 129.195 ;
        RECT 23.825 128.945 24.165 129.195 ;
        RECT 24.335 128.865 24.625 129.195 ;
        RECT 24.335 128.775 24.505 128.865 ;
        RECT 21.625 128.125 21.795 128.505 ;
        RECT 21.975 127.955 22.305 128.335 ;
        RECT 22.485 128.125 22.745 128.630 ;
        RECT 23.115 128.585 24.505 128.775 ;
        RECT 23.115 128.225 23.445 128.585 ;
        RECT 24.795 128.415 25.045 129.785 ;
        RECT 25.305 129.835 25.475 130.335 ;
        RECT 25.645 130.005 25.975 130.505 ;
        RECT 25.305 129.665 25.970 129.835 ;
        RECT 25.220 128.845 25.570 129.495 ;
        RECT 25.740 128.675 25.970 129.665 ;
        RECT 24.065 127.955 24.315 128.415 ;
        RECT 24.485 128.125 25.045 128.415 ;
        RECT 25.305 128.505 25.970 128.675 ;
        RECT 25.305 128.215 25.475 128.505 ;
        RECT 25.645 127.955 25.975 128.335 ;
        RECT 26.145 128.215 26.370 130.335 ;
        RECT 26.585 130.005 26.915 130.505 ;
        RECT 27.085 129.835 27.255 130.335 ;
        RECT 27.490 130.120 28.320 130.290 ;
        RECT 28.560 130.125 28.940 130.505 ;
        RECT 26.560 129.665 27.255 129.835 ;
        RECT 26.560 128.695 26.730 129.665 ;
        RECT 26.900 128.875 27.310 129.495 ;
        RECT 27.480 129.445 27.980 129.825 ;
        RECT 26.560 128.505 27.255 128.695 ;
        RECT 27.480 128.575 27.700 129.445 ;
        RECT 28.150 129.275 28.320 130.120 ;
        RECT 29.120 129.955 29.290 130.245 ;
        RECT 29.460 130.125 29.790 130.505 ;
        RECT 30.260 130.035 30.890 130.285 ;
        RECT 31.070 130.125 31.490 130.505 ;
        RECT 30.720 129.955 30.890 130.035 ;
        RECT 31.690 129.955 31.930 130.245 ;
        RECT 28.490 129.705 29.860 129.955 ;
        RECT 28.490 129.445 28.740 129.705 ;
        RECT 29.250 129.275 29.500 129.435 ;
        RECT 28.150 129.105 29.500 129.275 ;
        RECT 28.150 129.065 28.570 129.105 ;
        RECT 27.880 128.515 28.230 128.885 ;
        RECT 26.585 127.955 26.915 128.335 ;
        RECT 27.085 128.175 27.255 128.505 ;
        RECT 28.400 128.335 28.570 129.065 ;
        RECT 29.670 128.935 29.860 129.705 ;
        RECT 28.740 128.605 29.150 128.935 ;
        RECT 29.440 128.595 29.860 128.935 ;
        RECT 30.030 129.525 30.550 129.835 ;
        RECT 30.720 129.785 31.930 129.955 ;
        RECT 32.160 129.815 32.490 130.505 ;
        RECT 30.030 128.765 30.200 129.525 ;
        RECT 30.370 128.935 30.550 129.345 ;
        RECT 30.720 129.275 30.890 129.785 ;
        RECT 32.660 129.635 32.830 130.245 ;
        RECT 33.100 129.785 33.430 130.295 ;
        RECT 32.660 129.615 32.980 129.635 ;
        RECT 31.060 129.445 32.980 129.615 ;
        RECT 30.720 129.105 32.620 129.275 ;
        RECT 30.950 128.765 31.280 128.885 ;
        RECT 30.030 128.595 31.280 128.765 ;
        RECT 27.555 128.135 28.570 128.335 ;
        RECT 28.740 127.955 29.150 128.395 ;
        RECT 29.440 128.165 29.690 128.595 ;
        RECT 29.890 127.955 30.210 128.415 ;
        RECT 31.450 128.345 31.620 129.105 ;
        RECT 32.290 129.045 32.620 129.105 ;
        RECT 31.810 128.875 32.140 128.935 ;
        RECT 31.810 128.605 32.470 128.875 ;
        RECT 32.790 128.550 32.980 129.445 ;
        RECT 30.770 128.175 31.620 128.345 ;
        RECT 31.820 127.955 32.480 128.435 ;
        RECT 32.660 128.220 32.980 128.550 ;
        RECT 33.180 129.195 33.430 129.785 ;
        RECT 33.610 129.705 33.895 130.505 ;
        RECT 34.075 130.165 34.330 130.195 ;
        RECT 34.075 129.995 34.415 130.165 ;
        RECT 34.075 129.525 34.330 129.995 ;
        RECT 33.180 128.865 33.980 129.195 ;
        RECT 33.180 128.215 33.430 128.865 ;
        RECT 34.150 128.665 34.330 129.525 ;
        RECT 35.795 129.340 36.085 130.505 ;
        RECT 36.295 129.365 36.525 130.505 ;
        RECT 36.695 129.355 37.025 130.335 ;
        RECT 37.195 129.365 37.405 130.505 ;
        RECT 37.835 129.835 38.115 130.505 ;
        RECT 38.285 129.615 38.585 130.165 ;
        RECT 38.785 129.785 39.115 130.505 ;
        RECT 39.305 129.785 39.765 130.335 ;
        RECT 40.135 129.835 40.415 130.505 ;
        RECT 36.275 128.945 36.605 129.195 ;
        RECT 33.610 127.955 33.895 128.415 ;
        RECT 34.075 128.135 34.330 128.665 ;
        RECT 35.795 127.955 36.085 128.680 ;
        RECT 36.295 127.955 36.525 128.775 ;
        RECT 36.775 128.755 37.025 129.355 ;
        RECT 37.650 129.195 37.915 129.555 ;
        RECT 38.285 129.445 39.225 129.615 ;
        RECT 39.055 129.195 39.225 129.445 ;
        RECT 37.650 128.945 38.325 129.195 ;
        RECT 38.545 128.945 38.885 129.195 ;
        RECT 39.055 128.865 39.345 129.195 ;
        RECT 39.055 128.775 39.225 128.865 ;
        RECT 36.695 128.125 37.025 128.755 ;
        RECT 37.195 127.955 37.405 128.775 ;
        RECT 37.835 128.585 39.225 128.775 ;
        RECT 37.835 128.225 38.165 128.585 ;
        RECT 39.515 128.415 39.765 129.785 ;
        RECT 40.585 129.615 40.885 130.165 ;
        RECT 41.085 129.785 41.415 130.505 ;
        RECT 41.605 129.785 42.065 130.335 ;
        RECT 39.950 129.195 40.215 129.555 ;
        RECT 40.585 129.445 41.525 129.615 ;
        RECT 41.355 129.195 41.525 129.445 ;
        RECT 39.950 128.945 40.625 129.195 ;
        RECT 40.845 128.945 41.185 129.195 ;
        RECT 41.355 128.865 41.645 129.195 ;
        RECT 41.355 128.775 41.525 128.865 ;
        RECT 38.785 127.955 39.035 128.415 ;
        RECT 39.205 128.125 39.765 128.415 ;
        RECT 40.135 128.585 41.525 128.775 ;
        RECT 40.135 128.225 40.465 128.585 ;
        RECT 41.815 128.415 42.065 129.785 ;
        RECT 42.290 129.635 42.575 130.505 ;
        RECT 42.745 129.875 43.005 130.335 ;
        RECT 43.180 130.045 43.435 130.505 ;
        RECT 43.605 129.875 43.865 130.335 ;
        RECT 42.745 129.705 43.865 129.875 ;
        RECT 44.035 129.705 44.345 130.505 ;
        RECT 42.745 129.455 43.005 129.705 ;
        RECT 44.515 129.535 44.825 130.335 ;
        RECT 42.250 129.285 43.005 129.455 ;
        RECT 43.795 129.365 44.825 129.535 ;
        RECT 42.250 128.775 42.655 129.285 ;
        RECT 43.795 129.115 43.965 129.365 ;
        RECT 42.825 128.945 43.965 129.115 ;
        RECT 42.250 128.605 43.900 128.775 ;
        RECT 44.135 128.625 44.485 129.195 ;
        RECT 41.085 127.955 41.335 128.415 ;
        RECT 41.505 128.125 42.065 128.415 ;
        RECT 42.295 127.955 42.575 128.435 ;
        RECT 42.745 128.215 43.005 128.605 ;
        RECT 43.180 127.955 43.435 128.435 ;
        RECT 43.605 128.215 43.900 128.605 ;
        RECT 44.655 128.455 44.825 129.365 ;
        RECT 45.145 129.355 45.475 130.505 ;
        RECT 45.645 129.485 45.815 130.335 ;
        RECT 45.985 129.705 46.315 130.505 ;
        RECT 46.485 129.485 46.655 130.335 ;
        RECT 46.835 129.705 47.075 130.505 ;
        RECT 47.245 129.525 47.575 130.335 ;
        RECT 45.645 129.315 46.655 129.485 ;
        RECT 46.860 129.355 47.575 129.525 ;
        RECT 48.215 129.415 49.885 130.505 ;
        RECT 45.645 128.805 46.140 129.315 ;
        RECT 46.860 129.115 47.030 129.355 ;
        RECT 46.530 128.945 47.030 129.115 ;
        RECT 47.200 128.945 47.580 129.185 ;
        RECT 45.645 128.775 46.145 128.805 ;
        RECT 46.860 128.775 47.030 128.945 ;
        RECT 48.215 128.895 48.965 129.415 ;
        RECT 50.095 129.365 50.325 130.505 ;
        RECT 50.495 129.355 50.825 130.335 ;
        RECT 50.995 129.365 51.205 130.505 ;
        RECT 51.810 130.165 52.065 130.195 ;
        RECT 51.725 129.995 52.065 130.165 ;
        RECT 51.810 129.525 52.065 129.995 ;
        RECT 52.245 129.705 52.530 130.505 ;
        RECT 52.710 129.785 53.040 130.295 ;
        RECT 44.080 127.955 44.355 128.435 ;
        RECT 44.525 128.125 44.825 128.455 ;
        RECT 45.145 127.955 45.475 128.755 ;
        RECT 45.645 128.605 46.655 128.775 ;
        RECT 46.860 128.605 47.495 128.775 ;
        RECT 49.135 128.725 49.885 129.245 ;
        RECT 50.075 128.945 50.405 129.195 ;
        RECT 45.645 128.125 45.815 128.605 ;
        RECT 45.985 127.955 46.315 128.435 ;
        RECT 46.485 128.125 46.655 128.605 ;
        RECT 46.905 127.955 47.145 128.435 ;
        RECT 47.325 128.125 47.495 128.605 ;
        RECT 48.215 127.955 49.885 128.725 ;
        RECT 50.095 127.955 50.325 128.775 ;
        RECT 50.575 128.755 50.825 129.355 ;
        RECT 50.495 128.125 50.825 128.755 ;
        RECT 50.995 127.955 51.205 128.775 ;
        RECT 51.810 128.665 51.990 129.525 ;
        RECT 52.710 129.195 52.960 129.785 ;
        RECT 53.310 129.635 53.480 130.245 ;
        RECT 53.650 129.815 53.980 130.505 ;
        RECT 54.210 129.955 54.450 130.245 ;
        RECT 54.650 130.125 55.070 130.505 ;
        RECT 55.250 130.035 55.880 130.285 ;
        RECT 56.350 130.125 56.680 130.505 ;
        RECT 55.250 129.955 55.420 130.035 ;
        RECT 56.850 129.955 57.020 130.245 ;
        RECT 57.200 130.125 57.580 130.505 ;
        RECT 57.820 130.120 58.650 130.290 ;
        RECT 54.210 129.785 55.420 129.955 ;
        RECT 52.160 128.865 52.960 129.195 ;
        RECT 51.810 128.135 52.065 128.665 ;
        RECT 52.245 127.955 52.530 128.415 ;
        RECT 52.710 128.215 52.960 128.865 ;
        RECT 53.160 129.615 53.480 129.635 ;
        RECT 53.160 129.445 55.080 129.615 ;
        RECT 53.160 128.550 53.350 129.445 ;
        RECT 55.250 129.275 55.420 129.785 ;
        RECT 55.590 129.525 56.110 129.835 ;
        RECT 53.520 129.105 55.420 129.275 ;
        RECT 53.520 129.045 53.850 129.105 ;
        RECT 54.000 128.875 54.330 128.935 ;
        RECT 53.670 128.605 54.330 128.875 ;
        RECT 53.160 128.220 53.480 128.550 ;
        RECT 53.660 127.955 54.320 128.435 ;
        RECT 54.520 128.345 54.690 129.105 ;
        RECT 55.590 128.935 55.770 129.345 ;
        RECT 54.860 128.765 55.190 128.885 ;
        RECT 55.940 128.765 56.110 129.525 ;
        RECT 54.860 128.595 56.110 128.765 ;
        RECT 56.280 129.705 57.650 129.955 ;
        RECT 56.280 128.935 56.470 129.705 ;
        RECT 57.400 129.445 57.650 129.705 ;
        RECT 56.640 129.275 56.890 129.435 ;
        RECT 57.820 129.275 57.990 130.120 ;
        RECT 58.885 129.835 59.055 130.335 ;
        RECT 59.225 130.005 59.555 130.505 ;
        RECT 58.160 129.445 58.660 129.825 ;
        RECT 58.885 129.665 59.580 129.835 ;
        RECT 56.640 129.105 57.990 129.275 ;
        RECT 57.570 129.065 57.990 129.105 ;
        RECT 56.280 128.595 56.700 128.935 ;
        RECT 56.990 128.605 57.400 128.935 ;
        RECT 54.520 128.175 55.370 128.345 ;
        RECT 55.930 127.955 56.250 128.415 ;
        RECT 56.450 128.165 56.700 128.595 ;
        RECT 56.990 127.955 57.400 128.395 ;
        RECT 57.570 128.335 57.740 129.065 ;
        RECT 57.910 128.515 58.260 128.885 ;
        RECT 58.440 128.575 58.660 129.445 ;
        RECT 58.830 128.875 59.240 129.495 ;
        RECT 59.410 128.695 59.580 129.665 ;
        RECT 58.885 128.505 59.580 128.695 ;
        RECT 57.570 128.135 58.585 128.335 ;
        RECT 58.885 128.175 59.055 128.505 ;
        RECT 59.225 127.955 59.555 128.335 ;
        RECT 59.770 128.215 59.995 130.335 ;
        RECT 60.165 130.005 60.495 130.505 ;
        RECT 60.665 129.835 60.835 130.335 ;
        RECT 60.170 129.665 60.835 129.835 ;
        RECT 60.170 128.675 60.400 129.665 ;
        RECT 60.570 128.845 60.920 129.495 ;
        RECT 61.555 129.340 61.845 130.505 ;
        RECT 62.015 129.415 63.225 130.505 ;
        RECT 63.395 129.535 63.705 130.335 ;
        RECT 63.875 129.705 64.185 130.505 ;
        RECT 64.355 129.875 64.615 130.335 ;
        RECT 64.785 130.045 65.040 130.505 ;
        RECT 65.215 129.875 65.475 130.335 ;
        RECT 64.355 129.705 65.475 129.875 ;
        RECT 62.015 128.875 62.535 129.415 ;
        RECT 63.395 129.365 64.425 129.535 ;
        RECT 62.705 128.705 63.225 129.245 ;
        RECT 60.170 128.505 60.835 128.675 ;
        RECT 60.165 127.955 60.495 128.335 ;
        RECT 60.665 128.215 60.835 128.505 ;
        RECT 61.555 127.955 61.845 128.680 ;
        RECT 62.015 127.955 63.225 128.705 ;
        RECT 63.395 128.455 63.565 129.365 ;
        RECT 63.735 128.625 64.085 129.195 ;
        RECT 64.255 129.115 64.425 129.365 ;
        RECT 65.215 129.455 65.475 129.705 ;
        RECT 65.645 129.635 65.930 130.505 ;
        RECT 65.215 129.285 65.970 129.455 ;
        RECT 64.255 128.945 65.395 129.115 ;
        RECT 65.565 128.775 65.970 129.285 ;
        RECT 66.155 129.415 67.365 130.505 ;
        RECT 67.735 129.835 68.015 130.505 ;
        RECT 68.185 129.615 68.485 130.165 ;
        RECT 68.685 129.785 69.015 130.505 ;
        RECT 69.205 129.785 69.665 130.335 ;
        RECT 66.155 128.875 66.675 129.415 ;
        RECT 64.320 128.605 65.970 128.775 ;
        RECT 66.845 128.705 67.365 129.245 ;
        RECT 67.550 129.195 67.815 129.555 ;
        RECT 68.185 129.445 69.125 129.615 ;
        RECT 68.955 129.195 69.125 129.445 ;
        RECT 67.550 128.945 68.225 129.195 ;
        RECT 68.445 128.945 68.785 129.195 ;
        RECT 68.955 128.865 69.245 129.195 ;
        RECT 68.955 128.775 69.125 128.865 ;
        RECT 63.395 128.125 63.695 128.455 ;
        RECT 63.865 127.955 64.140 128.435 ;
        RECT 64.320 128.215 64.615 128.605 ;
        RECT 64.785 127.955 65.040 128.435 ;
        RECT 65.215 128.215 65.475 128.605 ;
        RECT 65.645 127.955 65.925 128.435 ;
        RECT 66.155 127.955 67.365 128.705 ;
        RECT 67.735 128.585 69.125 128.775 ;
        RECT 67.735 128.225 68.065 128.585 ;
        RECT 69.415 128.415 69.665 129.785 ;
        RECT 68.685 127.955 68.935 128.415 ;
        RECT 69.105 128.125 69.665 128.415 ;
        RECT 69.835 129.785 70.295 130.335 ;
        RECT 70.485 129.785 70.815 130.505 ;
        RECT 69.835 128.415 70.085 129.785 ;
        RECT 71.015 129.615 71.315 130.165 ;
        RECT 71.485 129.835 71.765 130.505 ;
        RECT 70.375 129.445 71.315 129.615 ;
        RECT 72.135 129.745 72.650 130.155 ;
        RECT 72.885 129.745 73.055 130.505 ;
        RECT 73.225 130.165 75.255 130.335 ;
        RECT 70.375 129.195 70.545 129.445 ;
        RECT 71.685 129.195 71.950 129.555 ;
        RECT 70.255 128.865 70.545 129.195 ;
        RECT 70.715 128.945 71.055 129.195 ;
        RECT 71.275 128.945 71.950 129.195 ;
        RECT 70.375 128.775 70.545 128.865 ;
        RECT 72.135 128.935 72.475 129.745 ;
        RECT 73.225 129.500 73.395 130.165 ;
        RECT 73.790 129.825 74.915 129.995 ;
        RECT 72.645 129.310 73.395 129.500 ;
        RECT 73.565 129.485 74.575 129.655 ;
        RECT 70.375 128.585 71.765 128.775 ;
        RECT 72.135 128.765 73.365 128.935 ;
        RECT 69.835 128.125 70.395 128.415 ;
        RECT 70.565 127.955 70.815 128.415 ;
        RECT 71.435 128.225 71.765 128.585 ;
        RECT 72.410 128.160 72.655 128.765 ;
        RECT 72.875 127.955 73.385 128.490 ;
        RECT 73.565 128.125 73.755 129.485 ;
        RECT 73.925 129.145 74.200 129.285 ;
        RECT 73.925 128.975 74.205 129.145 ;
        RECT 73.925 128.125 74.200 128.975 ;
        RECT 74.405 128.685 74.575 129.485 ;
        RECT 74.745 128.695 74.915 129.825 ;
        RECT 75.085 129.195 75.255 130.165 ;
        RECT 75.425 129.365 75.595 130.505 ;
        RECT 75.765 129.365 76.100 130.335 ;
        RECT 75.085 128.865 75.280 129.195 ;
        RECT 75.505 128.865 75.760 129.195 ;
        RECT 75.505 128.695 75.675 128.865 ;
        RECT 75.930 128.695 76.100 129.365 ;
        RECT 76.275 129.415 77.485 130.505 ;
        RECT 76.275 128.875 76.795 129.415 ;
        RECT 77.695 129.365 77.925 130.505 ;
        RECT 78.095 129.355 78.425 130.335 ;
        RECT 78.595 129.365 78.805 130.505 ;
        RECT 79.095 129.365 79.305 130.505 ;
        RECT 76.965 128.705 77.485 129.245 ;
        RECT 77.675 128.945 78.005 129.195 ;
        RECT 74.745 128.525 75.675 128.695 ;
        RECT 74.745 128.490 74.920 128.525 ;
        RECT 74.390 128.125 74.920 128.490 ;
        RECT 75.345 127.955 75.675 128.355 ;
        RECT 75.845 128.125 76.100 128.695 ;
        RECT 76.275 127.955 77.485 128.705 ;
        RECT 77.695 127.955 77.925 128.775 ;
        RECT 78.175 128.755 78.425 129.355 ;
        RECT 79.475 129.355 79.805 130.335 ;
        RECT 79.975 129.365 80.205 130.505 ;
        RECT 81.395 129.670 81.650 130.505 ;
        RECT 81.820 129.500 82.080 130.305 ;
        RECT 82.250 129.670 82.510 130.505 ;
        RECT 82.680 129.500 82.935 130.305 ;
        RECT 78.095 128.125 78.425 128.755 ;
        RECT 78.595 127.955 78.805 128.775 ;
        RECT 79.095 127.955 79.305 128.775 ;
        RECT 79.475 128.755 79.725 129.355 ;
        RECT 81.335 129.330 82.935 129.500 ;
        RECT 83.175 129.415 84.845 130.505 ;
        RECT 85.215 129.835 85.495 130.505 ;
        RECT 85.665 129.615 85.965 130.165 ;
        RECT 86.165 129.785 86.495 130.505 ;
        RECT 86.685 129.785 87.145 130.335 ;
        RECT 79.895 128.945 80.225 129.195 ;
        RECT 79.475 128.125 79.805 128.755 ;
        RECT 79.975 127.955 80.205 128.775 ;
        RECT 81.335 128.765 81.615 129.330 ;
        RECT 81.785 128.935 83.005 129.160 ;
        RECT 83.175 128.895 83.925 129.415 ;
        RECT 81.335 128.595 82.065 128.765 ;
        RECT 84.095 128.725 84.845 129.245 ;
        RECT 85.030 129.195 85.295 129.555 ;
        RECT 85.665 129.445 86.605 129.615 ;
        RECT 86.435 129.195 86.605 129.445 ;
        RECT 85.030 128.945 85.705 129.195 ;
        RECT 85.925 128.945 86.265 129.195 ;
        RECT 86.435 128.865 86.725 129.195 ;
        RECT 86.435 128.775 86.605 128.865 ;
        RECT 81.340 127.955 81.670 128.425 ;
        RECT 81.840 128.150 82.065 128.595 ;
        RECT 82.235 127.955 82.530 128.480 ;
        RECT 83.175 127.955 84.845 128.725 ;
        RECT 85.215 128.585 86.605 128.775 ;
        RECT 85.215 128.225 85.545 128.585 ;
        RECT 86.895 128.415 87.145 129.785 ;
        RECT 87.315 129.340 87.605 130.505 ;
        RECT 87.785 129.695 88.080 130.505 ;
        RECT 88.260 129.195 88.505 130.335 ;
        RECT 88.680 129.695 88.940 130.505 ;
        RECT 89.540 130.500 95.815 130.505 ;
        RECT 89.120 129.195 89.370 130.330 ;
        RECT 89.540 129.705 89.800 130.500 ;
        RECT 89.970 129.605 90.230 130.330 ;
        RECT 90.400 129.775 90.660 130.500 ;
        RECT 90.830 129.605 91.090 130.330 ;
        RECT 91.260 129.775 91.520 130.500 ;
        RECT 91.690 129.605 91.950 130.330 ;
        RECT 92.120 129.775 92.380 130.500 ;
        RECT 92.550 129.605 92.810 130.330 ;
        RECT 92.980 129.775 93.225 130.500 ;
        RECT 93.395 129.605 93.655 130.330 ;
        RECT 93.840 129.775 94.085 130.500 ;
        RECT 94.255 129.605 94.515 130.330 ;
        RECT 94.700 129.775 94.945 130.500 ;
        RECT 95.115 129.605 95.375 130.330 ;
        RECT 95.560 129.775 95.815 130.500 ;
        RECT 89.970 129.590 95.375 129.605 ;
        RECT 95.985 129.590 96.275 130.330 ;
        RECT 96.445 129.760 96.715 130.505 ;
        RECT 97.895 129.745 98.410 130.155 ;
        RECT 98.645 129.745 98.815 130.505 ;
        RECT 98.985 130.165 101.015 130.335 ;
        RECT 89.970 129.485 96.715 129.590 ;
        RECT 89.970 129.365 96.745 129.485 ;
        RECT 95.550 129.315 96.745 129.365 ;
        RECT 86.165 127.955 86.415 128.415 ;
        RECT 86.585 128.125 87.145 128.415 ;
        RECT 87.315 127.955 87.605 128.680 ;
        RECT 87.775 128.635 88.090 129.195 ;
        RECT 88.260 128.945 95.380 129.195 ;
        RECT 87.775 127.955 88.080 128.465 ;
        RECT 88.260 128.135 88.510 128.945 ;
        RECT 88.680 127.955 88.940 128.480 ;
        RECT 89.120 128.135 89.370 128.945 ;
        RECT 95.550 128.775 96.715 129.315 ;
        RECT 89.970 128.605 96.715 128.775 ;
        RECT 97.895 128.935 98.235 129.745 ;
        RECT 98.985 129.500 99.155 130.165 ;
        RECT 99.550 129.825 100.675 129.995 ;
        RECT 98.405 129.310 99.155 129.500 ;
        RECT 99.325 129.485 100.335 129.655 ;
        RECT 97.895 128.765 99.125 128.935 ;
        RECT 89.540 127.955 89.800 128.515 ;
        RECT 89.970 128.150 90.230 128.605 ;
        RECT 90.400 127.955 90.660 128.435 ;
        RECT 90.830 128.150 91.090 128.605 ;
        RECT 91.260 127.955 91.520 128.435 ;
        RECT 91.690 128.150 91.950 128.605 ;
        RECT 92.120 127.955 92.365 128.435 ;
        RECT 92.535 128.150 92.810 128.605 ;
        RECT 92.980 127.955 93.225 128.435 ;
        RECT 93.395 128.150 93.655 128.605 ;
        RECT 93.835 127.955 94.085 128.435 ;
        RECT 94.255 128.150 94.515 128.605 ;
        RECT 94.695 127.955 94.945 128.435 ;
        RECT 95.115 128.150 95.375 128.605 ;
        RECT 95.555 127.955 95.815 128.435 ;
        RECT 95.985 128.150 96.245 128.605 ;
        RECT 96.415 127.955 96.715 128.435 ;
        RECT 98.170 128.160 98.415 128.765 ;
        RECT 98.635 127.955 99.145 128.490 ;
        RECT 99.325 128.125 99.515 129.485 ;
        RECT 99.685 128.465 99.960 129.285 ;
        RECT 100.165 128.685 100.335 129.485 ;
        RECT 100.505 128.695 100.675 129.825 ;
        RECT 100.845 129.195 101.015 130.165 ;
        RECT 101.185 129.365 101.355 130.505 ;
        RECT 101.525 129.365 101.860 130.335 ;
        RECT 100.845 128.865 101.040 129.195 ;
        RECT 101.265 128.865 101.520 129.195 ;
        RECT 101.265 128.695 101.435 128.865 ;
        RECT 101.690 128.695 101.860 129.365 ;
        RECT 100.505 128.525 101.435 128.695 ;
        RECT 100.505 128.490 100.680 128.525 ;
        RECT 99.685 128.295 99.965 128.465 ;
        RECT 99.685 128.125 99.960 128.295 ;
        RECT 100.150 128.125 100.680 128.490 ;
        RECT 101.105 127.955 101.435 128.355 ;
        RECT 101.605 128.125 101.860 128.695 ;
        RECT 102.410 129.525 102.665 130.195 ;
        RECT 102.845 129.705 103.130 130.505 ;
        RECT 103.310 129.785 103.640 130.295 ;
        RECT 102.410 128.665 102.590 129.525 ;
        RECT 103.310 129.195 103.560 129.785 ;
        RECT 103.910 129.635 104.080 130.245 ;
        RECT 104.250 129.815 104.580 130.505 ;
        RECT 104.810 129.955 105.050 130.245 ;
        RECT 105.250 130.125 105.670 130.505 ;
        RECT 105.850 130.035 106.480 130.285 ;
        RECT 106.950 130.125 107.280 130.505 ;
        RECT 105.850 129.955 106.020 130.035 ;
        RECT 107.450 129.955 107.620 130.245 ;
        RECT 107.800 130.125 108.180 130.505 ;
        RECT 108.420 130.120 109.250 130.290 ;
        RECT 104.810 129.785 106.020 129.955 ;
        RECT 102.760 128.865 103.560 129.195 ;
        RECT 102.410 128.465 102.665 128.665 ;
        RECT 102.325 128.295 102.665 128.465 ;
        RECT 102.410 128.135 102.665 128.295 ;
        RECT 102.845 127.955 103.130 128.415 ;
        RECT 103.310 128.215 103.560 128.865 ;
        RECT 103.760 129.615 104.080 129.635 ;
        RECT 103.760 129.445 105.680 129.615 ;
        RECT 103.760 128.550 103.950 129.445 ;
        RECT 105.850 129.275 106.020 129.785 ;
        RECT 106.190 129.525 106.710 129.835 ;
        RECT 104.120 129.105 106.020 129.275 ;
        RECT 104.120 129.045 104.450 129.105 ;
        RECT 104.600 128.875 104.930 128.935 ;
        RECT 104.270 128.605 104.930 128.875 ;
        RECT 103.760 128.220 104.080 128.550 ;
        RECT 104.260 127.955 104.920 128.435 ;
        RECT 105.120 128.345 105.290 129.105 ;
        RECT 106.190 128.935 106.370 129.345 ;
        RECT 105.460 128.765 105.790 128.885 ;
        RECT 106.540 128.765 106.710 129.525 ;
        RECT 105.460 128.595 106.710 128.765 ;
        RECT 106.880 129.705 108.250 129.955 ;
        RECT 106.880 128.935 107.070 129.705 ;
        RECT 108.000 129.445 108.250 129.705 ;
        RECT 107.240 129.275 107.490 129.435 ;
        RECT 108.420 129.275 108.590 130.120 ;
        RECT 109.485 129.835 109.655 130.335 ;
        RECT 109.825 130.005 110.155 130.505 ;
        RECT 108.760 129.445 109.260 129.825 ;
        RECT 109.485 129.665 110.180 129.835 ;
        RECT 107.240 129.105 108.590 129.275 ;
        RECT 108.170 129.065 108.590 129.105 ;
        RECT 106.880 128.595 107.300 128.935 ;
        RECT 107.590 128.605 108.000 128.935 ;
        RECT 105.120 128.175 105.970 128.345 ;
        RECT 106.530 127.955 106.850 128.415 ;
        RECT 107.050 128.165 107.300 128.595 ;
        RECT 107.590 127.955 108.000 128.395 ;
        RECT 108.170 128.335 108.340 129.065 ;
        RECT 108.510 128.515 108.860 128.885 ;
        RECT 109.040 128.575 109.260 129.445 ;
        RECT 109.430 128.875 109.840 129.495 ;
        RECT 110.010 128.695 110.180 129.665 ;
        RECT 109.485 128.505 110.180 128.695 ;
        RECT 108.170 128.135 109.185 128.335 ;
        RECT 109.485 128.175 109.655 128.505 ;
        RECT 109.825 127.955 110.155 128.335 ;
        RECT 110.370 128.215 110.595 130.335 ;
        RECT 110.765 130.005 111.095 130.505 ;
        RECT 111.265 129.835 111.435 130.335 ;
        RECT 110.770 129.665 111.435 129.835 ;
        RECT 110.770 128.675 111.000 129.665 ;
        RECT 111.170 128.845 111.520 129.495 ;
        RECT 112.155 129.415 113.365 130.505 ;
        RECT 112.155 128.875 112.675 129.415 ;
        RECT 112.845 128.705 113.365 129.245 ;
        RECT 110.770 128.505 111.435 128.675 ;
        RECT 110.765 127.955 111.095 128.335 ;
        RECT 111.265 128.215 111.435 128.505 ;
        RECT 112.155 127.955 113.365 128.705 ;
        RECT 11.330 127.785 113.450 127.955 ;
        RECT 11.415 127.035 12.625 127.785 ;
        RECT 11.415 126.495 11.935 127.035 ;
        RECT 12.855 126.965 13.065 127.785 ;
        RECT 13.235 126.985 13.565 127.615 ;
        RECT 12.105 126.325 12.625 126.865 ;
        RECT 13.235 126.385 13.485 126.985 ;
        RECT 13.735 126.965 13.965 127.785 ;
        RECT 14.215 126.965 14.445 127.785 ;
        RECT 14.615 126.985 14.945 127.615 ;
        RECT 13.655 126.545 13.985 126.795 ;
        RECT 14.195 126.545 14.525 126.795 ;
        RECT 14.695 126.385 14.945 126.985 ;
        RECT 15.115 126.965 15.325 127.785 ;
        RECT 15.645 127.235 15.815 127.615 ;
        RECT 15.995 127.405 16.325 127.785 ;
        RECT 15.645 127.065 16.310 127.235 ;
        RECT 16.505 127.110 16.765 127.615 ;
        RECT 15.575 126.515 15.905 126.885 ;
        RECT 16.140 126.810 16.310 127.065 ;
        RECT 11.415 125.235 12.625 126.325 ;
        RECT 12.855 125.235 13.065 126.375 ;
        RECT 13.235 125.405 13.565 126.385 ;
        RECT 13.735 125.235 13.965 126.375 ;
        RECT 14.215 125.235 14.445 126.375 ;
        RECT 14.615 125.405 14.945 126.385 ;
        RECT 16.140 126.480 16.425 126.810 ;
        RECT 15.115 125.235 15.325 126.375 ;
        RECT 16.140 126.335 16.310 126.480 ;
        RECT 15.645 126.165 16.310 126.335 ;
        RECT 16.595 126.310 16.765 127.110 ;
        RECT 15.645 125.405 15.815 126.165 ;
        RECT 15.995 125.235 16.325 125.995 ;
        RECT 16.495 125.405 16.765 126.310 ;
        RECT 16.940 127.045 17.195 127.615 ;
        RECT 17.365 127.385 17.695 127.785 ;
        RECT 18.120 127.250 18.650 127.615 ;
        RECT 18.120 127.215 18.295 127.250 ;
        RECT 17.365 127.045 18.295 127.215 ;
        RECT 16.940 126.375 17.110 127.045 ;
        RECT 17.365 126.875 17.535 127.045 ;
        RECT 17.280 126.545 17.535 126.875 ;
        RECT 17.760 126.545 17.955 126.875 ;
        RECT 16.940 125.405 17.275 126.375 ;
        RECT 17.445 125.235 17.615 126.375 ;
        RECT 17.785 125.575 17.955 126.545 ;
        RECT 18.125 125.915 18.295 127.045 ;
        RECT 18.465 126.255 18.635 127.055 ;
        RECT 18.840 126.765 19.115 127.615 ;
        RECT 18.835 126.595 19.115 126.765 ;
        RECT 18.840 126.455 19.115 126.595 ;
        RECT 19.285 126.255 19.475 127.615 ;
        RECT 19.655 127.250 20.165 127.785 ;
        RECT 20.385 126.975 20.630 127.580 ;
        RECT 19.675 126.805 20.905 126.975 ;
        RECT 21.575 126.965 21.805 127.785 ;
        RECT 21.975 126.985 22.305 127.615 ;
        RECT 18.465 126.085 19.475 126.255 ;
        RECT 19.645 126.240 20.395 126.430 ;
        RECT 18.125 125.745 19.250 125.915 ;
        RECT 19.645 125.575 19.815 126.240 ;
        RECT 20.565 125.995 20.905 126.805 ;
        RECT 21.555 126.545 21.885 126.795 ;
        RECT 22.055 126.385 22.305 126.985 ;
        RECT 22.475 126.965 22.685 127.785 ;
        RECT 22.915 127.060 23.205 127.785 ;
        RECT 23.375 127.280 23.660 127.785 ;
        RECT 23.830 127.110 24.155 127.615 ;
        RECT 23.375 126.580 24.155 127.110 ;
        RECT 17.785 125.405 19.815 125.575 ;
        RECT 19.985 125.235 20.155 125.995 ;
        RECT 20.390 125.585 20.905 125.995 ;
        RECT 21.575 125.235 21.805 126.375 ;
        RECT 21.975 125.405 22.305 126.385 ;
        RECT 22.475 125.235 22.685 126.375 ;
        RECT 22.915 125.235 23.205 126.400 ;
        RECT 23.375 125.235 23.655 126.205 ;
        RECT 23.825 125.405 24.155 126.580 ;
        RECT 24.345 126.545 24.585 127.495 ;
        RECT 24.845 127.235 25.015 127.615 ;
        RECT 25.195 127.405 25.525 127.785 ;
        RECT 24.845 127.065 25.510 127.235 ;
        RECT 25.705 127.110 25.965 127.615 ;
        RECT 24.775 126.515 25.105 126.885 ;
        RECT 25.340 126.810 25.510 127.065 ;
        RECT 25.340 126.480 25.625 126.810 ;
        RECT 25.340 126.335 25.510 126.480 ;
        RECT 24.325 125.235 24.585 126.205 ;
        RECT 24.845 126.165 25.510 126.335 ;
        RECT 25.795 126.310 25.965 127.110 ;
        RECT 24.845 125.405 25.015 126.165 ;
        RECT 25.195 125.235 25.525 125.995 ;
        RECT 25.695 125.405 25.965 126.310 ;
        RECT 26.140 127.045 26.395 127.615 ;
        RECT 26.565 127.385 26.895 127.785 ;
        RECT 27.320 127.250 27.850 127.615 ;
        RECT 28.040 127.445 28.315 127.615 ;
        RECT 28.035 127.275 28.315 127.445 ;
        RECT 27.320 127.215 27.495 127.250 ;
        RECT 26.565 127.045 27.495 127.215 ;
        RECT 26.140 126.375 26.310 127.045 ;
        RECT 26.565 126.875 26.735 127.045 ;
        RECT 26.480 126.545 26.735 126.875 ;
        RECT 26.960 126.545 27.155 126.875 ;
        RECT 26.140 125.405 26.475 126.375 ;
        RECT 26.645 125.235 26.815 126.375 ;
        RECT 26.985 125.575 27.155 126.545 ;
        RECT 27.325 125.915 27.495 127.045 ;
        RECT 27.665 126.255 27.835 127.055 ;
        RECT 28.040 126.455 28.315 127.275 ;
        RECT 28.485 126.255 28.675 127.615 ;
        RECT 28.855 127.250 29.365 127.785 ;
        RECT 29.585 126.975 29.830 127.580 ;
        RECT 31.010 126.975 31.255 127.580 ;
        RECT 31.475 127.250 31.985 127.785 ;
        RECT 28.875 126.805 30.105 126.975 ;
        RECT 27.665 126.085 28.675 126.255 ;
        RECT 28.845 126.240 29.595 126.430 ;
        RECT 27.325 125.745 28.450 125.915 ;
        RECT 28.845 125.575 29.015 126.240 ;
        RECT 29.765 125.995 30.105 126.805 ;
        RECT 26.985 125.405 29.015 125.575 ;
        RECT 29.185 125.235 29.355 125.995 ;
        RECT 29.590 125.585 30.105 125.995 ;
        RECT 30.735 126.805 31.965 126.975 ;
        RECT 30.735 125.995 31.075 126.805 ;
        RECT 31.245 126.240 31.995 126.430 ;
        RECT 30.735 125.585 31.250 125.995 ;
        RECT 31.485 125.235 31.655 125.995 ;
        RECT 31.825 125.575 31.995 126.240 ;
        RECT 32.165 126.255 32.355 127.615 ;
        RECT 32.525 127.105 32.800 127.615 ;
        RECT 32.990 127.250 33.520 127.615 ;
        RECT 33.945 127.385 34.275 127.785 ;
        RECT 33.345 127.215 33.520 127.250 ;
        RECT 32.525 126.935 32.805 127.105 ;
        RECT 32.525 126.455 32.800 126.935 ;
        RECT 33.005 126.255 33.175 127.055 ;
        RECT 32.165 126.085 33.175 126.255 ;
        RECT 33.345 127.045 34.275 127.215 ;
        RECT 34.445 127.045 34.700 127.615 ;
        RECT 33.345 125.915 33.515 127.045 ;
        RECT 34.105 126.875 34.275 127.045 ;
        RECT 32.390 125.745 33.515 125.915 ;
        RECT 33.685 126.545 33.880 126.875 ;
        RECT 34.105 126.545 34.360 126.875 ;
        RECT 33.685 125.575 33.855 126.545 ;
        RECT 34.530 126.375 34.700 127.045 ;
        RECT 35.150 126.975 35.395 127.580 ;
        RECT 35.615 127.250 36.125 127.785 ;
        RECT 31.825 125.405 33.855 125.575 ;
        RECT 34.025 125.235 34.195 126.375 ;
        RECT 34.365 125.405 34.700 126.375 ;
        RECT 34.875 126.805 36.105 126.975 ;
        RECT 34.875 125.995 35.215 126.805 ;
        RECT 35.385 126.240 36.135 126.430 ;
        RECT 34.875 125.585 35.390 125.995 ;
        RECT 35.625 125.235 35.795 125.995 ;
        RECT 35.965 125.575 36.135 126.240 ;
        RECT 36.305 126.255 36.495 127.615 ;
        RECT 36.665 126.765 36.940 127.615 ;
        RECT 37.130 127.250 37.660 127.615 ;
        RECT 38.085 127.385 38.415 127.785 ;
        RECT 37.485 127.215 37.660 127.250 ;
        RECT 36.665 126.595 36.945 126.765 ;
        RECT 36.665 126.455 36.940 126.595 ;
        RECT 37.145 126.255 37.315 127.055 ;
        RECT 36.305 126.085 37.315 126.255 ;
        RECT 37.485 127.045 38.415 127.215 ;
        RECT 38.585 127.045 38.840 127.615 ;
        RECT 39.105 127.305 39.405 127.785 ;
        RECT 39.575 127.135 39.835 127.590 ;
        RECT 40.005 127.305 40.265 127.785 ;
        RECT 40.445 127.135 40.705 127.590 ;
        RECT 40.875 127.305 41.125 127.785 ;
        RECT 41.305 127.135 41.565 127.590 ;
        RECT 41.735 127.305 41.985 127.785 ;
        RECT 42.165 127.135 42.425 127.590 ;
        RECT 42.595 127.305 42.840 127.785 ;
        RECT 43.010 127.135 43.285 127.590 ;
        RECT 43.455 127.305 43.700 127.785 ;
        RECT 43.870 127.135 44.130 127.590 ;
        RECT 44.300 127.305 44.560 127.785 ;
        RECT 44.730 127.135 44.990 127.590 ;
        RECT 45.160 127.305 45.420 127.785 ;
        RECT 45.590 127.135 45.850 127.590 ;
        RECT 46.020 127.225 46.280 127.785 ;
        RECT 37.485 125.915 37.655 127.045 ;
        RECT 38.245 126.875 38.415 127.045 ;
        RECT 36.530 125.745 37.655 125.915 ;
        RECT 37.825 126.545 38.020 126.875 ;
        RECT 38.245 126.545 38.500 126.875 ;
        RECT 37.825 125.575 37.995 126.545 ;
        RECT 38.670 126.375 38.840 127.045 ;
        RECT 35.965 125.405 37.995 125.575 ;
        RECT 38.165 125.235 38.335 126.375 ;
        RECT 38.505 125.405 38.840 126.375 ;
        RECT 39.105 126.965 45.850 127.135 ;
        RECT 39.105 126.375 40.270 126.965 ;
        RECT 46.450 126.795 46.700 127.605 ;
        RECT 46.880 127.260 47.140 127.785 ;
        RECT 47.310 126.795 47.560 127.605 ;
        RECT 47.740 127.275 48.045 127.785 ;
        RECT 40.440 126.545 47.560 126.795 ;
        RECT 47.730 126.545 48.045 127.105 ;
        RECT 48.675 127.060 48.965 127.785 ;
        RECT 49.635 126.965 49.865 127.785 ;
        RECT 50.035 126.985 50.365 127.615 ;
        RECT 49.615 126.545 49.945 126.795 ;
        RECT 39.105 126.150 45.850 126.375 ;
        RECT 39.105 125.235 39.375 125.980 ;
        RECT 39.545 125.410 39.835 126.150 ;
        RECT 40.445 126.135 45.850 126.150 ;
        RECT 40.005 125.240 40.260 125.965 ;
        RECT 40.445 125.410 40.705 126.135 ;
        RECT 40.875 125.240 41.120 125.965 ;
        RECT 41.305 125.410 41.565 126.135 ;
        RECT 41.735 125.240 41.980 125.965 ;
        RECT 42.165 125.410 42.425 126.135 ;
        RECT 42.595 125.240 42.840 125.965 ;
        RECT 43.010 125.410 43.270 126.135 ;
        RECT 43.440 125.240 43.700 125.965 ;
        RECT 43.870 125.410 44.130 126.135 ;
        RECT 44.300 125.240 44.560 125.965 ;
        RECT 44.730 125.410 44.990 126.135 ;
        RECT 45.160 125.240 45.420 125.965 ;
        RECT 45.590 125.410 45.850 126.135 ;
        RECT 46.020 125.240 46.280 126.035 ;
        RECT 46.450 125.410 46.700 126.545 ;
        RECT 40.005 125.235 46.280 125.240 ;
        RECT 46.880 125.235 47.140 126.045 ;
        RECT 47.315 125.405 47.560 126.545 ;
        RECT 47.740 125.235 48.035 126.045 ;
        RECT 48.675 125.235 48.965 126.400 ;
        RECT 50.115 126.385 50.365 126.985 ;
        RECT 50.535 126.965 50.745 127.785 ;
        RECT 51.250 126.975 51.495 127.580 ;
        RECT 51.715 127.250 52.225 127.785 ;
        RECT 49.635 125.235 49.865 126.375 ;
        RECT 50.035 125.405 50.365 126.385 ;
        RECT 50.975 126.805 52.205 126.975 ;
        RECT 50.535 125.235 50.745 126.375 ;
        RECT 50.975 125.995 51.315 126.805 ;
        RECT 51.485 126.240 52.235 126.430 ;
        RECT 50.975 125.585 51.490 125.995 ;
        RECT 51.725 125.235 51.895 125.995 ;
        RECT 52.065 125.575 52.235 126.240 ;
        RECT 52.405 126.255 52.595 127.615 ;
        RECT 52.765 127.105 53.040 127.615 ;
        RECT 53.230 127.250 53.760 127.615 ;
        RECT 54.185 127.385 54.515 127.785 ;
        RECT 53.585 127.215 53.760 127.250 ;
        RECT 52.765 126.935 53.045 127.105 ;
        RECT 52.765 126.455 53.040 126.935 ;
        RECT 53.245 126.255 53.415 127.055 ;
        RECT 52.405 126.085 53.415 126.255 ;
        RECT 53.585 127.045 54.515 127.215 ;
        RECT 54.685 127.045 54.940 127.615 ;
        RECT 55.205 127.235 55.375 127.615 ;
        RECT 55.555 127.405 55.885 127.785 ;
        RECT 55.205 127.065 55.870 127.235 ;
        RECT 56.065 127.110 56.325 127.615 ;
        RECT 53.585 125.915 53.755 127.045 ;
        RECT 54.345 126.875 54.515 127.045 ;
        RECT 52.630 125.745 53.755 125.915 ;
        RECT 53.925 126.545 54.120 126.875 ;
        RECT 54.345 126.545 54.600 126.875 ;
        RECT 53.925 125.575 54.095 126.545 ;
        RECT 54.770 126.375 54.940 127.045 ;
        RECT 55.135 126.515 55.465 126.885 ;
        RECT 55.700 126.810 55.870 127.065 ;
        RECT 52.065 125.405 54.095 125.575 ;
        RECT 54.265 125.235 54.435 126.375 ;
        RECT 54.605 125.405 54.940 126.375 ;
        RECT 55.700 126.480 55.985 126.810 ;
        RECT 55.700 126.335 55.870 126.480 ;
        RECT 55.205 126.165 55.870 126.335 ;
        RECT 56.155 126.310 56.325 127.110 ;
        RECT 57.415 127.015 60.925 127.785 ;
        RECT 61.100 127.240 66.445 127.785 ;
        RECT 66.615 127.325 67.175 127.615 ;
        RECT 67.345 127.325 67.595 127.785 ;
        RECT 55.205 125.405 55.375 126.165 ;
        RECT 55.555 125.235 55.885 125.995 ;
        RECT 56.055 125.405 56.325 126.310 ;
        RECT 57.415 126.325 59.105 126.845 ;
        RECT 59.275 126.495 60.925 127.015 ;
        RECT 57.415 125.235 60.925 126.325 ;
        RECT 62.690 125.670 63.040 126.920 ;
        RECT 64.520 126.410 64.860 127.240 ;
        RECT 66.615 125.955 66.865 127.325 ;
        RECT 68.215 127.155 68.545 127.515 ;
        RECT 67.155 126.965 68.545 127.155 ;
        RECT 69.190 126.975 69.435 127.580 ;
        RECT 69.655 127.250 70.165 127.785 ;
        RECT 67.155 126.875 67.325 126.965 ;
        RECT 67.035 126.545 67.325 126.875 ;
        RECT 68.915 126.805 70.145 126.975 ;
        RECT 67.495 126.545 67.835 126.795 ;
        RECT 68.055 126.545 68.730 126.795 ;
        RECT 67.155 126.295 67.325 126.545 ;
        RECT 67.155 126.125 68.095 126.295 ;
        RECT 68.465 126.185 68.730 126.545 ;
        RECT 61.100 125.235 66.445 125.670 ;
        RECT 66.615 125.405 67.075 125.955 ;
        RECT 67.265 125.235 67.595 125.955 ;
        RECT 67.795 125.575 68.095 126.125 ;
        RECT 68.915 125.995 69.255 126.805 ;
        RECT 69.425 126.240 70.175 126.430 ;
        RECT 68.265 125.235 68.545 125.905 ;
        RECT 68.915 125.585 69.430 125.995 ;
        RECT 69.665 125.235 69.835 125.995 ;
        RECT 70.005 125.575 70.175 126.240 ;
        RECT 70.345 126.255 70.535 127.615 ;
        RECT 70.705 127.105 70.980 127.615 ;
        RECT 71.170 127.250 71.700 127.615 ;
        RECT 72.125 127.385 72.455 127.785 ;
        RECT 71.525 127.215 71.700 127.250 ;
        RECT 70.705 126.935 70.985 127.105 ;
        RECT 70.705 126.455 70.980 126.935 ;
        RECT 71.185 126.255 71.355 127.055 ;
        RECT 70.345 126.085 71.355 126.255 ;
        RECT 71.525 127.045 72.455 127.215 ;
        RECT 72.625 127.045 72.880 127.615 ;
        RECT 71.525 125.915 71.695 127.045 ;
        RECT 72.285 126.875 72.455 127.045 ;
        RECT 70.570 125.745 71.695 125.915 ;
        RECT 71.865 126.545 72.060 126.875 ;
        RECT 72.285 126.545 72.540 126.875 ;
        RECT 71.865 125.575 72.035 126.545 ;
        RECT 72.710 126.375 72.880 127.045 ;
        RECT 73.055 127.035 74.265 127.785 ;
        RECT 74.435 127.060 74.725 127.785 ;
        RECT 74.985 127.305 75.285 127.785 ;
        RECT 75.455 127.135 75.715 127.590 ;
        RECT 75.885 127.305 76.145 127.785 ;
        RECT 76.325 127.135 76.585 127.590 ;
        RECT 76.755 127.305 77.005 127.785 ;
        RECT 77.185 127.135 77.445 127.590 ;
        RECT 77.615 127.305 77.865 127.785 ;
        RECT 78.045 127.135 78.305 127.590 ;
        RECT 78.475 127.305 78.720 127.785 ;
        RECT 78.890 127.135 79.165 127.590 ;
        RECT 79.335 127.305 79.580 127.785 ;
        RECT 79.750 127.135 80.010 127.590 ;
        RECT 80.180 127.305 80.440 127.785 ;
        RECT 80.610 127.135 80.870 127.590 ;
        RECT 81.040 127.305 81.300 127.785 ;
        RECT 81.470 127.135 81.730 127.590 ;
        RECT 81.900 127.225 82.160 127.785 ;
        RECT 70.005 125.405 72.035 125.575 ;
        RECT 72.205 125.235 72.375 126.375 ;
        RECT 72.545 125.405 72.880 126.375 ;
        RECT 73.055 126.325 73.575 126.865 ;
        RECT 73.745 126.495 74.265 127.035 ;
        RECT 74.985 126.965 81.730 127.135 ;
        RECT 73.055 125.235 74.265 126.325 ;
        RECT 74.435 125.235 74.725 126.400 ;
        RECT 74.985 126.375 76.150 126.965 ;
        RECT 82.330 126.795 82.580 127.605 ;
        RECT 82.760 127.260 83.020 127.785 ;
        RECT 83.190 126.795 83.440 127.605 ;
        RECT 83.620 127.275 83.925 127.785 ;
        RECT 76.320 126.545 83.440 126.795 ;
        RECT 83.610 126.545 83.925 127.105 ;
        RECT 84.095 127.015 85.765 127.785 ;
        RECT 74.985 126.150 81.730 126.375 ;
        RECT 74.985 125.235 75.255 125.980 ;
        RECT 75.425 125.410 75.715 126.150 ;
        RECT 76.325 126.135 81.730 126.150 ;
        RECT 75.885 125.240 76.140 125.965 ;
        RECT 76.325 125.410 76.585 126.135 ;
        RECT 76.755 125.240 77.000 125.965 ;
        RECT 77.185 125.410 77.445 126.135 ;
        RECT 77.615 125.240 77.860 125.965 ;
        RECT 78.045 125.410 78.305 126.135 ;
        RECT 78.475 125.240 78.720 125.965 ;
        RECT 78.890 125.410 79.150 126.135 ;
        RECT 79.320 125.240 79.580 125.965 ;
        RECT 79.750 125.410 80.010 126.135 ;
        RECT 80.180 125.240 80.440 125.965 ;
        RECT 80.610 125.410 80.870 126.135 ;
        RECT 81.040 125.240 81.300 125.965 ;
        RECT 81.470 125.410 81.730 126.135 ;
        RECT 81.900 125.240 82.160 126.035 ;
        RECT 82.330 125.410 82.580 126.545 ;
        RECT 75.885 125.235 82.160 125.240 ;
        RECT 82.760 125.235 83.020 126.045 ;
        RECT 83.195 125.405 83.440 126.545 ;
        RECT 84.095 126.325 84.845 126.845 ;
        RECT 85.015 126.495 85.765 127.015 ;
        RECT 86.210 126.975 86.455 127.580 ;
        RECT 86.675 127.250 87.185 127.785 ;
        RECT 85.935 126.805 87.165 126.975 ;
        RECT 83.620 125.235 83.915 126.045 ;
        RECT 84.095 125.235 85.765 126.325 ;
        RECT 85.935 125.995 86.275 126.805 ;
        RECT 86.445 126.240 87.195 126.430 ;
        RECT 85.935 125.585 86.450 125.995 ;
        RECT 86.685 125.235 86.855 125.995 ;
        RECT 87.025 125.575 87.195 126.240 ;
        RECT 87.365 126.255 87.555 127.615 ;
        RECT 87.725 126.765 88.000 127.615 ;
        RECT 88.190 127.250 88.720 127.615 ;
        RECT 89.145 127.385 89.475 127.785 ;
        RECT 88.545 127.215 88.720 127.250 ;
        RECT 87.725 126.595 88.005 126.765 ;
        RECT 87.725 126.455 88.000 126.595 ;
        RECT 88.205 126.255 88.375 127.055 ;
        RECT 87.365 126.085 88.375 126.255 ;
        RECT 88.545 127.045 89.475 127.215 ;
        RECT 89.645 127.045 89.900 127.615 ;
        RECT 88.545 125.915 88.715 127.045 ;
        RECT 89.305 126.875 89.475 127.045 ;
        RECT 87.590 125.745 88.715 125.915 ;
        RECT 88.885 126.545 89.080 126.875 ;
        RECT 89.305 126.545 89.560 126.875 ;
        RECT 88.885 125.575 89.055 126.545 ;
        RECT 89.730 126.375 89.900 127.045 ;
        RECT 90.115 126.965 90.345 127.785 ;
        RECT 90.515 126.985 90.845 127.615 ;
        RECT 90.095 126.545 90.425 126.795 ;
        RECT 90.595 126.385 90.845 126.985 ;
        RECT 91.015 126.965 91.225 127.785 ;
        RECT 91.655 127.155 91.985 127.515 ;
        RECT 92.605 127.325 92.855 127.785 ;
        RECT 93.025 127.325 93.585 127.615 ;
        RECT 91.655 126.965 93.045 127.155 ;
        RECT 92.875 126.875 93.045 126.965 ;
        RECT 87.025 125.405 89.055 125.575 ;
        RECT 89.225 125.235 89.395 126.375 ;
        RECT 89.565 125.405 89.900 126.375 ;
        RECT 90.115 125.235 90.345 126.375 ;
        RECT 90.515 125.405 90.845 126.385 ;
        RECT 91.470 126.545 92.145 126.795 ;
        RECT 92.365 126.545 92.705 126.795 ;
        RECT 92.875 126.545 93.165 126.875 ;
        RECT 91.015 125.235 91.225 126.375 ;
        RECT 91.470 126.185 91.735 126.545 ;
        RECT 92.875 126.295 93.045 126.545 ;
        RECT 92.105 126.125 93.045 126.295 ;
        RECT 91.655 125.235 91.935 125.905 ;
        RECT 92.105 125.575 92.405 126.125 ;
        RECT 93.335 125.955 93.585 127.325 ;
        RECT 94.030 126.975 94.275 127.580 ;
        RECT 94.495 127.250 95.005 127.785 ;
        RECT 92.605 125.235 92.935 125.955 ;
        RECT 93.125 125.405 93.585 125.955 ;
        RECT 93.755 126.805 94.985 126.975 ;
        RECT 93.755 125.995 94.095 126.805 ;
        RECT 94.265 126.240 95.015 126.430 ;
        RECT 93.755 125.585 94.270 125.995 ;
        RECT 94.505 125.235 94.675 125.995 ;
        RECT 94.845 125.575 95.015 126.240 ;
        RECT 95.185 126.255 95.375 127.615 ;
        RECT 95.545 126.765 95.820 127.615 ;
        RECT 96.010 127.250 96.540 127.615 ;
        RECT 96.965 127.385 97.295 127.785 ;
        RECT 96.365 127.215 96.540 127.250 ;
        RECT 95.545 126.595 95.825 126.765 ;
        RECT 95.545 126.455 95.820 126.595 ;
        RECT 96.025 126.255 96.195 127.055 ;
        RECT 95.185 126.085 96.195 126.255 ;
        RECT 96.365 127.045 97.295 127.215 ;
        RECT 97.465 127.045 97.720 127.615 ;
        RECT 96.365 125.915 96.535 127.045 ;
        RECT 97.125 126.875 97.295 127.045 ;
        RECT 95.410 125.745 96.535 125.915 ;
        RECT 96.705 126.545 96.900 126.875 ;
        RECT 97.125 126.545 97.380 126.875 ;
        RECT 96.705 125.575 96.875 126.545 ;
        RECT 97.550 126.375 97.720 127.045 ;
        RECT 98.855 126.965 99.085 127.785 ;
        RECT 99.255 126.985 99.585 127.615 ;
        RECT 98.835 126.545 99.165 126.795 ;
        RECT 99.335 126.385 99.585 126.985 ;
        RECT 99.755 126.965 99.965 127.785 ;
        RECT 100.195 127.060 100.485 127.785 ;
        RECT 101.490 127.075 101.745 127.605 ;
        RECT 101.925 127.325 102.210 127.785 ;
        RECT 94.845 125.405 96.875 125.575 ;
        RECT 97.045 125.235 97.215 126.375 ;
        RECT 97.385 125.405 97.720 126.375 ;
        RECT 98.855 125.235 99.085 126.375 ;
        RECT 99.255 125.405 99.585 126.385 ;
        RECT 99.755 125.235 99.965 126.375 ;
        RECT 100.195 125.235 100.485 126.400 ;
        RECT 101.490 126.215 101.670 127.075 ;
        RECT 102.390 126.875 102.640 127.525 ;
        RECT 101.840 126.545 102.640 126.875 ;
        RECT 101.490 125.745 101.745 126.215 ;
        RECT 101.405 125.575 101.745 125.745 ;
        RECT 101.490 125.545 101.745 125.575 ;
        RECT 101.925 125.235 102.210 126.035 ;
        RECT 102.390 125.955 102.640 126.545 ;
        RECT 102.840 127.190 103.160 127.520 ;
        RECT 103.340 127.305 104.000 127.785 ;
        RECT 104.200 127.395 105.050 127.565 ;
        RECT 102.840 126.295 103.030 127.190 ;
        RECT 103.350 126.865 104.010 127.135 ;
        RECT 103.680 126.805 104.010 126.865 ;
        RECT 103.200 126.635 103.530 126.695 ;
        RECT 104.200 126.635 104.370 127.395 ;
        RECT 105.610 127.325 105.930 127.785 ;
        RECT 106.130 127.145 106.380 127.575 ;
        RECT 106.670 127.345 107.080 127.785 ;
        RECT 107.250 127.405 108.265 127.605 ;
        RECT 104.540 126.975 105.790 127.145 ;
        RECT 104.540 126.855 104.870 126.975 ;
        RECT 103.200 126.465 105.100 126.635 ;
        RECT 102.840 126.125 104.760 126.295 ;
        RECT 102.840 126.105 103.160 126.125 ;
        RECT 102.390 125.445 102.720 125.955 ;
        RECT 102.990 125.495 103.160 126.105 ;
        RECT 104.930 125.955 105.100 126.465 ;
        RECT 105.270 126.395 105.450 126.805 ;
        RECT 105.620 126.215 105.790 126.975 ;
        RECT 103.330 125.235 103.660 125.925 ;
        RECT 103.890 125.785 105.100 125.955 ;
        RECT 105.270 125.905 105.790 126.215 ;
        RECT 105.960 126.805 106.380 127.145 ;
        RECT 106.670 126.805 107.080 127.135 ;
        RECT 105.960 126.035 106.150 126.805 ;
        RECT 107.250 126.675 107.420 127.405 ;
        RECT 108.565 127.235 108.735 127.565 ;
        RECT 108.905 127.405 109.235 127.785 ;
        RECT 107.590 126.855 107.940 127.225 ;
        RECT 107.250 126.635 107.670 126.675 ;
        RECT 106.320 126.465 107.670 126.635 ;
        RECT 106.320 126.305 106.570 126.465 ;
        RECT 107.080 126.035 107.330 126.295 ;
        RECT 105.960 125.785 107.330 126.035 ;
        RECT 103.890 125.495 104.130 125.785 ;
        RECT 104.930 125.705 105.100 125.785 ;
        RECT 104.330 125.235 104.750 125.615 ;
        RECT 104.930 125.455 105.560 125.705 ;
        RECT 106.030 125.235 106.360 125.615 ;
        RECT 106.530 125.495 106.700 125.785 ;
        RECT 107.500 125.620 107.670 126.465 ;
        RECT 108.120 126.295 108.340 127.165 ;
        RECT 108.565 127.045 109.260 127.235 ;
        RECT 107.840 125.915 108.340 126.295 ;
        RECT 108.510 126.245 108.920 126.865 ;
        RECT 109.090 126.075 109.260 127.045 ;
        RECT 108.565 125.905 109.260 126.075 ;
        RECT 106.880 125.235 107.260 125.615 ;
        RECT 107.500 125.450 108.330 125.620 ;
        RECT 108.565 125.405 108.735 125.905 ;
        RECT 108.905 125.235 109.235 125.735 ;
        RECT 109.450 125.405 109.675 127.525 ;
        RECT 109.845 127.405 110.175 127.785 ;
        RECT 110.345 127.235 110.515 127.525 ;
        RECT 109.850 127.065 110.515 127.235 ;
        RECT 109.850 126.075 110.080 127.065 ;
        RECT 110.775 127.035 111.985 127.785 ;
        RECT 112.155 127.035 113.365 127.785 ;
        RECT 110.250 126.245 110.600 126.895 ;
        RECT 110.775 126.325 111.295 126.865 ;
        RECT 111.465 126.495 111.985 127.035 ;
        RECT 112.155 126.325 112.675 126.865 ;
        RECT 112.845 126.495 113.365 127.035 ;
        RECT 109.850 125.905 110.515 126.075 ;
        RECT 109.845 125.235 110.175 125.735 ;
        RECT 110.345 125.405 110.515 125.905 ;
        RECT 110.775 125.235 111.985 126.325 ;
        RECT 112.155 125.235 113.365 126.325 ;
        RECT 11.330 125.065 113.450 125.235 ;
        RECT 11.415 123.975 12.625 125.065 ;
        RECT 13.630 124.725 13.885 124.755 ;
        RECT 13.545 124.555 13.885 124.725 ;
        RECT 11.415 123.265 11.935 123.805 ;
        RECT 12.105 123.435 12.625 123.975 ;
        RECT 13.630 124.085 13.885 124.555 ;
        RECT 14.065 124.265 14.350 125.065 ;
        RECT 14.530 124.345 14.860 124.855 ;
        RECT 11.415 122.515 12.625 123.265 ;
        RECT 13.630 123.225 13.810 124.085 ;
        RECT 14.530 123.755 14.780 124.345 ;
        RECT 15.130 124.195 15.300 124.805 ;
        RECT 15.470 124.375 15.800 125.065 ;
        RECT 16.030 124.515 16.270 124.805 ;
        RECT 16.470 124.685 16.890 125.065 ;
        RECT 17.070 124.595 17.700 124.845 ;
        RECT 18.170 124.685 18.500 125.065 ;
        RECT 17.070 124.515 17.240 124.595 ;
        RECT 18.670 124.515 18.840 124.805 ;
        RECT 19.020 124.685 19.400 125.065 ;
        RECT 19.640 124.680 20.470 124.850 ;
        RECT 16.030 124.345 17.240 124.515 ;
        RECT 13.980 123.425 14.780 123.755 ;
        RECT 13.630 122.695 13.885 123.225 ;
        RECT 14.065 122.515 14.350 122.975 ;
        RECT 14.530 122.775 14.780 123.425 ;
        RECT 14.980 124.175 15.300 124.195 ;
        RECT 14.980 124.005 16.900 124.175 ;
        RECT 14.980 123.110 15.170 124.005 ;
        RECT 17.070 123.835 17.240 124.345 ;
        RECT 17.410 124.085 17.930 124.395 ;
        RECT 15.340 123.665 17.240 123.835 ;
        RECT 15.340 123.605 15.670 123.665 ;
        RECT 15.820 123.435 16.150 123.495 ;
        RECT 15.490 123.165 16.150 123.435 ;
        RECT 14.980 122.780 15.300 123.110 ;
        RECT 15.480 122.515 16.140 122.995 ;
        RECT 16.340 122.905 16.510 123.665 ;
        RECT 17.410 123.495 17.590 123.905 ;
        RECT 16.680 123.325 17.010 123.445 ;
        RECT 17.760 123.325 17.930 124.085 ;
        RECT 16.680 123.155 17.930 123.325 ;
        RECT 18.100 124.265 19.470 124.515 ;
        RECT 18.100 123.495 18.290 124.265 ;
        RECT 19.220 124.005 19.470 124.265 ;
        RECT 18.460 123.835 18.710 123.995 ;
        RECT 19.640 123.835 19.810 124.680 ;
        RECT 20.705 124.395 20.875 124.895 ;
        RECT 21.045 124.565 21.375 125.065 ;
        RECT 19.980 124.005 20.480 124.385 ;
        RECT 20.705 124.225 21.400 124.395 ;
        RECT 18.460 123.665 19.810 123.835 ;
        RECT 19.390 123.625 19.810 123.665 ;
        RECT 18.100 123.155 18.520 123.495 ;
        RECT 18.810 123.165 19.220 123.495 ;
        RECT 16.340 122.735 17.190 122.905 ;
        RECT 17.750 122.515 18.070 122.975 ;
        RECT 18.270 122.725 18.520 123.155 ;
        RECT 18.810 122.515 19.220 122.955 ;
        RECT 19.390 122.895 19.560 123.625 ;
        RECT 19.730 123.075 20.080 123.445 ;
        RECT 20.260 123.135 20.480 124.005 ;
        RECT 20.650 123.435 21.060 124.055 ;
        RECT 21.230 123.255 21.400 124.225 ;
        RECT 20.705 123.065 21.400 123.255 ;
        RECT 19.390 122.695 20.405 122.895 ;
        RECT 20.705 122.735 20.875 123.065 ;
        RECT 21.045 122.515 21.375 122.895 ;
        RECT 21.590 122.775 21.815 124.895 ;
        RECT 21.985 124.565 22.315 125.065 ;
        RECT 22.485 124.395 22.655 124.895 ;
        RECT 21.990 124.225 22.655 124.395 ;
        RECT 23.925 124.320 24.195 125.065 ;
        RECT 24.825 125.060 31.100 125.065 ;
        RECT 21.990 123.235 22.220 124.225 ;
        RECT 24.365 124.150 24.655 124.890 ;
        RECT 24.825 124.335 25.080 125.060 ;
        RECT 25.265 124.165 25.525 124.890 ;
        RECT 25.695 124.335 25.940 125.060 ;
        RECT 26.125 124.165 26.385 124.890 ;
        RECT 26.555 124.335 26.800 125.060 ;
        RECT 26.985 124.165 27.245 124.890 ;
        RECT 27.415 124.335 27.660 125.060 ;
        RECT 27.830 124.165 28.090 124.890 ;
        RECT 28.260 124.335 28.520 125.060 ;
        RECT 28.690 124.165 28.950 124.890 ;
        RECT 29.120 124.335 29.380 125.060 ;
        RECT 29.550 124.165 29.810 124.890 ;
        RECT 29.980 124.335 30.240 125.060 ;
        RECT 30.410 124.165 30.670 124.890 ;
        RECT 30.840 124.265 31.100 125.060 ;
        RECT 25.265 124.150 30.670 124.165 ;
        RECT 22.390 123.405 22.740 124.055 ;
        RECT 23.925 123.925 30.670 124.150 ;
        RECT 23.925 123.335 25.090 123.925 ;
        RECT 31.270 123.755 31.520 124.890 ;
        RECT 31.700 124.255 31.960 125.065 ;
        RECT 32.135 123.755 32.380 124.895 ;
        RECT 32.560 124.255 32.855 125.065 ;
        RECT 33.695 124.395 33.975 125.065 ;
        RECT 34.145 124.175 34.445 124.725 ;
        RECT 34.645 124.345 34.975 125.065 ;
        RECT 35.165 124.345 35.625 124.895 ;
        RECT 33.510 123.755 33.775 124.115 ;
        RECT 34.145 124.005 35.085 124.175 ;
        RECT 34.915 123.755 35.085 124.005 ;
        RECT 25.260 123.505 32.380 123.755 ;
        RECT 21.990 123.065 22.655 123.235 ;
        RECT 23.925 123.165 30.670 123.335 ;
        RECT 21.985 122.515 22.315 122.895 ;
        RECT 22.485 122.775 22.655 123.065 ;
        RECT 23.925 122.515 24.225 122.995 ;
        RECT 24.395 122.710 24.655 123.165 ;
        RECT 24.825 122.515 25.085 122.995 ;
        RECT 25.265 122.710 25.525 123.165 ;
        RECT 25.695 122.515 25.945 122.995 ;
        RECT 26.125 122.710 26.385 123.165 ;
        RECT 26.555 122.515 26.805 122.995 ;
        RECT 26.985 122.710 27.245 123.165 ;
        RECT 27.415 122.515 27.660 122.995 ;
        RECT 27.830 122.710 28.105 123.165 ;
        RECT 28.275 122.515 28.520 122.995 ;
        RECT 28.690 122.710 28.950 123.165 ;
        RECT 29.120 122.515 29.380 122.995 ;
        RECT 29.550 122.710 29.810 123.165 ;
        RECT 29.980 122.515 30.240 122.995 ;
        RECT 30.410 122.710 30.670 123.165 ;
        RECT 30.840 122.515 31.100 123.075 ;
        RECT 31.270 122.695 31.520 123.505 ;
        RECT 31.700 122.515 31.960 123.040 ;
        RECT 32.130 122.695 32.380 123.505 ;
        RECT 32.550 123.195 32.865 123.755 ;
        RECT 33.510 123.505 34.185 123.755 ;
        RECT 34.405 123.505 34.745 123.755 ;
        RECT 34.915 123.425 35.205 123.755 ;
        RECT 34.915 123.335 35.085 123.425 ;
        RECT 33.695 123.145 35.085 123.335 ;
        RECT 32.560 122.515 32.865 123.025 ;
        RECT 33.695 122.785 34.025 123.145 ;
        RECT 35.375 122.975 35.625 124.345 ;
        RECT 35.795 123.900 36.085 125.065 ;
        RECT 37.285 124.265 37.455 125.065 ;
        RECT 37.625 124.045 37.955 124.895 ;
        RECT 38.125 124.265 38.295 125.065 ;
        RECT 38.465 124.045 38.795 124.895 ;
        RECT 38.965 124.265 39.135 125.065 ;
        RECT 39.305 124.045 39.635 124.895 ;
        RECT 39.805 124.265 39.975 125.065 ;
        RECT 40.145 124.045 40.475 124.895 ;
        RECT 40.645 124.265 40.815 125.065 ;
        RECT 40.985 124.045 41.315 124.895 ;
        RECT 41.485 124.265 41.655 125.065 ;
        RECT 41.825 124.045 42.155 124.895 ;
        RECT 42.325 124.265 42.495 125.065 ;
        RECT 42.665 124.045 42.995 124.895 ;
        RECT 43.165 124.265 43.335 125.065 ;
        RECT 43.505 124.045 43.835 124.895 ;
        RECT 44.005 124.265 44.175 125.065 ;
        RECT 44.345 124.045 44.675 124.895 ;
        RECT 44.845 124.265 45.015 125.065 ;
        RECT 45.185 124.045 45.515 124.895 ;
        RECT 45.685 124.265 45.855 125.065 ;
        RECT 46.025 124.045 46.355 124.895 ;
        RECT 46.525 124.215 46.695 125.065 ;
        RECT 46.865 124.045 47.195 124.895 ;
        RECT 47.365 124.215 47.535 125.065 ;
        RECT 47.705 124.045 48.035 124.895 ;
        RECT 48.590 124.725 48.845 124.755 ;
        RECT 48.505 124.555 48.845 124.725 ;
        RECT 37.175 123.875 43.835 124.045 ;
        RECT 44.005 123.875 46.355 124.045 ;
        RECT 46.525 123.875 48.035 124.045 ;
        RECT 48.590 124.085 48.845 124.555 ;
        RECT 49.025 124.265 49.310 125.065 ;
        RECT 49.490 124.345 49.820 124.855 ;
        RECT 37.175 123.335 37.450 123.875 ;
        RECT 44.005 123.705 44.180 123.875 ;
        RECT 46.525 123.705 46.695 123.875 ;
        RECT 37.620 123.505 44.180 123.705 ;
        RECT 44.385 123.505 46.695 123.705 ;
        RECT 46.865 123.505 48.040 123.705 ;
        RECT 44.005 123.335 44.180 123.505 ;
        RECT 46.525 123.335 46.695 123.505 ;
        RECT 34.645 122.515 34.895 122.975 ;
        RECT 35.065 122.685 35.625 122.975 ;
        RECT 35.795 122.515 36.085 123.240 ;
        RECT 37.175 123.165 43.835 123.335 ;
        RECT 44.005 123.165 46.355 123.335 ;
        RECT 46.525 123.165 48.035 123.335 ;
        RECT 37.285 122.515 37.455 122.995 ;
        RECT 37.625 122.690 37.955 123.165 ;
        RECT 38.125 122.515 38.295 122.995 ;
        RECT 38.465 122.690 38.795 123.165 ;
        RECT 38.965 122.515 39.135 122.995 ;
        RECT 39.305 122.690 39.635 123.165 ;
        RECT 39.805 122.515 39.975 122.995 ;
        RECT 40.145 122.690 40.475 123.165 ;
        RECT 40.645 122.515 40.815 122.995 ;
        RECT 40.985 122.690 41.315 123.165 ;
        RECT 41.485 122.515 41.655 122.995 ;
        RECT 41.825 122.690 42.155 123.165 ;
        RECT 41.905 122.685 42.075 122.690 ;
        RECT 42.325 122.515 42.495 122.995 ;
        RECT 42.665 122.690 42.995 123.165 ;
        RECT 42.745 122.685 42.915 122.690 ;
        RECT 43.165 122.515 43.335 122.995 ;
        RECT 43.505 122.690 43.835 123.165 ;
        RECT 43.585 122.685 43.835 122.690 ;
        RECT 44.005 122.515 44.175 122.995 ;
        RECT 44.345 122.690 44.675 123.165 ;
        RECT 44.845 122.515 45.015 122.995 ;
        RECT 45.185 122.690 45.515 123.165 ;
        RECT 45.685 122.515 45.855 122.995 ;
        RECT 46.025 122.690 46.355 123.165 ;
        RECT 46.525 122.515 46.695 122.995 ;
        RECT 46.865 122.690 47.195 123.165 ;
        RECT 47.365 122.515 47.535 122.995 ;
        RECT 47.705 122.690 48.035 123.165 ;
        RECT 48.590 123.225 48.770 124.085 ;
        RECT 49.490 123.755 49.740 124.345 ;
        RECT 50.090 124.195 50.260 124.805 ;
        RECT 50.430 124.375 50.760 125.065 ;
        RECT 50.990 124.515 51.230 124.805 ;
        RECT 51.430 124.685 51.850 125.065 ;
        RECT 52.030 124.595 52.660 124.845 ;
        RECT 53.130 124.685 53.460 125.065 ;
        RECT 52.030 124.515 52.200 124.595 ;
        RECT 53.630 124.515 53.800 124.805 ;
        RECT 53.980 124.685 54.360 125.065 ;
        RECT 54.600 124.680 55.430 124.850 ;
        RECT 50.990 124.345 52.200 124.515 ;
        RECT 48.940 123.425 49.740 123.755 ;
        RECT 48.590 122.695 48.845 123.225 ;
        RECT 49.025 122.515 49.310 122.975 ;
        RECT 49.490 122.775 49.740 123.425 ;
        RECT 49.940 124.175 50.260 124.195 ;
        RECT 49.940 124.005 51.860 124.175 ;
        RECT 49.940 123.110 50.130 124.005 ;
        RECT 52.030 123.835 52.200 124.345 ;
        RECT 52.370 124.085 52.890 124.395 ;
        RECT 50.300 123.665 52.200 123.835 ;
        RECT 50.300 123.605 50.630 123.665 ;
        RECT 50.780 123.435 51.110 123.495 ;
        RECT 50.450 123.165 51.110 123.435 ;
        RECT 49.940 122.780 50.260 123.110 ;
        RECT 50.440 122.515 51.100 122.995 ;
        RECT 51.300 122.905 51.470 123.665 ;
        RECT 52.370 123.495 52.550 123.905 ;
        RECT 51.640 123.325 51.970 123.445 ;
        RECT 52.720 123.325 52.890 124.085 ;
        RECT 51.640 123.155 52.890 123.325 ;
        RECT 53.060 124.265 54.430 124.515 ;
        RECT 53.060 123.495 53.250 124.265 ;
        RECT 54.180 124.005 54.430 124.265 ;
        RECT 53.420 123.835 53.670 123.995 ;
        RECT 54.600 123.835 54.770 124.680 ;
        RECT 55.665 124.395 55.835 124.895 ;
        RECT 56.005 124.565 56.335 125.065 ;
        RECT 54.940 124.005 55.440 124.385 ;
        RECT 55.665 124.225 56.360 124.395 ;
        RECT 53.420 123.665 54.770 123.835 ;
        RECT 54.350 123.625 54.770 123.665 ;
        RECT 53.060 123.155 53.480 123.495 ;
        RECT 53.770 123.165 54.180 123.495 ;
        RECT 51.300 122.735 52.150 122.905 ;
        RECT 52.710 122.515 53.030 122.975 ;
        RECT 53.230 122.725 53.480 123.155 ;
        RECT 53.770 122.515 54.180 122.955 ;
        RECT 54.350 122.895 54.520 123.625 ;
        RECT 54.690 123.075 55.040 123.445 ;
        RECT 55.220 123.135 55.440 124.005 ;
        RECT 55.610 123.435 56.020 124.055 ;
        RECT 56.190 123.255 56.360 124.225 ;
        RECT 55.665 123.065 56.360 123.255 ;
        RECT 54.350 122.695 55.365 122.895 ;
        RECT 55.665 122.735 55.835 123.065 ;
        RECT 56.005 122.515 56.335 122.895 ;
        RECT 56.550 122.775 56.775 124.895 ;
        RECT 56.945 124.565 57.275 125.065 ;
        RECT 57.445 124.395 57.615 124.895 ;
        RECT 56.950 124.225 57.615 124.395 ;
        RECT 56.950 123.235 57.180 124.225 ;
        RECT 57.350 123.405 57.700 124.055 ;
        RECT 57.875 123.975 61.385 125.065 ;
        RECT 57.875 123.455 59.565 123.975 ;
        RECT 61.555 123.900 61.845 125.065 ;
        RECT 62.015 123.975 64.605 125.065 ;
        RECT 59.735 123.285 61.385 123.805 ;
        RECT 62.015 123.455 63.225 123.975 ;
        RECT 64.815 123.925 65.045 125.065 ;
        RECT 65.215 123.915 65.545 124.895 ;
        RECT 65.715 123.925 65.925 125.065 ;
        RECT 66.155 124.305 66.670 124.715 ;
        RECT 66.905 124.305 67.075 125.065 ;
        RECT 67.245 124.725 69.275 124.895 ;
        RECT 63.395 123.285 64.605 123.805 ;
        RECT 64.795 123.505 65.125 123.755 ;
        RECT 56.950 123.065 57.615 123.235 ;
        RECT 56.945 122.515 57.275 122.895 ;
        RECT 57.445 122.775 57.615 123.065 ;
        RECT 57.875 122.515 61.385 123.285 ;
        RECT 61.555 122.515 61.845 123.240 ;
        RECT 62.015 122.515 64.605 123.285 ;
        RECT 64.815 122.515 65.045 123.335 ;
        RECT 65.295 123.315 65.545 123.915 ;
        RECT 66.155 123.495 66.495 124.305 ;
        RECT 67.245 124.060 67.415 124.725 ;
        RECT 67.810 124.385 68.935 124.555 ;
        RECT 66.665 123.870 67.415 124.060 ;
        RECT 67.585 124.045 68.595 124.215 ;
        RECT 65.215 122.685 65.545 123.315 ;
        RECT 65.715 122.515 65.925 123.335 ;
        RECT 66.155 123.325 67.385 123.495 ;
        RECT 66.430 122.720 66.675 123.325 ;
        RECT 66.895 122.515 67.405 123.050 ;
        RECT 67.585 122.685 67.775 124.045 ;
        RECT 67.945 123.025 68.220 123.845 ;
        RECT 68.425 123.245 68.595 124.045 ;
        RECT 68.765 123.255 68.935 124.385 ;
        RECT 69.105 123.755 69.275 124.725 ;
        RECT 69.445 123.925 69.615 125.065 ;
        RECT 69.785 123.925 70.120 124.895 ;
        RECT 69.105 123.425 69.300 123.755 ;
        RECT 69.525 123.425 69.780 123.755 ;
        RECT 69.525 123.255 69.695 123.425 ;
        RECT 69.950 123.255 70.120 123.925 ;
        RECT 70.295 123.975 71.965 125.065 ;
        RECT 72.510 124.725 72.765 124.755 ;
        RECT 72.425 124.555 72.765 124.725 ;
        RECT 72.510 124.085 72.765 124.555 ;
        RECT 72.945 124.265 73.230 125.065 ;
        RECT 73.410 124.345 73.740 124.855 ;
        RECT 70.295 123.455 71.045 123.975 ;
        RECT 71.215 123.285 71.965 123.805 ;
        RECT 68.765 123.085 69.695 123.255 ;
        RECT 68.765 123.050 68.940 123.085 ;
        RECT 67.945 122.855 68.225 123.025 ;
        RECT 67.945 122.685 68.220 122.855 ;
        RECT 68.410 122.685 68.940 123.050 ;
        RECT 69.365 122.515 69.695 122.915 ;
        RECT 69.865 122.685 70.120 123.255 ;
        RECT 70.295 122.515 71.965 123.285 ;
        RECT 72.510 123.225 72.690 124.085 ;
        RECT 73.410 123.755 73.660 124.345 ;
        RECT 74.010 124.195 74.180 124.805 ;
        RECT 74.350 124.375 74.680 125.065 ;
        RECT 74.910 124.515 75.150 124.805 ;
        RECT 75.350 124.685 75.770 125.065 ;
        RECT 75.950 124.595 76.580 124.845 ;
        RECT 77.050 124.685 77.380 125.065 ;
        RECT 75.950 124.515 76.120 124.595 ;
        RECT 77.550 124.515 77.720 124.805 ;
        RECT 77.900 124.685 78.280 125.065 ;
        RECT 78.520 124.680 79.350 124.850 ;
        RECT 74.910 124.345 76.120 124.515 ;
        RECT 72.860 123.425 73.660 123.755 ;
        RECT 72.510 122.695 72.765 123.225 ;
        RECT 72.945 122.515 73.230 122.975 ;
        RECT 73.410 122.775 73.660 123.425 ;
        RECT 73.860 124.175 74.180 124.195 ;
        RECT 73.860 124.005 75.780 124.175 ;
        RECT 73.860 123.110 74.050 124.005 ;
        RECT 75.950 123.835 76.120 124.345 ;
        RECT 76.290 124.085 76.810 124.395 ;
        RECT 74.220 123.665 76.120 123.835 ;
        RECT 74.220 123.605 74.550 123.665 ;
        RECT 74.700 123.435 75.030 123.495 ;
        RECT 74.370 123.165 75.030 123.435 ;
        RECT 73.860 122.780 74.180 123.110 ;
        RECT 74.360 122.515 75.020 122.995 ;
        RECT 75.220 122.905 75.390 123.665 ;
        RECT 76.290 123.495 76.470 123.905 ;
        RECT 75.560 123.325 75.890 123.445 ;
        RECT 76.640 123.325 76.810 124.085 ;
        RECT 75.560 123.155 76.810 123.325 ;
        RECT 76.980 124.265 78.350 124.515 ;
        RECT 76.980 123.495 77.170 124.265 ;
        RECT 78.100 124.005 78.350 124.265 ;
        RECT 77.340 123.835 77.590 123.995 ;
        RECT 78.520 123.835 78.690 124.680 ;
        RECT 79.585 124.395 79.755 124.895 ;
        RECT 79.925 124.565 80.255 125.065 ;
        RECT 78.860 124.005 79.360 124.385 ;
        RECT 79.585 124.225 80.280 124.395 ;
        RECT 77.340 123.665 78.690 123.835 ;
        RECT 78.270 123.625 78.690 123.665 ;
        RECT 76.980 123.155 77.400 123.495 ;
        RECT 77.690 123.165 78.100 123.495 ;
        RECT 75.220 122.735 76.070 122.905 ;
        RECT 76.630 122.515 76.950 122.975 ;
        RECT 77.150 122.725 77.400 123.155 ;
        RECT 77.690 122.515 78.100 122.955 ;
        RECT 78.270 122.895 78.440 123.625 ;
        RECT 78.610 123.075 78.960 123.445 ;
        RECT 79.140 123.135 79.360 124.005 ;
        RECT 79.530 123.435 79.940 124.055 ;
        RECT 80.110 123.255 80.280 124.225 ;
        RECT 79.585 123.065 80.280 123.255 ;
        RECT 78.270 122.695 79.285 122.895 ;
        RECT 79.585 122.735 79.755 123.065 ;
        RECT 79.925 122.515 80.255 122.895 ;
        RECT 80.470 122.775 80.695 124.895 ;
        RECT 80.865 124.565 81.195 125.065 ;
        RECT 81.365 124.395 81.535 124.895 ;
        RECT 80.870 124.225 81.535 124.395 ;
        RECT 81.795 124.305 82.310 124.715 ;
        RECT 82.545 124.305 82.715 125.065 ;
        RECT 82.885 124.725 84.915 124.895 ;
        RECT 80.870 123.235 81.100 124.225 ;
        RECT 81.270 123.405 81.620 124.055 ;
        RECT 81.795 123.495 82.135 124.305 ;
        RECT 82.885 124.060 83.055 124.725 ;
        RECT 83.450 124.385 84.575 124.555 ;
        RECT 82.305 123.870 83.055 124.060 ;
        RECT 83.225 124.045 84.235 124.215 ;
        RECT 81.795 123.325 83.025 123.495 ;
        RECT 80.870 123.065 81.535 123.235 ;
        RECT 80.865 122.515 81.195 122.895 ;
        RECT 81.365 122.775 81.535 123.065 ;
        RECT 82.070 122.720 82.315 123.325 ;
        RECT 82.535 122.515 83.045 123.050 ;
        RECT 83.225 122.685 83.415 124.045 ;
        RECT 83.585 123.365 83.860 123.845 ;
        RECT 83.585 123.195 83.865 123.365 ;
        RECT 84.065 123.245 84.235 124.045 ;
        RECT 84.405 123.255 84.575 124.385 ;
        RECT 84.745 123.755 84.915 124.725 ;
        RECT 85.085 123.925 85.255 125.065 ;
        RECT 85.425 123.925 85.760 124.895 ;
        RECT 84.745 123.425 84.940 123.755 ;
        RECT 85.165 123.425 85.420 123.755 ;
        RECT 85.165 123.255 85.335 123.425 ;
        RECT 85.590 123.255 85.760 123.925 ;
        RECT 85.935 123.975 87.145 125.065 ;
        RECT 85.935 123.435 86.455 123.975 ;
        RECT 87.315 123.900 87.605 125.065 ;
        RECT 88.610 124.725 88.865 124.755 ;
        RECT 88.525 124.555 88.865 124.725 ;
        RECT 88.610 124.085 88.865 124.555 ;
        RECT 89.045 124.265 89.330 125.065 ;
        RECT 89.510 124.345 89.840 124.855 ;
        RECT 86.625 123.265 87.145 123.805 ;
        RECT 83.585 122.685 83.860 123.195 ;
        RECT 84.405 123.085 85.335 123.255 ;
        RECT 84.405 123.050 84.580 123.085 ;
        RECT 84.050 122.685 84.580 123.050 ;
        RECT 85.005 122.515 85.335 122.915 ;
        RECT 85.505 122.685 85.760 123.255 ;
        RECT 85.935 122.515 87.145 123.265 ;
        RECT 87.315 122.515 87.605 123.240 ;
        RECT 88.610 123.225 88.790 124.085 ;
        RECT 89.510 123.755 89.760 124.345 ;
        RECT 90.110 124.195 90.280 124.805 ;
        RECT 90.450 124.375 90.780 125.065 ;
        RECT 91.010 124.515 91.250 124.805 ;
        RECT 91.450 124.685 91.870 125.065 ;
        RECT 92.050 124.595 92.680 124.845 ;
        RECT 93.150 124.685 93.480 125.065 ;
        RECT 92.050 124.515 92.220 124.595 ;
        RECT 93.650 124.515 93.820 124.805 ;
        RECT 94.000 124.685 94.380 125.065 ;
        RECT 94.620 124.680 95.450 124.850 ;
        RECT 91.010 124.345 92.220 124.515 ;
        RECT 88.960 123.425 89.760 123.755 ;
        RECT 88.610 122.695 88.865 123.225 ;
        RECT 89.045 122.515 89.330 122.975 ;
        RECT 89.510 122.775 89.760 123.425 ;
        RECT 89.960 124.175 90.280 124.195 ;
        RECT 89.960 124.005 91.880 124.175 ;
        RECT 89.960 123.110 90.150 124.005 ;
        RECT 92.050 123.835 92.220 124.345 ;
        RECT 92.390 124.085 92.910 124.395 ;
        RECT 90.320 123.665 92.220 123.835 ;
        RECT 90.320 123.605 90.650 123.665 ;
        RECT 90.800 123.435 91.130 123.495 ;
        RECT 90.470 123.165 91.130 123.435 ;
        RECT 89.960 122.780 90.280 123.110 ;
        RECT 90.460 122.515 91.120 122.995 ;
        RECT 91.320 122.905 91.490 123.665 ;
        RECT 92.390 123.495 92.570 123.905 ;
        RECT 91.660 123.325 91.990 123.445 ;
        RECT 92.740 123.325 92.910 124.085 ;
        RECT 91.660 123.155 92.910 123.325 ;
        RECT 93.080 124.265 94.450 124.515 ;
        RECT 93.080 123.495 93.270 124.265 ;
        RECT 94.200 124.005 94.450 124.265 ;
        RECT 93.440 123.835 93.690 123.995 ;
        RECT 94.620 123.835 94.790 124.680 ;
        RECT 95.685 124.395 95.855 124.895 ;
        RECT 96.025 124.565 96.355 125.065 ;
        RECT 94.960 124.005 95.460 124.385 ;
        RECT 95.685 124.225 96.380 124.395 ;
        RECT 93.440 123.665 94.790 123.835 ;
        RECT 94.370 123.625 94.790 123.665 ;
        RECT 93.080 123.155 93.500 123.495 ;
        RECT 93.790 123.165 94.200 123.495 ;
        RECT 91.320 122.735 92.170 122.905 ;
        RECT 92.730 122.515 93.050 122.975 ;
        RECT 93.250 122.725 93.500 123.155 ;
        RECT 93.790 122.515 94.200 122.955 ;
        RECT 94.370 122.895 94.540 123.625 ;
        RECT 94.710 123.075 95.060 123.445 ;
        RECT 95.240 123.135 95.460 124.005 ;
        RECT 95.630 123.435 96.040 124.055 ;
        RECT 96.210 123.255 96.380 124.225 ;
        RECT 95.685 123.065 96.380 123.255 ;
        RECT 94.370 122.695 95.385 122.895 ;
        RECT 95.685 122.735 95.855 123.065 ;
        RECT 96.025 122.515 96.355 122.895 ;
        RECT 96.570 122.775 96.795 124.895 ;
        RECT 96.965 124.565 97.295 125.065 ;
        RECT 97.465 124.395 97.635 124.895 ;
        RECT 96.970 124.225 97.635 124.395 ;
        RECT 96.970 123.235 97.200 124.225 ;
        RECT 97.370 123.405 97.720 124.055 ;
        RECT 97.895 123.990 98.165 124.895 ;
        RECT 98.335 124.305 98.665 125.065 ;
        RECT 98.845 124.135 99.015 124.895 ;
        RECT 96.970 123.065 97.635 123.235 ;
        RECT 96.965 122.515 97.295 122.895 ;
        RECT 97.465 122.775 97.635 123.065 ;
        RECT 97.895 123.190 98.065 123.990 ;
        RECT 98.350 123.965 99.015 124.135 ;
        RECT 99.275 123.975 100.485 125.065 ;
        RECT 100.655 124.305 101.170 124.715 ;
        RECT 101.405 124.305 101.575 125.065 ;
        RECT 101.745 124.725 103.775 124.895 ;
        RECT 98.350 123.820 98.520 123.965 ;
        RECT 98.235 123.490 98.520 123.820 ;
        RECT 98.350 123.235 98.520 123.490 ;
        RECT 98.755 123.415 99.085 123.785 ;
        RECT 99.275 123.435 99.795 123.975 ;
        RECT 99.965 123.265 100.485 123.805 ;
        RECT 100.655 123.495 100.995 124.305 ;
        RECT 101.745 124.060 101.915 124.725 ;
        RECT 102.310 124.385 103.435 124.555 ;
        RECT 101.165 123.870 101.915 124.060 ;
        RECT 102.085 124.045 103.095 124.215 ;
        RECT 100.655 123.325 101.885 123.495 ;
        RECT 97.895 122.685 98.155 123.190 ;
        RECT 98.350 123.065 99.015 123.235 ;
        RECT 98.335 122.515 98.665 122.895 ;
        RECT 98.845 122.685 99.015 123.065 ;
        RECT 99.275 122.515 100.485 123.265 ;
        RECT 100.930 122.720 101.175 123.325 ;
        RECT 101.395 122.515 101.905 123.050 ;
        RECT 102.085 122.685 102.275 124.045 ;
        RECT 102.445 123.705 102.720 123.845 ;
        RECT 102.445 123.535 102.725 123.705 ;
        RECT 102.445 122.685 102.720 123.535 ;
        RECT 102.925 123.245 103.095 124.045 ;
        RECT 103.265 123.255 103.435 124.385 ;
        RECT 103.605 123.755 103.775 124.725 ;
        RECT 103.945 123.925 104.115 125.065 ;
        RECT 104.285 123.925 104.620 124.895 ;
        RECT 103.605 123.425 103.800 123.755 ;
        RECT 104.025 123.425 104.280 123.755 ;
        RECT 104.025 123.255 104.195 123.425 ;
        RECT 104.450 123.255 104.620 123.925 ;
        RECT 104.795 123.975 106.005 125.065 ;
        RECT 106.265 124.135 106.435 124.895 ;
        RECT 106.615 124.305 106.945 125.065 ;
        RECT 104.795 123.435 105.315 123.975 ;
        RECT 106.265 123.965 106.930 124.135 ;
        RECT 107.115 123.990 107.385 124.895 ;
        RECT 106.760 123.820 106.930 123.965 ;
        RECT 105.485 123.265 106.005 123.805 ;
        RECT 106.195 123.415 106.525 123.785 ;
        RECT 106.760 123.490 107.045 123.820 ;
        RECT 103.265 123.085 104.195 123.255 ;
        RECT 103.265 123.050 103.440 123.085 ;
        RECT 102.910 122.685 103.440 123.050 ;
        RECT 103.865 122.515 104.195 122.915 ;
        RECT 104.365 122.685 104.620 123.255 ;
        RECT 104.795 122.515 106.005 123.265 ;
        RECT 106.760 123.235 106.930 123.490 ;
        RECT 106.265 123.065 106.930 123.235 ;
        RECT 107.215 123.190 107.385 123.990 ;
        RECT 108.475 123.975 111.985 125.065 ;
        RECT 112.155 123.975 113.365 125.065 ;
        RECT 108.475 123.455 110.165 123.975 ;
        RECT 110.335 123.285 111.985 123.805 ;
        RECT 112.155 123.435 112.675 123.975 ;
        RECT 106.265 122.685 106.435 123.065 ;
        RECT 106.615 122.515 106.945 122.895 ;
        RECT 107.125 122.685 107.385 123.190 ;
        RECT 108.475 122.515 111.985 123.285 ;
        RECT 112.845 123.265 113.365 123.805 ;
        RECT 112.155 122.515 113.365 123.265 ;
        RECT 11.330 122.345 113.450 122.515 ;
        RECT 11.415 121.595 12.625 122.345 ;
        RECT 13.170 121.635 13.425 122.165 ;
        RECT 13.605 121.885 13.890 122.345 ;
        RECT 11.415 121.055 11.935 121.595 ;
        RECT 12.105 120.885 12.625 121.425 ;
        RECT 11.415 119.795 12.625 120.885 ;
        RECT 13.170 120.775 13.350 121.635 ;
        RECT 14.070 121.435 14.320 122.085 ;
        RECT 13.520 121.105 14.320 121.435 ;
        RECT 13.170 120.305 13.425 120.775 ;
        RECT 13.085 120.135 13.425 120.305 ;
        RECT 13.170 120.105 13.425 120.135 ;
        RECT 13.605 119.795 13.890 120.595 ;
        RECT 14.070 120.515 14.320 121.105 ;
        RECT 14.520 121.750 14.840 122.080 ;
        RECT 15.020 121.865 15.680 122.345 ;
        RECT 15.880 121.955 16.730 122.125 ;
        RECT 14.520 120.855 14.710 121.750 ;
        RECT 15.030 121.425 15.690 121.695 ;
        RECT 15.360 121.365 15.690 121.425 ;
        RECT 14.880 121.195 15.210 121.255 ;
        RECT 15.880 121.195 16.050 121.955 ;
        RECT 17.290 121.885 17.610 122.345 ;
        RECT 17.810 121.705 18.060 122.135 ;
        RECT 18.350 121.905 18.760 122.345 ;
        RECT 18.930 121.965 19.945 122.165 ;
        RECT 16.220 121.535 17.470 121.705 ;
        RECT 16.220 121.415 16.550 121.535 ;
        RECT 14.880 121.025 16.780 121.195 ;
        RECT 14.520 120.685 16.440 120.855 ;
        RECT 14.520 120.665 14.840 120.685 ;
        RECT 14.070 120.005 14.400 120.515 ;
        RECT 14.670 120.055 14.840 120.665 ;
        RECT 16.610 120.515 16.780 121.025 ;
        RECT 16.950 120.955 17.130 121.365 ;
        RECT 17.300 120.775 17.470 121.535 ;
        RECT 15.010 119.795 15.340 120.485 ;
        RECT 15.570 120.345 16.780 120.515 ;
        RECT 16.950 120.465 17.470 120.775 ;
        RECT 17.640 121.365 18.060 121.705 ;
        RECT 18.350 121.365 18.760 121.695 ;
        RECT 17.640 120.595 17.830 121.365 ;
        RECT 18.930 121.235 19.100 121.965 ;
        RECT 20.245 121.795 20.415 122.125 ;
        RECT 20.585 121.965 20.915 122.345 ;
        RECT 19.270 121.415 19.620 121.785 ;
        RECT 18.930 121.195 19.350 121.235 ;
        RECT 18.000 121.025 19.350 121.195 ;
        RECT 18.000 120.865 18.250 121.025 ;
        RECT 18.760 120.595 19.010 120.855 ;
        RECT 17.640 120.345 19.010 120.595 ;
        RECT 15.570 120.055 15.810 120.345 ;
        RECT 16.610 120.265 16.780 120.345 ;
        RECT 16.010 119.795 16.430 120.175 ;
        RECT 16.610 120.015 17.240 120.265 ;
        RECT 17.710 119.795 18.040 120.175 ;
        RECT 18.210 120.055 18.380 120.345 ;
        RECT 19.180 120.180 19.350 121.025 ;
        RECT 19.800 120.855 20.020 121.725 ;
        RECT 20.245 121.605 20.940 121.795 ;
        RECT 19.520 120.475 20.020 120.855 ;
        RECT 20.190 120.805 20.600 121.425 ;
        RECT 20.770 120.635 20.940 121.605 ;
        RECT 20.245 120.465 20.940 120.635 ;
        RECT 18.560 119.795 18.940 120.175 ;
        RECT 19.180 120.010 20.010 120.180 ;
        RECT 20.245 119.965 20.415 120.465 ;
        RECT 20.585 119.795 20.915 120.295 ;
        RECT 21.130 119.965 21.355 122.085 ;
        RECT 21.525 121.965 21.855 122.345 ;
        RECT 22.025 121.795 22.195 122.085 ;
        RECT 21.530 121.625 22.195 121.795 ;
        RECT 21.530 120.635 21.760 121.625 ;
        RECT 22.915 121.620 23.205 122.345 ;
        RECT 23.465 121.795 23.635 122.085 ;
        RECT 23.805 121.965 24.135 122.345 ;
        RECT 23.465 121.625 24.130 121.795 ;
        RECT 21.930 120.805 22.280 121.455 ;
        RECT 21.530 120.465 22.195 120.635 ;
        RECT 21.525 119.795 21.855 120.295 ;
        RECT 22.025 119.965 22.195 120.465 ;
        RECT 22.915 119.795 23.205 120.960 ;
        RECT 23.380 120.805 23.730 121.455 ;
        RECT 23.900 120.635 24.130 121.625 ;
        RECT 23.465 120.465 24.130 120.635 ;
        RECT 23.465 119.965 23.635 120.465 ;
        RECT 23.805 119.795 24.135 120.295 ;
        RECT 24.305 119.965 24.530 122.085 ;
        RECT 24.745 121.965 25.075 122.345 ;
        RECT 25.245 121.795 25.415 122.125 ;
        RECT 25.715 121.965 26.730 122.165 ;
        RECT 24.720 121.605 25.415 121.795 ;
        RECT 24.720 120.635 24.890 121.605 ;
        RECT 25.060 120.805 25.470 121.425 ;
        RECT 25.640 120.855 25.860 121.725 ;
        RECT 26.040 121.415 26.390 121.785 ;
        RECT 26.560 121.235 26.730 121.965 ;
        RECT 26.900 121.905 27.310 122.345 ;
        RECT 27.600 121.705 27.850 122.135 ;
        RECT 28.050 121.885 28.370 122.345 ;
        RECT 28.930 121.955 29.780 122.125 ;
        RECT 26.900 121.365 27.310 121.695 ;
        RECT 27.600 121.365 28.020 121.705 ;
        RECT 26.310 121.195 26.730 121.235 ;
        RECT 26.310 121.025 27.660 121.195 ;
        RECT 24.720 120.465 25.415 120.635 ;
        RECT 25.640 120.475 26.140 120.855 ;
        RECT 24.745 119.795 25.075 120.295 ;
        RECT 25.245 119.965 25.415 120.465 ;
        RECT 26.310 120.180 26.480 121.025 ;
        RECT 27.410 120.865 27.660 121.025 ;
        RECT 26.650 120.595 26.900 120.855 ;
        RECT 27.830 120.595 28.020 121.365 ;
        RECT 26.650 120.345 28.020 120.595 ;
        RECT 28.190 121.535 29.440 121.705 ;
        RECT 28.190 120.775 28.360 121.535 ;
        RECT 29.110 121.415 29.440 121.535 ;
        RECT 28.530 120.955 28.710 121.365 ;
        RECT 29.610 121.195 29.780 121.955 ;
        RECT 29.980 121.865 30.640 122.345 ;
        RECT 30.820 121.750 31.140 122.080 ;
        RECT 29.970 121.425 30.630 121.695 ;
        RECT 29.970 121.365 30.300 121.425 ;
        RECT 30.450 121.195 30.780 121.255 ;
        RECT 28.880 121.025 30.780 121.195 ;
        RECT 28.190 120.465 28.710 120.775 ;
        RECT 28.880 120.515 29.050 121.025 ;
        RECT 30.950 120.855 31.140 121.750 ;
        RECT 29.220 120.685 31.140 120.855 ;
        RECT 30.820 120.665 31.140 120.685 ;
        RECT 31.340 121.435 31.590 122.085 ;
        RECT 31.770 121.885 32.055 122.345 ;
        RECT 32.235 122.005 32.490 122.165 ;
        RECT 32.235 121.835 32.575 122.005 ;
        RECT 32.235 121.635 32.490 121.835 ;
        RECT 31.340 121.105 32.140 121.435 ;
        RECT 28.880 120.345 30.090 120.515 ;
        RECT 25.650 120.010 26.480 120.180 ;
        RECT 26.720 119.795 27.100 120.175 ;
        RECT 27.280 120.055 27.450 120.345 ;
        RECT 28.880 120.265 29.050 120.345 ;
        RECT 27.620 119.795 27.950 120.175 ;
        RECT 28.420 120.015 29.050 120.265 ;
        RECT 29.230 119.795 29.650 120.175 ;
        RECT 29.850 120.055 30.090 120.345 ;
        RECT 30.320 119.795 30.650 120.485 ;
        RECT 30.820 120.055 30.990 120.665 ;
        RECT 31.340 120.515 31.590 121.105 ;
        RECT 32.310 120.775 32.490 121.635 ;
        RECT 33.410 121.635 33.665 122.165 ;
        RECT 33.845 121.885 34.130 122.345 ;
        RECT 33.410 121.325 33.590 121.635 ;
        RECT 34.310 121.435 34.560 122.085 ;
        RECT 33.325 121.155 33.590 121.325 ;
        RECT 31.260 120.005 31.590 120.515 ;
        RECT 31.770 119.795 32.055 120.595 ;
        RECT 32.235 120.105 32.490 120.775 ;
        RECT 33.410 120.775 33.590 121.155 ;
        RECT 33.760 121.105 34.560 121.435 ;
        RECT 33.410 120.105 33.665 120.775 ;
        RECT 33.845 119.795 34.130 120.595 ;
        RECT 34.310 120.515 34.560 121.105 ;
        RECT 34.760 121.750 35.080 122.080 ;
        RECT 35.260 121.865 35.920 122.345 ;
        RECT 36.120 121.955 36.970 122.125 ;
        RECT 34.760 120.855 34.950 121.750 ;
        RECT 35.270 121.425 35.930 121.695 ;
        RECT 35.600 121.365 35.930 121.425 ;
        RECT 35.120 121.195 35.450 121.255 ;
        RECT 36.120 121.195 36.290 121.955 ;
        RECT 37.530 121.885 37.850 122.345 ;
        RECT 38.050 121.705 38.300 122.135 ;
        RECT 38.590 121.905 39.000 122.345 ;
        RECT 39.170 121.965 40.185 122.165 ;
        RECT 36.460 121.535 37.710 121.705 ;
        RECT 36.460 121.415 36.790 121.535 ;
        RECT 35.120 121.025 37.020 121.195 ;
        RECT 34.760 120.685 36.680 120.855 ;
        RECT 34.760 120.665 35.080 120.685 ;
        RECT 34.310 120.005 34.640 120.515 ;
        RECT 34.910 120.055 35.080 120.665 ;
        RECT 36.850 120.515 37.020 121.025 ;
        RECT 37.190 120.955 37.370 121.365 ;
        RECT 37.540 120.775 37.710 121.535 ;
        RECT 35.250 119.795 35.580 120.485 ;
        RECT 35.810 120.345 37.020 120.515 ;
        RECT 37.190 120.465 37.710 120.775 ;
        RECT 37.880 121.365 38.300 121.705 ;
        RECT 38.590 121.365 39.000 121.695 ;
        RECT 37.880 120.595 38.070 121.365 ;
        RECT 39.170 121.235 39.340 121.965 ;
        RECT 40.485 121.795 40.655 122.125 ;
        RECT 40.825 121.965 41.155 122.345 ;
        RECT 39.510 121.415 39.860 121.785 ;
        RECT 39.170 121.195 39.590 121.235 ;
        RECT 38.240 121.025 39.590 121.195 ;
        RECT 38.240 120.865 38.490 121.025 ;
        RECT 39.000 120.595 39.250 120.855 ;
        RECT 37.880 120.345 39.250 120.595 ;
        RECT 35.810 120.055 36.050 120.345 ;
        RECT 36.850 120.265 37.020 120.345 ;
        RECT 36.250 119.795 36.670 120.175 ;
        RECT 36.850 120.015 37.480 120.265 ;
        RECT 37.950 119.795 38.280 120.175 ;
        RECT 38.450 120.055 38.620 120.345 ;
        RECT 39.420 120.180 39.590 121.025 ;
        RECT 40.040 120.855 40.260 121.725 ;
        RECT 40.485 121.605 41.180 121.795 ;
        RECT 39.760 120.475 40.260 120.855 ;
        RECT 40.430 120.805 40.840 121.425 ;
        RECT 41.010 120.635 41.180 121.605 ;
        RECT 40.485 120.465 41.180 120.635 ;
        RECT 38.800 119.795 39.180 120.175 ;
        RECT 39.420 120.010 40.250 120.180 ;
        RECT 40.485 119.965 40.655 120.465 ;
        RECT 40.825 119.795 41.155 120.295 ;
        RECT 41.370 119.965 41.595 122.085 ;
        RECT 41.765 121.965 42.095 122.345 ;
        RECT 42.265 121.795 42.435 122.085 ;
        RECT 41.770 121.625 42.435 121.795 ;
        RECT 41.770 120.635 42.000 121.625 ;
        RECT 42.970 121.535 43.215 122.140 ;
        RECT 43.435 121.810 43.945 122.345 ;
        RECT 42.170 120.805 42.520 121.455 ;
        RECT 42.695 121.365 43.925 121.535 ;
        RECT 41.770 120.465 42.435 120.635 ;
        RECT 41.765 119.795 42.095 120.295 ;
        RECT 42.265 119.965 42.435 120.465 ;
        RECT 42.695 120.555 43.035 121.365 ;
        RECT 43.205 120.800 43.955 120.990 ;
        RECT 42.695 120.145 43.210 120.555 ;
        RECT 43.445 119.795 43.615 120.555 ;
        RECT 43.785 120.135 43.955 120.800 ;
        RECT 44.125 120.815 44.315 122.175 ;
        RECT 44.485 121.325 44.760 122.175 ;
        RECT 44.950 121.810 45.480 122.175 ;
        RECT 45.905 121.945 46.235 122.345 ;
        RECT 45.305 121.775 45.480 121.810 ;
        RECT 44.485 121.155 44.765 121.325 ;
        RECT 44.485 121.015 44.760 121.155 ;
        RECT 44.965 120.815 45.135 121.615 ;
        RECT 44.125 120.645 45.135 120.815 ;
        RECT 45.305 121.605 46.235 121.775 ;
        RECT 46.405 121.605 46.660 122.175 ;
        RECT 46.925 121.795 47.095 122.175 ;
        RECT 47.275 121.965 47.605 122.345 ;
        RECT 46.925 121.625 47.590 121.795 ;
        RECT 47.785 121.670 48.045 122.175 ;
        RECT 45.305 120.475 45.475 121.605 ;
        RECT 46.065 121.435 46.235 121.605 ;
        RECT 44.350 120.305 45.475 120.475 ;
        RECT 45.645 121.105 45.840 121.435 ;
        RECT 46.065 121.105 46.320 121.435 ;
        RECT 45.645 120.135 45.815 121.105 ;
        RECT 46.490 120.935 46.660 121.605 ;
        RECT 46.855 121.075 47.185 121.445 ;
        RECT 47.420 121.370 47.590 121.625 ;
        RECT 43.785 119.965 45.815 120.135 ;
        RECT 45.985 119.795 46.155 120.935 ;
        RECT 46.325 119.965 46.660 120.935 ;
        RECT 47.420 121.040 47.705 121.370 ;
        RECT 47.420 120.895 47.590 121.040 ;
        RECT 46.925 120.725 47.590 120.895 ;
        RECT 47.875 120.870 48.045 121.670 ;
        RECT 48.675 121.620 48.965 122.345 ;
        RECT 49.135 121.575 50.805 122.345 ;
        RECT 46.925 119.965 47.095 120.725 ;
        RECT 47.275 119.795 47.605 120.555 ;
        RECT 47.775 119.965 48.045 120.870 ;
        RECT 48.675 119.795 48.965 120.960 ;
        RECT 49.135 120.885 49.885 121.405 ;
        RECT 50.055 121.055 50.805 121.575 ;
        RECT 50.980 121.605 51.235 122.175 ;
        RECT 51.405 121.945 51.735 122.345 ;
        RECT 52.160 121.810 52.690 122.175 ;
        RECT 52.880 122.005 53.155 122.175 ;
        RECT 52.875 121.835 53.155 122.005 ;
        RECT 52.160 121.775 52.335 121.810 ;
        RECT 51.405 121.605 52.335 121.775 ;
        RECT 50.980 120.935 51.150 121.605 ;
        RECT 51.405 121.435 51.575 121.605 ;
        RECT 51.320 121.105 51.575 121.435 ;
        RECT 51.800 121.105 51.995 121.435 ;
        RECT 49.135 119.795 50.805 120.885 ;
        RECT 50.980 119.965 51.315 120.935 ;
        RECT 51.485 119.795 51.655 120.935 ;
        RECT 51.825 120.135 51.995 121.105 ;
        RECT 52.165 120.475 52.335 121.605 ;
        RECT 52.505 120.815 52.675 121.615 ;
        RECT 52.880 121.015 53.155 121.835 ;
        RECT 53.325 120.815 53.515 122.175 ;
        RECT 53.695 121.810 54.205 122.345 ;
        RECT 54.425 121.535 54.670 122.140 ;
        RECT 55.390 121.535 55.635 122.140 ;
        RECT 55.855 121.810 56.365 122.345 ;
        RECT 53.715 121.365 54.945 121.535 ;
        RECT 52.505 120.645 53.515 120.815 ;
        RECT 53.685 120.800 54.435 120.990 ;
        RECT 52.165 120.305 53.290 120.475 ;
        RECT 53.685 120.135 53.855 120.800 ;
        RECT 54.605 120.555 54.945 121.365 ;
        RECT 51.825 119.965 53.855 120.135 ;
        RECT 54.025 119.795 54.195 120.555 ;
        RECT 54.430 120.145 54.945 120.555 ;
        RECT 55.115 121.365 56.345 121.535 ;
        RECT 55.115 120.555 55.455 121.365 ;
        RECT 55.625 120.800 56.375 120.990 ;
        RECT 55.115 120.145 55.630 120.555 ;
        RECT 55.865 119.795 56.035 120.555 ;
        RECT 56.205 120.135 56.375 120.800 ;
        RECT 56.545 120.815 56.735 122.175 ;
        RECT 56.905 121.325 57.180 122.175 ;
        RECT 57.370 121.810 57.900 122.175 ;
        RECT 58.325 121.945 58.655 122.345 ;
        RECT 57.725 121.775 57.900 121.810 ;
        RECT 56.905 121.155 57.185 121.325 ;
        RECT 56.905 121.015 57.180 121.155 ;
        RECT 57.385 120.815 57.555 121.615 ;
        RECT 56.545 120.645 57.555 120.815 ;
        RECT 57.725 121.605 58.655 121.775 ;
        RECT 58.825 121.605 59.080 122.175 ;
        RECT 59.345 121.795 59.515 122.175 ;
        RECT 59.695 121.965 60.025 122.345 ;
        RECT 59.345 121.625 60.010 121.795 ;
        RECT 60.205 121.670 60.465 122.175 ;
        RECT 57.725 120.475 57.895 121.605 ;
        RECT 58.485 121.435 58.655 121.605 ;
        RECT 56.770 120.305 57.895 120.475 ;
        RECT 58.065 121.105 58.260 121.435 ;
        RECT 58.485 121.105 58.740 121.435 ;
        RECT 58.065 120.135 58.235 121.105 ;
        RECT 58.910 120.935 59.080 121.605 ;
        RECT 59.275 121.075 59.605 121.445 ;
        RECT 59.840 121.370 60.010 121.625 ;
        RECT 56.205 119.965 58.235 120.135 ;
        RECT 58.405 119.795 58.575 120.935 ;
        RECT 58.745 119.965 59.080 120.935 ;
        RECT 59.840 121.040 60.125 121.370 ;
        RECT 59.840 120.895 60.010 121.040 ;
        RECT 59.345 120.725 60.010 120.895 ;
        RECT 60.295 120.870 60.465 121.670 ;
        RECT 60.675 121.525 60.905 122.345 ;
        RECT 61.075 121.545 61.405 122.175 ;
        RECT 60.655 121.105 60.985 121.355 ;
        RECT 61.155 120.945 61.405 121.545 ;
        RECT 61.575 121.525 61.785 122.345 ;
        RECT 62.390 122.005 62.645 122.165 ;
        RECT 62.305 121.835 62.645 122.005 ;
        RECT 62.825 121.885 63.110 122.345 ;
        RECT 62.390 121.635 62.645 121.835 ;
        RECT 59.345 119.965 59.515 120.725 ;
        RECT 59.695 119.795 60.025 120.555 ;
        RECT 60.195 119.965 60.465 120.870 ;
        RECT 60.675 119.795 60.905 120.935 ;
        RECT 61.075 119.965 61.405 120.945 ;
        RECT 61.575 119.795 61.785 120.935 ;
        RECT 62.390 120.775 62.570 121.635 ;
        RECT 63.290 121.435 63.540 122.085 ;
        RECT 62.740 121.105 63.540 121.435 ;
        RECT 62.390 120.105 62.645 120.775 ;
        RECT 62.825 119.795 63.110 120.595 ;
        RECT 63.290 120.515 63.540 121.105 ;
        RECT 63.740 121.750 64.060 122.080 ;
        RECT 64.240 121.865 64.900 122.345 ;
        RECT 65.100 121.955 65.950 122.125 ;
        RECT 63.740 120.855 63.930 121.750 ;
        RECT 64.250 121.425 64.910 121.695 ;
        RECT 64.580 121.365 64.910 121.425 ;
        RECT 64.100 121.195 64.430 121.255 ;
        RECT 65.100 121.195 65.270 121.955 ;
        RECT 66.510 121.885 66.830 122.345 ;
        RECT 67.030 121.705 67.280 122.135 ;
        RECT 67.570 121.905 67.980 122.345 ;
        RECT 68.150 121.965 69.165 122.165 ;
        RECT 65.440 121.535 66.690 121.705 ;
        RECT 65.440 121.415 65.770 121.535 ;
        RECT 64.100 121.025 66.000 121.195 ;
        RECT 63.740 120.685 65.660 120.855 ;
        RECT 63.740 120.665 64.060 120.685 ;
        RECT 63.290 120.005 63.620 120.515 ;
        RECT 63.890 120.055 64.060 120.665 ;
        RECT 65.830 120.515 66.000 121.025 ;
        RECT 66.170 120.955 66.350 121.365 ;
        RECT 66.520 120.775 66.690 121.535 ;
        RECT 64.230 119.795 64.560 120.485 ;
        RECT 64.790 120.345 66.000 120.515 ;
        RECT 66.170 120.465 66.690 120.775 ;
        RECT 66.860 121.365 67.280 121.705 ;
        RECT 67.570 121.365 67.980 121.695 ;
        RECT 66.860 120.595 67.050 121.365 ;
        RECT 68.150 121.235 68.320 121.965 ;
        RECT 69.465 121.795 69.635 122.125 ;
        RECT 69.805 121.965 70.135 122.345 ;
        RECT 68.490 121.415 68.840 121.785 ;
        RECT 68.150 121.195 68.570 121.235 ;
        RECT 67.220 121.025 68.570 121.195 ;
        RECT 67.220 120.865 67.470 121.025 ;
        RECT 67.980 120.595 68.230 120.855 ;
        RECT 66.860 120.345 68.230 120.595 ;
        RECT 64.790 120.055 65.030 120.345 ;
        RECT 65.830 120.265 66.000 120.345 ;
        RECT 65.230 119.795 65.650 120.175 ;
        RECT 65.830 120.015 66.460 120.265 ;
        RECT 66.930 119.795 67.260 120.175 ;
        RECT 67.430 120.055 67.600 120.345 ;
        RECT 68.400 120.180 68.570 121.025 ;
        RECT 69.020 120.855 69.240 121.725 ;
        RECT 69.465 121.605 70.160 121.795 ;
        RECT 68.740 120.475 69.240 120.855 ;
        RECT 69.410 120.805 69.820 121.425 ;
        RECT 69.990 120.635 70.160 121.605 ;
        RECT 69.465 120.465 70.160 120.635 ;
        RECT 67.780 119.795 68.160 120.175 ;
        RECT 68.400 120.010 69.230 120.180 ;
        RECT 69.465 119.965 69.635 120.465 ;
        RECT 69.805 119.795 70.135 120.295 ;
        RECT 70.350 119.965 70.575 122.085 ;
        RECT 70.745 121.965 71.075 122.345 ;
        RECT 71.245 121.795 71.415 122.085 ;
        RECT 70.750 121.625 71.415 121.795 ;
        RECT 71.675 121.670 71.935 122.175 ;
        RECT 72.115 121.965 72.445 122.345 ;
        RECT 72.625 121.795 72.795 122.175 ;
        RECT 70.750 120.635 70.980 121.625 ;
        RECT 71.150 120.805 71.500 121.455 ;
        RECT 71.675 120.870 71.845 121.670 ;
        RECT 72.130 121.625 72.795 121.795 ;
        RECT 73.055 121.670 73.315 122.175 ;
        RECT 73.495 121.965 73.825 122.345 ;
        RECT 74.005 121.795 74.175 122.175 ;
        RECT 72.130 121.370 72.300 121.625 ;
        RECT 72.015 121.040 72.300 121.370 ;
        RECT 72.535 121.075 72.865 121.445 ;
        RECT 72.130 120.895 72.300 121.040 ;
        RECT 70.750 120.465 71.415 120.635 ;
        RECT 70.745 119.795 71.075 120.295 ;
        RECT 71.245 119.965 71.415 120.465 ;
        RECT 71.675 119.965 71.945 120.870 ;
        RECT 72.130 120.725 72.795 120.895 ;
        RECT 72.115 119.795 72.445 120.555 ;
        RECT 72.625 119.965 72.795 120.725 ;
        RECT 73.055 120.870 73.225 121.670 ;
        RECT 73.510 121.625 74.175 121.795 ;
        RECT 73.510 121.370 73.680 121.625 ;
        RECT 74.435 121.620 74.725 122.345 ;
        RECT 74.935 121.525 75.165 122.345 ;
        RECT 75.335 121.545 75.665 122.175 ;
        RECT 73.395 121.040 73.680 121.370 ;
        RECT 73.915 121.075 74.245 121.445 ;
        RECT 74.915 121.105 75.245 121.355 ;
        RECT 73.510 120.895 73.680 121.040 ;
        RECT 73.055 119.965 73.325 120.870 ;
        RECT 73.510 120.725 74.175 120.895 ;
        RECT 73.495 119.795 73.825 120.555 ;
        RECT 74.005 119.965 74.175 120.725 ;
        RECT 74.435 119.795 74.725 120.960 ;
        RECT 75.415 120.945 75.665 121.545 ;
        RECT 75.835 121.525 76.045 122.345 ;
        RECT 76.650 121.635 76.905 122.165 ;
        RECT 77.085 121.885 77.370 122.345 ;
        RECT 74.935 119.795 75.165 120.935 ;
        RECT 75.335 119.965 75.665 120.945 ;
        RECT 75.835 119.795 76.045 120.935 ;
        RECT 76.650 120.775 76.830 121.635 ;
        RECT 77.550 121.435 77.800 122.085 ;
        RECT 77.000 121.105 77.800 121.435 ;
        RECT 76.650 120.305 76.905 120.775 ;
        RECT 76.565 120.135 76.905 120.305 ;
        RECT 76.650 120.105 76.905 120.135 ;
        RECT 77.085 119.795 77.370 120.595 ;
        RECT 77.550 120.515 77.800 121.105 ;
        RECT 78.000 121.750 78.320 122.080 ;
        RECT 78.500 121.865 79.160 122.345 ;
        RECT 79.360 121.955 80.210 122.125 ;
        RECT 78.000 120.855 78.190 121.750 ;
        RECT 78.510 121.425 79.170 121.695 ;
        RECT 78.840 121.365 79.170 121.425 ;
        RECT 78.360 121.195 78.690 121.255 ;
        RECT 79.360 121.195 79.530 121.955 ;
        RECT 80.770 121.885 81.090 122.345 ;
        RECT 81.290 121.705 81.540 122.135 ;
        RECT 81.830 121.905 82.240 122.345 ;
        RECT 82.410 121.965 83.425 122.165 ;
        RECT 79.700 121.535 80.950 121.705 ;
        RECT 79.700 121.415 80.030 121.535 ;
        RECT 78.360 121.025 80.260 121.195 ;
        RECT 78.000 120.685 79.920 120.855 ;
        RECT 78.000 120.665 78.320 120.685 ;
        RECT 77.550 120.005 77.880 120.515 ;
        RECT 78.150 120.055 78.320 120.665 ;
        RECT 80.090 120.515 80.260 121.025 ;
        RECT 80.430 120.955 80.610 121.365 ;
        RECT 80.780 120.775 80.950 121.535 ;
        RECT 78.490 119.795 78.820 120.485 ;
        RECT 79.050 120.345 80.260 120.515 ;
        RECT 80.430 120.465 80.950 120.775 ;
        RECT 81.120 121.365 81.540 121.705 ;
        RECT 81.830 121.365 82.240 121.695 ;
        RECT 81.120 120.595 81.310 121.365 ;
        RECT 82.410 121.235 82.580 121.965 ;
        RECT 83.725 121.795 83.895 122.125 ;
        RECT 84.065 121.965 84.395 122.345 ;
        RECT 82.750 121.415 83.100 121.785 ;
        RECT 82.410 121.195 82.830 121.235 ;
        RECT 81.480 121.025 82.830 121.195 ;
        RECT 81.480 120.865 81.730 121.025 ;
        RECT 82.240 120.595 82.490 120.855 ;
        RECT 81.120 120.345 82.490 120.595 ;
        RECT 79.050 120.055 79.290 120.345 ;
        RECT 80.090 120.265 80.260 120.345 ;
        RECT 79.490 119.795 79.910 120.175 ;
        RECT 80.090 120.015 80.720 120.265 ;
        RECT 81.190 119.795 81.520 120.175 ;
        RECT 81.690 120.055 81.860 120.345 ;
        RECT 82.660 120.180 82.830 121.025 ;
        RECT 83.280 120.855 83.500 121.725 ;
        RECT 83.725 121.605 84.420 121.795 ;
        RECT 83.000 120.475 83.500 120.855 ;
        RECT 83.670 120.805 84.080 121.425 ;
        RECT 84.250 120.635 84.420 121.605 ;
        RECT 83.725 120.465 84.420 120.635 ;
        RECT 82.040 119.795 82.420 120.175 ;
        RECT 82.660 120.010 83.490 120.180 ;
        RECT 83.725 119.965 83.895 120.465 ;
        RECT 84.065 119.795 84.395 120.295 ;
        RECT 84.610 119.965 84.835 122.085 ;
        RECT 85.005 121.965 85.335 122.345 ;
        RECT 85.505 121.795 85.675 122.085 ;
        RECT 85.010 121.625 85.675 121.795 ;
        RECT 85.010 120.635 85.240 121.625 ;
        RECT 85.975 121.525 86.205 122.345 ;
        RECT 86.375 121.545 86.705 122.175 ;
        RECT 85.410 120.805 85.760 121.455 ;
        RECT 85.955 121.105 86.285 121.355 ;
        RECT 86.455 120.945 86.705 121.545 ;
        RECT 86.875 121.525 87.085 122.345 ;
        RECT 87.315 121.670 87.575 122.175 ;
        RECT 87.755 121.965 88.085 122.345 ;
        RECT 88.265 121.795 88.435 122.175 ;
        RECT 85.010 120.465 85.675 120.635 ;
        RECT 85.005 119.795 85.335 120.295 ;
        RECT 85.505 119.965 85.675 120.465 ;
        RECT 85.975 119.795 86.205 120.935 ;
        RECT 86.375 119.965 86.705 120.945 ;
        RECT 86.875 119.795 87.085 120.935 ;
        RECT 87.315 120.870 87.485 121.670 ;
        RECT 87.770 121.625 88.435 121.795 ;
        RECT 88.695 121.670 88.955 122.175 ;
        RECT 89.135 121.965 89.465 122.345 ;
        RECT 89.645 121.795 89.815 122.175 ;
        RECT 87.770 121.370 87.940 121.625 ;
        RECT 87.655 121.040 87.940 121.370 ;
        RECT 88.175 121.075 88.505 121.445 ;
        RECT 87.770 120.895 87.940 121.040 ;
        RECT 87.315 119.965 87.585 120.870 ;
        RECT 87.770 120.725 88.435 120.895 ;
        RECT 87.755 119.795 88.085 120.555 ;
        RECT 88.265 119.965 88.435 120.725 ;
        RECT 88.695 120.870 88.865 121.670 ;
        RECT 89.150 121.625 89.815 121.795 ;
        RECT 89.150 121.370 89.320 121.625 ;
        RECT 90.115 121.525 90.345 122.345 ;
        RECT 90.515 121.545 90.845 122.175 ;
        RECT 89.035 121.040 89.320 121.370 ;
        RECT 89.555 121.075 89.885 121.445 ;
        RECT 90.095 121.105 90.425 121.355 ;
        RECT 89.150 120.895 89.320 121.040 ;
        RECT 90.595 120.945 90.845 121.545 ;
        RECT 91.015 121.525 91.225 122.345 ;
        RECT 91.730 121.535 91.975 122.140 ;
        RECT 92.195 121.810 92.705 122.345 ;
        RECT 88.695 119.965 88.965 120.870 ;
        RECT 89.150 120.725 89.815 120.895 ;
        RECT 89.135 119.795 89.465 120.555 ;
        RECT 89.645 119.965 89.815 120.725 ;
        RECT 90.115 119.795 90.345 120.935 ;
        RECT 90.515 119.965 90.845 120.945 ;
        RECT 91.455 121.365 92.685 121.535 ;
        RECT 91.015 119.795 91.225 120.935 ;
        RECT 91.455 120.555 91.795 121.365 ;
        RECT 91.965 120.800 92.715 120.990 ;
        RECT 91.455 120.145 91.970 120.555 ;
        RECT 92.205 119.795 92.375 120.555 ;
        RECT 92.545 120.135 92.715 120.800 ;
        RECT 92.885 120.815 93.075 122.175 ;
        RECT 93.245 121.665 93.520 122.175 ;
        RECT 93.710 121.810 94.240 122.175 ;
        RECT 94.665 121.945 94.995 122.345 ;
        RECT 94.065 121.775 94.240 121.810 ;
        RECT 93.245 121.495 93.525 121.665 ;
        RECT 93.245 121.015 93.520 121.495 ;
        RECT 93.725 120.815 93.895 121.615 ;
        RECT 92.885 120.645 93.895 120.815 ;
        RECT 94.065 121.605 94.995 121.775 ;
        RECT 95.165 121.605 95.420 122.175 ;
        RECT 94.065 120.475 94.235 121.605 ;
        RECT 94.825 121.435 94.995 121.605 ;
        RECT 93.110 120.305 94.235 120.475 ;
        RECT 94.405 121.105 94.600 121.435 ;
        RECT 94.825 121.105 95.080 121.435 ;
        RECT 94.405 120.135 94.575 121.105 ;
        RECT 95.250 120.935 95.420 121.605 ;
        RECT 96.330 121.535 96.575 122.140 ;
        RECT 96.795 121.810 97.305 122.345 ;
        RECT 92.545 119.965 94.575 120.135 ;
        RECT 94.745 119.795 94.915 120.935 ;
        RECT 95.085 119.965 95.420 120.935 ;
        RECT 96.055 121.365 97.285 121.535 ;
        RECT 96.055 120.555 96.395 121.365 ;
        RECT 96.565 120.800 97.315 120.990 ;
        RECT 96.055 120.145 96.570 120.555 ;
        RECT 96.805 119.795 96.975 120.555 ;
        RECT 97.145 120.135 97.315 120.800 ;
        RECT 97.485 120.815 97.675 122.175 ;
        RECT 97.845 122.005 98.120 122.175 ;
        RECT 97.845 121.835 98.125 122.005 ;
        RECT 97.845 121.015 98.120 121.835 ;
        RECT 98.310 121.810 98.840 122.175 ;
        RECT 99.265 121.945 99.595 122.345 ;
        RECT 98.665 121.775 98.840 121.810 ;
        RECT 98.325 120.815 98.495 121.615 ;
        RECT 97.485 120.645 98.495 120.815 ;
        RECT 98.665 121.605 99.595 121.775 ;
        RECT 99.765 121.605 100.020 122.175 ;
        RECT 100.195 121.620 100.485 122.345 ;
        RECT 101.030 122.005 101.285 122.165 ;
        RECT 100.945 121.835 101.285 122.005 ;
        RECT 101.465 121.885 101.750 122.345 ;
        RECT 101.030 121.635 101.285 121.835 ;
        RECT 98.665 120.475 98.835 121.605 ;
        RECT 99.425 121.435 99.595 121.605 ;
        RECT 97.710 120.305 98.835 120.475 ;
        RECT 99.005 121.105 99.200 121.435 ;
        RECT 99.425 121.105 99.680 121.435 ;
        RECT 99.005 120.135 99.175 121.105 ;
        RECT 99.850 120.935 100.020 121.605 ;
        RECT 97.145 119.965 99.175 120.135 ;
        RECT 99.345 119.795 99.515 120.935 ;
        RECT 99.685 119.965 100.020 120.935 ;
        RECT 100.195 119.795 100.485 120.960 ;
        RECT 101.030 120.775 101.210 121.635 ;
        RECT 101.930 121.435 102.180 122.085 ;
        RECT 101.380 121.105 102.180 121.435 ;
        RECT 101.030 120.105 101.285 120.775 ;
        RECT 101.465 119.795 101.750 120.595 ;
        RECT 101.930 120.515 102.180 121.105 ;
        RECT 102.380 121.750 102.700 122.080 ;
        RECT 102.880 121.865 103.540 122.345 ;
        RECT 103.740 121.955 104.590 122.125 ;
        RECT 102.380 120.855 102.570 121.750 ;
        RECT 102.890 121.425 103.550 121.695 ;
        RECT 103.220 121.365 103.550 121.425 ;
        RECT 102.740 121.195 103.070 121.255 ;
        RECT 103.740 121.195 103.910 121.955 ;
        RECT 105.150 121.885 105.470 122.345 ;
        RECT 105.670 121.705 105.920 122.135 ;
        RECT 106.210 121.905 106.620 122.345 ;
        RECT 106.790 121.965 107.805 122.165 ;
        RECT 104.080 121.535 105.330 121.705 ;
        RECT 104.080 121.415 104.410 121.535 ;
        RECT 102.740 121.025 104.640 121.195 ;
        RECT 102.380 120.685 104.300 120.855 ;
        RECT 102.380 120.665 102.700 120.685 ;
        RECT 101.930 120.005 102.260 120.515 ;
        RECT 102.530 120.055 102.700 120.665 ;
        RECT 104.470 120.515 104.640 121.025 ;
        RECT 104.810 120.955 104.990 121.365 ;
        RECT 105.160 120.775 105.330 121.535 ;
        RECT 102.870 119.795 103.200 120.485 ;
        RECT 103.430 120.345 104.640 120.515 ;
        RECT 104.810 120.465 105.330 120.775 ;
        RECT 105.500 121.365 105.920 121.705 ;
        RECT 106.210 121.365 106.620 121.695 ;
        RECT 105.500 120.595 105.690 121.365 ;
        RECT 106.790 121.235 106.960 121.965 ;
        RECT 108.105 121.795 108.275 122.125 ;
        RECT 108.445 121.965 108.775 122.345 ;
        RECT 107.130 121.415 107.480 121.785 ;
        RECT 106.790 121.195 107.210 121.235 ;
        RECT 105.860 121.025 107.210 121.195 ;
        RECT 105.860 120.865 106.110 121.025 ;
        RECT 106.620 120.595 106.870 120.855 ;
        RECT 105.500 120.345 106.870 120.595 ;
        RECT 103.430 120.055 103.670 120.345 ;
        RECT 104.470 120.265 104.640 120.345 ;
        RECT 103.870 119.795 104.290 120.175 ;
        RECT 104.470 120.015 105.100 120.265 ;
        RECT 105.570 119.795 105.900 120.175 ;
        RECT 106.070 120.055 106.240 120.345 ;
        RECT 107.040 120.180 107.210 121.025 ;
        RECT 107.660 120.855 107.880 121.725 ;
        RECT 108.105 121.605 108.800 121.795 ;
        RECT 107.380 120.475 107.880 120.855 ;
        RECT 108.050 120.805 108.460 121.425 ;
        RECT 108.630 120.635 108.800 121.605 ;
        RECT 108.105 120.465 108.800 120.635 ;
        RECT 106.420 119.795 106.800 120.175 ;
        RECT 107.040 120.010 107.870 120.180 ;
        RECT 108.105 119.965 108.275 120.465 ;
        RECT 108.445 119.795 108.775 120.295 ;
        RECT 108.990 119.965 109.215 122.085 ;
        RECT 109.385 121.965 109.715 122.345 ;
        RECT 109.885 121.795 110.055 122.085 ;
        RECT 109.390 121.625 110.055 121.795 ;
        RECT 109.390 120.635 109.620 121.625 ;
        RECT 110.315 121.575 111.985 122.345 ;
        RECT 112.155 121.595 113.365 122.345 ;
        RECT 109.790 120.805 110.140 121.455 ;
        RECT 110.315 120.885 111.065 121.405 ;
        RECT 111.235 121.055 111.985 121.575 ;
        RECT 112.155 120.885 112.675 121.425 ;
        RECT 112.845 121.055 113.365 121.595 ;
        RECT 109.390 120.465 110.055 120.635 ;
        RECT 109.385 119.795 109.715 120.295 ;
        RECT 109.885 119.965 110.055 120.465 ;
        RECT 110.315 119.795 111.985 120.885 ;
        RECT 112.155 119.795 113.365 120.885 ;
        RECT 11.330 119.625 113.450 119.795 ;
        RECT 11.415 118.535 12.625 119.625 ;
        RECT 13.105 118.785 13.275 119.625 ;
        RECT 13.485 118.615 13.735 119.455 ;
        RECT 13.945 118.785 14.115 119.625 ;
        RECT 14.285 118.615 14.575 119.455 ;
        RECT 11.415 117.825 11.935 118.365 ;
        RECT 12.105 117.995 12.625 118.535 ;
        RECT 12.850 118.445 14.575 118.615 ;
        RECT 14.785 118.565 14.955 119.625 ;
        RECT 15.250 119.245 15.580 119.625 ;
        RECT 15.760 119.075 15.930 119.365 ;
        RECT 16.100 119.165 16.350 119.625 ;
        RECT 15.130 118.905 15.930 119.075 ;
        RECT 16.520 119.115 17.390 119.455 ;
        RECT 12.850 117.895 13.260 118.445 ;
        RECT 15.130 118.285 15.300 118.905 ;
        RECT 16.520 118.735 16.690 119.115 ;
        RECT 17.625 118.995 17.795 119.455 ;
        RECT 17.965 119.165 18.335 119.625 ;
        RECT 18.630 119.025 18.800 119.365 ;
        RECT 18.970 119.195 19.300 119.625 ;
        RECT 19.535 119.025 19.705 119.365 ;
        RECT 15.470 118.565 16.690 118.735 ;
        RECT 16.860 118.655 17.320 118.945 ;
        RECT 17.625 118.825 18.185 118.995 ;
        RECT 18.630 118.855 19.705 119.025 ;
        RECT 19.875 119.125 20.555 119.455 ;
        RECT 20.770 119.125 21.020 119.455 ;
        RECT 21.190 119.165 21.440 119.625 ;
        RECT 18.015 118.685 18.185 118.825 ;
        RECT 16.860 118.645 17.825 118.655 ;
        RECT 16.520 118.475 16.690 118.565 ;
        RECT 17.150 118.485 17.825 118.645 ;
        RECT 15.130 118.275 15.475 118.285 ;
        RECT 13.445 118.065 15.475 118.275 ;
        RECT 11.415 117.075 12.625 117.825 ;
        RECT 12.850 117.725 14.615 117.895 ;
        RECT 13.105 117.075 13.275 117.545 ;
        RECT 13.445 117.245 13.775 117.725 ;
        RECT 13.945 117.075 14.115 117.545 ;
        RECT 14.285 117.245 14.615 117.725 ;
        RECT 14.785 117.075 14.955 117.885 ;
        RECT 15.150 117.810 15.475 118.065 ;
        RECT 15.155 117.455 15.475 117.810 ;
        RECT 15.645 118.025 16.185 118.395 ;
        RECT 16.520 118.305 16.925 118.475 ;
        RECT 15.645 117.625 15.885 118.025 ;
        RECT 16.365 117.855 16.585 118.135 ;
        RECT 16.055 117.685 16.585 117.855 ;
        RECT 16.055 117.455 16.225 117.685 ;
        RECT 16.755 117.525 16.925 118.305 ;
        RECT 17.095 117.695 17.445 118.315 ;
        RECT 17.615 117.695 17.825 118.485 ;
        RECT 18.015 118.515 19.515 118.685 ;
        RECT 18.015 117.825 18.185 118.515 ;
        RECT 19.875 118.345 20.045 119.125 ;
        RECT 20.850 118.995 21.020 119.125 ;
        RECT 18.355 118.175 20.045 118.345 ;
        RECT 20.215 118.565 20.680 118.955 ;
        RECT 20.850 118.825 21.245 118.995 ;
        RECT 18.355 117.995 18.525 118.175 ;
        RECT 15.155 117.285 16.225 117.455 ;
        RECT 16.395 117.075 16.585 117.515 ;
        RECT 16.755 117.245 17.705 117.525 ;
        RECT 18.015 117.435 18.275 117.825 ;
        RECT 18.695 117.755 19.485 118.005 ;
        RECT 17.925 117.265 18.275 117.435 ;
        RECT 18.485 117.075 18.815 117.535 ;
        RECT 19.690 117.465 19.860 118.175 ;
        RECT 20.215 117.975 20.385 118.565 ;
        RECT 20.030 117.755 20.385 117.975 ;
        RECT 20.555 117.755 20.905 118.375 ;
        RECT 21.075 117.465 21.245 118.825 ;
        RECT 21.610 118.655 21.935 119.440 ;
        RECT 21.415 117.605 21.875 118.655 ;
        RECT 19.690 117.295 20.545 117.465 ;
        RECT 20.750 117.295 21.245 117.465 ;
        RECT 21.415 117.075 21.745 117.435 ;
        RECT 22.105 117.335 22.275 119.455 ;
        RECT 22.445 119.125 22.775 119.625 ;
        RECT 22.945 118.955 23.200 119.455 ;
        RECT 22.450 118.785 23.200 118.955 ;
        RECT 23.465 118.955 23.635 119.455 ;
        RECT 23.805 119.125 24.135 119.625 ;
        RECT 23.465 118.785 24.130 118.955 ;
        RECT 22.450 117.795 22.680 118.785 ;
        RECT 22.850 117.965 23.200 118.615 ;
        RECT 23.380 117.965 23.730 118.615 ;
        RECT 23.900 117.795 24.130 118.785 ;
        RECT 22.450 117.625 23.200 117.795 ;
        RECT 22.445 117.075 22.775 117.455 ;
        RECT 22.945 117.335 23.200 117.625 ;
        RECT 23.465 117.625 24.130 117.795 ;
        RECT 23.465 117.335 23.635 117.625 ;
        RECT 23.805 117.075 24.135 117.455 ;
        RECT 24.305 117.335 24.530 119.455 ;
        RECT 24.745 119.125 25.075 119.625 ;
        RECT 25.245 118.955 25.415 119.455 ;
        RECT 25.650 119.240 26.480 119.410 ;
        RECT 26.720 119.245 27.100 119.625 ;
        RECT 24.720 118.785 25.415 118.955 ;
        RECT 24.720 117.815 24.890 118.785 ;
        RECT 25.060 117.995 25.470 118.615 ;
        RECT 25.640 118.565 26.140 118.945 ;
        RECT 24.720 117.625 25.415 117.815 ;
        RECT 25.640 117.695 25.860 118.565 ;
        RECT 26.310 118.395 26.480 119.240 ;
        RECT 27.280 119.075 27.450 119.365 ;
        RECT 27.620 119.245 27.950 119.625 ;
        RECT 28.420 119.155 29.050 119.405 ;
        RECT 29.230 119.245 29.650 119.625 ;
        RECT 28.880 119.075 29.050 119.155 ;
        RECT 29.850 119.075 30.090 119.365 ;
        RECT 26.650 118.825 28.020 119.075 ;
        RECT 26.650 118.565 26.900 118.825 ;
        RECT 27.410 118.395 27.660 118.555 ;
        RECT 26.310 118.225 27.660 118.395 ;
        RECT 26.310 118.185 26.730 118.225 ;
        RECT 26.040 117.635 26.390 118.005 ;
        RECT 24.745 117.075 25.075 117.455 ;
        RECT 25.245 117.295 25.415 117.625 ;
        RECT 26.560 117.455 26.730 118.185 ;
        RECT 27.830 118.055 28.020 118.825 ;
        RECT 26.900 117.725 27.310 118.055 ;
        RECT 27.600 117.715 28.020 118.055 ;
        RECT 28.190 118.645 28.710 118.955 ;
        RECT 28.880 118.905 30.090 119.075 ;
        RECT 30.320 118.935 30.650 119.625 ;
        RECT 28.190 117.885 28.360 118.645 ;
        RECT 28.530 118.055 28.710 118.465 ;
        RECT 28.880 118.395 29.050 118.905 ;
        RECT 30.820 118.755 30.990 119.365 ;
        RECT 31.260 118.905 31.590 119.415 ;
        RECT 30.820 118.735 31.140 118.755 ;
        RECT 29.220 118.565 31.140 118.735 ;
        RECT 28.880 118.225 30.780 118.395 ;
        RECT 29.110 117.885 29.440 118.005 ;
        RECT 28.190 117.715 29.440 117.885 ;
        RECT 25.715 117.255 26.730 117.455 ;
        RECT 26.900 117.075 27.310 117.515 ;
        RECT 27.600 117.285 27.850 117.715 ;
        RECT 28.050 117.075 28.370 117.535 ;
        RECT 29.610 117.465 29.780 118.225 ;
        RECT 30.450 118.165 30.780 118.225 ;
        RECT 29.970 117.995 30.300 118.055 ;
        RECT 29.970 117.725 30.630 117.995 ;
        RECT 30.950 117.670 31.140 118.565 ;
        RECT 28.930 117.295 29.780 117.465 ;
        RECT 29.980 117.075 30.640 117.555 ;
        RECT 30.820 117.340 31.140 117.670 ;
        RECT 31.340 118.315 31.590 118.905 ;
        RECT 31.770 118.825 32.055 119.625 ;
        RECT 32.235 119.285 32.490 119.315 ;
        RECT 32.235 119.115 32.575 119.285 ;
        RECT 32.235 118.645 32.490 119.115 ;
        RECT 31.340 117.985 32.140 118.315 ;
        RECT 31.340 117.335 31.590 117.985 ;
        RECT 32.310 117.785 32.490 118.645 ;
        RECT 31.770 117.075 32.055 117.535 ;
        RECT 32.235 117.255 32.490 117.785 ;
        RECT 33.955 118.550 34.225 119.455 ;
        RECT 34.395 118.865 34.725 119.625 ;
        RECT 34.905 118.695 35.075 119.455 ;
        RECT 33.955 117.750 34.125 118.550 ;
        RECT 34.410 118.525 35.075 118.695 ;
        RECT 34.410 118.380 34.580 118.525 ;
        RECT 35.795 118.460 36.085 119.625 ;
        RECT 36.255 118.535 37.925 119.625 ;
        RECT 38.185 118.695 38.355 119.455 ;
        RECT 38.535 118.865 38.865 119.625 ;
        RECT 34.295 118.050 34.580 118.380 ;
        RECT 34.410 117.795 34.580 118.050 ;
        RECT 34.815 117.975 35.145 118.345 ;
        RECT 36.255 118.015 37.005 118.535 ;
        RECT 38.185 118.525 38.850 118.695 ;
        RECT 39.035 118.550 39.305 119.455 ;
        RECT 38.680 118.380 38.850 118.525 ;
        RECT 37.175 117.845 37.925 118.365 ;
        RECT 38.115 117.975 38.445 118.345 ;
        RECT 38.680 118.050 38.965 118.380 ;
        RECT 33.955 117.245 34.215 117.750 ;
        RECT 34.410 117.625 35.075 117.795 ;
        RECT 34.395 117.075 34.725 117.455 ;
        RECT 34.905 117.245 35.075 117.625 ;
        RECT 35.795 117.075 36.085 117.800 ;
        RECT 36.255 117.075 37.925 117.845 ;
        RECT 38.680 117.795 38.850 118.050 ;
        RECT 38.185 117.625 38.850 117.795 ;
        RECT 39.135 117.750 39.305 118.550 ;
        RECT 39.850 118.645 40.105 119.315 ;
        RECT 40.285 118.825 40.570 119.625 ;
        RECT 40.750 118.905 41.080 119.415 ;
        RECT 39.850 118.265 40.030 118.645 ;
        RECT 40.750 118.315 41.000 118.905 ;
        RECT 41.350 118.755 41.520 119.365 ;
        RECT 41.690 118.935 42.020 119.625 ;
        RECT 42.250 119.075 42.490 119.365 ;
        RECT 42.690 119.245 43.110 119.625 ;
        RECT 43.290 119.155 43.920 119.405 ;
        RECT 44.390 119.245 44.720 119.625 ;
        RECT 43.290 119.075 43.460 119.155 ;
        RECT 44.890 119.075 45.060 119.365 ;
        RECT 45.240 119.245 45.620 119.625 ;
        RECT 45.860 119.240 46.690 119.410 ;
        RECT 42.250 118.905 43.460 119.075 ;
        RECT 39.765 118.095 40.030 118.265 ;
        RECT 38.185 117.245 38.355 117.625 ;
        RECT 38.535 117.075 38.865 117.455 ;
        RECT 39.045 117.245 39.305 117.750 ;
        RECT 39.850 117.785 40.030 118.095 ;
        RECT 40.200 117.985 41.000 118.315 ;
        RECT 39.850 117.255 40.105 117.785 ;
        RECT 40.285 117.075 40.570 117.535 ;
        RECT 40.750 117.335 41.000 117.985 ;
        RECT 41.200 118.735 41.520 118.755 ;
        RECT 41.200 118.565 43.120 118.735 ;
        RECT 41.200 117.670 41.390 118.565 ;
        RECT 43.290 118.395 43.460 118.905 ;
        RECT 43.630 118.645 44.150 118.955 ;
        RECT 41.560 118.225 43.460 118.395 ;
        RECT 41.560 118.165 41.890 118.225 ;
        RECT 42.040 117.995 42.370 118.055 ;
        RECT 41.710 117.725 42.370 117.995 ;
        RECT 41.200 117.340 41.520 117.670 ;
        RECT 41.700 117.075 42.360 117.555 ;
        RECT 42.560 117.465 42.730 118.225 ;
        RECT 43.630 118.055 43.810 118.465 ;
        RECT 42.900 117.885 43.230 118.005 ;
        RECT 43.980 117.885 44.150 118.645 ;
        RECT 42.900 117.715 44.150 117.885 ;
        RECT 44.320 118.825 45.690 119.075 ;
        RECT 44.320 118.055 44.510 118.825 ;
        RECT 45.440 118.565 45.690 118.825 ;
        RECT 44.680 118.395 44.930 118.555 ;
        RECT 45.860 118.395 46.030 119.240 ;
        RECT 46.925 118.955 47.095 119.455 ;
        RECT 47.265 119.125 47.595 119.625 ;
        RECT 46.200 118.565 46.700 118.945 ;
        RECT 46.925 118.785 47.620 118.955 ;
        RECT 44.680 118.225 46.030 118.395 ;
        RECT 45.610 118.185 46.030 118.225 ;
        RECT 44.320 117.715 44.740 118.055 ;
        RECT 45.030 117.725 45.440 118.055 ;
        RECT 42.560 117.295 43.410 117.465 ;
        RECT 43.970 117.075 44.290 117.535 ;
        RECT 44.490 117.285 44.740 117.715 ;
        RECT 45.030 117.075 45.440 117.515 ;
        RECT 45.610 117.455 45.780 118.185 ;
        RECT 45.950 117.635 46.300 118.005 ;
        RECT 46.480 117.695 46.700 118.565 ;
        RECT 46.870 117.995 47.280 118.615 ;
        RECT 47.450 117.815 47.620 118.785 ;
        RECT 46.925 117.625 47.620 117.815 ;
        RECT 45.610 117.255 46.625 117.455 ;
        RECT 46.925 117.295 47.095 117.625 ;
        RECT 47.265 117.075 47.595 117.455 ;
        RECT 47.810 117.335 48.035 119.455 ;
        RECT 48.205 119.125 48.535 119.625 ;
        RECT 48.705 118.955 48.875 119.455 ;
        RECT 48.210 118.785 48.875 118.955 ;
        RECT 48.210 117.795 48.440 118.785 ;
        RECT 48.610 117.965 48.960 118.615 ;
        RECT 49.135 118.535 50.345 119.625 ;
        RECT 50.515 118.550 50.785 119.455 ;
        RECT 50.955 118.865 51.285 119.625 ;
        RECT 51.465 118.695 51.635 119.455 ;
        RECT 49.135 117.995 49.655 118.535 ;
        RECT 49.825 117.825 50.345 118.365 ;
        RECT 48.210 117.625 48.875 117.795 ;
        RECT 48.205 117.075 48.535 117.455 ;
        RECT 48.705 117.335 48.875 117.625 ;
        RECT 49.135 117.075 50.345 117.825 ;
        RECT 50.515 117.750 50.685 118.550 ;
        RECT 50.970 118.525 51.635 118.695 ;
        RECT 52.270 118.645 52.525 119.315 ;
        RECT 52.705 118.825 52.990 119.625 ;
        RECT 53.170 118.905 53.500 119.415 ;
        RECT 50.970 118.380 51.140 118.525 ;
        RECT 50.855 118.050 51.140 118.380 ;
        RECT 50.970 117.795 51.140 118.050 ;
        RECT 51.375 117.975 51.705 118.345 ;
        RECT 52.270 118.265 52.450 118.645 ;
        RECT 53.170 118.315 53.420 118.905 ;
        RECT 53.770 118.755 53.940 119.365 ;
        RECT 54.110 118.935 54.440 119.625 ;
        RECT 54.670 119.075 54.910 119.365 ;
        RECT 55.110 119.245 55.530 119.625 ;
        RECT 55.710 119.155 56.340 119.405 ;
        RECT 56.810 119.245 57.140 119.625 ;
        RECT 55.710 119.075 55.880 119.155 ;
        RECT 57.310 119.075 57.480 119.365 ;
        RECT 57.660 119.245 58.040 119.625 ;
        RECT 58.280 119.240 59.110 119.410 ;
        RECT 54.670 118.905 55.880 119.075 ;
        RECT 52.185 118.095 52.450 118.265 ;
        RECT 50.515 117.245 50.775 117.750 ;
        RECT 50.970 117.625 51.635 117.795 ;
        RECT 50.955 117.075 51.285 117.455 ;
        RECT 51.465 117.245 51.635 117.625 ;
        RECT 52.270 117.785 52.450 118.095 ;
        RECT 52.620 117.985 53.420 118.315 ;
        RECT 52.270 117.255 52.525 117.785 ;
        RECT 52.705 117.075 52.990 117.535 ;
        RECT 53.170 117.335 53.420 117.985 ;
        RECT 53.620 118.735 53.940 118.755 ;
        RECT 53.620 118.565 55.540 118.735 ;
        RECT 53.620 117.670 53.810 118.565 ;
        RECT 55.710 118.395 55.880 118.905 ;
        RECT 56.050 118.645 56.570 118.955 ;
        RECT 53.980 118.225 55.880 118.395 ;
        RECT 53.980 118.165 54.310 118.225 ;
        RECT 54.460 117.995 54.790 118.055 ;
        RECT 54.130 117.725 54.790 117.995 ;
        RECT 53.620 117.340 53.940 117.670 ;
        RECT 54.120 117.075 54.780 117.555 ;
        RECT 54.980 117.465 55.150 118.225 ;
        RECT 56.050 118.055 56.230 118.465 ;
        RECT 55.320 117.885 55.650 118.005 ;
        RECT 56.400 117.885 56.570 118.645 ;
        RECT 55.320 117.715 56.570 117.885 ;
        RECT 56.740 118.825 58.110 119.075 ;
        RECT 56.740 118.055 56.930 118.825 ;
        RECT 57.860 118.565 58.110 118.825 ;
        RECT 57.100 118.395 57.350 118.555 ;
        RECT 58.280 118.395 58.450 119.240 ;
        RECT 59.345 118.955 59.515 119.455 ;
        RECT 59.685 119.125 60.015 119.625 ;
        RECT 58.620 118.565 59.120 118.945 ;
        RECT 59.345 118.785 60.040 118.955 ;
        RECT 57.100 118.225 58.450 118.395 ;
        RECT 58.030 118.185 58.450 118.225 ;
        RECT 56.740 117.715 57.160 118.055 ;
        RECT 57.450 117.725 57.860 118.055 ;
        RECT 54.980 117.295 55.830 117.465 ;
        RECT 56.390 117.075 56.710 117.535 ;
        RECT 56.910 117.285 57.160 117.715 ;
        RECT 57.450 117.075 57.860 117.515 ;
        RECT 58.030 117.455 58.200 118.185 ;
        RECT 58.370 117.635 58.720 118.005 ;
        RECT 58.900 117.695 59.120 118.565 ;
        RECT 59.290 117.995 59.700 118.615 ;
        RECT 59.870 117.815 60.040 118.785 ;
        RECT 59.345 117.625 60.040 117.815 ;
        RECT 58.030 117.255 59.045 117.455 ;
        RECT 59.345 117.295 59.515 117.625 ;
        RECT 59.685 117.075 60.015 117.455 ;
        RECT 60.230 117.335 60.455 119.455 ;
        RECT 60.625 119.125 60.955 119.625 ;
        RECT 61.125 118.955 61.295 119.455 ;
        RECT 60.630 118.785 61.295 118.955 ;
        RECT 60.630 117.795 60.860 118.785 ;
        RECT 61.030 117.965 61.380 118.615 ;
        RECT 61.555 118.460 61.845 119.625 ;
        RECT 62.075 118.485 62.285 119.625 ;
        RECT 62.455 118.475 62.785 119.455 ;
        RECT 62.955 118.485 63.185 119.625 ;
        RECT 63.395 118.535 64.605 119.625 ;
        RECT 65.150 119.285 65.405 119.315 ;
        RECT 65.065 119.115 65.405 119.285 ;
        RECT 65.150 118.645 65.405 119.115 ;
        RECT 65.585 118.825 65.870 119.625 ;
        RECT 66.050 118.905 66.380 119.415 ;
        RECT 60.630 117.625 61.295 117.795 ;
        RECT 60.625 117.075 60.955 117.455 ;
        RECT 61.125 117.335 61.295 117.625 ;
        RECT 61.555 117.075 61.845 117.800 ;
        RECT 62.075 117.075 62.285 117.895 ;
        RECT 62.455 117.875 62.705 118.475 ;
        RECT 62.875 118.065 63.205 118.315 ;
        RECT 63.395 117.995 63.915 118.535 ;
        RECT 62.455 117.245 62.785 117.875 ;
        RECT 62.955 117.075 63.185 117.895 ;
        RECT 64.085 117.825 64.605 118.365 ;
        RECT 63.395 117.075 64.605 117.825 ;
        RECT 65.150 117.785 65.330 118.645 ;
        RECT 66.050 118.315 66.300 118.905 ;
        RECT 66.650 118.755 66.820 119.365 ;
        RECT 66.990 118.935 67.320 119.625 ;
        RECT 67.550 119.075 67.790 119.365 ;
        RECT 67.990 119.245 68.410 119.625 ;
        RECT 68.590 119.155 69.220 119.405 ;
        RECT 69.690 119.245 70.020 119.625 ;
        RECT 68.590 119.075 68.760 119.155 ;
        RECT 70.190 119.075 70.360 119.365 ;
        RECT 70.540 119.245 70.920 119.625 ;
        RECT 71.160 119.240 71.990 119.410 ;
        RECT 67.550 118.905 68.760 119.075 ;
        RECT 65.500 117.985 66.300 118.315 ;
        RECT 65.150 117.255 65.405 117.785 ;
        RECT 65.585 117.075 65.870 117.535 ;
        RECT 66.050 117.335 66.300 117.985 ;
        RECT 66.500 118.735 66.820 118.755 ;
        RECT 66.500 118.565 68.420 118.735 ;
        RECT 66.500 117.670 66.690 118.565 ;
        RECT 68.590 118.395 68.760 118.905 ;
        RECT 68.930 118.645 69.450 118.955 ;
        RECT 66.860 118.225 68.760 118.395 ;
        RECT 66.860 118.165 67.190 118.225 ;
        RECT 67.340 117.995 67.670 118.055 ;
        RECT 67.010 117.725 67.670 117.995 ;
        RECT 66.500 117.340 66.820 117.670 ;
        RECT 67.000 117.075 67.660 117.555 ;
        RECT 67.860 117.465 68.030 118.225 ;
        RECT 68.930 118.055 69.110 118.465 ;
        RECT 68.200 117.885 68.530 118.005 ;
        RECT 69.280 117.885 69.450 118.645 ;
        RECT 68.200 117.715 69.450 117.885 ;
        RECT 69.620 118.825 70.990 119.075 ;
        RECT 69.620 118.055 69.810 118.825 ;
        RECT 70.740 118.565 70.990 118.825 ;
        RECT 69.980 118.395 70.230 118.555 ;
        RECT 71.160 118.395 71.330 119.240 ;
        RECT 72.225 118.955 72.395 119.455 ;
        RECT 72.565 119.125 72.895 119.625 ;
        RECT 71.500 118.565 72.000 118.945 ;
        RECT 72.225 118.785 72.920 118.955 ;
        RECT 69.980 118.225 71.330 118.395 ;
        RECT 70.910 118.185 71.330 118.225 ;
        RECT 69.620 117.715 70.040 118.055 ;
        RECT 70.330 117.725 70.740 118.055 ;
        RECT 67.860 117.295 68.710 117.465 ;
        RECT 69.270 117.075 69.590 117.535 ;
        RECT 69.790 117.285 70.040 117.715 ;
        RECT 70.330 117.075 70.740 117.515 ;
        RECT 70.910 117.455 71.080 118.185 ;
        RECT 71.250 117.635 71.600 118.005 ;
        RECT 71.780 117.695 72.000 118.565 ;
        RECT 72.170 117.995 72.580 118.615 ;
        RECT 72.750 117.815 72.920 118.785 ;
        RECT 72.225 117.625 72.920 117.815 ;
        RECT 70.910 117.255 71.925 117.455 ;
        RECT 72.225 117.295 72.395 117.625 ;
        RECT 72.565 117.075 72.895 117.455 ;
        RECT 73.110 117.335 73.335 119.455 ;
        RECT 73.505 119.125 73.835 119.625 ;
        RECT 74.005 118.955 74.175 119.455 ;
        RECT 73.510 118.785 74.175 118.955 ;
        RECT 73.510 117.795 73.740 118.785 ;
        RECT 73.910 117.965 74.260 118.615 ;
        RECT 74.435 118.535 76.105 119.625 ;
        RECT 76.365 118.695 76.535 119.455 ;
        RECT 76.715 118.865 77.045 119.625 ;
        RECT 74.435 118.015 75.185 118.535 ;
        RECT 76.365 118.525 77.030 118.695 ;
        RECT 77.215 118.550 77.485 119.455 ;
        RECT 77.745 118.955 77.915 119.455 ;
        RECT 78.085 119.125 78.415 119.625 ;
        RECT 77.745 118.785 78.410 118.955 ;
        RECT 76.860 118.380 77.030 118.525 ;
        RECT 75.355 117.845 76.105 118.365 ;
        RECT 76.295 117.975 76.625 118.345 ;
        RECT 76.860 118.050 77.145 118.380 ;
        RECT 73.510 117.625 74.175 117.795 ;
        RECT 73.505 117.075 73.835 117.455 ;
        RECT 74.005 117.335 74.175 117.625 ;
        RECT 74.435 117.075 76.105 117.845 ;
        RECT 76.860 117.795 77.030 118.050 ;
        RECT 76.365 117.625 77.030 117.795 ;
        RECT 77.315 117.750 77.485 118.550 ;
        RECT 77.660 117.965 78.010 118.615 ;
        RECT 78.180 117.795 78.410 118.785 ;
        RECT 76.365 117.245 76.535 117.625 ;
        RECT 76.715 117.075 77.045 117.455 ;
        RECT 77.225 117.245 77.485 117.750 ;
        RECT 77.745 117.625 78.410 117.795 ;
        RECT 77.745 117.335 77.915 117.625 ;
        RECT 78.085 117.075 78.415 117.455 ;
        RECT 78.585 117.335 78.810 119.455 ;
        RECT 79.025 119.125 79.355 119.625 ;
        RECT 79.525 118.955 79.695 119.455 ;
        RECT 79.930 119.240 80.760 119.410 ;
        RECT 81.000 119.245 81.380 119.625 ;
        RECT 79.000 118.785 79.695 118.955 ;
        RECT 79.000 117.815 79.170 118.785 ;
        RECT 79.340 117.995 79.750 118.615 ;
        RECT 79.920 118.565 80.420 118.945 ;
        RECT 79.000 117.625 79.695 117.815 ;
        RECT 79.920 117.695 80.140 118.565 ;
        RECT 80.590 118.395 80.760 119.240 ;
        RECT 81.560 119.075 81.730 119.365 ;
        RECT 81.900 119.245 82.230 119.625 ;
        RECT 82.700 119.155 83.330 119.405 ;
        RECT 83.510 119.245 83.930 119.625 ;
        RECT 83.160 119.075 83.330 119.155 ;
        RECT 84.130 119.075 84.370 119.365 ;
        RECT 80.930 118.825 82.300 119.075 ;
        RECT 80.930 118.565 81.180 118.825 ;
        RECT 81.690 118.395 81.940 118.555 ;
        RECT 80.590 118.225 81.940 118.395 ;
        RECT 80.590 118.185 81.010 118.225 ;
        RECT 80.320 117.635 80.670 118.005 ;
        RECT 79.025 117.075 79.355 117.455 ;
        RECT 79.525 117.295 79.695 117.625 ;
        RECT 80.840 117.455 81.010 118.185 ;
        RECT 82.110 118.055 82.300 118.825 ;
        RECT 81.180 117.725 81.590 118.055 ;
        RECT 81.880 117.715 82.300 118.055 ;
        RECT 82.470 118.645 82.990 118.955 ;
        RECT 83.160 118.905 84.370 119.075 ;
        RECT 84.600 118.935 84.930 119.625 ;
        RECT 82.470 117.885 82.640 118.645 ;
        RECT 82.810 118.055 82.990 118.465 ;
        RECT 83.160 118.395 83.330 118.905 ;
        RECT 85.100 118.755 85.270 119.365 ;
        RECT 85.540 118.905 85.870 119.415 ;
        RECT 85.100 118.735 85.420 118.755 ;
        RECT 83.500 118.565 85.420 118.735 ;
        RECT 83.160 118.225 85.060 118.395 ;
        RECT 83.390 117.885 83.720 118.005 ;
        RECT 82.470 117.715 83.720 117.885 ;
        RECT 79.995 117.255 81.010 117.455 ;
        RECT 81.180 117.075 81.590 117.515 ;
        RECT 81.880 117.285 82.130 117.715 ;
        RECT 82.330 117.075 82.650 117.535 ;
        RECT 83.890 117.465 84.060 118.225 ;
        RECT 84.730 118.165 85.060 118.225 ;
        RECT 84.250 117.995 84.580 118.055 ;
        RECT 84.250 117.725 84.910 117.995 ;
        RECT 85.230 117.670 85.420 118.565 ;
        RECT 83.210 117.295 84.060 117.465 ;
        RECT 84.260 117.075 84.920 117.555 ;
        RECT 85.100 117.340 85.420 117.670 ;
        RECT 85.620 118.315 85.870 118.905 ;
        RECT 86.050 118.825 86.335 119.625 ;
        RECT 86.515 119.285 86.770 119.315 ;
        RECT 86.515 119.115 86.855 119.285 ;
        RECT 86.515 118.645 86.770 119.115 ;
        RECT 85.620 117.985 86.420 118.315 ;
        RECT 85.620 117.335 85.870 117.985 ;
        RECT 86.590 117.785 86.770 118.645 ;
        RECT 87.315 118.460 87.605 119.625 ;
        RECT 88.235 118.535 90.825 119.625 ;
        RECT 91.370 119.285 91.625 119.315 ;
        RECT 91.285 119.115 91.625 119.285 ;
        RECT 91.370 118.645 91.625 119.115 ;
        RECT 91.805 118.825 92.090 119.625 ;
        RECT 92.270 118.905 92.600 119.415 ;
        RECT 88.235 118.015 89.445 118.535 ;
        RECT 89.615 117.845 90.825 118.365 ;
        RECT 86.050 117.075 86.335 117.535 ;
        RECT 86.515 117.255 86.770 117.785 ;
        RECT 87.315 117.075 87.605 117.800 ;
        RECT 88.235 117.075 90.825 117.845 ;
        RECT 91.370 117.785 91.550 118.645 ;
        RECT 92.270 118.315 92.520 118.905 ;
        RECT 92.870 118.755 93.040 119.365 ;
        RECT 93.210 118.935 93.540 119.625 ;
        RECT 93.770 119.075 94.010 119.365 ;
        RECT 94.210 119.245 94.630 119.625 ;
        RECT 94.810 119.155 95.440 119.405 ;
        RECT 95.910 119.245 96.240 119.625 ;
        RECT 94.810 119.075 94.980 119.155 ;
        RECT 96.410 119.075 96.580 119.365 ;
        RECT 96.760 119.245 97.140 119.625 ;
        RECT 97.380 119.240 98.210 119.410 ;
        RECT 93.770 118.905 94.980 119.075 ;
        RECT 91.720 117.985 92.520 118.315 ;
        RECT 91.370 117.255 91.625 117.785 ;
        RECT 91.805 117.075 92.090 117.535 ;
        RECT 92.270 117.335 92.520 117.985 ;
        RECT 92.720 118.735 93.040 118.755 ;
        RECT 92.720 118.565 94.640 118.735 ;
        RECT 92.720 117.670 92.910 118.565 ;
        RECT 94.810 118.395 94.980 118.905 ;
        RECT 95.150 118.645 95.670 118.955 ;
        RECT 93.080 118.225 94.980 118.395 ;
        RECT 93.080 118.165 93.410 118.225 ;
        RECT 93.560 117.995 93.890 118.055 ;
        RECT 93.230 117.725 93.890 117.995 ;
        RECT 92.720 117.340 93.040 117.670 ;
        RECT 93.220 117.075 93.880 117.555 ;
        RECT 94.080 117.465 94.250 118.225 ;
        RECT 95.150 118.055 95.330 118.465 ;
        RECT 94.420 117.885 94.750 118.005 ;
        RECT 95.500 117.885 95.670 118.645 ;
        RECT 94.420 117.715 95.670 117.885 ;
        RECT 95.840 118.825 97.210 119.075 ;
        RECT 95.840 118.055 96.030 118.825 ;
        RECT 96.960 118.565 97.210 118.825 ;
        RECT 96.200 118.395 96.450 118.555 ;
        RECT 97.380 118.395 97.550 119.240 ;
        RECT 98.445 118.955 98.615 119.455 ;
        RECT 98.785 119.125 99.115 119.625 ;
        RECT 97.720 118.565 98.220 118.945 ;
        RECT 98.445 118.785 99.140 118.955 ;
        RECT 96.200 118.225 97.550 118.395 ;
        RECT 97.130 118.185 97.550 118.225 ;
        RECT 95.840 117.715 96.260 118.055 ;
        RECT 96.550 117.725 96.960 118.055 ;
        RECT 94.080 117.295 94.930 117.465 ;
        RECT 95.490 117.075 95.810 117.535 ;
        RECT 96.010 117.285 96.260 117.715 ;
        RECT 96.550 117.075 96.960 117.515 ;
        RECT 97.130 117.455 97.300 118.185 ;
        RECT 97.470 117.635 97.820 118.005 ;
        RECT 98.000 117.695 98.220 118.565 ;
        RECT 98.390 117.995 98.800 118.615 ;
        RECT 98.970 117.815 99.140 118.785 ;
        RECT 98.445 117.625 99.140 117.815 ;
        RECT 97.130 117.255 98.145 117.455 ;
        RECT 98.445 117.295 98.615 117.625 ;
        RECT 98.785 117.075 99.115 117.455 ;
        RECT 99.330 117.335 99.555 119.455 ;
        RECT 99.725 119.125 100.055 119.625 ;
        RECT 100.225 118.955 100.395 119.455 ;
        RECT 99.730 118.785 100.395 118.955 ;
        RECT 99.730 117.795 99.960 118.785 ;
        RECT 100.130 117.965 100.480 118.615 ;
        RECT 101.115 118.535 103.705 119.625 ;
        RECT 101.115 118.015 102.325 118.535 ;
        RECT 103.915 118.485 104.145 119.625 ;
        RECT 104.315 118.475 104.645 119.455 ;
        RECT 104.815 118.485 105.025 119.625 ;
        RECT 105.345 118.695 105.515 119.455 ;
        RECT 105.695 118.865 106.025 119.625 ;
        RECT 105.345 118.525 106.010 118.695 ;
        RECT 106.195 118.550 106.465 119.455 ;
        RECT 106.640 119.190 111.985 119.625 ;
        RECT 102.495 117.845 103.705 118.365 ;
        RECT 103.895 118.065 104.225 118.315 ;
        RECT 99.730 117.625 100.395 117.795 ;
        RECT 99.725 117.075 100.055 117.455 ;
        RECT 100.225 117.335 100.395 117.625 ;
        RECT 101.115 117.075 103.705 117.845 ;
        RECT 103.915 117.075 104.145 117.895 ;
        RECT 104.395 117.875 104.645 118.475 ;
        RECT 105.840 118.380 106.010 118.525 ;
        RECT 105.275 117.975 105.605 118.345 ;
        RECT 105.840 118.050 106.125 118.380 ;
        RECT 104.315 117.245 104.645 117.875 ;
        RECT 104.815 117.075 105.025 117.895 ;
        RECT 105.840 117.795 106.010 118.050 ;
        RECT 105.345 117.625 106.010 117.795 ;
        RECT 106.295 117.750 106.465 118.550 ;
        RECT 108.230 117.940 108.580 119.190 ;
        RECT 112.155 118.535 113.365 119.625 ;
        RECT 105.345 117.245 105.515 117.625 ;
        RECT 105.695 117.075 106.025 117.455 ;
        RECT 106.205 117.245 106.465 117.750 ;
        RECT 110.060 117.620 110.400 118.450 ;
        RECT 112.155 117.995 112.675 118.535 ;
        RECT 112.845 117.825 113.365 118.365 ;
        RECT 106.640 117.075 111.985 117.620 ;
        RECT 112.155 117.075 113.365 117.825 ;
        RECT 11.330 116.905 113.450 117.075 ;
        RECT 11.415 116.155 12.625 116.905 ;
        RECT 11.415 115.615 11.935 116.155 ;
        RECT 12.795 116.135 15.385 116.905 ;
        RECT 15.645 116.355 15.815 116.735 ;
        RECT 15.995 116.525 16.325 116.905 ;
        RECT 15.645 116.185 16.310 116.355 ;
        RECT 16.505 116.230 16.765 116.735 ;
        RECT 12.105 115.445 12.625 115.985 ;
        RECT 11.415 114.355 12.625 115.445 ;
        RECT 12.795 115.445 14.005 115.965 ;
        RECT 14.175 115.615 15.385 116.135 ;
        RECT 15.575 115.635 15.905 116.005 ;
        RECT 16.140 115.930 16.310 116.185 ;
        RECT 16.140 115.600 16.425 115.930 ;
        RECT 16.140 115.455 16.310 115.600 ;
        RECT 12.795 114.355 15.385 115.445 ;
        RECT 15.645 115.285 16.310 115.455 ;
        RECT 16.595 115.430 16.765 116.230 ;
        RECT 15.645 114.525 15.815 115.285 ;
        RECT 15.995 114.355 16.325 115.115 ;
        RECT 16.495 114.525 16.765 115.430 ;
        RECT 16.940 116.165 17.195 116.735 ;
        RECT 17.365 116.505 17.695 116.905 ;
        RECT 18.120 116.370 18.650 116.735 ;
        RECT 18.120 116.335 18.295 116.370 ;
        RECT 17.365 116.165 18.295 116.335 ;
        RECT 18.840 116.225 19.115 116.735 ;
        RECT 16.940 115.495 17.110 116.165 ;
        RECT 17.365 115.995 17.535 116.165 ;
        RECT 17.280 115.665 17.535 115.995 ;
        RECT 17.760 115.665 17.955 115.995 ;
        RECT 16.940 114.525 17.275 115.495 ;
        RECT 17.445 114.355 17.615 115.495 ;
        RECT 17.785 114.695 17.955 115.665 ;
        RECT 18.125 115.035 18.295 116.165 ;
        RECT 18.465 115.375 18.635 116.175 ;
        RECT 18.835 116.055 19.115 116.225 ;
        RECT 18.840 115.575 19.115 116.055 ;
        RECT 19.285 115.375 19.475 116.735 ;
        RECT 19.655 116.370 20.165 116.905 ;
        RECT 20.385 116.095 20.630 116.700 ;
        RECT 21.075 116.135 22.745 116.905 ;
        RECT 22.915 116.180 23.205 116.905 ;
        RECT 23.375 116.155 24.585 116.905 ;
        RECT 24.760 116.360 30.105 116.905 ;
        RECT 19.675 115.925 20.905 116.095 ;
        RECT 18.465 115.205 19.475 115.375 ;
        RECT 19.645 115.360 20.395 115.550 ;
        RECT 18.125 114.865 19.250 115.035 ;
        RECT 19.645 114.695 19.815 115.360 ;
        RECT 20.565 115.115 20.905 115.925 ;
        RECT 17.785 114.525 19.815 114.695 ;
        RECT 19.985 114.355 20.155 115.115 ;
        RECT 20.390 114.705 20.905 115.115 ;
        RECT 21.075 115.445 21.825 115.965 ;
        RECT 21.995 115.615 22.745 116.135 ;
        RECT 21.075 114.355 22.745 115.445 ;
        RECT 22.915 114.355 23.205 115.520 ;
        RECT 23.375 115.445 23.895 115.985 ;
        RECT 24.065 115.615 24.585 116.155 ;
        RECT 23.375 114.355 24.585 115.445 ;
        RECT 26.350 114.790 26.700 116.040 ;
        RECT 28.180 115.530 28.520 116.360 ;
        RECT 30.335 116.085 30.545 116.905 ;
        RECT 30.715 116.105 31.045 116.735 ;
        RECT 30.715 115.505 30.965 116.105 ;
        RECT 31.215 116.085 31.445 116.905 ;
        RECT 32.120 116.360 37.465 116.905 ;
        RECT 37.640 116.360 42.985 116.905 ;
        RECT 31.135 115.665 31.465 115.915 ;
        RECT 24.760 114.355 30.105 114.790 ;
        RECT 30.335 114.355 30.545 115.495 ;
        RECT 30.715 114.525 31.045 115.505 ;
        RECT 31.215 114.355 31.445 115.495 ;
        RECT 33.710 114.790 34.060 116.040 ;
        RECT 35.540 115.530 35.880 116.360 ;
        RECT 39.230 114.790 39.580 116.040 ;
        RECT 41.060 115.530 41.400 116.360 ;
        RECT 43.215 116.085 43.425 116.905 ;
        RECT 43.595 116.105 43.925 116.735 ;
        RECT 43.595 115.505 43.845 116.105 ;
        RECT 44.095 116.085 44.325 116.905 ;
        RECT 44.995 116.135 48.505 116.905 ;
        RECT 48.675 116.180 48.965 116.905 ;
        RECT 49.225 116.355 49.395 116.645 ;
        RECT 49.565 116.525 49.895 116.905 ;
        RECT 49.225 116.185 49.890 116.355 ;
        RECT 44.015 115.665 44.345 115.915 ;
        RECT 32.120 114.355 37.465 114.790 ;
        RECT 37.640 114.355 42.985 114.790 ;
        RECT 43.215 114.355 43.425 115.495 ;
        RECT 43.595 114.525 43.925 115.505 ;
        RECT 44.095 114.355 44.325 115.495 ;
        RECT 44.995 115.445 46.685 115.965 ;
        RECT 46.855 115.615 48.505 116.135 ;
        RECT 44.995 114.355 48.505 115.445 ;
        RECT 48.675 114.355 48.965 115.520 ;
        RECT 49.140 115.365 49.490 116.015 ;
        RECT 49.660 115.195 49.890 116.185 ;
        RECT 49.225 115.025 49.890 115.195 ;
        RECT 49.225 114.525 49.395 115.025 ;
        RECT 49.565 114.355 49.895 114.855 ;
        RECT 50.065 114.525 50.290 116.645 ;
        RECT 50.505 116.525 50.835 116.905 ;
        RECT 51.005 116.355 51.175 116.685 ;
        RECT 51.475 116.525 52.490 116.725 ;
        RECT 50.480 116.165 51.175 116.355 ;
        RECT 50.480 115.195 50.650 116.165 ;
        RECT 50.820 115.365 51.230 115.985 ;
        RECT 51.400 115.415 51.620 116.285 ;
        RECT 51.800 115.975 52.150 116.345 ;
        RECT 52.320 115.795 52.490 116.525 ;
        RECT 52.660 116.465 53.070 116.905 ;
        RECT 53.360 116.265 53.610 116.695 ;
        RECT 53.810 116.445 54.130 116.905 ;
        RECT 54.690 116.515 55.540 116.685 ;
        RECT 52.660 115.925 53.070 116.255 ;
        RECT 53.360 115.925 53.780 116.265 ;
        RECT 52.070 115.755 52.490 115.795 ;
        RECT 52.070 115.585 53.420 115.755 ;
        RECT 50.480 115.025 51.175 115.195 ;
        RECT 51.400 115.035 51.900 115.415 ;
        RECT 50.505 114.355 50.835 114.855 ;
        RECT 51.005 114.525 51.175 115.025 ;
        RECT 52.070 114.740 52.240 115.585 ;
        RECT 53.170 115.425 53.420 115.585 ;
        RECT 52.410 115.155 52.660 115.415 ;
        RECT 53.590 115.155 53.780 115.925 ;
        RECT 52.410 114.905 53.780 115.155 ;
        RECT 53.950 116.095 55.200 116.265 ;
        RECT 53.950 115.335 54.120 116.095 ;
        RECT 54.870 115.975 55.200 116.095 ;
        RECT 54.290 115.515 54.470 115.925 ;
        RECT 55.370 115.755 55.540 116.515 ;
        RECT 55.740 116.425 56.400 116.905 ;
        RECT 56.580 116.310 56.900 116.640 ;
        RECT 55.730 115.985 56.390 116.255 ;
        RECT 55.730 115.925 56.060 115.985 ;
        RECT 56.210 115.755 56.540 115.815 ;
        RECT 54.640 115.585 56.540 115.755 ;
        RECT 53.950 115.025 54.470 115.335 ;
        RECT 54.640 115.075 54.810 115.585 ;
        RECT 56.710 115.415 56.900 116.310 ;
        RECT 54.980 115.245 56.900 115.415 ;
        RECT 56.580 115.225 56.900 115.245 ;
        RECT 57.100 115.995 57.350 116.645 ;
        RECT 57.530 116.445 57.815 116.905 ;
        RECT 57.995 116.565 58.250 116.725 ;
        RECT 57.995 116.395 58.335 116.565 ;
        RECT 57.995 116.195 58.250 116.395 ;
        RECT 57.100 115.665 57.900 115.995 ;
        RECT 54.640 114.905 55.850 115.075 ;
        RECT 51.410 114.570 52.240 114.740 ;
        RECT 52.480 114.355 52.860 114.735 ;
        RECT 53.040 114.615 53.210 114.905 ;
        RECT 54.640 114.825 54.810 114.905 ;
        RECT 53.380 114.355 53.710 114.735 ;
        RECT 54.180 114.575 54.810 114.825 ;
        RECT 54.990 114.355 55.410 114.735 ;
        RECT 55.610 114.615 55.850 114.905 ;
        RECT 56.080 114.355 56.410 115.045 ;
        RECT 56.580 114.615 56.750 115.225 ;
        RECT 57.100 115.075 57.350 115.665 ;
        RECT 58.070 115.335 58.250 116.195 ;
        RECT 59.715 116.135 63.225 116.905 ;
        RECT 63.400 116.360 68.745 116.905 ;
        RECT 68.920 116.360 74.265 116.905 ;
        RECT 57.020 114.565 57.350 115.075 ;
        RECT 57.530 114.355 57.815 115.155 ;
        RECT 57.995 114.665 58.250 115.335 ;
        RECT 59.715 115.445 61.405 115.965 ;
        RECT 61.575 115.615 63.225 116.135 ;
        RECT 59.715 114.355 63.225 115.445 ;
        RECT 64.990 114.790 65.340 116.040 ;
        RECT 66.820 115.530 67.160 116.360 ;
        RECT 70.510 114.790 70.860 116.040 ;
        RECT 72.340 115.530 72.680 116.360 ;
        RECT 74.435 116.180 74.725 116.905 ;
        RECT 75.815 116.135 79.325 116.905 ;
        RECT 79.500 116.360 84.845 116.905 ;
        RECT 85.020 116.360 90.365 116.905 ;
        RECT 90.540 116.360 95.885 116.905 ;
        RECT 63.400 114.355 68.745 114.790 ;
        RECT 68.920 114.355 74.265 114.790 ;
        RECT 74.435 114.355 74.725 115.520 ;
        RECT 75.815 115.445 77.505 115.965 ;
        RECT 77.675 115.615 79.325 116.135 ;
        RECT 75.815 114.355 79.325 115.445 ;
        RECT 81.090 114.790 81.440 116.040 ;
        RECT 82.920 115.530 83.260 116.360 ;
        RECT 86.610 114.790 86.960 116.040 ;
        RECT 88.440 115.530 88.780 116.360 ;
        RECT 92.130 114.790 92.480 116.040 ;
        RECT 93.960 115.530 94.300 116.360 ;
        RECT 96.145 116.355 96.315 116.735 ;
        RECT 96.495 116.525 96.825 116.905 ;
        RECT 96.145 116.185 96.810 116.355 ;
        RECT 97.005 116.230 97.265 116.735 ;
        RECT 96.075 115.635 96.405 116.005 ;
        RECT 96.640 115.930 96.810 116.185 ;
        RECT 96.640 115.600 96.925 115.930 ;
        RECT 96.640 115.455 96.810 115.600 ;
        RECT 96.145 115.285 96.810 115.455 ;
        RECT 97.095 115.430 97.265 116.230 ;
        RECT 97.435 116.135 100.025 116.905 ;
        RECT 100.195 116.180 100.485 116.905 ;
        RECT 100.655 116.135 104.165 116.905 ;
        RECT 79.500 114.355 84.845 114.790 ;
        RECT 85.020 114.355 90.365 114.790 ;
        RECT 90.540 114.355 95.885 114.790 ;
        RECT 96.145 114.525 96.315 115.285 ;
        RECT 96.495 114.355 96.825 115.115 ;
        RECT 96.995 114.525 97.265 115.430 ;
        RECT 97.435 115.445 98.645 115.965 ;
        RECT 98.815 115.615 100.025 116.135 ;
        RECT 97.435 114.355 100.025 115.445 ;
        RECT 100.195 114.355 100.485 115.520 ;
        RECT 100.655 115.445 102.345 115.965 ;
        RECT 102.515 115.615 104.165 116.135 ;
        RECT 104.335 116.230 104.595 116.735 ;
        RECT 104.775 116.525 105.105 116.905 ;
        RECT 105.285 116.355 105.455 116.735 ;
        RECT 100.655 114.355 104.165 115.445 ;
        RECT 104.335 115.430 104.505 116.230 ;
        RECT 104.790 116.185 105.455 116.355 ;
        RECT 104.790 115.930 104.960 116.185 ;
        RECT 105.755 116.085 105.985 116.905 ;
        RECT 106.155 116.105 106.485 116.735 ;
        RECT 104.675 115.600 104.960 115.930 ;
        RECT 105.195 115.635 105.525 116.005 ;
        RECT 105.735 115.665 106.065 115.915 ;
        RECT 104.790 115.455 104.960 115.600 ;
        RECT 106.235 115.505 106.485 116.105 ;
        RECT 106.655 116.085 106.865 116.905 ;
        RECT 108.015 116.230 108.275 116.735 ;
        RECT 108.455 116.525 108.785 116.905 ;
        RECT 108.965 116.355 109.135 116.735 ;
        RECT 104.335 114.525 104.605 115.430 ;
        RECT 104.790 115.285 105.455 115.455 ;
        RECT 104.775 114.355 105.105 115.115 ;
        RECT 105.285 114.525 105.455 115.285 ;
        RECT 105.755 114.355 105.985 115.495 ;
        RECT 106.155 114.525 106.485 115.505 ;
        RECT 106.655 114.355 106.865 115.495 ;
        RECT 108.015 115.430 108.185 116.230 ;
        RECT 108.470 116.185 109.135 116.355 ;
        RECT 108.470 115.930 108.640 116.185 ;
        RECT 109.395 116.135 111.985 116.905 ;
        RECT 112.155 116.155 113.365 116.905 ;
        RECT 108.355 115.600 108.640 115.930 ;
        RECT 108.875 115.635 109.205 116.005 ;
        RECT 108.470 115.455 108.640 115.600 ;
        RECT 108.015 114.525 108.285 115.430 ;
        RECT 108.470 115.285 109.135 115.455 ;
        RECT 108.455 114.355 108.785 115.115 ;
        RECT 108.965 114.525 109.135 115.285 ;
        RECT 109.395 115.445 110.605 115.965 ;
        RECT 110.775 115.615 111.985 116.135 ;
        RECT 112.155 115.445 112.675 115.985 ;
        RECT 112.845 115.615 113.365 116.155 ;
        RECT 109.395 114.355 111.985 115.445 ;
        RECT 112.155 114.355 113.365 115.445 ;
        RECT 11.330 114.185 113.450 114.355 ;
        RECT 11.415 113.095 12.625 114.185 ;
        RECT 11.415 112.385 11.935 112.925 ;
        RECT 12.105 112.555 12.625 113.095 ;
        RECT 12.795 113.095 14.005 114.185 ;
        RECT 14.485 113.345 14.655 114.185 ;
        RECT 14.865 113.175 15.115 114.015 ;
        RECT 15.325 113.345 15.495 114.185 ;
        RECT 15.665 113.175 15.955 114.015 ;
        RECT 12.795 112.555 13.315 113.095 ;
        RECT 14.230 113.005 15.955 113.175 ;
        RECT 16.165 113.125 16.335 114.185 ;
        RECT 16.630 113.805 16.960 114.185 ;
        RECT 17.140 113.635 17.310 113.925 ;
        RECT 17.480 113.725 17.730 114.185 ;
        RECT 16.510 113.465 17.310 113.635 ;
        RECT 17.900 113.675 18.770 114.015 ;
        RECT 13.485 112.385 14.005 112.925 ;
        RECT 11.415 111.635 12.625 112.385 ;
        RECT 12.795 111.635 14.005 112.385 ;
        RECT 14.230 112.455 14.640 113.005 ;
        RECT 16.510 112.845 16.680 113.465 ;
        RECT 17.900 113.295 18.070 113.675 ;
        RECT 19.005 113.555 19.175 114.015 ;
        RECT 19.345 113.725 19.715 114.185 ;
        RECT 20.010 113.585 20.180 113.925 ;
        RECT 20.350 113.755 20.680 114.185 ;
        RECT 20.915 113.585 21.085 113.925 ;
        RECT 16.850 113.125 18.070 113.295 ;
        RECT 18.240 113.215 18.700 113.505 ;
        RECT 19.005 113.385 19.565 113.555 ;
        RECT 20.010 113.415 21.085 113.585 ;
        RECT 21.255 113.685 21.935 114.015 ;
        RECT 22.150 113.685 22.400 114.015 ;
        RECT 22.570 113.725 22.820 114.185 ;
        RECT 19.395 113.245 19.565 113.385 ;
        RECT 18.240 113.205 19.205 113.215 ;
        RECT 17.900 113.035 18.070 113.125 ;
        RECT 18.530 113.045 19.205 113.205 ;
        RECT 16.510 112.835 16.855 112.845 ;
        RECT 14.825 112.625 16.855 112.835 ;
        RECT 14.230 112.285 15.995 112.455 ;
        RECT 14.485 111.635 14.655 112.105 ;
        RECT 14.825 111.805 15.155 112.285 ;
        RECT 15.325 111.635 15.495 112.105 ;
        RECT 15.665 111.805 15.995 112.285 ;
        RECT 16.165 111.635 16.335 112.445 ;
        RECT 16.530 112.370 16.855 112.625 ;
        RECT 16.535 112.015 16.855 112.370 ;
        RECT 17.025 112.585 17.565 112.955 ;
        RECT 17.900 112.865 18.305 113.035 ;
        RECT 17.025 112.185 17.265 112.585 ;
        RECT 17.745 112.415 17.965 112.695 ;
        RECT 17.435 112.245 17.965 112.415 ;
        RECT 17.435 112.015 17.605 112.245 ;
        RECT 18.135 112.085 18.305 112.865 ;
        RECT 18.475 112.255 18.825 112.875 ;
        RECT 18.995 112.255 19.205 113.045 ;
        RECT 19.395 113.075 20.895 113.245 ;
        RECT 19.395 112.385 19.565 113.075 ;
        RECT 21.255 112.905 21.425 113.685 ;
        RECT 22.230 113.555 22.400 113.685 ;
        RECT 19.735 112.735 21.425 112.905 ;
        RECT 21.595 113.125 22.060 113.515 ;
        RECT 22.230 113.385 22.625 113.555 ;
        RECT 19.735 112.555 19.905 112.735 ;
        RECT 16.535 111.845 17.605 112.015 ;
        RECT 17.775 111.635 17.965 112.075 ;
        RECT 18.135 111.805 19.085 112.085 ;
        RECT 19.395 111.995 19.655 112.385 ;
        RECT 20.075 112.315 20.865 112.565 ;
        RECT 19.305 111.825 19.655 111.995 ;
        RECT 19.865 111.635 20.195 112.095 ;
        RECT 21.070 112.025 21.240 112.735 ;
        RECT 21.595 112.535 21.765 113.125 ;
        RECT 21.410 112.315 21.765 112.535 ;
        RECT 21.935 112.315 22.285 112.935 ;
        RECT 22.455 112.025 22.625 113.385 ;
        RECT 22.990 113.215 23.315 114.000 ;
        RECT 22.795 112.165 23.255 113.215 ;
        RECT 21.070 111.855 21.925 112.025 ;
        RECT 22.130 111.855 22.625 112.025 ;
        RECT 22.795 111.635 23.125 111.995 ;
        RECT 23.485 111.895 23.655 114.015 ;
        RECT 23.825 113.685 24.155 114.185 ;
        RECT 24.325 113.515 24.580 114.015 ;
        RECT 23.830 113.345 24.580 113.515 ;
        RECT 23.830 112.355 24.060 113.345 ;
        RECT 24.230 112.525 24.580 113.175 ;
        RECT 24.755 113.095 27.345 114.185 ;
        RECT 24.755 112.575 25.965 113.095 ;
        RECT 27.575 113.045 27.785 114.185 ;
        RECT 27.955 113.035 28.285 114.015 ;
        RECT 28.455 113.045 28.685 114.185 ;
        RECT 28.895 113.095 30.105 114.185 ;
        RECT 30.280 113.750 35.625 114.185 ;
        RECT 26.135 112.405 27.345 112.925 ;
        RECT 23.830 112.185 24.580 112.355 ;
        RECT 23.825 111.635 24.155 112.015 ;
        RECT 24.325 111.895 24.580 112.185 ;
        RECT 24.755 111.635 27.345 112.405 ;
        RECT 27.575 111.635 27.785 112.455 ;
        RECT 27.955 112.435 28.205 113.035 ;
        RECT 28.375 112.625 28.705 112.875 ;
        RECT 28.895 112.555 29.415 113.095 ;
        RECT 27.955 111.805 28.285 112.435 ;
        RECT 28.455 111.635 28.685 112.455 ;
        RECT 29.585 112.385 30.105 112.925 ;
        RECT 31.870 112.500 32.220 113.750 ;
        RECT 35.795 113.020 36.085 114.185 ;
        RECT 36.255 113.110 36.525 114.015 ;
        RECT 36.695 113.425 37.025 114.185 ;
        RECT 37.205 113.255 37.375 114.015 ;
        RECT 28.895 111.635 30.105 112.385 ;
        RECT 33.700 112.180 34.040 113.010 ;
        RECT 30.280 111.635 35.625 112.180 ;
        RECT 35.795 111.635 36.085 112.360 ;
        RECT 36.255 112.310 36.425 113.110 ;
        RECT 36.710 113.085 37.375 113.255 ;
        RECT 38.095 113.095 39.765 114.185 ;
        RECT 39.935 113.110 40.205 114.015 ;
        RECT 40.375 113.425 40.705 114.185 ;
        RECT 40.885 113.255 41.055 114.015 ;
        RECT 36.710 112.940 36.880 113.085 ;
        RECT 36.595 112.610 36.880 112.940 ;
        RECT 36.710 112.355 36.880 112.610 ;
        RECT 37.115 112.535 37.445 112.905 ;
        RECT 38.095 112.575 38.845 113.095 ;
        RECT 39.015 112.405 39.765 112.925 ;
        RECT 36.255 111.805 36.515 112.310 ;
        RECT 36.710 112.185 37.375 112.355 ;
        RECT 36.695 111.635 37.025 112.015 ;
        RECT 37.205 111.805 37.375 112.185 ;
        RECT 38.095 111.635 39.765 112.405 ;
        RECT 39.935 112.310 40.105 113.110 ;
        RECT 40.390 113.085 41.055 113.255 ;
        RECT 41.315 113.095 43.905 114.185 ;
        RECT 44.165 113.255 44.335 114.015 ;
        RECT 44.515 113.425 44.845 114.185 ;
        RECT 40.390 112.940 40.560 113.085 ;
        RECT 40.275 112.610 40.560 112.940 ;
        RECT 40.390 112.355 40.560 112.610 ;
        RECT 40.795 112.535 41.125 112.905 ;
        RECT 41.315 112.575 42.525 113.095 ;
        RECT 44.165 113.085 44.830 113.255 ;
        RECT 45.015 113.110 45.285 114.015 ;
        RECT 44.660 112.940 44.830 113.085 ;
        RECT 42.695 112.405 43.905 112.925 ;
        RECT 44.095 112.535 44.425 112.905 ;
        RECT 44.660 112.610 44.945 112.940 ;
        RECT 39.935 111.805 40.195 112.310 ;
        RECT 40.390 112.185 41.055 112.355 ;
        RECT 40.375 111.635 40.705 112.015 ;
        RECT 40.885 111.805 41.055 112.185 ;
        RECT 41.315 111.635 43.905 112.405 ;
        RECT 44.660 112.355 44.830 112.610 ;
        RECT 44.165 112.185 44.830 112.355 ;
        RECT 45.115 112.310 45.285 113.110 ;
        RECT 46.375 113.095 49.885 114.185 ;
        RECT 46.375 112.575 48.065 113.095 ;
        RECT 50.095 113.045 50.325 114.185 ;
        RECT 50.495 113.035 50.825 114.015 ;
        RECT 50.995 113.045 51.205 114.185 ;
        RECT 51.445 113.205 51.775 114.015 ;
        RECT 51.945 113.385 52.185 114.185 ;
        RECT 51.445 113.035 52.160 113.205 ;
        RECT 48.235 112.405 49.885 112.925 ;
        RECT 50.075 112.625 50.405 112.875 ;
        RECT 44.165 111.805 44.335 112.185 ;
        RECT 44.515 111.635 44.845 112.015 ;
        RECT 45.025 111.805 45.285 112.310 ;
        RECT 46.375 111.635 49.885 112.405 ;
        RECT 50.095 111.635 50.325 112.455 ;
        RECT 50.575 112.435 50.825 113.035 ;
        RECT 51.440 112.625 51.820 112.865 ;
        RECT 51.990 112.795 52.160 113.035 ;
        RECT 52.365 113.165 52.535 114.015 ;
        RECT 52.705 113.385 53.035 114.185 ;
        RECT 53.205 113.165 53.375 114.015 ;
        RECT 52.365 112.995 53.375 113.165 ;
        RECT 53.545 113.035 53.875 114.185 ;
        RECT 54.195 113.095 56.785 114.185 ;
        RECT 57.045 113.255 57.215 114.015 ;
        RECT 57.395 113.425 57.725 114.185 ;
        RECT 51.990 112.625 52.490 112.795 ;
        RECT 51.990 112.455 52.160 112.625 ;
        RECT 52.880 112.485 53.375 112.995 ;
        RECT 54.195 112.575 55.405 113.095 ;
        RECT 57.045 113.085 57.710 113.255 ;
        RECT 57.895 113.110 58.165 114.015 ;
        RECT 57.540 112.940 57.710 113.085 ;
        RECT 52.875 112.455 53.375 112.485 ;
        RECT 50.495 111.805 50.825 112.435 ;
        RECT 50.995 111.635 51.205 112.455 ;
        RECT 51.525 112.285 52.160 112.455 ;
        RECT 52.365 112.285 53.375 112.455 ;
        RECT 51.525 111.805 51.695 112.285 ;
        RECT 51.875 111.635 52.115 112.115 ;
        RECT 52.365 111.805 52.535 112.285 ;
        RECT 52.705 111.635 53.035 112.115 ;
        RECT 53.205 111.805 53.375 112.285 ;
        RECT 53.545 111.635 53.875 112.435 ;
        RECT 55.575 112.405 56.785 112.925 ;
        RECT 56.975 112.535 57.305 112.905 ;
        RECT 57.540 112.610 57.825 112.940 ;
        RECT 54.195 111.635 56.785 112.405 ;
        RECT 57.540 112.355 57.710 112.610 ;
        RECT 57.045 112.185 57.710 112.355 ;
        RECT 57.995 112.310 58.165 113.110 ;
        RECT 58.335 113.095 60.005 114.185 ;
        RECT 60.265 113.255 60.435 114.015 ;
        RECT 60.615 113.425 60.945 114.185 ;
        RECT 58.335 112.575 59.085 113.095 ;
        RECT 60.265 113.085 60.930 113.255 ;
        RECT 61.115 113.110 61.385 114.015 ;
        RECT 60.760 112.940 60.930 113.085 ;
        RECT 59.255 112.405 60.005 112.925 ;
        RECT 60.195 112.535 60.525 112.905 ;
        RECT 60.760 112.610 61.045 112.940 ;
        RECT 57.045 111.805 57.215 112.185 ;
        RECT 57.395 111.635 57.725 112.015 ;
        RECT 57.905 111.805 58.165 112.310 ;
        RECT 58.335 111.635 60.005 112.405 ;
        RECT 60.760 112.355 60.930 112.610 ;
        RECT 60.265 112.185 60.930 112.355 ;
        RECT 61.215 112.310 61.385 113.110 ;
        RECT 61.555 113.020 61.845 114.185 ;
        RECT 62.935 113.095 66.445 114.185 ;
        RECT 62.935 112.575 64.625 113.095 ;
        RECT 66.675 113.045 66.885 114.185 ;
        RECT 67.055 113.035 67.385 114.015 ;
        RECT 67.555 113.045 67.785 114.185 ;
        RECT 67.995 113.110 68.265 114.015 ;
        RECT 68.435 113.425 68.765 114.185 ;
        RECT 68.945 113.255 69.115 114.015 ;
        RECT 64.795 112.405 66.445 112.925 ;
        RECT 60.265 111.805 60.435 112.185 ;
        RECT 60.615 111.635 60.945 112.015 ;
        RECT 61.125 111.805 61.385 112.310 ;
        RECT 61.555 111.635 61.845 112.360 ;
        RECT 62.935 111.635 66.445 112.405 ;
        RECT 66.675 111.635 66.885 112.455 ;
        RECT 67.055 112.435 67.305 113.035 ;
        RECT 67.475 112.625 67.805 112.875 ;
        RECT 67.055 111.805 67.385 112.435 ;
        RECT 67.555 111.635 67.785 112.455 ;
        RECT 67.995 112.310 68.165 113.110 ;
        RECT 68.450 113.085 69.115 113.255 ;
        RECT 68.450 112.940 68.620 113.085 ;
        RECT 69.435 113.045 69.645 114.185 ;
        RECT 68.335 112.610 68.620 112.940 ;
        RECT 69.815 113.035 70.145 114.015 ;
        RECT 70.315 113.045 70.545 114.185 ;
        RECT 70.765 113.205 71.095 114.015 ;
        RECT 71.265 113.385 71.505 114.185 ;
        RECT 70.765 113.035 71.480 113.205 ;
        RECT 68.450 112.355 68.620 112.610 ;
        RECT 68.855 112.535 69.185 112.905 ;
        RECT 67.995 111.805 68.255 112.310 ;
        RECT 68.450 112.185 69.115 112.355 ;
        RECT 68.435 111.635 68.765 112.015 ;
        RECT 68.945 111.805 69.115 112.185 ;
        RECT 69.435 111.635 69.645 112.455 ;
        RECT 69.815 112.435 70.065 113.035 ;
        RECT 70.235 112.625 70.565 112.875 ;
        RECT 70.760 112.625 71.140 112.865 ;
        RECT 71.310 112.795 71.480 113.035 ;
        RECT 71.685 113.165 71.855 114.015 ;
        RECT 72.025 113.385 72.355 114.185 ;
        RECT 72.525 113.165 72.695 114.015 ;
        RECT 71.685 112.995 72.695 113.165 ;
        RECT 72.865 113.035 73.195 114.185 ;
        RECT 73.975 113.095 77.485 114.185 ;
        RECT 77.660 113.750 83.005 114.185 ;
        RECT 71.310 112.625 71.810 112.795 ;
        RECT 71.310 112.455 71.480 112.625 ;
        RECT 72.200 112.455 72.695 112.995 ;
        RECT 73.975 112.575 75.665 113.095 ;
        RECT 69.815 111.805 70.145 112.435 ;
        RECT 70.315 111.635 70.545 112.455 ;
        RECT 70.845 112.285 71.480 112.455 ;
        RECT 71.685 112.285 72.695 112.455 ;
        RECT 70.845 111.805 71.015 112.285 ;
        RECT 71.195 111.635 71.435 112.115 ;
        RECT 71.685 111.805 71.855 112.285 ;
        RECT 72.025 111.635 72.355 112.115 ;
        RECT 72.525 111.805 72.695 112.285 ;
        RECT 72.865 111.635 73.195 112.435 ;
        RECT 75.835 112.405 77.485 112.925 ;
        RECT 79.250 112.500 79.600 113.750 ;
        RECT 83.265 113.255 83.435 114.015 ;
        RECT 83.615 113.425 83.945 114.185 ;
        RECT 83.265 113.085 83.930 113.255 ;
        RECT 84.115 113.110 84.385 114.015 ;
        RECT 73.975 111.635 77.485 112.405 ;
        RECT 81.080 112.180 81.420 113.010 ;
        RECT 83.760 112.940 83.930 113.085 ;
        RECT 83.195 112.535 83.525 112.905 ;
        RECT 83.760 112.610 84.045 112.940 ;
        RECT 83.760 112.355 83.930 112.610 ;
        RECT 83.265 112.185 83.930 112.355 ;
        RECT 84.215 112.310 84.385 113.110 ;
        RECT 84.555 113.095 87.145 114.185 ;
        RECT 84.555 112.575 85.765 113.095 ;
        RECT 87.315 113.020 87.605 114.185 ;
        RECT 88.325 113.255 88.495 114.015 ;
        RECT 88.675 113.425 89.005 114.185 ;
        RECT 88.325 113.085 88.990 113.255 ;
        RECT 89.175 113.110 89.445 114.015 ;
        RECT 88.820 112.940 88.990 113.085 ;
        RECT 85.935 112.405 87.145 112.925 ;
        RECT 88.255 112.535 88.585 112.905 ;
        RECT 88.820 112.610 89.105 112.940 ;
        RECT 77.660 111.635 83.005 112.180 ;
        RECT 83.265 111.805 83.435 112.185 ;
        RECT 83.615 111.635 83.945 112.015 ;
        RECT 84.125 111.805 84.385 112.310 ;
        RECT 84.555 111.635 87.145 112.405 ;
        RECT 87.315 111.635 87.605 112.360 ;
        RECT 88.820 112.355 88.990 112.610 ;
        RECT 88.325 112.185 88.990 112.355 ;
        RECT 89.275 112.310 89.445 113.110 ;
        RECT 90.075 113.095 93.585 114.185 ;
        RECT 93.845 113.255 94.015 114.015 ;
        RECT 94.195 113.425 94.525 114.185 ;
        RECT 90.075 112.575 91.765 113.095 ;
        RECT 93.845 113.085 94.510 113.255 ;
        RECT 94.695 113.110 94.965 114.015 ;
        RECT 94.340 112.940 94.510 113.085 ;
        RECT 91.935 112.405 93.585 112.925 ;
        RECT 93.775 112.535 94.105 112.905 ;
        RECT 94.340 112.610 94.625 112.940 ;
        RECT 88.325 111.805 88.495 112.185 ;
        RECT 88.675 111.635 89.005 112.015 ;
        RECT 89.185 111.805 89.445 112.310 ;
        RECT 90.075 111.635 93.585 112.405 ;
        RECT 94.340 112.355 94.510 112.610 ;
        RECT 93.845 112.185 94.510 112.355 ;
        RECT 94.795 112.310 94.965 113.110 ;
        RECT 96.145 113.255 96.315 114.015 ;
        RECT 96.495 113.425 96.825 114.185 ;
        RECT 96.145 113.085 96.810 113.255 ;
        RECT 96.995 113.110 97.265 114.015 ;
        RECT 96.640 112.940 96.810 113.085 ;
        RECT 96.075 112.535 96.405 112.905 ;
        RECT 96.640 112.610 96.925 112.940 ;
        RECT 96.640 112.355 96.810 112.610 ;
        RECT 93.845 111.805 94.015 112.185 ;
        RECT 94.195 111.635 94.525 112.015 ;
        RECT 94.705 111.805 94.965 112.310 ;
        RECT 96.145 112.185 96.810 112.355 ;
        RECT 97.095 112.310 97.265 113.110 ;
        RECT 96.145 111.805 96.315 112.185 ;
        RECT 96.495 111.635 96.825 112.015 ;
        RECT 97.005 111.805 97.265 112.310 ;
        RECT 97.435 113.110 97.705 114.015 ;
        RECT 97.875 113.425 98.205 114.185 ;
        RECT 98.385 113.255 98.555 114.015 ;
        RECT 97.435 112.310 97.605 113.110 ;
        RECT 97.890 113.085 98.555 113.255 ;
        RECT 98.815 113.095 101.405 114.185 ;
        RECT 101.580 113.515 101.835 114.015 ;
        RECT 102.005 113.685 102.335 114.185 ;
        RECT 101.580 113.345 102.330 113.515 ;
        RECT 97.890 112.940 98.060 113.085 ;
        RECT 97.775 112.610 98.060 112.940 ;
        RECT 97.890 112.355 98.060 112.610 ;
        RECT 98.295 112.535 98.625 112.905 ;
        RECT 98.815 112.575 100.025 113.095 ;
        RECT 100.195 112.405 101.405 112.925 ;
        RECT 101.580 112.525 101.930 113.175 ;
        RECT 97.435 111.805 97.695 112.310 ;
        RECT 97.890 112.185 98.555 112.355 ;
        RECT 97.875 111.635 98.205 112.015 ;
        RECT 98.385 111.805 98.555 112.185 ;
        RECT 98.815 111.635 101.405 112.405 ;
        RECT 102.100 112.355 102.330 113.345 ;
        RECT 101.580 112.185 102.330 112.355 ;
        RECT 101.580 111.895 101.835 112.185 ;
        RECT 102.005 111.635 102.335 112.015 ;
        RECT 102.505 111.895 102.675 114.015 ;
        RECT 102.845 113.215 103.170 114.000 ;
        RECT 103.340 113.725 103.590 114.185 ;
        RECT 103.760 113.685 104.010 114.015 ;
        RECT 104.225 113.685 104.905 114.015 ;
        RECT 103.760 113.555 103.930 113.685 ;
        RECT 103.535 113.385 103.930 113.555 ;
        RECT 102.905 112.165 103.365 113.215 ;
        RECT 103.535 112.025 103.705 113.385 ;
        RECT 104.100 113.125 104.565 113.515 ;
        RECT 103.875 112.315 104.225 112.935 ;
        RECT 104.395 112.535 104.565 113.125 ;
        RECT 104.735 112.905 104.905 113.685 ;
        RECT 105.075 113.585 105.245 113.925 ;
        RECT 105.480 113.755 105.810 114.185 ;
        RECT 105.980 113.585 106.150 113.925 ;
        RECT 106.445 113.725 106.815 114.185 ;
        RECT 105.075 113.415 106.150 113.585 ;
        RECT 106.985 113.555 107.155 114.015 ;
        RECT 107.390 113.675 108.260 114.015 ;
        RECT 108.430 113.725 108.680 114.185 ;
        RECT 106.595 113.385 107.155 113.555 ;
        RECT 106.595 113.245 106.765 113.385 ;
        RECT 105.265 113.075 106.765 113.245 ;
        RECT 107.460 113.215 107.920 113.505 ;
        RECT 104.735 112.735 106.425 112.905 ;
        RECT 104.395 112.315 104.750 112.535 ;
        RECT 104.920 112.025 105.090 112.735 ;
        RECT 105.295 112.315 106.085 112.565 ;
        RECT 106.255 112.555 106.425 112.735 ;
        RECT 106.595 112.385 106.765 113.075 ;
        RECT 103.035 111.635 103.365 111.995 ;
        RECT 103.535 111.855 104.030 112.025 ;
        RECT 104.235 111.855 105.090 112.025 ;
        RECT 105.965 111.635 106.295 112.095 ;
        RECT 106.505 111.995 106.765 112.385 ;
        RECT 106.955 113.205 107.920 113.215 ;
        RECT 108.090 113.295 108.260 113.675 ;
        RECT 108.850 113.635 109.020 113.925 ;
        RECT 109.200 113.805 109.530 114.185 ;
        RECT 108.850 113.465 109.650 113.635 ;
        RECT 106.955 113.045 107.630 113.205 ;
        RECT 108.090 113.125 109.310 113.295 ;
        RECT 106.955 112.255 107.165 113.045 ;
        RECT 108.090 113.035 108.260 113.125 ;
        RECT 107.335 112.255 107.685 112.875 ;
        RECT 107.855 112.865 108.260 113.035 ;
        RECT 107.855 112.085 108.025 112.865 ;
        RECT 108.195 112.415 108.415 112.695 ;
        RECT 108.595 112.585 109.135 112.955 ;
        RECT 109.480 112.845 109.650 113.465 ;
        RECT 109.825 113.125 109.995 114.185 ;
        RECT 110.205 113.175 110.495 114.015 ;
        RECT 110.665 113.345 110.835 114.185 ;
        RECT 111.045 113.175 111.295 114.015 ;
        RECT 111.505 113.345 111.675 114.185 ;
        RECT 110.205 113.005 111.930 113.175 ;
        RECT 108.195 112.245 108.725 112.415 ;
        RECT 106.505 111.825 106.855 111.995 ;
        RECT 107.075 111.805 108.025 112.085 ;
        RECT 108.195 111.635 108.385 112.075 ;
        RECT 108.555 112.015 108.725 112.245 ;
        RECT 108.895 112.185 109.135 112.585 ;
        RECT 109.305 112.835 109.650 112.845 ;
        RECT 109.305 112.625 111.335 112.835 ;
        RECT 109.305 112.370 109.630 112.625 ;
        RECT 111.520 112.455 111.930 113.005 ;
        RECT 112.155 113.095 113.365 114.185 ;
        RECT 112.155 112.555 112.675 113.095 ;
        RECT 109.305 112.015 109.625 112.370 ;
        RECT 108.555 111.845 109.625 112.015 ;
        RECT 109.825 111.635 109.995 112.445 ;
        RECT 110.165 112.285 111.930 112.455 ;
        RECT 112.845 112.385 113.365 112.925 ;
        RECT 110.165 111.805 110.495 112.285 ;
        RECT 110.665 111.635 110.835 112.105 ;
        RECT 111.005 111.805 111.335 112.285 ;
        RECT 111.505 111.635 111.675 112.105 ;
        RECT 112.155 111.635 113.365 112.385 ;
        RECT 11.330 111.465 113.450 111.635 ;
        RECT 11.415 110.715 12.625 111.465 ;
        RECT 12.800 110.920 18.145 111.465 ;
        RECT 11.415 110.175 11.935 110.715 ;
        RECT 12.105 110.005 12.625 110.545 ;
        RECT 11.415 108.915 12.625 110.005 ;
        RECT 14.390 109.350 14.740 110.600 ;
        RECT 16.220 110.090 16.560 110.920 ;
        RECT 18.375 110.645 18.585 111.465 ;
        RECT 18.755 110.665 19.085 111.295 ;
        RECT 18.755 110.065 19.005 110.665 ;
        RECT 19.255 110.645 19.485 111.465 ;
        RECT 19.695 110.695 21.365 111.465 ;
        RECT 19.175 110.225 19.505 110.475 ;
        RECT 12.800 108.915 18.145 109.350 ;
        RECT 18.375 108.915 18.585 110.055 ;
        RECT 18.755 109.085 19.085 110.065 ;
        RECT 19.255 108.915 19.485 110.055 ;
        RECT 19.695 110.005 20.445 110.525 ;
        RECT 20.615 110.175 21.365 110.695 ;
        RECT 21.535 110.790 21.795 111.295 ;
        RECT 21.975 111.085 22.305 111.465 ;
        RECT 22.485 110.915 22.655 111.295 ;
        RECT 19.695 108.915 21.365 110.005 ;
        RECT 21.535 109.990 21.705 110.790 ;
        RECT 21.990 110.745 22.655 110.915 ;
        RECT 21.990 110.490 22.160 110.745 ;
        RECT 22.915 110.740 23.205 111.465 ;
        RECT 23.375 110.790 23.635 111.295 ;
        RECT 23.815 111.085 24.145 111.465 ;
        RECT 24.325 110.915 24.495 111.295 ;
        RECT 21.875 110.160 22.160 110.490 ;
        RECT 22.395 110.195 22.725 110.565 ;
        RECT 21.990 110.015 22.160 110.160 ;
        RECT 21.535 109.085 21.805 109.990 ;
        RECT 21.990 109.845 22.655 110.015 ;
        RECT 21.975 108.915 22.305 109.675 ;
        RECT 22.485 109.085 22.655 109.845 ;
        RECT 22.915 108.915 23.205 110.080 ;
        RECT 23.375 109.990 23.545 110.790 ;
        RECT 23.830 110.745 24.495 110.915 ;
        RECT 24.755 110.790 25.015 111.295 ;
        RECT 25.195 111.085 25.525 111.465 ;
        RECT 25.705 110.915 25.875 111.295 ;
        RECT 23.830 110.490 24.000 110.745 ;
        RECT 23.715 110.160 24.000 110.490 ;
        RECT 24.235 110.195 24.565 110.565 ;
        RECT 23.830 110.015 24.000 110.160 ;
        RECT 23.375 109.085 23.645 109.990 ;
        RECT 23.830 109.845 24.495 110.015 ;
        RECT 23.815 108.915 24.145 109.675 ;
        RECT 24.325 109.085 24.495 109.845 ;
        RECT 24.755 109.990 24.925 110.790 ;
        RECT 25.210 110.745 25.875 110.915 ;
        RECT 26.225 110.915 26.395 111.295 ;
        RECT 26.575 111.085 26.905 111.465 ;
        RECT 26.225 110.745 26.890 110.915 ;
        RECT 27.085 110.790 27.345 111.295 ;
        RECT 27.825 110.995 27.995 111.465 ;
        RECT 28.165 110.815 28.495 111.295 ;
        RECT 28.665 110.995 28.835 111.465 ;
        RECT 29.005 110.815 29.335 111.295 ;
        RECT 25.210 110.490 25.380 110.745 ;
        RECT 25.095 110.160 25.380 110.490 ;
        RECT 25.615 110.195 25.945 110.565 ;
        RECT 26.155 110.195 26.485 110.565 ;
        RECT 26.720 110.490 26.890 110.745 ;
        RECT 25.210 110.015 25.380 110.160 ;
        RECT 26.720 110.160 27.005 110.490 ;
        RECT 26.720 110.015 26.890 110.160 ;
        RECT 24.755 109.085 25.025 109.990 ;
        RECT 25.210 109.845 25.875 110.015 ;
        RECT 25.195 108.915 25.525 109.675 ;
        RECT 25.705 109.085 25.875 109.845 ;
        RECT 26.225 109.845 26.890 110.015 ;
        RECT 27.175 109.990 27.345 110.790 ;
        RECT 26.225 109.085 26.395 109.845 ;
        RECT 26.575 108.915 26.905 109.675 ;
        RECT 27.075 109.085 27.345 109.990 ;
        RECT 27.570 110.645 29.335 110.815 ;
        RECT 29.505 110.655 29.675 111.465 ;
        RECT 29.875 111.085 30.945 111.255 ;
        RECT 29.875 110.730 30.195 111.085 ;
        RECT 27.570 110.095 27.980 110.645 ;
        RECT 29.870 110.475 30.195 110.730 ;
        RECT 28.165 110.265 30.195 110.475 ;
        RECT 29.850 110.255 30.195 110.265 ;
        RECT 30.365 110.515 30.605 110.915 ;
        RECT 30.775 110.855 30.945 111.085 ;
        RECT 31.115 111.025 31.305 111.465 ;
        RECT 31.475 111.015 32.425 111.295 ;
        RECT 32.645 111.105 32.995 111.275 ;
        RECT 30.775 110.685 31.305 110.855 ;
        RECT 27.570 109.925 29.295 110.095 ;
        RECT 27.825 108.915 27.995 109.755 ;
        RECT 28.205 109.085 28.455 109.925 ;
        RECT 28.665 108.915 28.835 109.755 ;
        RECT 29.005 109.085 29.295 109.925 ;
        RECT 29.505 108.915 29.675 109.975 ;
        RECT 29.850 109.635 30.020 110.255 ;
        RECT 30.365 110.145 30.905 110.515 ;
        RECT 31.085 110.405 31.305 110.685 ;
        RECT 31.475 110.235 31.645 111.015 ;
        RECT 31.240 110.065 31.645 110.235 ;
        RECT 31.815 110.225 32.165 110.845 ;
        RECT 31.240 109.975 31.410 110.065 ;
        RECT 32.335 110.055 32.545 110.845 ;
        RECT 30.190 109.805 31.410 109.975 ;
        RECT 31.870 109.895 32.545 110.055 ;
        RECT 29.850 109.465 30.650 109.635 ;
        RECT 29.970 108.915 30.300 109.295 ;
        RECT 30.480 109.175 30.650 109.465 ;
        RECT 31.240 109.425 31.410 109.805 ;
        RECT 31.580 109.885 32.545 109.895 ;
        RECT 32.735 110.715 32.995 111.105 ;
        RECT 33.205 111.005 33.535 111.465 ;
        RECT 34.410 111.075 35.265 111.245 ;
        RECT 35.470 111.075 35.965 111.245 ;
        RECT 36.135 111.105 36.465 111.465 ;
        RECT 32.735 110.025 32.905 110.715 ;
        RECT 33.075 110.365 33.245 110.545 ;
        RECT 33.415 110.535 34.205 110.785 ;
        RECT 34.410 110.365 34.580 111.075 ;
        RECT 34.750 110.565 35.105 110.785 ;
        RECT 33.075 110.195 34.765 110.365 ;
        RECT 31.580 109.595 32.040 109.885 ;
        RECT 32.735 109.855 34.235 110.025 ;
        RECT 32.735 109.715 32.905 109.855 ;
        RECT 32.345 109.545 32.905 109.715 ;
        RECT 30.820 108.915 31.070 109.375 ;
        RECT 31.240 109.085 32.110 109.425 ;
        RECT 32.345 109.085 32.515 109.545 ;
        RECT 33.350 109.515 34.425 109.685 ;
        RECT 32.685 108.915 33.055 109.375 ;
        RECT 33.350 109.175 33.520 109.515 ;
        RECT 33.690 108.915 34.020 109.345 ;
        RECT 34.255 109.175 34.425 109.515 ;
        RECT 34.595 109.415 34.765 110.195 ;
        RECT 34.935 109.975 35.105 110.565 ;
        RECT 35.275 110.165 35.625 110.785 ;
        RECT 34.935 109.585 35.400 109.975 ;
        RECT 35.795 109.715 35.965 111.075 ;
        RECT 36.135 109.885 36.595 110.935 ;
        RECT 35.570 109.545 35.965 109.715 ;
        RECT 35.570 109.415 35.740 109.545 ;
        RECT 34.595 109.085 35.275 109.415 ;
        RECT 35.490 109.085 35.740 109.415 ;
        RECT 35.910 108.915 36.160 109.375 ;
        RECT 36.330 109.100 36.655 109.885 ;
        RECT 36.825 109.085 36.995 111.205 ;
        RECT 37.165 111.085 37.495 111.465 ;
        RECT 37.665 110.915 37.920 111.205 ;
        RECT 38.405 110.995 38.575 111.465 ;
        RECT 37.170 110.745 37.920 110.915 ;
        RECT 38.745 110.815 39.075 111.295 ;
        RECT 39.245 110.995 39.415 111.465 ;
        RECT 39.585 110.815 39.915 111.295 ;
        RECT 37.170 109.755 37.400 110.745 ;
        RECT 38.150 110.645 39.915 110.815 ;
        RECT 40.085 110.655 40.255 111.465 ;
        RECT 40.455 111.085 41.525 111.255 ;
        RECT 40.455 110.730 40.775 111.085 ;
        RECT 37.570 109.925 37.920 110.575 ;
        RECT 38.150 110.095 38.560 110.645 ;
        RECT 40.450 110.475 40.775 110.730 ;
        RECT 38.745 110.265 40.775 110.475 ;
        RECT 40.430 110.255 40.775 110.265 ;
        RECT 40.945 110.515 41.185 110.915 ;
        RECT 41.355 110.855 41.525 111.085 ;
        RECT 41.695 111.025 41.885 111.465 ;
        RECT 42.055 111.015 43.005 111.295 ;
        RECT 43.225 111.105 43.575 111.275 ;
        RECT 41.355 110.685 41.885 110.855 ;
        RECT 38.150 109.925 39.875 110.095 ;
        RECT 37.170 109.585 37.920 109.755 ;
        RECT 37.165 108.915 37.495 109.415 ;
        RECT 37.665 109.085 37.920 109.585 ;
        RECT 38.405 108.915 38.575 109.755 ;
        RECT 38.785 109.085 39.035 109.925 ;
        RECT 39.245 108.915 39.415 109.755 ;
        RECT 39.585 109.085 39.875 109.925 ;
        RECT 40.085 108.915 40.255 109.975 ;
        RECT 40.430 109.635 40.600 110.255 ;
        RECT 40.945 110.145 41.485 110.515 ;
        RECT 41.665 110.405 41.885 110.685 ;
        RECT 42.055 110.235 42.225 111.015 ;
        RECT 41.820 110.065 42.225 110.235 ;
        RECT 42.395 110.225 42.745 110.845 ;
        RECT 41.820 109.975 41.990 110.065 ;
        RECT 42.915 110.055 43.125 110.845 ;
        RECT 40.770 109.805 41.990 109.975 ;
        RECT 42.450 109.895 43.125 110.055 ;
        RECT 40.430 109.465 41.230 109.635 ;
        RECT 40.550 108.915 40.880 109.295 ;
        RECT 41.060 109.175 41.230 109.465 ;
        RECT 41.820 109.425 41.990 109.805 ;
        RECT 42.160 109.885 43.125 109.895 ;
        RECT 43.315 110.715 43.575 111.105 ;
        RECT 43.785 111.005 44.115 111.465 ;
        RECT 44.990 111.075 45.845 111.245 ;
        RECT 46.050 111.075 46.545 111.245 ;
        RECT 46.715 111.105 47.045 111.465 ;
        RECT 43.315 110.025 43.485 110.715 ;
        RECT 43.655 110.365 43.825 110.545 ;
        RECT 43.995 110.535 44.785 110.785 ;
        RECT 44.990 110.365 45.160 111.075 ;
        RECT 45.330 110.565 45.685 110.785 ;
        RECT 43.655 110.195 45.345 110.365 ;
        RECT 42.160 109.595 42.620 109.885 ;
        RECT 43.315 109.855 44.815 110.025 ;
        RECT 43.315 109.715 43.485 109.855 ;
        RECT 42.925 109.545 43.485 109.715 ;
        RECT 41.400 108.915 41.650 109.375 ;
        RECT 41.820 109.085 42.690 109.425 ;
        RECT 42.925 109.085 43.095 109.545 ;
        RECT 43.930 109.515 45.005 109.685 ;
        RECT 43.265 108.915 43.635 109.375 ;
        RECT 43.930 109.175 44.100 109.515 ;
        RECT 44.270 108.915 44.600 109.345 ;
        RECT 44.835 109.175 45.005 109.515 ;
        RECT 45.175 109.415 45.345 110.195 ;
        RECT 45.515 109.975 45.685 110.565 ;
        RECT 45.855 110.165 46.205 110.785 ;
        RECT 45.515 109.585 45.980 109.975 ;
        RECT 46.375 109.715 46.545 111.075 ;
        RECT 46.715 109.885 47.175 110.935 ;
        RECT 46.150 109.545 46.545 109.715 ;
        RECT 46.150 109.415 46.320 109.545 ;
        RECT 45.175 109.085 45.855 109.415 ;
        RECT 46.070 109.085 46.320 109.415 ;
        RECT 46.490 108.915 46.740 109.375 ;
        RECT 46.910 109.100 47.235 109.885 ;
        RECT 47.405 109.085 47.575 111.205 ;
        RECT 47.745 111.085 48.075 111.465 ;
        RECT 48.245 110.915 48.500 111.205 ;
        RECT 47.750 110.745 48.500 110.915 ;
        RECT 47.750 109.755 47.980 110.745 ;
        RECT 48.675 110.740 48.965 111.465 ;
        RECT 49.225 110.915 49.395 111.295 ;
        RECT 49.575 111.085 49.905 111.465 ;
        RECT 49.225 110.745 49.890 110.915 ;
        RECT 50.085 110.790 50.345 111.295 ;
        RECT 51.745 110.995 51.915 111.465 ;
        RECT 52.085 110.815 52.415 111.295 ;
        RECT 52.585 110.995 52.755 111.465 ;
        RECT 52.925 110.815 53.255 111.295 ;
        RECT 48.150 109.925 48.500 110.575 ;
        RECT 49.155 110.195 49.485 110.565 ;
        RECT 49.720 110.490 49.890 110.745 ;
        RECT 49.720 110.160 50.005 110.490 ;
        RECT 47.750 109.585 48.500 109.755 ;
        RECT 47.745 108.915 48.075 109.415 ;
        RECT 48.245 109.085 48.500 109.585 ;
        RECT 48.675 108.915 48.965 110.080 ;
        RECT 49.720 110.015 49.890 110.160 ;
        RECT 49.225 109.845 49.890 110.015 ;
        RECT 50.175 109.990 50.345 110.790 ;
        RECT 49.225 109.085 49.395 109.845 ;
        RECT 49.575 108.915 49.905 109.675 ;
        RECT 50.075 109.085 50.345 109.990 ;
        RECT 51.490 110.645 53.255 110.815 ;
        RECT 53.425 110.655 53.595 111.465 ;
        RECT 53.795 111.085 54.865 111.255 ;
        RECT 53.795 110.730 54.115 111.085 ;
        RECT 51.490 110.095 51.900 110.645 ;
        RECT 53.790 110.475 54.115 110.730 ;
        RECT 52.085 110.265 54.115 110.475 ;
        RECT 53.770 110.255 54.115 110.265 ;
        RECT 54.285 110.515 54.525 110.915 ;
        RECT 54.695 110.855 54.865 111.085 ;
        RECT 55.035 111.025 55.225 111.465 ;
        RECT 55.395 111.015 56.345 111.295 ;
        RECT 56.565 111.105 56.915 111.275 ;
        RECT 54.695 110.685 55.225 110.855 ;
        RECT 51.490 109.925 53.215 110.095 ;
        RECT 51.745 108.915 51.915 109.755 ;
        RECT 52.125 109.085 52.375 109.925 ;
        RECT 52.585 108.915 52.755 109.755 ;
        RECT 52.925 109.085 53.215 109.925 ;
        RECT 53.425 108.915 53.595 109.975 ;
        RECT 53.770 109.635 53.940 110.255 ;
        RECT 54.285 110.145 54.825 110.515 ;
        RECT 55.005 110.405 55.225 110.685 ;
        RECT 55.395 110.235 55.565 111.015 ;
        RECT 55.160 110.065 55.565 110.235 ;
        RECT 55.735 110.225 56.085 110.845 ;
        RECT 55.160 109.975 55.330 110.065 ;
        RECT 56.255 110.055 56.465 110.845 ;
        RECT 54.110 109.805 55.330 109.975 ;
        RECT 55.790 109.895 56.465 110.055 ;
        RECT 53.770 109.465 54.570 109.635 ;
        RECT 53.890 108.915 54.220 109.295 ;
        RECT 54.400 109.175 54.570 109.465 ;
        RECT 55.160 109.425 55.330 109.805 ;
        RECT 55.500 109.885 56.465 109.895 ;
        RECT 56.655 110.715 56.915 111.105 ;
        RECT 57.125 111.005 57.455 111.465 ;
        RECT 58.330 111.075 59.185 111.245 ;
        RECT 59.390 111.075 59.885 111.245 ;
        RECT 60.055 111.105 60.385 111.465 ;
        RECT 56.655 110.025 56.825 110.715 ;
        RECT 56.995 110.365 57.165 110.545 ;
        RECT 57.335 110.535 58.125 110.785 ;
        RECT 58.330 110.365 58.500 111.075 ;
        RECT 58.670 110.565 59.025 110.785 ;
        RECT 56.995 110.195 58.685 110.365 ;
        RECT 55.500 109.595 55.960 109.885 ;
        RECT 56.655 109.855 58.155 110.025 ;
        RECT 56.655 109.715 56.825 109.855 ;
        RECT 56.265 109.545 56.825 109.715 ;
        RECT 54.740 108.915 54.990 109.375 ;
        RECT 55.160 109.085 56.030 109.425 ;
        RECT 56.265 109.085 56.435 109.545 ;
        RECT 57.270 109.515 58.345 109.685 ;
        RECT 56.605 108.915 56.975 109.375 ;
        RECT 57.270 109.175 57.440 109.515 ;
        RECT 57.610 108.915 57.940 109.345 ;
        RECT 58.175 109.175 58.345 109.515 ;
        RECT 58.515 109.415 58.685 110.195 ;
        RECT 58.855 109.975 59.025 110.565 ;
        RECT 59.195 110.165 59.545 110.785 ;
        RECT 58.855 109.585 59.320 109.975 ;
        RECT 59.715 109.715 59.885 111.075 ;
        RECT 60.055 109.885 60.515 110.935 ;
        RECT 59.490 109.545 59.885 109.715 ;
        RECT 59.490 109.415 59.660 109.545 ;
        RECT 58.515 109.085 59.195 109.415 ;
        RECT 59.410 109.085 59.660 109.415 ;
        RECT 59.830 108.915 60.080 109.375 ;
        RECT 60.250 109.100 60.575 109.885 ;
        RECT 60.745 109.085 60.915 111.205 ;
        RECT 61.085 111.085 61.415 111.465 ;
        RECT 61.585 110.915 61.840 111.205 ;
        RECT 63.245 110.995 63.415 111.465 ;
        RECT 61.090 110.745 61.840 110.915 ;
        RECT 63.585 110.815 63.915 111.295 ;
        RECT 64.085 110.995 64.255 111.465 ;
        RECT 64.425 110.815 64.755 111.295 ;
        RECT 61.090 109.755 61.320 110.745 ;
        RECT 62.990 110.645 64.755 110.815 ;
        RECT 64.925 110.655 65.095 111.465 ;
        RECT 65.295 111.085 66.365 111.255 ;
        RECT 65.295 110.730 65.615 111.085 ;
        RECT 61.490 109.925 61.840 110.575 ;
        RECT 62.990 110.095 63.400 110.645 ;
        RECT 65.290 110.475 65.615 110.730 ;
        RECT 63.585 110.265 65.615 110.475 ;
        RECT 65.270 110.255 65.615 110.265 ;
        RECT 65.785 110.515 66.025 110.915 ;
        RECT 66.195 110.855 66.365 111.085 ;
        RECT 66.535 111.025 66.725 111.465 ;
        RECT 66.895 111.015 67.845 111.295 ;
        RECT 68.065 111.105 68.415 111.275 ;
        RECT 66.195 110.685 66.725 110.855 ;
        RECT 62.990 109.925 64.715 110.095 ;
        RECT 61.090 109.585 61.840 109.755 ;
        RECT 61.085 108.915 61.415 109.415 ;
        RECT 61.585 109.085 61.840 109.585 ;
        RECT 63.245 108.915 63.415 109.755 ;
        RECT 63.625 109.085 63.875 109.925 ;
        RECT 64.085 108.915 64.255 109.755 ;
        RECT 64.425 109.085 64.715 109.925 ;
        RECT 64.925 108.915 65.095 109.975 ;
        RECT 65.270 109.635 65.440 110.255 ;
        RECT 65.785 110.145 66.325 110.515 ;
        RECT 66.505 110.405 66.725 110.685 ;
        RECT 66.895 110.235 67.065 111.015 ;
        RECT 66.660 110.065 67.065 110.235 ;
        RECT 67.235 110.225 67.585 110.845 ;
        RECT 66.660 109.975 66.830 110.065 ;
        RECT 67.755 110.055 67.965 110.845 ;
        RECT 65.610 109.805 66.830 109.975 ;
        RECT 67.290 109.895 67.965 110.055 ;
        RECT 65.270 109.465 66.070 109.635 ;
        RECT 65.390 108.915 65.720 109.295 ;
        RECT 65.900 109.175 66.070 109.465 ;
        RECT 66.660 109.425 66.830 109.805 ;
        RECT 67.000 109.885 67.965 109.895 ;
        RECT 68.155 110.715 68.415 111.105 ;
        RECT 68.625 111.005 68.955 111.465 ;
        RECT 69.830 111.075 70.685 111.245 ;
        RECT 70.890 111.075 71.385 111.245 ;
        RECT 71.555 111.105 71.885 111.465 ;
        RECT 68.155 110.025 68.325 110.715 ;
        RECT 68.495 110.365 68.665 110.545 ;
        RECT 68.835 110.535 69.625 110.785 ;
        RECT 69.830 110.365 70.000 111.075 ;
        RECT 70.170 110.565 70.525 110.785 ;
        RECT 68.495 110.195 70.185 110.365 ;
        RECT 67.000 109.595 67.460 109.885 ;
        RECT 68.155 109.855 69.655 110.025 ;
        RECT 68.155 109.715 68.325 109.855 ;
        RECT 67.765 109.545 68.325 109.715 ;
        RECT 66.240 108.915 66.490 109.375 ;
        RECT 66.660 109.085 67.530 109.425 ;
        RECT 67.765 109.085 67.935 109.545 ;
        RECT 68.770 109.515 69.845 109.685 ;
        RECT 68.105 108.915 68.475 109.375 ;
        RECT 68.770 109.175 68.940 109.515 ;
        RECT 69.110 108.915 69.440 109.345 ;
        RECT 69.675 109.175 69.845 109.515 ;
        RECT 70.015 109.415 70.185 110.195 ;
        RECT 70.355 109.975 70.525 110.565 ;
        RECT 70.695 110.165 71.045 110.785 ;
        RECT 70.355 109.585 70.820 109.975 ;
        RECT 71.215 109.715 71.385 111.075 ;
        RECT 71.555 109.885 72.015 110.935 ;
        RECT 70.990 109.545 71.385 109.715 ;
        RECT 70.990 109.415 71.160 109.545 ;
        RECT 70.015 109.085 70.695 109.415 ;
        RECT 70.910 109.085 71.160 109.415 ;
        RECT 71.330 108.915 71.580 109.375 ;
        RECT 71.750 109.100 72.075 109.885 ;
        RECT 72.245 109.085 72.415 111.205 ;
        RECT 72.585 111.085 72.915 111.465 ;
        RECT 73.085 110.915 73.340 111.205 ;
        RECT 72.590 110.745 73.340 110.915 ;
        RECT 72.590 109.755 72.820 110.745 ;
        RECT 74.435 110.740 74.725 111.465 ;
        RECT 74.895 110.790 75.155 111.295 ;
        RECT 75.335 111.085 75.665 111.465 ;
        RECT 75.845 110.915 76.015 111.295 ;
        RECT 72.990 109.925 73.340 110.575 ;
        RECT 72.590 109.585 73.340 109.755 ;
        RECT 72.585 108.915 72.915 109.415 ;
        RECT 73.085 109.085 73.340 109.585 ;
        RECT 74.435 108.915 74.725 110.080 ;
        RECT 74.895 109.990 75.065 110.790 ;
        RECT 75.350 110.745 76.015 110.915 ;
        RECT 76.825 110.915 76.995 111.295 ;
        RECT 77.175 111.085 77.505 111.465 ;
        RECT 76.825 110.745 77.490 110.915 ;
        RECT 77.685 110.790 77.945 111.295 ;
        RECT 78.425 110.995 78.595 111.465 ;
        RECT 78.765 110.815 79.095 111.295 ;
        RECT 79.265 110.995 79.435 111.465 ;
        RECT 79.605 110.815 79.935 111.295 ;
        RECT 75.350 110.490 75.520 110.745 ;
        RECT 75.235 110.160 75.520 110.490 ;
        RECT 75.755 110.195 76.085 110.565 ;
        RECT 76.755 110.195 77.085 110.565 ;
        RECT 77.320 110.490 77.490 110.745 ;
        RECT 75.350 110.015 75.520 110.160 ;
        RECT 77.320 110.160 77.605 110.490 ;
        RECT 77.320 110.015 77.490 110.160 ;
        RECT 74.895 109.085 75.165 109.990 ;
        RECT 75.350 109.845 76.015 110.015 ;
        RECT 75.335 108.915 75.665 109.675 ;
        RECT 75.845 109.085 76.015 109.845 ;
        RECT 76.825 109.845 77.490 110.015 ;
        RECT 77.775 109.990 77.945 110.790 ;
        RECT 76.825 109.085 76.995 109.845 ;
        RECT 77.175 108.915 77.505 109.675 ;
        RECT 77.675 109.085 77.945 109.990 ;
        RECT 78.170 110.645 79.935 110.815 ;
        RECT 80.105 110.655 80.275 111.465 ;
        RECT 80.475 111.085 81.545 111.255 ;
        RECT 80.475 110.730 80.795 111.085 ;
        RECT 78.170 110.095 78.580 110.645 ;
        RECT 80.470 110.475 80.795 110.730 ;
        RECT 78.765 110.265 80.795 110.475 ;
        RECT 80.450 110.255 80.795 110.265 ;
        RECT 80.965 110.515 81.205 110.915 ;
        RECT 81.375 110.855 81.545 111.085 ;
        RECT 81.715 111.025 81.905 111.465 ;
        RECT 82.075 111.015 83.025 111.295 ;
        RECT 83.245 111.105 83.595 111.275 ;
        RECT 81.375 110.685 81.905 110.855 ;
        RECT 78.170 109.925 79.895 110.095 ;
        RECT 78.425 108.915 78.595 109.755 ;
        RECT 78.805 109.085 79.055 109.925 ;
        RECT 79.265 108.915 79.435 109.755 ;
        RECT 79.605 109.085 79.895 109.925 ;
        RECT 80.105 108.915 80.275 109.975 ;
        RECT 80.450 109.635 80.620 110.255 ;
        RECT 80.965 110.145 81.505 110.515 ;
        RECT 81.685 110.405 81.905 110.685 ;
        RECT 82.075 110.235 82.245 111.015 ;
        RECT 81.840 110.065 82.245 110.235 ;
        RECT 82.415 110.225 82.765 110.845 ;
        RECT 81.840 109.975 82.010 110.065 ;
        RECT 82.935 110.055 83.145 110.845 ;
        RECT 80.790 109.805 82.010 109.975 ;
        RECT 82.470 109.895 83.145 110.055 ;
        RECT 80.450 109.465 81.250 109.635 ;
        RECT 80.570 108.915 80.900 109.295 ;
        RECT 81.080 109.175 81.250 109.465 ;
        RECT 81.840 109.425 82.010 109.805 ;
        RECT 82.180 109.885 83.145 109.895 ;
        RECT 83.335 110.715 83.595 111.105 ;
        RECT 83.805 111.005 84.135 111.465 ;
        RECT 85.010 111.075 85.865 111.245 ;
        RECT 86.070 111.075 86.565 111.245 ;
        RECT 86.735 111.105 87.065 111.465 ;
        RECT 83.335 110.025 83.505 110.715 ;
        RECT 83.675 110.365 83.845 110.545 ;
        RECT 84.015 110.535 84.805 110.785 ;
        RECT 85.010 110.365 85.180 111.075 ;
        RECT 85.350 110.565 85.705 110.785 ;
        RECT 83.675 110.195 85.365 110.365 ;
        RECT 82.180 109.595 82.640 109.885 ;
        RECT 83.335 109.855 84.835 110.025 ;
        RECT 83.335 109.715 83.505 109.855 ;
        RECT 82.945 109.545 83.505 109.715 ;
        RECT 81.420 108.915 81.670 109.375 ;
        RECT 81.840 109.085 82.710 109.425 ;
        RECT 82.945 109.085 83.115 109.545 ;
        RECT 83.950 109.515 85.025 109.685 ;
        RECT 83.285 108.915 83.655 109.375 ;
        RECT 83.950 109.175 84.120 109.515 ;
        RECT 84.290 108.915 84.620 109.345 ;
        RECT 84.855 109.175 85.025 109.515 ;
        RECT 85.195 109.415 85.365 110.195 ;
        RECT 85.535 109.975 85.705 110.565 ;
        RECT 85.875 110.165 86.225 110.785 ;
        RECT 85.535 109.585 86.000 109.975 ;
        RECT 86.395 109.715 86.565 111.075 ;
        RECT 86.735 109.885 87.195 110.935 ;
        RECT 86.170 109.545 86.565 109.715 ;
        RECT 86.170 109.415 86.340 109.545 ;
        RECT 85.195 109.085 85.875 109.415 ;
        RECT 86.090 109.085 86.340 109.415 ;
        RECT 86.510 108.915 86.760 109.375 ;
        RECT 86.930 109.100 87.255 109.885 ;
        RECT 87.425 109.085 87.595 111.205 ;
        RECT 87.765 111.085 88.095 111.465 ;
        RECT 88.265 110.915 88.520 111.205 ;
        RECT 89.005 110.995 89.175 111.465 ;
        RECT 87.770 110.745 88.520 110.915 ;
        RECT 89.345 110.815 89.675 111.295 ;
        RECT 89.845 110.995 90.015 111.465 ;
        RECT 90.185 110.815 90.515 111.295 ;
        RECT 87.770 109.755 88.000 110.745 ;
        RECT 88.750 110.645 90.515 110.815 ;
        RECT 90.685 110.655 90.855 111.465 ;
        RECT 91.055 111.085 92.125 111.255 ;
        RECT 91.055 110.730 91.375 111.085 ;
        RECT 88.170 109.925 88.520 110.575 ;
        RECT 88.750 110.095 89.160 110.645 ;
        RECT 91.050 110.475 91.375 110.730 ;
        RECT 89.345 110.265 91.375 110.475 ;
        RECT 91.030 110.255 91.375 110.265 ;
        RECT 91.545 110.515 91.785 110.915 ;
        RECT 91.955 110.855 92.125 111.085 ;
        RECT 92.295 111.025 92.485 111.465 ;
        RECT 92.655 111.015 93.605 111.295 ;
        RECT 93.825 111.105 94.175 111.275 ;
        RECT 91.955 110.685 92.485 110.855 ;
        RECT 88.750 109.925 90.475 110.095 ;
        RECT 87.770 109.585 88.520 109.755 ;
        RECT 87.765 108.915 88.095 109.415 ;
        RECT 88.265 109.085 88.520 109.585 ;
        RECT 89.005 108.915 89.175 109.755 ;
        RECT 89.385 109.085 89.635 109.925 ;
        RECT 89.845 108.915 90.015 109.755 ;
        RECT 90.185 109.085 90.475 109.925 ;
        RECT 90.685 108.915 90.855 109.975 ;
        RECT 91.030 109.635 91.200 110.255 ;
        RECT 91.545 110.145 92.085 110.515 ;
        RECT 92.265 110.405 92.485 110.685 ;
        RECT 92.655 110.235 92.825 111.015 ;
        RECT 92.420 110.065 92.825 110.235 ;
        RECT 92.995 110.225 93.345 110.845 ;
        RECT 92.420 109.975 92.590 110.065 ;
        RECT 93.515 110.055 93.725 110.845 ;
        RECT 91.370 109.805 92.590 109.975 ;
        RECT 93.050 109.895 93.725 110.055 ;
        RECT 91.030 109.465 91.830 109.635 ;
        RECT 91.150 108.915 91.480 109.295 ;
        RECT 91.660 109.175 91.830 109.465 ;
        RECT 92.420 109.425 92.590 109.805 ;
        RECT 92.760 109.885 93.725 109.895 ;
        RECT 93.915 110.715 94.175 111.105 ;
        RECT 94.385 111.005 94.715 111.465 ;
        RECT 95.590 111.075 96.445 111.245 ;
        RECT 96.650 111.075 97.145 111.245 ;
        RECT 97.315 111.105 97.645 111.465 ;
        RECT 93.915 110.025 94.085 110.715 ;
        RECT 94.255 110.365 94.425 110.545 ;
        RECT 94.595 110.535 95.385 110.785 ;
        RECT 95.590 110.365 95.760 111.075 ;
        RECT 95.930 110.565 96.285 110.785 ;
        RECT 94.255 110.195 95.945 110.365 ;
        RECT 92.760 109.595 93.220 109.885 ;
        RECT 93.915 109.855 95.415 110.025 ;
        RECT 93.915 109.715 94.085 109.855 ;
        RECT 93.525 109.545 94.085 109.715 ;
        RECT 92.000 108.915 92.250 109.375 ;
        RECT 92.420 109.085 93.290 109.425 ;
        RECT 93.525 109.085 93.695 109.545 ;
        RECT 94.530 109.515 95.605 109.685 ;
        RECT 93.865 108.915 94.235 109.375 ;
        RECT 94.530 109.175 94.700 109.515 ;
        RECT 94.870 108.915 95.200 109.345 ;
        RECT 95.435 109.175 95.605 109.515 ;
        RECT 95.775 109.415 95.945 110.195 ;
        RECT 96.115 109.975 96.285 110.565 ;
        RECT 96.455 110.165 96.805 110.785 ;
        RECT 96.115 109.585 96.580 109.975 ;
        RECT 96.975 109.715 97.145 111.075 ;
        RECT 97.315 109.885 97.775 110.935 ;
        RECT 96.750 109.545 97.145 109.715 ;
        RECT 96.750 109.415 96.920 109.545 ;
        RECT 95.775 109.085 96.455 109.415 ;
        RECT 96.670 109.085 96.920 109.415 ;
        RECT 97.090 108.915 97.340 109.375 ;
        RECT 97.510 109.100 97.835 109.885 ;
        RECT 98.005 109.085 98.175 111.205 ;
        RECT 98.345 111.085 98.675 111.465 ;
        RECT 98.845 110.915 99.100 111.205 ;
        RECT 98.350 110.745 99.100 110.915 ;
        RECT 98.350 109.755 98.580 110.745 ;
        RECT 100.195 110.740 100.485 111.465 ;
        RECT 101.580 110.915 101.835 111.205 ;
        RECT 102.005 111.085 102.335 111.465 ;
        RECT 101.580 110.745 102.330 110.915 ;
        RECT 98.750 109.925 99.100 110.575 ;
        RECT 98.350 109.585 99.100 109.755 ;
        RECT 98.345 108.915 98.675 109.415 ;
        RECT 98.845 109.085 99.100 109.585 ;
        RECT 100.195 108.915 100.485 110.080 ;
        RECT 101.580 109.925 101.930 110.575 ;
        RECT 102.100 109.755 102.330 110.745 ;
        RECT 101.580 109.585 102.330 109.755 ;
        RECT 101.580 109.085 101.835 109.585 ;
        RECT 102.005 108.915 102.335 109.415 ;
        RECT 102.505 109.085 102.675 111.205 ;
        RECT 103.035 111.105 103.365 111.465 ;
        RECT 103.535 111.075 104.030 111.245 ;
        RECT 104.235 111.075 105.090 111.245 ;
        RECT 102.905 109.885 103.365 110.935 ;
        RECT 102.845 109.100 103.170 109.885 ;
        RECT 103.535 109.715 103.705 111.075 ;
        RECT 103.875 110.165 104.225 110.785 ;
        RECT 104.395 110.565 104.750 110.785 ;
        RECT 104.395 109.975 104.565 110.565 ;
        RECT 104.920 110.365 105.090 111.075 ;
        RECT 105.965 111.005 106.295 111.465 ;
        RECT 106.505 111.105 106.855 111.275 ;
        RECT 105.295 110.535 106.085 110.785 ;
        RECT 106.505 110.715 106.765 111.105 ;
        RECT 107.075 111.015 108.025 111.295 ;
        RECT 108.195 111.025 108.385 111.465 ;
        RECT 108.555 111.085 109.625 111.255 ;
        RECT 106.255 110.365 106.425 110.545 ;
        RECT 103.535 109.545 103.930 109.715 ;
        RECT 104.100 109.585 104.565 109.975 ;
        RECT 104.735 110.195 106.425 110.365 ;
        RECT 103.760 109.415 103.930 109.545 ;
        RECT 104.735 109.415 104.905 110.195 ;
        RECT 106.595 110.025 106.765 110.715 ;
        RECT 105.265 109.855 106.765 110.025 ;
        RECT 106.955 110.055 107.165 110.845 ;
        RECT 107.335 110.225 107.685 110.845 ;
        RECT 107.855 110.235 108.025 111.015 ;
        RECT 108.555 110.855 108.725 111.085 ;
        RECT 108.195 110.685 108.725 110.855 ;
        RECT 108.195 110.405 108.415 110.685 ;
        RECT 108.895 110.515 109.135 110.915 ;
        RECT 107.855 110.065 108.260 110.235 ;
        RECT 108.595 110.145 109.135 110.515 ;
        RECT 109.305 110.730 109.625 111.085 ;
        RECT 109.305 110.475 109.630 110.730 ;
        RECT 109.825 110.655 109.995 111.465 ;
        RECT 110.165 110.815 110.495 111.295 ;
        RECT 110.665 110.995 110.835 111.465 ;
        RECT 111.005 110.815 111.335 111.295 ;
        RECT 111.505 110.995 111.675 111.465 ;
        RECT 110.165 110.645 111.930 110.815 ;
        RECT 112.155 110.715 113.365 111.465 ;
        RECT 109.305 110.265 111.335 110.475 ;
        RECT 109.305 110.255 109.650 110.265 ;
        RECT 106.955 109.895 107.630 110.055 ;
        RECT 108.090 109.975 108.260 110.065 ;
        RECT 106.955 109.885 107.920 109.895 ;
        RECT 106.595 109.715 106.765 109.855 ;
        RECT 103.340 108.915 103.590 109.375 ;
        RECT 103.760 109.085 104.010 109.415 ;
        RECT 104.225 109.085 104.905 109.415 ;
        RECT 105.075 109.515 106.150 109.685 ;
        RECT 106.595 109.545 107.155 109.715 ;
        RECT 107.460 109.595 107.920 109.885 ;
        RECT 108.090 109.805 109.310 109.975 ;
        RECT 105.075 109.175 105.245 109.515 ;
        RECT 105.480 108.915 105.810 109.345 ;
        RECT 105.980 109.175 106.150 109.515 ;
        RECT 106.445 108.915 106.815 109.375 ;
        RECT 106.985 109.085 107.155 109.545 ;
        RECT 108.090 109.425 108.260 109.805 ;
        RECT 109.480 109.635 109.650 110.255 ;
        RECT 111.520 110.095 111.930 110.645 ;
        RECT 107.390 109.085 108.260 109.425 ;
        RECT 108.850 109.465 109.650 109.635 ;
        RECT 108.430 108.915 108.680 109.375 ;
        RECT 108.850 109.175 109.020 109.465 ;
        RECT 109.200 108.915 109.530 109.295 ;
        RECT 109.825 108.915 109.995 109.975 ;
        RECT 110.205 109.925 111.930 110.095 ;
        RECT 112.155 110.005 112.675 110.545 ;
        RECT 112.845 110.175 113.365 110.715 ;
        RECT 110.205 109.085 110.495 109.925 ;
        RECT 110.665 108.915 110.835 109.755 ;
        RECT 111.045 109.085 111.295 109.925 ;
        RECT 111.505 108.915 111.675 109.755 ;
        RECT 112.155 108.915 113.365 110.005 ;
        RECT 11.330 108.745 113.450 108.915 ;
        RECT 11.415 107.655 12.625 108.745 ;
        RECT 11.415 106.945 11.935 107.485 ;
        RECT 12.105 107.115 12.625 107.655 ;
        RECT 13.315 107.605 13.525 108.745 ;
        RECT 13.695 107.595 14.025 108.575 ;
        RECT 14.195 107.605 14.425 108.745 ;
        RECT 14.945 107.905 15.115 108.745 ;
        RECT 15.325 107.735 15.575 108.575 ;
        RECT 15.785 107.905 15.955 108.745 ;
        RECT 16.125 107.735 16.415 108.575 ;
        RECT 11.415 106.195 12.625 106.945 ;
        RECT 13.315 106.195 13.525 107.015 ;
        RECT 13.695 106.995 13.945 107.595 ;
        RECT 14.690 107.565 16.415 107.735 ;
        RECT 16.625 107.685 16.795 108.745 ;
        RECT 17.090 108.365 17.420 108.745 ;
        RECT 17.600 108.195 17.770 108.485 ;
        RECT 17.940 108.285 18.190 108.745 ;
        RECT 16.970 108.025 17.770 108.195 ;
        RECT 18.360 108.235 19.230 108.575 ;
        RECT 14.115 107.185 14.445 107.435 ;
        RECT 14.690 107.015 15.100 107.565 ;
        RECT 16.970 107.405 17.140 108.025 ;
        RECT 18.360 107.855 18.530 108.235 ;
        RECT 19.465 108.115 19.635 108.575 ;
        RECT 19.805 108.285 20.175 108.745 ;
        RECT 20.470 108.145 20.640 108.485 ;
        RECT 20.810 108.315 21.140 108.745 ;
        RECT 21.375 108.145 21.545 108.485 ;
        RECT 17.310 107.685 18.530 107.855 ;
        RECT 18.700 107.775 19.160 108.065 ;
        RECT 19.465 107.945 20.025 108.115 ;
        RECT 20.470 107.975 21.545 108.145 ;
        RECT 21.715 108.245 22.395 108.575 ;
        RECT 22.610 108.245 22.860 108.575 ;
        RECT 23.030 108.285 23.280 108.745 ;
        RECT 19.855 107.805 20.025 107.945 ;
        RECT 18.700 107.765 19.665 107.775 ;
        RECT 18.360 107.595 18.530 107.685 ;
        RECT 18.990 107.605 19.665 107.765 ;
        RECT 16.970 107.395 17.315 107.405 ;
        RECT 15.285 107.185 17.315 107.395 ;
        RECT 13.695 106.365 14.025 106.995 ;
        RECT 14.195 106.195 14.425 107.015 ;
        RECT 14.690 106.845 16.455 107.015 ;
        RECT 14.945 106.195 15.115 106.665 ;
        RECT 15.285 106.365 15.615 106.845 ;
        RECT 15.785 106.195 15.955 106.665 ;
        RECT 16.125 106.365 16.455 106.845 ;
        RECT 16.625 106.195 16.795 107.005 ;
        RECT 16.990 106.930 17.315 107.185 ;
        RECT 16.995 106.575 17.315 106.930 ;
        RECT 17.485 107.145 18.025 107.515 ;
        RECT 18.360 107.425 18.765 107.595 ;
        RECT 17.485 106.745 17.725 107.145 ;
        RECT 18.205 106.975 18.425 107.255 ;
        RECT 17.895 106.805 18.425 106.975 ;
        RECT 17.895 106.575 18.065 106.805 ;
        RECT 18.595 106.645 18.765 107.425 ;
        RECT 18.935 106.815 19.285 107.435 ;
        RECT 19.455 106.815 19.665 107.605 ;
        RECT 19.855 107.635 21.355 107.805 ;
        RECT 19.855 106.945 20.025 107.635 ;
        RECT 21.715 107.465 21.885 108.245 ;
        RECT 22.690 108.115 22.860 108.245 ;
        RECT 20.195 107.295 21.885 107.465 ;
        RECT 22.055 107.685 22.520 108.075 ;
        RECT 22.690 107.945 23.085 108.115 ;
        RECT 20.195 107.115 20.365 107.295 ;
        RECT 16.995 106.405 18.065 106.575 ;
        RECT 18.235 106.195 18.425 106.635 ;
        RECT 18.595 106.365 19.545 106.645 ;
        RECT 19.855 106.555 20.115 106.945 ;
        RECT 20.535 106.875 21.325 107.125 ;
        RECT 19.765 106.385 20.115 106.555 ;
        RECT 20.325 106.195 20.655 106.655 ;
        RECT 21.530 106.585 21.700 107.295 ;
        RECT 22.055 107.095 22.225 107.685 ;
        RECT 21.870 106.875 22.225 107.095 ;
        RECT 22.395 106.875 22.745 107.495 ;
        RECT 22.915 106.585 23.085 107.945 ;
        RECT 23.450 107.775 23.775 108.560 ;
        RECT 23.255 106.725 23.715 107.775 ;
        RECT 21.530 106.415 22.385 106.585 ;
        RECT 22.590 106.415 23.085 106.585 ;
        RECT 23.255 106.195 23.585 106.555 ;
        RECT 23.945 106.455 24.115 108.575 ;
        RECT 24.285 108.245 24.615 108.745 ;
        RECT 24.785 108.075 25.040 108.575 ;
        RECT 24.290 107.905 25.040 108.075 ;
        RECT 25.220 108.075 25.475 108.575 ;
        RECT 25.645 108.245 25.975 108.745 ;
        RECT 25.220 107.905 25.970 108.075 ;
        RECT 24.290 106.915 24.520 107.905 ;
        RECT 24.690 107.085 25.040 107.735 ;
        RECT 25.220 107.085 25.570 107.735 ;
        RECT 25.740 106.915 25.970 107.905 ;
        RECT 24.290 106.745 25.040 106.915 ;
        RECT 24.285 106.195 24.615 106.575 ;
        RECT 24.785 106.455 25.040 106.745 ;
        RECT 25.220 106.745 25.970 106.915 ;
        RECT 25.220 106.455 25.475 106.745 ;
        RECT 25.645 106.195 25.975 106.575 ;
        RECT 26.145 106.455 26.315 108.575 ;
        RECT 26.485 107.775 26.810 108.560 ;
        RECT 26.980 108.285 27.230 108.745 ;
        RECT 27.400 108.245 27.650 108.575 ;
        RECT 27.865 108.245 28.545 108.575 ;
        RECT 27.400 108.115 27.570 108.245 ;
        RECT 27.175 107.945 27.570 108.115 ;
        RECT 26.545 106.725 27.005 107.775 ;
        RECT 27.175 106.585 27.345 107.945 ;
        RECT 27.740 107.685 28.205 108.075 ;
        RECT 27.515 106.875 27.865 107.495 ;
        RECT 28.035 107.095 28.205 107.685 ;
        RECT 28.375 107.465 28.545 108.245 ;
        RECT 28.715 108.145 28.885 108.485 ;
        RECT 29.120 108.315 29.450 108.745 ;
        RECT 29.620 108.145 29.790 108.485 ;
        RECT 30.085 108.285 30.455 108.745 ;
        RECT 28.715 107.975 29.790 108.145 ;
        RECT 30.625 108.115 30.795 108.575 ;
        RECT 31.030 108.235 31.900 108.575 ;
        RECT 32.070 108.285 32.320 108.745 ;
        RECT 30.235 107.945 30.795 108.115 ;
        RECT 30.235 107.805 30.405 107.945 ;
        RECT 28.905 107.635 30.405 107.805 ;
        RECT 31.100 107.775 31.560 108.065 ;
        RECT 28.375 107.295 30.065 107.465 ;
        RECT 28.035 106.875 28.390 107.095 ;
        RECT 28.560 106.585 28.730 107.295 ;
        RECT 28.935 106.875 29.725 107.125 ;
        RECT 29.895 107.115 30.065 107.295 ;
        RECT 30.235 106.945 30.405 107.635 ;
        RECT 26.675 106.195 27.005 106.555 ;
        RECT 27.175 106.415 27.670 106.585 ;
        RECT 27.875 106.415 28.730 106.585 ;
        RECT 29.605 106.195 29.935 106.655 ;
        RECT 30.145 106.555 30.405 106.945 ;
        RECT 30.595 107.765 31.560 107.775 ;
        RECT 31.730 107.855 31.900 108.235 ;
        RECT 32.490 108.195 32.660 108.485 ;
        RECT 32.840 108.365 33.170 108.745 ;
        RECT 32.490 108.025 33.290 108.195 ;
        RECT 30.595 107.605 31.270 107.765 ;
        RECT 31.730 107.685 32.950 107.855 ;
        RECT 30.595 106.815 30.805 107.605 ;
        RECT 31.730 107.595 31.900 107.685 ;
        RECT 30.975 106.815 31.325 107.435 ;
        RECT 31.495 107.425 31.900 107.595 ;
        RECT 31.495 106.645 31.665 107.425 ;
        RECT 31.835 106.975 32.055 107.255 ;
        RECT 32.235 107.145 32.775 107.515 ;
        RECT 33.120 107.405 33.290 108.025 ;
        RECT 33.465 107.685 33.635 108.745 ;
        RECT 33.845 107.735 34.135 108.575 ;
        RECT 34.305 107.905 34.475 108.745 ;
        RECT 34.685 107.735 34.935 108.575 ;
        RECT 35.145 107.905 35.315 108.745 ;
        RECT 33.845 107.565 35.570 107.735 ;
        RECT 35.795 107.580 36.085 108.745 ;
        RECT 36.315 107.605 36.525 108.745 ;
        RECT 36.695 107.595 37.025 108.575 ;
        RECT 37.195 107.605 37.425 108.745 ;
        RECT 38.155 107.605 38.365 108.745 ;
        RECT 38.535 107.595 38.865 108.575 ;
        RECT 39.035 107.605 39.265 108.745 ;
        RECT 39.935 107.655 43.445 108.745 ;
        RECT 31.835 106.805 32.365 106.975 ;
        RECT 30.145 106.385 30.495 106.555 ;
        RECT 30.715 106.365 31.665 106.645 ;
        RECT 31.835 106.195 32.025 106.635 ;
        RECT 32.195 106.575 32.365 106.805 ;
        RECT 32.535 106.745 32.775 107.145 ;
        RECT 32.945 107.395 33.290 107.405 ;
        RECT 32.945 107.185 34.975 107.395 ;
        RECT 32.945 106.930 33.270 107.185 ;
        RECT 35.160 107.015 35.570 107.565 ;
        RECT 32.945 106.575 33.265 106.930 ;
        RECT 32.195 106.405 33.265 106.575 ;
        RECT 33.465 106.195 33.635 107.005 ;
        RECT 33.805 106.845 35.570 107.015 ;
        RECT 33.805 106.365 34.135 106.845 ;
        RECT 34.305 106.195 34.475 106.665 ;
        RECT 34.645 106.365 34.975 106.845 ;
        RECT 35.145 106.195 35.315 106.665 ;
        RECT 35.795 106.195 36.085 106.920 ;
        RECT 36.315 106.195 36.525 107.015 ;
        RECT 36.695 106.995 36.945 107.595 ;
        RECT 37.115 107.185 37.445 107.435 ;
        RECT 36.695 106.365 37.025 106.995 ;
        RECT 37.195 106.195 37.425 107.015 ;
        RECT 38.155 106.195 38.365 107.015 ;
        RECT 38.535 106.995 38.785 107.595 ;
        RECT 38.955 107.185 39.285 107.435 ;
        RECT 39.935 107.135 41.625 107.655 ;
        RECT 43.675 107.605 43.885 108.745 ;
        RECT 44.055 107.595 44.385 108.575 ;
        RECT 44.555 107.605 44.785 108.745 ;
        RECT 45.305 107.905 45.475 108.745 ;
        RECT 45.685 107.735 45.935 108.575 ;
        RECT 46.145 107.905 46.315 108.745 ;
        RECT 46.485 107.735 46.775 108.575 ;
        RECT 38.535 106.365 38.865 106.995 ;
        RECT 39.035 106.195 39.265 107.015 ;
        RECT 41.795 106.965 43.445 107.485 ;
        RECT 39.935 106.195 43.445 106.965 ;
        RECT 43.675 106.195 43.885 107.015 ;
        RECT 44.055 106.995 44.305 107.595 ;
        RECT 45.050 107.565 46.775 107.735 ;
        RECT 46.985 107.685 47.155 108.745 ;
        RECT 47.450 108.365 47.780 108.745 ;
        RECT 47.960 108.195 48.130 108.485 ;
        RECT 48.300 108.285 48.550 108.745 ;
        RECT 47.330 108.025 48.130 108.195 ;
        RECT 48.720 108.235 49.590 108.575 ;
        RECT 44.475 107.185 44.805 107.435 ;
        RECT 45.050 107.015 45.460 107.565 ;
        RECT 47.330 107.405 47.500 108.025 ;
        RECT 48.720 107.855 48.890 108.235 ;
        RECT 49.825 108.115 49.995 108.575 ;
        RECT 50.165 108.285 50.535 108.745 ;
        RECT 50.830 108.145 51.000 108.485 ;
        RECT 51.170 108.315 51.500 108.745 ;
        RECT 51.735 108.145 51.905 108.485 ;
        RECT 47.670 107.685 48.890 107.855 ;
        RECT 49.060 107.775 49.520 108.065 ;
        RECT 49.825 107.945 50.385 108.115 ;
        RECT 50.830 107.975 51.905 108.145 ;
        RECT 52.075 108.245 52.755 108.575 ;
        RECT 52.970 108.245 53.220 108.575 ;
        RECT 53.390 108.285 53.640 108.745 ;
        RECT 50.215 107.805 50.385 107.945 ;
        RECT 49.060 107.765 50.025 107.775 ;
        RECT 48.720 107.595 48.890 107.685 ;
        RECT 49.350 107.605 50.025 107.765 ;
        RECT 47.330 107.395 47.675 107.405 ;
        RECT 45.645 107.185 47.675 107.395 ;
        RECT 44.055 106.365 44.385 106.995 ;
        RECT 44.555 106.195 44.785 107.015 ;
        RECT 45.050 106.845 46.815 107.015 ;
        RECT 45.305 106.195 45.475 106.665 ;
        RECT 45.645 106.365 45.975 106.845 ;
        RECT 46.145 106.195 46.315 106.665 ;
        RECT 46.485 106.365 46.815 106.845 ;
        RECT 46.985 106.195 47.155 107.005 ;
        RECT 47.350 106.930 47.675 107.185 ;
        RECT 47.355 106.575 47.675 106.930 ;
        RECT 47.845 107.145 48.385 107.515 ;
        RECT 48.720 107.425 49.125 107.595 ;
        RECT 47.845 106.745 48.085 107.145 ;
        RECT 48.565 106.975 48.785 107.255 ;
        RECT 48.255 106.805 48.785 106.975 ;
        RECT 48.255 106.575 48.425 106.805 ;
        RECT 48.955 106.645 49.125 107.425 ;
        RECT 49.295 106.815 49.645 107.435 ;
        RECT 49.815 106.815 50.025 107.605 ;
        RECT 50.215 107.635 51.715 107.805 ;
        RECT 50.215 106.945 50.385 107.635 ;
        RECT 52.075 107.465 52.245 108.245 ;
        RECT 53.050 108.115 53.220 108.245 ;
        RECT 50.555 107.295 52.245 107.465 ;
        RECT 52.415 107.685 52.880 108.075 ;
        RECT 53.050 107.945 53.445 108.115 ;
        RECT 50.555 107.115 50.725 107.295 ;
        RECT 47.355 106.405 48.425 106.575 ;
        RECT 48.595 106.195 48.785 106.635 ;
        RECT 48.955 106.365 49.905 106.645 ;
        RECT 50.215 106.555 50.475 106.945 ;
        RECT 50.895 106.875 51.685 107.125 ;
        RECT 50.125 106.385 50.475 106.555 ;
        RECT 50.685 106.195 51.015 106.655 ;
        RECT 51.890 106.585 52.060 107.295 ;
        RECT 52.415 107.095 52.585 107.685 ;
        RECT 52.230 106.875 52.585 107.095 ;
        RECT 52.755 106.875 53.105 107.495 ;
        RECT 53.275 106.585 53.445 107.945 ;
        RECT 53.810 107.775 54.135 108.560 ;
        RECT 53.615 106.725 54.075 107.775 ;
        RECT 51.890 106.415 52.745 106.585 ;
        RECT 52.950 106.415 53.445 106.585 ;
        RECT 53.615 106.195 53.945 106.555 ;
        RECT 54.305 106.455 54.475 108.575 ;
        RECT 54.645 108.245 54.975 108.745 ;
        RECT 55.145 108.075 55.400 108.575 ;
        RECT 54.650 107.905 55.400 108.075 ;
        RECT 54.650 106.915 54.880 107.905 ;
        RECT 55.050 107.085 55.400 107.735 ;
        RECT 55.635 107.605 55.845 108.745 ;
        RECT 56.015 107.595 56.345 108.575 ;
        RECT 56.515 107.605 56.745 108.745 ;
        RECT 57.455 107.605 57.685 108.745 ;
        RECT 57.855 107.595 58.185 108.575 ;
        RECT 58.355 107.605 58.565 108.745 ;
        RECT 58.795 107.655 61.385 108.745 ;
        RECT 54.650 106.745 55.400 106.915 ;
        RECT 54.645 106.195 54.975 106.575 ;
        RECT 55.145 106.455 55.400 106.745 ;
        RECT 55.635 106.195 55.845 107.015 ;
        RECT 56.015 106.995 56.265 107.595 ;
        RECT 56.435 107.185 56.765 107.435 ;
        RECT 57.435 107.185 57.765 107.435 ;
        RECT 56.015 106.365 56.345 106.995 ;
        RECT 56.515 106.195 56.745 107.015 ;
        RECT 57.455 106.195 57.685 107.015 ;
        RECT 57.935 106.995 58.185 107.595 ;
        RECT 58.795 107.135 60.005 107.655 ;
        RECT 61.555 107.580 61.845 108.745 ;
        RECT 62.325 107.905 62.495 108.745 ;
        RECT 62.705 107.735 62.955 108.575 ;
        RECT 63.165 107.905 63.335 108.745 ;
        RECT 63.505 107.735 63.795 108.575 ;
        RECT 62.070 107.565 63.795 107.735 ;
        RECT 64.005 107.685 64.175 108.745 ;
        RECT 64.470 108.365 64.800 108.745 ;
        RECT 64.980 108.195 65.150 108.485 ;
        RECT 65.320 108.285 65.570 108.745 ;
        RECT 64.350 108.025 65.150 108.195 ;
        RECT 65.740 108.235 66.610 108.575 ;
        RECT 57.855 106.365 58.185 106.995 ;
        RECT 58.355 106.195 58.565 107.015 ;
        RECT 60.175 106.965 61.385 107.485 ;
        RECT 58.795 106.195 61.385 106.965 ;
        RECT 62.070 107.015 62.480 107.565 ;
        RECT 64.350 107.405 64.520 108.025 ;
        RECT 65.740 107.855 65.910 108.235 ;
        RECT 66.845 108.115 67.015 108.575 ;
        RECT 67.185 108.285 67.555 108.745 ;
        RECT 67.850 108.145 68.020 108.485 ;
        RECT 68.190 108.315 68.520 108.745 ;
        RECT 68.755 108.145 68.925 108.485 ;
        RECT 64.690 107.685 65.910 107.855 ;
        RECT 66.080 107.775 66.540 108.065 ;
        RECT 66.845 107.945 67.405 108.115 ;
        RECT 67.850 107.975 68.925 108.145 ;
        RECT 69.095 108.245 69.775 108.575 ;
        RECT 69.990 108.245 70.240 108.575 ;
        RECT 70.410 108.285 70.660 108.745 ;
        RECT 67.235 107.805 67.405 107.945 ;
        RECT 66.080 107.765 67.045 107.775 ;
        RECT 65.740 107.595 65.910 107.685 ;
        RECT 66.370 107.605 67.045 107.765 ;
        RECT 64.350 107.395 64.695 107.405 ;
        RECT 62.665 107.185 64.695 107.395 ;
        RECT 61.555 106.195 61.845 106.920 ;
        RECT 62.070 106.845 63.835 107.015 ;
        RECT 62.325 106.195 62.495 106.665 ;
        RECT 62.665 106.365 62.995 106.845 ;
        RECT 63.165 106.195 63.335 106.665 ;
        RECT 63.505 106.365 63.835 106.845 ;
        RECT 64.005 106.195 64.175 107.005 ;
        RECT 64.370 106.930 64.695 107.185 ;
        RECT 64.375 106.575 64.695 106.930 ;
        RECT 64.865 107.145 65.405 107.515 ;
        RECT 65.740 107.425 66.145 107.595 ;
        RECT 64.865 106.745 65.105 107.145 ;
        RECT 65.585 106.975 65.805 107.255 ;
        RECT 65.275 106.805 65.805 106.975 ;
        RECT 65.275 106.575 65.445 106.805 ;
        RECT 65.975 106.645 66.145 107.425 ;
        RECT 66.315 106.815 66.665 107.435 ;
        RECT 66.835 106.815 67.045 107.605 ;
        RECT 67.235 107.635 68.735 107.805 ;
        RECT 67.235 106.945 67.405 107.635 ;
        RECT 69.095 107.465 69.265 108.245 ;
        RECT 70.070 108.115 70.240 108.245 ;
        RECT 67.575 107.295 69.265 107.465 ;
        RECT 69.435 107.685 69.900 108.075 ;
        RECT 70.070 107.945 70.465 108.115 ;
        RECT 67.575 107.115 67.745 107.295 ;
        RECT 64.375 106.405 65.445 106.575 ;
        RECT 65.615 106.195 65.805 106.635 ;
        RECT 65.975 106.365 66.925 106.645 ;
        RECT 67.235 106.555 67.495 106.945 ;
        RECT 67.915 106.875 68.705 107.125 ;
        RECT 67.145 106.385 67.495 106.555 ;
        RECT 67.705 106.195 68.035 106.655 ;
        RECT 68.910 106.585 69.080 107.295 ;
        RECT 69.435 107.095 69.605 107.685 ;
        RECT 69.250 106.875 69.605 107.095 ;
        RECT 69.775 106.875 70.125 107.495 ;
        RECT 70.295 106.585 70.465 107.945 ;
        RECT 70.830 107.775 71.155 108.560 ;
        RECT 70.635 106.725 71.095 107.775 ;
        RECT 68.910 106.415 69.765 106.585 ;
        RECT 69.970 106.415 70.465 106.585 ;
        RECT 70.635 106.195 70.965 106.555 ;
        RECT 71.325 106.455 71.495 108.575 ;
        RECT 71.665 108.245 71.995 108.745 ;
        RECT 72.165 108.075 72.420 108.575 ;
        RECT 71.670 107.905 72.420 108.075 ;
        RECT 73.825 107.905 73.995 108.745 ;
        RECT 71.670 106.915 71.900 107.905 ;
        RECT 74.205 107.735 74.455 108.575 ;
        RECT 74.665 107.905 74.835 108.745 ;
        RECT 75.005 107.735 75.295 108.575 ;
        RECT 72.070 107.085 72.420 107.735 ;
        RECT 73.570 107.565 75.295 107.735 ;
        RECT 75.505 107.685 75.675 108.745 ;
        RECT 75.970 108.365 76.300 108.745 ;
        RECT 76.480 108.195 76.650 108.485 ;
        RECT 76.820 108.285 77.070 108.745 ;
        RECT 75.850 108.025 76.650 108.195 ;
        RECT 77.240 108.235 78.110 108.575 ;
        RECT 73.570 107.015 73.980 107.565 ;
        RECT 75.850 107.405 76.020 108.025 ;
        RECT 77.240 107.855 77.410 108.235 ;
        RECT 78.345 108.115 78.515 108.575 ;
        RECT 78.685 108.285 79.055 108.745 ;
        RECT 79.350 108.145 79.520 108.485 ;
        RECT 79.690 108.315 80.020 108.745 ;
        RECT 80.255 108.145 80.425 108.485 ;
        RECT 76.190 107.685 77.410 107.855 ;
        RECT 77.580 107.775 78.040 108.065 ;
        RECT 78.345 107.945 78.905 108.115 ;
        RECT 79.350 107.975 80.425 108.145 ;
        RECT 80.595 108.245 81.275 108.575 ;
        RECT 81.490 108.245 81.740 108.575 ;
        RECT 81.910 108.285 82.160 108.745 ;
        RECT 78.735 107.805 78.905 107.945 ;
        RECT 77.580 107.765 78.545 107.775 ;
        RECT 77.240 107.595 77.410 107.685 ;
        RECT 77.870 107.605 78.545 107.765 ;
        RECT 75.850 107.395 76.195 107.405 ;
        RECT 74.165 107.185 76.195 107.395 ;
        RECT 71.670 106.745 72.420 106.915 ;
        RECT 73.570 106.845 75.335 107.015 ;
        RECT 71.665 106.195 71.995 106.575 ;
        RECT 72.165 106.455 72.420 106.745 ;
        RECT 73.825 106.195 73.995 106.665 ;
        RECT 74.165 106.365 74.495 106.845 ;
        RECT 74.665 106.195 74.835 106.665 ;
        RECT 75.005 106.365 75.335 106.845 ;
        RECT 75.505 106.195 75.675 107.005 ;
        RECT 75.870 106.930 76.195 107.185 ;
        RECT 75.875 106.575 76.195 106.930 ;
        RECT 76.365 107.145 76.905 107.515 ;
        RECT 77.240 107.425 77.645 107.595 ;
        RECT 76.365 106.745 76.605 107.145 ;
        RECT 77.085 106.975 77.305 107.255 ;
        RECT 76.775 106.805 77.305 106.975 ;
        RECT 76.775 106.575 76.945 106.805 ;
        RECT 77.475 106.645 77.645 107.425 ;
        RECT 77.815 106.815 78.165 107.435 ;
        RECT 78.335 106.815 78.545 107.605 ;
        RECT 78.735 107.635 80.235 107.805 ;
        RECT 78.735 106.945 78.905 107.635 ;
        RECT 80.595 107.465 80.765 108.245 ;
        RECT 81.570 108.115 81.740 108.245 ;
        RECT 79.075 107.295 80.765 107.465 ;
        RECT 80.935 107.685 81.400 108.075 ;
        RECT 81.570 107.945 81.965 108.115 ;
        RECT 79.075 107.115 79.245 107.295 ;
        RECT 75.875 106.405 76.945 106.575 ;
        RECT 77.115 106.195 77.305 106.635 ;
        RECT 77.475 106.365 78.425 106.645 ;
        RECT 78.735 106.555 78.995 106.945 ;
        RECT 79.415 106.875 80.205 107.125 ;
        RECT 78.645 106.385 78.995 106.555 ;
        RECT 79.205 106.195 79.535 106.655 ;
        RECT 80.410 106.585 80.580 107.295 ;
        RECT 80.935 107.095 81.105 107.685 ;
        RECT 80.750 106.875 81.105 107.095 ;
        RECT 81.275 106.875 81.625 107.495 ;
        RECT 81.795 106.585 81.965 107.945 ;
        RECT 82.330 107.775 82.655 108.560 ;
        RECT 82.135 106.725 82.595 107.775 ;
        RECT 80.410 106.415 81.265 106.585 ;
        RECT 81.470 106.415 81.965 106.585 ;
        RECT 82.135 106.195 82.465 106.555 ;
        RECT 82.825 106.455 82.995 108.575 ;
        RECT 83.165 108.245 83.495 108.745 ;
        RECT 83.665 108.075 83.920 108.575 ;
        RECT 83.170 107.905 83.920 108.075 ;
        RECT 83.170 106.915 83.400 107.905 ;
        RECT 83.570 107.085 83.920 107.735 ;
        RECT 84.155 107.605 84.365 108.745 ;
        RECT 84.535 107.595 84.865 108.575 ;
        RECT 85.035 107.605 85.265 108.745 ;
        RECT 85.975 107.605 86.205 108.745 ;
        RECT 86.375 107.595 86.705 108.575 ;
        RECT 86.875 107.605 87.085 108.745 ;
        RECT 83.170 106.745 83.920 106.915 ;
        RECT 83.165 106.195 83.495 106.575 ;
        RECT 83.665 106.455 83.920 106.745 ;
        RECT 84.155 106.195 84.365 107.015 ;
        RECT 84.535 106.995 84.785 107.595 ;
        RECT 84.955 107.185 85.285 107.435 ;
        RECT 85.955 107.185 86.285 107.435 ;
        RECT 84.535 106.365 84.865 106.995 ;
        RECT 85.035 106.195 85.265 107.015 ;
        RECT 85.975 106.195 86.205 107.015 ;
        RECT 86.455 106.995 86.705 107.595 ;
        RECT 87.315 107.580 87.605 108.745 ;
        RECT 88.085 107.905 88.255 108.745 ;
        RECT 88.465 107.735 88.715 108.575 ;
        RECT 88.925 107.905 89.095 108.745 ;
        RECT 89.265 107.735 89.555 108.575 ;
        RECT 87.830 107.565 89.555 107.735 ;
        RECT 89.765 107.685 89.935 108.745 ;
        RECT 90.230 108.365 90.560 108.745 ;
        RECT 90.740 108.195 90.910 108.485 ;
        RECT 91.080 108.285 91.330 108.745 ;
        RECT 90.110 108.025 90.910 108.195 ;
        RECT 91.500 108.235 92.370 108.575 ;
        RECT 87.830 107.015 88.240 107.565 ;
        RECT 90.110 107.405 90.280 108.025 ;
        RECT 91.500 107.855 91.670 108.235 ;
        RECT 92.605 108.115 92.775 108.575 ;
        RECT 92.945 108.285 93.315 108.745 ;
        RECT 93.610 108.145 93.780 108.485 ;
        RECT 93.950 108.315 94.280 108.745 ;
        RECT 94.515 108.145 94.685 108.485 ;
        RECT 90.450 107.685 91.670 107.855 ;
        RECT 91.840 107.775 92.300 108.065 ;
        RECT 92.605 107.945 93.165 108.115 ;
        RECT 93.610 107.975 94.685 108.145 ;
        RECT 94.855 108.245 95.535 108.575 ;
        RECT 95.750 108.245 96.000 108.575 ;
        RECT 96.170 108.285 96.420 108.745 ;
        RECT 92.995 107.805 93.165 107.945 ;
        RECT 91.840 107.765 92.805 107.775 ;
        RECT 91.500 107.595 91.670 107.685 ;
        RECT 92.130 107.605 92.805 107.765 ;
        RECT 90.110 107.395 90.455 107.405 ;
        RECT 88.425 107.185 90.455 107.395 ;
        RECT 86.375 106.365 86.705 106.995 ;
        RECT 86.875 106.195 87.085 107.015 ;
        RECT 87.315 106.195 87.605 106.920 ;
        RECT 87.830 106.845 89.595 107.015 ;
        RECT 88.085 106.195 88.255 106.665 ;
        RECT 88.425 106.365 88.755 106.845 ;
        RECT 88.925 106.195 89.095 106.665 ;
        RECT 89.265 106.365 89.595 106.845 ;
        RECT 89.765 106.195 89.935 107.005 ;
        RECT 90.130 106.930 90.455 107.185 ;
        RECT 90.135 106.575 90.455 106.930 ;
        RECT 90.625 107.145 91.165 107.515 ;
        RECT 91.500 107.425 91.905 107.595 ;
        RECT 90.625 106.745 90.865 107.145 ;
        RECT 91.345 106.975 91.565 107.255 ;
        RECT 91.035 106.805 91.565 106.975 ;
        RECT 91.035 106.575 91.205 106.805 ;
        RECT 91.735 106.645 91.905 107.425 ;
        RECT 92.075 106.815 92.425 107.435 ;
        RECT 92.595 106.815 92.805 107.605 ;
        RECT 92.995 107.635 94.495 107.805 ;
        RECT 92.995 106.945 93.165 107.635 ;
        RECT 94.855 107.465 95.025 108.245 ;
        RECT 95.830 108.115 96.000 108.245 ;
        RECT 93.335 107.295 95.025 107.465 ;
        RECT 95.195 107.685 95.660 108.075 ;
        RECT 95.830 107.945 96.225 108.115 ;
        RECT 93.335 107.115 93.505 107.295 ;
        RECT 90.135 106.405 91.205 106.575 ;
        RECT 91.375 106.195 91.565 106.635 ;
        RECT 91.735 106.365 92.685 106.645 ;
        RECT 92.995 106.555 93.255 106.945 ;
        RECT 93.675 106.875 94.465 107.125 ;
        RECT 92.905 106.385 93.255 106.555 ;
        RECT 93.465 106.195 93.795 106.655 ;
        RECT 94.670 106.585 94.840 107.295 ;
        RECT 95.195 107.095 95.365 107.685 ;
        RECT 95.010 106.875 95.365 107.095 ;
        RECT 95.535 106.875 95.885 107.495 ;
        RECT 96.055 106.585 96.225 107.945 ;
        RECT 96.590 107.775 96.915 108.560 ;
        RECT 96.395 106.725 96.855 107.775 ;
        RECT 94.670 106.415 95.525 106.585 ;
        RECT 95.730 106.415 96.225 106.585 ;
        RECT 96.395 106.195 96.725 106.555 ;
        RECT 97.085 106.455 97.255 108.575 ;
        RECT 97.425 108.245 97.755 108.745 ;
        RECT 97.925 108.075 98.180 108.575 ;
        RECT 97.430 107.905 98.180 108.075 ;
        RECT 99.280 108.075 99.535 108.575 ;
        RECT 99.705 108.245 100.035 108.745 ;
        RECT 99.280 107.905 100.030 108.075 ;
        RECT 97.430 106.915 97.660 107.905 ;
        RECT 97.830 107.085 98.180 107.735 ;
        RECT 99.280 107.085 99.630 107.735 ;
        RECT 99.800 106.915 100.030 107.905 ;
        RECT 97.430 106.745 98.180 106.915 ;
        RECT 97.425 106.195 97.755 106.575 ;
        RECT 97.925 106.455 98.180 106.745 ;
        RECT 99.280 106.745 100.030 106.915 ;
        RECT 99.280 106.455 99.535 106.745 ;
        RECT 99.705 106.195 100.035 106.575 ;
        RECT 100.205 106.455 100.375 108.575 ;
        RECT 100.545 107.775 100.870 108.560 ;
        RECT 101.040 108.285 101.290 108.745 ;
        RECT 101.460 108.245 101.710 108.575 ;
        RECT 101.925 108.245 102.605 108.575 ;
        RECT 101.460 108.115 101.630 108.245 ;
        RECT 101.235 107.945 101.630 108.115 ;
        RECT 100.605 106.725 101.065 107.775 ;
        RECT 101.235 106.585 101.405 107.945 ;
        RECT 101.800 107.685 102.265 108.075 ;
        RECT 101.575 106.875 101.925 107.495 ;
        RECT 102.095 107.095 102.265 107.685 ;
        RECT 102.435 107.465 102.605 108.245 ;
        RECT 102.775 108.145 102.945 108.485 ;
        RECT 103.180 108.315 103.510 108.745 ;
        RECT 103.680 108.145 103.850 108.485 ;
        RECT 104.145 108.285 104.515 108.745 ;
        RECT 102.775 107.975 103.850 108.145 ;
        RECT 104.685 108.115 104.855 108.575 ;
        RECT 105.090 108.235 105.960 108.575 ;
        RECT 106.130 108.285 106.380 108.745 ;
        RECT 104.295 107.945 104.855 108.115 ;
        RECT 104.295 107.805 104.465 107.945 ;
        RECT 102.965 107.635 104.465 107.805 ;
        RECT 105.160 107.775 105.620 108.065 ;
        RECT 102.435 107.295 104.125 107.465 ;
        RECT 102.095 106.875 102.450 107.095 ;
        RECT 102.620 106.585 102.790 107.295 ;
        RECT 102.995 106.875 103.785 107.125 ;
        RECT 103.955 107.115 104.125 107.295 ;
        RECT 104.295 106.945 104.465 107.635 ;
        RECT 100.735 106.195 101.065 106.555 ;
        RECT 101.235 106.415 101.730 106.585 ;
        RECT 101.935 106.415 102.790 106.585 ;
        RECT 103.665 106.195 103.995 106.655 ;
        RECT 104.205 106.555 104.465 106.945 ;
        RECT 104.655 107.765 105.620 107.775 ;
        RECT 105.790 107.855 105.960 108.235 ;
        RECT 106.550 108.195 106.720 108.485 ;
        RECT 106.900 108.365 107.230 108.745 ;
        RECT 106.550 108.025 107.350 108.195 ;
        RECT 104.655 107.605 105.330 107.765 ;
        RECT 105.790 107.685 107.010 107.855 ;
        RECT 104.655 106.815 104.865 107.605 ;
        RECT 105.790 107.595 105.960 107.685 ;
        RECT 105.035 106.815 105.385 107.435 ;
        RECT 105.555 107.425 105.960 107.595 ;
        RECT 105.555 106.645 105.725 107.425 ;
        RECT 105.895 106.975 106.115 107.255 ;
        RECT 106.295 107.145 106.835 107.515 ;
        RECT 107.180 107.405 107.350 108.025 ;
        RECT 107.525 107.685 107.695 108.745 ;
        RECT 107.905 107.735 108.195 108.575 ;
        RECT 108.365 107.905 108.535 108.745 ;
        RECT 108.745 107.735 108.995 108.575 ;
        RECT 109.205 107.905 109.375 108.745 ;
        RECT 107.905 107.565 109.630 107.735 ;
        RECT 105.895 106.805 106.425 106.975 ;
        RECT 104.205 106.385 104.555 106.555 ;
        RECT 104.775 106.365 105.725 106.645 ;
        RECT 105.895 106.195 106.085 106.635 ;
        RECT 106.255 106.575 106.425 106.805 ;
        RECT 106.595 106.745 106.835 107.145 ;
        RECT 107.005 107.395 107.350 107.405 ;
        RECT 107.005 107.185 109.035 107.395 ;
        RECT 107.005 106.930 107.330 107.185 ;
        RECT 109.220 107.015 109.630 107.565 ;
        RECT 107.005 106.575 107.325 106.930 ;
        RECT 106.255 106.405 107.325 106.575 ;
        RECT 107.525 106.195 107.695 107.005 ;
        RECT 107.865 106.845 109.630 107.015 ;
        RECT 110.775 107.670 111.045 108.575 ;
        RECT 111.215 107.985 111.545 108.745 ;
        RECT 111.725 107.815 111.905 108.575 ;
        RECT 110.775 106.870 110.955 107.670 ;
        RECT 111.230 107.645 111.905 107.815 ;
        RECT 112.155 107.655 113.365 108.745 ;
        RECT 111.230 107.500 111.400 107.645 ;
        RECT 111.125 107.170 111.400 107.500 ;
        RECT 111.230 106.915 111.400 107.170 ;
        RECT 111.625 107.095 111.965 107.465 ;
        RECT 112.155 107.115 112.675 107.655 ;
        RECT 112.845 106.945 113.365 107.485 ;
        RECT 107.865 106.365 108.195 106.845 ;
        RECT 108.365 106.195 108.535 106.665 ;
        RECT 108.705 106.365 109.035 106.845 ;
        RECT 109.205 106.195 109.375 106.665 ;
        RECT 110.775 106.365 111.035 106.870 ;
        RECT 111.230 106.745 111.895 106.915 ;
        RECT 111.215 106.195 111.545 106.575 ;
        RECT 111.725 106.365 111.895 106.745 ;
        RECT 112.155 106.195 113.365 106.945 ;
        RECT 11.330 106.025 113.450 106.195 ;
        RECT 11.415 105.275 12.625 106.025 ;
        RECT 11.415 104.735 11.935 105.275 ;
        RECT 13.255 105.255 15.845 106.025 ;
        RECT 16.020 105.480 21.365 106.025 ;
        RECT 12.105 104.565 12.625 105.105 ;
        RECT 11.415 103.475 12.625 104.565 ;
        RECT 13.255 104.565 14.465 105.085 ;
        RECT 14.635 104.735 15.845 105.255 ;
        RECT 13.255 103.475 15.845 104.565 ;
        RECT 17.610 103.910 17.960 105.160 ;
        RECT 19.440 104.650 19.780 105.480 ;
        RECT 21.595 105.205 21.805 106.025 ;
        RECT 21.975 105.225 22.305 105.855 ;
        RECT 21.975 104.625 22.225 105.225 ;
        RECT 22.475 105.205 22.705 106.025 ;
        RECT 22.915 105.300 23.205 106.025 ;
        RECT 23.685 105.555 23.855 106.025 ;
        RECT 24.025 105.375 24.355 105.855 ;
        RECT 24.525 105.555 24.695 106.025 ;
        RECT 24.865 105.375 25.195 105.855 ;
        RECT 23.430 105.205 25.195 105.375 ;
        RECT 25.365 105.215 25.535 106.025 ;
        RECT 25.735 105.645 26.805 105.815 ;
        RECT 25.735 105.290 26.055 105.645 ;
        RECT 22.395 104.785 22.725 105.035 ;
        RECT 23.430 104.655 23.840 105.205 ;
        RECT 25.730 105.035 26.055 105.290 ;
        RECT 24.025 104.825 26.055 105.035 ;
        RECT 25.710 104.815 26.055 104.825 ;
        RECT 26.225 105.075 26.465 105.475 ;
        RECT 26.635 105.415 26.805 105.645 ;
        RECT 26.975 105.585 27.165 106.025 ;
        RECT 27.335 105.575 28.285 105.855 ;
        RECT 28.505 105.665 28.855 105.835 ;
        RECT 26.635 105.245 27.165 105.415 ;
        RECT 16.020 103.475 21.365 103.910 ;
        RECT 21.595 103.475 21.805 104.615 ;
        RECT 21.975 103.645 22.305 104.625 ;
        RECT 22.475 103.475 22.705 104.615 ;
        RECT 22.915 103.475 23.205 104.640 ;
        RECT 23.430 104.485 25.155 104.655 ;
        RECT 23.685 103.475 23.855 104.315 ;
        RECT 24.065 103.645 24.315 104.485 ;
        RECT 24.525 103.475 24.695 104.315 ;
        RECT 24.865 103.645 25.155 104.485 ;
        RECT 25.365 103.475 25.535 104.535 ;
        RECT 25.710 104.195 25.880 104.815 ;
        RECT 26.225 104.705 26.765 105.075 ;
        RECT 26.945 104.965 27.165 105.245 ;
        RECT 27.335 104.795 27.505 105.575 ;
        RECT 27.100 104.625 27.505 104.795 ;
        RECT 27.675 104.785 28.025 105.405 ;
        RECT 27.100 104.535 27.270 104.625 ;
        RECT 28.195 104.615 28.405 105.405 ;
        RECT 26.050 104.365 27.270 104.535 ;
        RECT 27.730 104.455 28.405 104.615 ;
        RECT 25.710 104.025 26.510 104.195 ;
        RECT 25.830 103.475 26.160 103.855 ;
        RECT 26.340 103.735 26.510 104.025 ;
        RECT 27.100 103.985 27.270 104.365 ;
        RECT 27.440 104.445 28.405 104.455 ;
        RECT 28.595 105.275 28.855 105.665 ;
        RECT 29.065 105.565 29.395 106.025 ;
        RECT 30.270 105.635 31.125 105.805 ;
        RECT 31.330 105.635 31.825 105.805 ;
        RECT 31.995 105.665 32.325 106.025 ;
        RECT 28.595 104.585 28.765 105.275 ;
        RECT 28.935 104.925 29.105 105.105 ;
        RECT 29.275 105.095 30.065 105.345 ;
        RECT 30.270 104.925 30.440 105.635 ;
        RECT 30.610 105.125 30.965 105.345 ;
        RECT 28.935 104.755 30.625 104.925 ;
        RECT 27.440 104.155 27.900 104.445 ;
        RECT 28.595 104.415 30.095 104.585 ;
        RECT 28.595 104.275 28.765 104.415 ;
        RECT 28.205 104.105 28.765 104.275 ;
        RECT 26.680 103.475 26.930 103.935 ;
        RECT 27.100 103.645 27.970 103.985 ;
        RECT 28.205 103.645 28.375 104.105 ;
        RECT 29.210 104.075 30.285 104.245 ;
        RECT 28.545 103.475 28.915 103.935 ;
        RECT 29.210 103.735 29.380 104.075 ;
        RECT 29.550 103.475 29.880 103.905 ;
        RECT 30.115 103.735 30.285 104.075 ;
        RECT 30.455 103.975 30.625 104.755 ;
        RECT 30.795 104.535 30.965 105.125 ;
        RECT 31.135 104.725 31.485 105.345 ;
        RECT 30.795 104.145 31.260 104.535 ;
        RECT 31.655 104.275 31.825 105.635 ;
        RECT 31.995 104.445 32.455 105.495 ;
        RECT 31.430 104.105 31.825 104.275 ;
        RECT 31.430 103.975 31.600 104.105 ;
        RECT 30.455 103.645 31.135 103.975 ;
        RECT 31.350 103.645 31.600 103.975 ;
        RECT 31.770 103.475 32.020 103.935 ;
        RECT 32.190 103.660 32.515 104.445 ;
        RECT 32.685 103.645 32.855 105.765 ;
        RECT 33.025 105.645 33.355 106.025 ;
        RECT 33.525 105.475 33.780 105.765 ;
        RECT 33.030 105.305 33.780 105.475 ;
        RECT 33.030 104.315 33.260 105.305 ;
        RECT 33.955 105.255 35.625 106.025 ;
        RECT 35.795 105.300 36.085 106.025 ;
        RECT 36.255 105.275 37.465 106.025 ;
        RECT 37.640 105.480 42.985 106.025 ;
        RECT 43.160 105.480 48.505 106.025 ;
        RECT 33.430 104.485 33.780 105.135 ;
        RECT 33.955 104.565 34.705 105.085 ;
        RECT 34.875 104.735 35.625 105.255 ;
        RECT 33.030 104.145 33.780 104.315 ;
        RECT 33.025 103.475 33.355 103.975 ;
        RECT 33.525 103.645 33.780 104.145 ;
        RECT 33.955 103.475 35.625 104.565 ;
        RECT 35.795 103.475 36.085 104.640 ;
        RECT 36.255 104.565 36.775 105.105 ;
        RECT 36.945 104.735 37.465 105.275 ;
        RECT 36.255 103.475 37.465 104.565 ;
        RECT 39.230 103.910 39.580 105.160 ;
        RECT 41.060 104.650 41.400 105.480 ;
        RECT 44.750 103.910 45.100 105.160 ;
        RECT 46.580 104.650 46.920 105.480 ;
        RECT 48.675 105.300 48.965 106.025 ;
        RECT 49.195 105.205 49.405 106.025 ;
        RECT 49.575 105.225 49.905 105.855 ;
        RECT 37.640 103.475 42.985 103.910 ;
        RECT 43.160 103.475 48.505 103.910 ;
        RECT 48.675 103.475 48.965 104.640 ;
        RECT 49.575 104.625 49.825 105.225 ;
        RECT 50.075 105.205 50.305 106.025 ;
        RECT 50.520 105.480 55.865 106.025 ;
        RECT 56.040 105.480 61.385 106.025 ;
        RECT 49.995 104.785 50.325 105.035 ;
        RECT 49.195 103.475 49.405 104.615 ;
        RECT 49.575 103.645 49.905 104.625 ;
        RECT 50.075 103.475 50.305 104.615 ;
        RECT 52.110 103.910 52.460 105.160 ;
        RECT 53.940 104.650 54.280 105.480 ;
        RECT 57.630 103.910 57.980 105.160 ;
        RECT 59.460 104.650 59.800 105.480 ;
        RECT 61.555 105.300 61.845 106.025 ;
        RECT 62.015 105.255 63.685 106.025 ;
        RECT 63.860 105.475 64.115 105.765 ;
        RECT 64.285 105.645 64.615 106.025 ;
        RECT 63.860 105.305 64.610 105.475 ;
        RECT 50.520 103.475 55.865 103.910 ;
        RECT 56.040 103.475 61.385 103.910 ;
        RECT 61.555 103.475 61.845 104.640 ;
        RECT 62.015 104.565 62.765 105.085 ;
        RECT 62.935 104.735 63.685 105.255 ;
        RECT 62.015 103.475 63.685 104.565 ;
        RECT 63.860 104.485 64.210 105.135 ;
        RECT 64.380 104.315 64.610 105.305 ;
        RECT 63.860 104.145 64.610 104.315 ;
        RECT 63.860 103.645 64.115 104.145 ;
        RECT 64.285 103.475 64.615 103.975 ;
        RECT 64.785 103.645 64.955 105.765 ;
        RECT 65.315 105.665 65.645 106.025 ;
        RECT 65.815 105.635 66.310 105.805 ;
        RECT 66.515 105.635 67.370 105.805 ;
        RECT 65.185 104.445 65.645 105.495 ;
        RECT 65.125 103.660 65.450 104.445 ;
        RECT 65.815 104.275 65.985 105.635 ;
        RECT 66.155 104.725 66.505 105.345 ;
        RECT 66.675 105.125 67.030 105.345 ;
        RECT 66.675 104.535 66.845 105.125 ;
        RECT 67.200 104.925 67.370 105.635 ;
        RECT 68.245 105.565 68.575 106.025 ;
        RECT 68.785 105.665 69.135 105.835 ;
        RECT 67.575 105.095 68.365 105.345 ;
        RECT 68.785 105.275 69.045 105.665 ;
        RECT 69.355 105.575 70.305 105.855 ;
        RECT 70.475 105.585 70.665 106.025 ;
        RECT 70.835 105.645 71.905 105.815 ;
        RECT 68.535 104.925 68.705 105.105 ;
        RECT 65.815 104.105 66.210 104.275 ;
        RECT 66.380 104.145 66.845 104.535 ;
        RECT 67.015 104.755 68.705 104.925 ;
        RECT 66.040 103.975 66.210 104.105 ;
        RECT 67.015 103.975 67.185 104.755 ;
        RECT 68.875 104.585 69.045 105.275 ;
        RECT 67.545 104.415 69.045 104.585 ;
        RECT 69.235 104.615 69.445 105.405 ;
        RECT 69.615 104.785 69.965 105.405 ;
        RECT 70.135 104.795 70.305 105.575 ;
        RECT 70.835 105.415 71.005 105.645 ;
        RECT 70.475 105.245 71.005 105.415 ;
        RECT 70.475 104.965 70.695 105.245 ;
        RECT 71.175 105.075 71.415 105.475 ;
        RECT 70.135 104.625 70.540 104.795 ;
        RECT 70.875 104.705 71.415 105.075 ;
        RECT 71.585 105.290 71.905 105.645 ;
        RECT 71.585 105.035 71.910 105.290 ;
        RECT 72.105 105.215 72.275 106.025 ;
        RECT 72.445 105.375 72.775 105.855 ;
        RECT 72.945 105.555 73.115 106.025 ;
        RECT 73.285 105.375 73.615 105.855 ;
        RECT 73.785 105.555 73.955 106.025 ;
        RECT 72.445 105.205 74.210 105.375 ;
        RECT 74.435 105.300 74.725 106.025 ;
        RECT 74.955 105.205 75.165 106.025 ;
        RECT 75.335 105.225 75.665 105.855 ;
        RECT 71.585 104.825 73.615 105.035 ;
        RECT 71.585 104.815 71.930 104.825 ;
        RECT 69.235 104.455 69.910 104.615 ;
        RECT 70.370 104.535 70.540 104.625 ;
        RECT 69.235 104.445 70.200 104.455 ;
        RECT 68.875 104.275 69.045 104.415 ;
        RECT 65.620 103.475 65.870 103.935 ;
        RECT 66.040 103.645 66.290 103.975 ;
        RECT 66.505 103.645 67.185 103.975 ;
        RECT 67.355 104.075 68.430 104.245 ;
        RECT 68.875 104.105 69.435 104.275 ;
        RECT 69.740 104.155 70.200 104.445 ;
        RECT 70.370 104.365 71.590 104.535 ;
        RECT 67.355 103.735 67.525 104.075 ;
        RECT 67.760 103.475 68.090 103.905 ;
        RECT 68.260 103.735 68.430 104.075 ;
        RECT 68.725 103.475 69.095 103.935 ;
        RECT 69.265 103.645 69.435 104.105 ;
        RECT 70.370 103.985 70.540 104.365 ;
        RECT 71.760 104.195 71.930 104.815 ;
        RECT 73.800 104.655 74.210 105.205 ;
        RECT 69.670 103.645 70.540 103.985 ;
        RECT 71.130 104.025 71.930 104.195 ;
        RECT 70.710 103.475 70.960 103.935 ;
        RECT 71.130 103.735 71.300 104.025 ;
        RECT 71.480 103.475 71.810 103.855 ;
        RECT 72.105 103.475 72.275 104.535 ;
        RECT 72.485 104.485 74.210 104.655 ;
        RECT 72.485 103.645 72.775 104.485 ;
        RECT 72.945 103.475 73.115 104.315 ;
        RECT 73.325 103.645 73.575 104.485 ;
        RECT 73.785 103.475 73.955 104.315 ;
        RECT 74.435 103.475 74.725 104.640 ;
        RECT 75.335 104.625 75.585 105.225 ;
        RECT 75.835 105.205 76.065 106.025 ;
        RECT 76.275 105.275 77.485 106.025 ;
        RECT 75.755 104.785 76.085 105.035 ;
        RECT 74.955 103.475 75.165 104.615 ;
        RECT 75.335 103.645 75.665 104.625 ;
        RECT 75.835 103.475 76.065 104.615 ;
        RECT 76.275 104.565 76.795 105.105 ;
        RECT 76.965 104.735 77.485 105.275 ;
        RECT 77.715 105.205 77.925 106.025 ;
        RECT 78.095 105.225 78.425 105.855 ;
        RECT 78.095 104.625 78.345 105.225 ;
        RECT 78.595 105.205 78.825 106.025 ;
        RECT 79.035 105.255 81.625 106.025 ;
        RECT 81.800 105.480 87.145 106.025 ;
        RECT 78.515 104.785 78.845 105.035 ;
        RECT 76.275 103.475 77.485 104.565 ;
        RECT 77.715 103.475 77.925 104.615 ;
        RECT 78.095 103.645 78.425 104.625 ;
        RECT 78.595 103.475 78.825 104.615 ;
        RECT 79.035 104.565 80.245 105.085 ;
        RECT 80.415 104.735 81.625 105.255 ;
        RECT 79.035 103.475 81.625 104.565 ;
        RECT 83.390 103.910 83.740 105.160 ;
        RECT 85.220 104.650 85.560 105.480 ;
        RECT 87.315 105.300 87.605 106.025 ;
        RECT 88.275 105.205 88.505 106.025 ;
        RECT 88.675 105.225 89.005 105.855 ;
        RECT 88.255 104.785 88.585 105.035 ;
        RECT 81.800 103.475 87.145 103.910 ;
        RECT 87.315 103.475 87.605 104.640 ;
        RECT 88.755 104.625 89.005 105.225 ;
        RECT 89.175 105.205 89.385 106.025 ;
        RECT 89.620 105.475 89.875 105.765 ;
        RECT 90.045 105.645 90.375 106.025 ;
        RECT 89.620 105.305 90.370 105.475 ;
        RECT 88.275 103.475 88.505 104.615 ;
        RECT 88.675 103.645 89.005 104.625 ;
        RECT 89.175 103.475 89.385 104.615 ;
        RECT 89.620 104.485 89.970 105.135 ;
        RECT 90.140 104.315 90.370 105.305 ;
        RECT 89.620 104.145 90.370 104.315 ;
        RECT 89.620 103.645 89.875 104.145 ;
        RECT 90.045 103.475 90.375 103.975 ;
        RECT 90.545 103.645 90.715 105.765 ;
        RECT 91.075 105.665 91.405 106.025 ;
        RECT 91.575 105.635 92.070 105.805 ;
        RECT 92.275 105.635 93.130 105.805 ;
        RECT 90.945 104.445 91.405 105.495 ;
        RECT 90.885 103.660 91.210 104.445 ;
        RECT 91.575 104.275 91.745 105.635 ;
        RECT 91.915 104.725 92.265 105.345 ;
        RECT 92.435 105.125 92.790 105.345 ;
        RECT 92.435 104.535 92.605 105.125 ;
        RECT 92.960 104.925 93.130 105.635 ;
        RECT 94.005 105.565 94.335 106.025 ;
        RECT 94.545 105.665 94.895 105.835 ;
        RECT 93.335 105.095 94.125 105.345 ;
        RECT 94.545 105.275 94.805 105.665 ;
        RECT 95.115 105.575 96.065 105.855 ;
        RECT 96.235 105.585 96.425 106.025 ;
        RECT 96.595 105.645 97.665 105.815 ;
        RECT 94.295 104.925 94.465 105.105 ;
        RECT 91.575 104.105 91.970 104.275 ;
        RECT 92.140 104.145 92.605 104.535 ;
        RECT 92.775 104.755 94.465 104.925 ;
        RECT 91.800 103.975 91.970 104.105 ;
        RECT 92.775 103.975 92.945 104.755 ;
        RECT 94.635 104.585 94.805 105.275 ;
        RECT 93.305 104.415 94.805 104.585 ;
        RECT 94.995 104.615 95.205 105.405 ;
        RECT 95.375 104.785 95.725 105.405 ;
        RECT 95.895 104.795 96.065 105.575 ;
        RECT 96.595 105.415 96.765 105.645 ;
        RECT 96.235 105.245 96.765 105.415 ;
        RECT 96.235 104.965 96.455 105.245 ;
        RECT 96.935 105.075 97.175 105.475 ;
        RECT 95.895 104.625 96.300 104.795 ;
        RECT 96.635 104.705 97.175 105.075 ;
        RECT 97.345 105.290 97.665 105.645 ;
        RECT 97.345 105.035 97.670 105.290 ;
        RECT 97.865 105.215 98.035 106.025 ;
        RECT 98.205 105.375 98.535 105.855 ;
        RECT 98.705 105.555 98.875 106.025 ;
        RECT 99.045 105.375 99.375 105.855 ;
        RECT 99.545 105.555 99.715 106.025 ;
        RECT 98.205 105.205 99.970 105.375 ;
        RECT 100.195 105.300 100.485 106.025 ;
        RECT 100.715 105.205 100.925 106.025 ;
        RECT 101.095 105.225 101.425 105.855 ;
        RECT 97.345 104.825 99.375 105.035 ;
        RECT 97.345 104.815 97.690 104.825 ;
        RECT 94.995 104.455 95.670 104.615 ;
        RECT 96.130 104.535 96.300 104.625 ;
        RECT 94.995 104.445 95.960 104.455 ;
        RECT 94.635 104.275 94.805 104.415 ;
        RECT 91.380 103.475 91.630 103.935 ;
        RECT 91.800 103.645 92.050 103.975 ;
        RECT 92.265 103.645 92.945 103.975 ;
        RECT 93.115 104.075 94.190 104.245 ;
        RECT 94.635 104.105 95.195 104.275 ;
        RECT 95.500 104.155 95.960 104.445 ;
        RECT 96.130 104.365 97.350 104.535 ;
        RECT 93.115 103.735 93.285 104.075 ;
        RECT 93.520 103.475 93.850 103.905 ;
        RECT 94.020 103.735 94.190 104.075 ;
        RECT 94.485 103.475 94.855 103.935 ;
        RECT 95.025 103.645 95.195 104.105 ;
        RECT 96.130 103.985 96.300 104.365 ;
        RECT 97.520 104.195 97.690 104.815 ;
        RECT 99.560 104.655 99.970 105.205 ;
        RECT 95.430 103.645 96.300 103.985 ;
        RECT 96.890 104.025 97.690 104.195 ;
        RECT 96.470 103.475 96.720 103.935 ;
        RECT 96.890 103.735 97.060 104.025 ;
        RECT 97.240 103.475 97.570 103.855 ;
        RECT 97.865 103.475 98.035 104.535 ;
        RECT 98.245 104.485 99.970 104.655 ;
        RECT 98.245 103.645 98.535 104.485 ;
        RECT 98.705 103.475 98.875 104.315 ;
        RECT 99.085 103.645 99.335 104.485 ;
        RECT 99.545 103.475 99.715 104.315 ;
        RECT 100.195 103.475 100.485 104.640 ;
        RECT 101.095 104.625 101.345 105.225 ;
        RECT 101.595 105.205 101.825 106.025 ;
        RECT 102.035 105.275 103.245 106.025 ;
        RECT 101.515 104.785 101.845 105.035 ;
        RECT 100.715 103.475 100.925 104.615 ;
        RECT 101.095 103.645 101.425 104.625 ;
        RECT 101.595 103.475 101.825 104.615 ;
        RECT 102.035 104.565 102.555 105.105 ;
        RECT 102.725 104.735 103.245 105.275 ;
        RECT 103.475 105.205 103.685 106.025 ;
        RECT 103.855 105.225 104.185 105.855 ;
        RECT 103.855 104.625 104.105 105.225 ;
        RECT 104.355 105.205 104.585 106.025 ;
        RECT 105.755 105.205 105.985 106.025 ;
        RECT 106.155 105.225 106.485 105.855 ;
        RECT 104.275 104.785 104.605 105.035 ;
        RECT 105.735 104.785 106.065 105.035 ;
        RECT 106.235 104.625 106.485 105.225 ;
        RECT 106.655 105.205 106.865 106.025 ;
        RECT 107.095 105.275 108.305 106.025 ;
        RECT 102.035 103.475 103.245 104.565 ;
        RECT 103.475 103.475 103.685 104.615 ;
        RECT 103.855 103.645 104.185 104.625 ;
        RECT 104.355 103.475 104.585 104.615 ;
        RECT 105.755 103.475 105.985 104.615 ;
        RECT 106.155 103.645 106.485 104.625 ;
        RECT 106.655 103.475 106.865 104.615 ;
        RECT 107.095 104.565 107.615 105.105 ;
        RECT 107.785 104.735 108.305 105.275 ;
        RECT 108.475 105.255 111.985 106.025 ;
        RECT 112.155 105.275 113.365 106.025 ;
        RECT 108.475 104.565 110.165 105.085 ;
        RECT 110.335 104.735 111.985 105.255 ;
        RECT 112.155 104.565 112.675 105.105 ;
        RECT 112.845 104.735 113.365 105.275 ;
        RECT 107.095 103.475 108.305 104.565 ;
        RECT 108.475 103.475 111.985 104.565 ;
        RECT 112.155 103.475 113.365 104.565 ;
        RECT 11.330 103.305 113.450 103.475 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 11.330 203.790 113.450 204.270 ;
        RECT 11.330 201.070 113.450 201.550 ;
        RECT 64.875 200.530 65.165 200.575 ;
        RECT 67.995 200.530 68.285 200.575 ;
        RECT 69.885 200.530 70.175 200.575 ;
        RECT 64.875 200.390 70.175 200.530 ;
        RECT 64.875 200.345 65.165 200.390 ;
        RECT 67.995 200.345 68.285 200.390 ;
        RECT 69.885 200.345 70.175 200.390 ;
        RECT 58.795 200.190 59.085 200.235 ;
        RECT 58.795 200.050 64.070 200.190 ;
        RECT 58.795 200.005 59.085 200.050 ;
        RECT 56.955 199.850 57.245 199.895 ;
        RECT 58.320 199.850 58.640 199.910 ;
        RECT 56.955 199.710 58.640 199.850 ;
        RECT 56.955 199.665 57.245 199.710 ;
        RECT 58.320 199.650 58.640 199.710 ;
        RECT 61.095 199.850 61.385 199.895 ;
        RECT 63.930 199.870 64.070 200.050 ;
        RECT 61.095 199.710 62.230 199.850 ;
        RECT 61.095 199.665 61.385 199.710 ;
        RECT 56.480 198.970 56.800 199.230 ;
        RECT 60.160 198.970 60.480 199.230 ;
        RECT 62.090 199.215 62.230 199.710 ;
        RECT 63.795 199.555 64.085 199.870 ;
        RECT 64.875 199.850 65.165 199.895 ;
        RECT 68.455 199.850 68.745 199.895 ;
        RECT 70.290 199.850 70.580 199.895 ;
        RECT 64.875 199.710 70.580 199.850 ;
        RECT 64.875 199.665 65.165 199.710 ;
        RECT 68.455 199.665 68.745 199.710 ;
        RECT 70.290 199.665 70.580 199.710 ;
        RECT 70.740 199.650 71.060 199.910 ;
        RECT 71.660 199.850 71.980 199.910 ;
        RECT 73.055 199.850 73.345 199.895 ;
        RECT 71.660 199.710 73.345 199.850 ;
        RECT 71.660 199.650 71.980 199.710 ;
        RECT 73.055 199.665 73.345 199.710 ;
        RECT 74.435 199.665 74.725 199.895 ;
        RECT 63.495 199.510 64.085 199.555 ;
        RECT 66.735 199.510 67.385 199.555 ;
        RECT 63.495 199.370 67.385 199.510 ;
        RECT 63.495 199.325 63.785 199.370 ;
        RECT 66.735 199.325 67.385 199.370 ;
        RECT 69.360 199.310 69.680 199.570 ;
        RECT 74.510 199.510 74.650 199.665 ;
        RECT 70.830 199.370 74.650 199.510 ;
        RECT 62.015 199.170 62.305 199.215 ;
        RECT 64.760 199.170 65.080 199.230 ;
        RECT 62.015 199.030 65.080 199.170 ;
        RECT 62.015 198.985 62.305 199.030 ;
        RECT 64.760 198.970 65.080 199.030 ;
        RECT 70.280 199.170 70.600 199.230 ;
        RECT 70.830 199.170 70.970 199.370 ;
        RECT 70.280 199.030 70.970 199.170 ;
        RECT 70.280 198.970 70.600 199.030 ;
        RECT 73.500 198.970 73.820 199.230 ;
        RECT 74.895 199.170 75.185 199.215 ;
        RECT 82.240 199.170 82.560 199.230 ;
        RECT 74.895 199.030 82.560 199.170 ;
        RECT 74.895 198.985 75.185 199.030 ;
        RECT 82.240 198.970 82.560 199.030 ;
        RECT 11.330 198.350 113.450 198.830 ;
        RECT 64.315 198.150 64.605 198.195 ;
        RECT 64.760 198.150 65.080 198.210 ;
        RECT 64.315 198.010 65.080 198.150 ;
        RECT 64.315 197.965 64.605 198.010 ;
        RECT 64.760 197.950 65.080 198.010 ;
        RECT 69.360 198.150 69.680 198.210 ;
        RECT 70.295 198.150 70.585 198.195 ;
        RECT 69.360 198.010 70.585 198.150 ;
        RECT 69.360 197.950 69.680 198.010 ;
        RECT 70.295 197.965 70.585 198.010 ;
        RECT 55.095 197.810 55.745 197.855 ;
        RECT 56.480 197.810 56.800 197.870 ;
        RECT 58.695 197.810 58.985 197.855 ;
        RECT 55.095 197.670 58.985 197.810 ;
        RECT 55.095 197.625 55.745 197.670 ;
        RECT 56.480 197.610 56.800 197.670 ;
        RECT 58.395 197.625 58.985 197.670 ;
        RECT 59.240 197.810 59.560 197.870 ;
        RECT 73.500 197.810 73.820 197.870 ;
        RECT 76.375 197.810 76.665 197.855 ;
        RECT 79.615 197.810 80.265 197.855 ;
        RECT 59.240 197.670 70.740 197.810 ;
        RECT 51.900 197.470 52.190 197.515 ;
        RECT 53.735 197.470 54.025 197.515 ;
        RECT 57.315 197.470 57.605 197.515 ;
        RECT 51.900 197.330 57.605 197.470 ;
        RECT 51.900 197.285 52.190 197.330 ;
        RECT 53.735 197.285 54.025 197.330 ;
        RECT 57.315 197.285 57.605 197.330 ;
        RECT 58.395 197.310 58.685 197.625 ;
        RECT 59.240 197.610 59.560 197.670 ;
        RECT 61.555 197.470 61.845 197.515 ;
        RECT 66.140 197.470 66.460 197.530 ;
        RECT 68.455 197.470 68.745 197.515 ;
        RECT 61.555 197.330 65.450 197.470 ;
        RECT 61.555 197.285 61.845 197.330 ;
        RECT 65.310 197.190 65.450 197.330 ;
        RECT 66.140 197.330 68.745 197.470 ;
        RECT 70.600 197.470 70.740 197.670 ;
        RECT 73.500 197.670 80.265 197.810 ;
        RECT 73.500 197.610 73.820 197.670 ;
        RECT 76.375 197.625 76.965 197.670 ;
        RECT 79.615 197.625 80.265 197.670 ;
        RECT 71.660 197.470 71.980 197.530 ;
        RECT 70.600 197.330 71.980 197.470 ;
        RECT 66.140 197.270 66.460 197.330 ;
        RECT 68.455 197.285 68.745 197.330 ;
        RECT 71.660 197.270 71.980 197.330 ;
        RECT 73.055 197.285 73.345 197.515 ;
        RECT 76.675 197.310 76.965 197.625 ;
        RECT 82.240 197.610 82.560 197.870 ;
        RECT 77.755 197.470 78.045 197.515 ;
        RECT 81.335 197.470 81.625 197.515 ;
        RECT 83.170 197.470 83.460 197.515 ;
        RECT 77.755 197.330 83.460 197.470 ;
        RECT 77.755 197.285 78.045 197.330 ;
        RECT 81.335 197.285 81.625 197.330 ;
        RECT 83.170 197.285 83.460 197.330 ;
        RECT 50.040 197.130 50.360 197.190 ;
        RECT 51.435 197.130 51.725 197.175 ;
        RECT 50.040 196.990 51.725 197.130 ;
        RECT 50.040 196.930 50.360 196.990 ;
        RECT 51.435 196.945 51.725 196.990 ;
        RECT 52.800 196.930 53.120 197.190 ;
        RECT 63.380 197.175 63.700 197.190 ;
        RECT 63.270 196.945 63.700 197.175 ;
        RECT 63.855 196.945 64.145 197.175 ;
        RECT 65.220 197.130 65.540 197.190 ;
        RECT 65.695 197.130 65.985 197.175 ;
        RECT 65.220 196.990 65.985 197.130 ;
        RECT 63.380 196.930 63.700 196.945 ;
        RECT 52.305 196.790 52.595 196.835 ;
        RECT 54.195 196.790 54.485 196.835 ;
        RECT 57.315 196.790 57.605 196.835 ;
        RECT 52.305 196.650 57.605 196.790 ;
        RECT 63.930 196.790 64.070 196.945 ;
        RECT 65.220 196.930 65.540 196.990 ;
        RECT 65.695 196.945 65.985 196.990 ;
        RECT 67.520 197.130 67.840 197.190 ;
        RECT 67.995 197.130 68.285 197.175 ;
        RECT 67.520 196.990 68.285 197.130 ;
        RECT 67.520 196.930 67.840 196.990 ;
        RECT 67.995 196.945 68.285 196.990 ;
        RECT 69.360 197.130 69.680 197.190 ;
        RECT 73.130 197.130 73.270 197.285 ;
        RECT 98.800 197.270 99.120 197.530 ;
        RECT 69.360 196.990 73.270 197.130 ;
        RECT 83.635 197.130 83.925 197.175 ;
        RECT 84.540 197.130 84.860 197.190 ;
        RECT 83.635 196.990 84.860 197.130 ;
        RECT 69.360 196.930 69.680 196.990 ;
        RECT 83.635 196.945 83.925 196.990 ;
        RECT 84.540 196.930 84.860 196.990 ;
        RECT 77.755 196.790 78.045 196.835 ;
        RECT 80.875 196.790 81.165 196.835 ;
        RECT 82.765 196.790 83.055 196.835 ;
        RECT 63.930 196.650 75.110 196.790 ;
        RECT 52.305 196.605 52.595 196.650 ;
        RECT 54.195 196.605 54.485 196.650 ;
        RECT 57.315 196.605 57.605 196.650 ;
        RECT 74.970 196.510 75.110 196.650 ;
        RECT 77.755 196.650 83.055 196.790 ;
        RECT 77.755 196.605 78.045 196.650 ;
        RECT 80.875 196.605 81.165 196.650 ;
        RECT 82.765 196.605 83.055 196.650 ;
        RECT 61.080 196.450 61.400 196.510 ;
        RECT 62.475 196.450 62.765 196.495 ;
        RECT 61.080 196.310 62.765 196.450 ;
        RECT 61.080 196.250 61.400 196.310 ;
        RECT 62.475 196.265 62.765 196.310 ;
        RECT 72.120 196.250 72.440 196.510 ;
        RECT 73.960 196.250 74.280 196.510 ;
        RECT 74.880 196.250 75.200 196.510 ;
        RECT 99.720 196.250 100.040 196.510 ;
        RECT 11.330 195.630 113.450 196.110 ;
        RECT 52.800 195.430 53.120 195.490 ;
        RECT 56.955 195.430 57.245 195.475 ;
        RECT 52.800 195.290 57.245 195.430 ;
        RECT 52.800 195.230 53.120 195.290 ;
        RECT 56.955 195.245 57.245 195.290 ;
        RECT 62.000 195.430 62.320 195.490 ;
        RECT 68.440 195.430 68.760 195.490 ;
        RECT 62.000 195.290 68.760 195.430 ;
        RECT 62.000 195.230 62.320 195.290 ;
        RECT 68.440 195.230 68.760 195.290 ;
        RECT 70.740 195.430 71.060 195.490 ;
        RECT 84.540 195.430 84.860 195.490 ;
        RECT 70.740 195.290 84.860 195.430 ;
        RECT 70.740 195.230 71.060 195.290 ;
        RECT 64.315 195.090 64.605 195.135 ;
        RECT 64.760 195.090 65.080 195.150 ;
        RECT 66.140 195.090 66.460 195.150 ;
        RECT 69.835 195.090 70.125 195.135 ;
        RECT 60.250 194.950 66.460 195.090 ;
        RECT 60.250 194.810 60.390 194.950 ;
        RECT 64.315 194.905 64.605 194.950 ;
        RECT 64.760 194.890 65.080 194.950 ;
        RECT 66.140 194.890 66.460 194.950 ;
        RECT 66.690 194.950 70.125 195.090 ;
        RECT 59.700 194.550 60.020 194.810 ;
        RECT 60.160 194.550 60.480 194.810 ;
        RECT 63.380 194.750 63.700 194.810 ;
        RECT 66.690 194.795 66.830 194.950 ;
        RECT 69.835 194.905 70.125 194.950 ;
        RECT 72.695 195.090 72.985 195.135 ;
        RECT 75.815 195.090 76.105 195.135 ;
        RECT 77.705 195.090 77.995 195.135 ;
        RECT 72.695 194.950 77.995 195.090 ;
        RECT 72.695 194.905 72.985 194.950 ;
        RECT 75.815 194.905 76.105 194.950 ;
        RECT 77.705 194.905 77.995 194.950 ;
        RECT 66.615 194.750 66.905 194.795 ;
        RECT 63.010 194.610 66.905 194.750 ;
        RECT 57.860 194.210 58.180 194.470 ;
        RECT 58.795 194.225 59.085 194.455 ;
        RECT 59.255 194.410 59.545 194.455 ;
        RECT 62.000 194.410 62.320 194.470 ;
        RECT 63.010 194.455 63.150 194.610 ;
        RECT 63.380 194.550 63.700 194.610 ;
        RECT 66.615 194.565 66.905 194.610 ;
        RECT 67.980 194.550 68.300 194.810 ;
        RECT 73.960 194.750 74.280 194.810 ;
        RECT 78.650 194.795 78.790 195.290 ;
        RECT 84.540 195.230 84.860 195.290 ;
        RECT 96.500 195.430 96.820 195.490 ;
        RECT 96.500 195.290 103.170 195.430 ;
        RECT 96.500 195.230 96.820 195.290 ;
        RECT 97.075 195.090 97.365 195.135 ;
        RECT 100.195 195.090 100.485 195.135 ;
        RECT 102.085 195.090 102.375 195.135 ;
        RECT 97.075 194.950 102.375 195.090 ;
        RECT 97.075 194.905 97.365 194.950 ;
        RECT 100.195 194.905 100.485 194.950 ;
        RECT 102.085 194.905 102.375 194.950 ;
        RECT 77.195 194.750 77.485 194.795 ;
        RECT 73.960 194.610 77.485 194.750 ;
        RECT 73.960 194.550 74.280 194.610 ;
        RECT 77.195 194.565 77.485 194.610 ;
        RECT 78.575 194.565 78.865 194.795 ;
        RECT 99.720 194.750 100.040 194.810 ;
        RECT 103.030 194.795 103.170 195.290 ;
        RECT 101.575 194.750 101.865 194.795 ;
        RECT 99.720 194.610 101.865 194.750 ;
        RECT 99.720 194.550 100.040 194.610 ;
        RECT 101.575 194.565 101.865 194.610 ;
        RECT 102.955 194.750 103.245 194.795 ;
        RECT 102.955 194.610 105.240 194.750 ;
        RECT 102.955 194.565 103.245 194.610 ;
        RECT 59.255 194.270 62.320 194.410 ;
        RECT 59.255 194.225 59.545 194.270 ;
        RECT 58.870 194.070 59.010 194.225 ;
        RECT 62.000 194.210 62.320 194.270 ;
        RECT 62.935 194.225 63.225 194.455 ;
        RECT 67.075 194.410 67.365 194.455 ;
        RECT 67.075 194.270 68.210 194.410 ;
        RECT 67.075 194.225 67.365 194.270 ;
        RECT 64.315 194.070 64.605 194.115 ;
        RECT 65.220 194.070 65.540 194.130 ;
        RECT 58.870 193.930 65.540 194.070 ;
        RECT 68.070 194.070 68.210 194.270 ;
        RECT 68.440 194.210 68.760 194.470 ;
        RECT 69.375 194.410 69.665 194.455 ;
        RECT 70.280 194.410 70.600 194.470 ;
        RECT 69.375 194.270 70.600 194.410 ;
        RECT 69.375 194.225 69.665 194.270 ;
        RECT 70.280 194.210 70.600 194.270 ;
        RECT 70.740 194.070 71.060 194.130 ;
        RECT 71.615 194.115 71.905 194.430 ;
        RECT 72.695 194.410 72.985 194.455 ;
        RECT 76.275 194.410 76.565 194.455 ;
        RECT 78.110 194.410 78.400 194.455 ;
        RECT 72.695 194.270 78.400 194.410 ;
        RECT 72.695 194.225 72.985 194.270 ;
        RECT 76.275 194.225 76.565 194.270 ;
        RECT 78.110 194.225 78.400 194.270 ;
        RECT 90.060 194.210 90.380 194.470 ;
        RECT 68.070 193.930 71.060 194.070 ;
        RECT 64.315 193.885 64.605 193.930 ;
        RECT 65.220 193.870 65.540 193.930 ;
        RECT 70.740 193.870 71.060 193.930 ;
        RECT 71.315 194.070 71.905 194.115 ;
        RECT 72.120 194.070 72.440 194.130 ;
        RECT 74.555 194.070 75.205 194.115 ;
        RECT 71.315 193.930 75.205 194.070 ;
        RECT 71.315 193.885 71.605 193.930 ;
        RECT 72.120 193.870 72.440 193.930 ;
        RECT 74.555 193.885 75.205 193.930 ;
        RECT 94.660 194.070 94.980 194.130 ;
        RECT 95.995 194.115 96.285 194.430 ;
        RECT 97.075 194.410 97.365 194.455 ;
        RECT 100.655 194.410 100.945 194.455 ;
        RECT 102.490 194.410 102.780 194.455 ;
        RECT 97.075 194.270 102.780 194.410 ;
        RECT 97.075 194.225 97.365 194.270 ;
        RECT 100.655 194.225 100.945 194.270 ;
        RECT 102.490 194.225 102.780 194.270 ;
        RECT 95.695 194.070 96.285 194.115 ;
        RECT 98.935 194.070 99.585 194.115 ;
        RECT 94.660 193.930 99.585 194.070 ;
        RECT 105.100 194.070 105.240 194.610 ;
        RECT 109.380 194.070 109.700 194.130 ;
        RECT 105.100 193.930 109.700 194.070 ;
        RECT 94.660 193.870 94.980 193.930 ;
        RECT 95.695 193.885 95.985 193.930 ;
        RECT 98.935 193.885 99.585 193.930 ;
        RECT 109.380 193.870 109.700 193.930 ;
        RECT 61.095 193.730 61.385 193.775 ;
        RECT 62.000 193.730 62.320 193.790 ;
        RECT 61.095 193.590 62.320 193.730 ;
        RECT 61.095 193.545 61.385 193.590 ;
        RECT 62.000 193.530 62.320 193.590 ;
        RECT 67.520 193.730 67.840 193.790 ;
        RECT 68.455 193.730 68.745 193.775 ;
        RECT 67.520 193.590 68.745 193.730 ;
        RECT 67.520 193.530 67.840 193.590 ;
        RECT 68.455 193.545 68.745 193.590 ;
        RECT 90.980 193.530 91.300 193.790 ;
        RECT 94.215 193.730 94.505 193.775 ;
        RECT 96.960 193.730 97.280 193.790 ;
        RECT 94.215 193.590 97.280 193.730 ;
        RECT 94.215 193.545 94.505 193.590 ;
        RECT 96.960 193.530 97.280 193.590 ;
        RECT 11.330 192.910 113.450 193.390 ;
        RECT 57.860 192.710 58.180 192.770 ;
        RECT 62.000 192.755 62.320 192.770 ;
        RECT 61.095 192.710 61.385 192.755 ;
        RECT 57.860 192.570 61.385 192.710 ;
        RECT 57.860 192.510 58.180 192.570 ;
        RECT 61.095 192.525 61.385 192.570 ;
        RECT 61.935 192.525 62.320 192.755 ;
        RECT 70.280 192.710 70.600 192.770 ;
        RECT 71.215 192.710 71.505 192.755 ;
        RECT 62.000 192.510 62.320 192.525 ;
        RECT 69.910 192.570 71.505 192.710 ;
        RECT 34.860 192.415 35.180 192.430 ;
        RECT 31.755 192.370 32.045 192.415 ;
        RECT 34.860 192.370 35.645 192.415 ;
        RECT 31.755 192.230 35.645 192.370 ;
        RECT 31.755 192.185 32.345 192.230 ;
        RECT 32.055 191.870 32.345 192.185 ;
        RECT 34.860 192.185 35.645 192.230 ;
        RECT 40.380 192.370 40.700 192.430 ;
        RECT 40.955 192.370 41.245 192.415 ;
        RECT 44.195 192.370 44.845 192.415 ;
        RECT 40.380 192.230 44.845 192.370 ;
        RECT 34.860 192.170 35.180 192.185 ;
        RECT 40.380 192.170 40.700 192.230 ;
        RECT 40.955 192.185 41.545 192.230 ;
        RECT 44.195 192.185 44.845 192.230 ;
        RECT 62.935 192.370 63.225 192.415 ;
        RECT 68.440 192.370 68.760 192.430 ;
        RECT 69.910 192.415 70.050 192.570 ;
        RECT 70.280 192.510 70.600 192.570 ;
        RECT 71.215 192.525 71.505 192.570 ;
        RECT 68.915 192.370 69.205 192.415 ;
        RECT 62.935 192.230 66.370 192.370 ;
        RECT 62.935 192.185 63.225 192.230 ;
        RECT 33.135 192.030 33.425 192.075 ;
        RECT 36.715 192.030 37.005 192.075 ;
        RECT 38.550 192.030 38.840 192.075 ;
        RECT 33.135 191.890 38.840 192.030 ;
        RECT 33.135 191.845 33.425 191.890 ;
        RECT 36.715 191.845 37.005 191.890 ;
        RECT 38.550 191.845 38.840 191.890 ;
        RECT 41.255 191.870 41.545 192.185 ;
        RECT 42.335 192.030 42.625 192.075 ;
        RECT 45.915 192.030 46.205 192.075 ;
        RECT 47.750 192.030 48.040 192.075 ;
        RECT 42.335 191.890 48.040 192.030 ;
        RECT 42.335 191.845 42.625 191.890 ;
        RECT 45.915 191.845 46.205 191.890 ;
        RECT 47.750 191.845 48.040 191.890 ;
        RECT 57.415 192.030 57.705 192.075 ;
        RECT 58.320 192.030 58.640 192.090 ;
        RECT 57.415 191.890 58.640 192.030 ;
        RECT 57.415 191.845 57.705 191.890 ;
        RECT 58.320 191.830 58.640 191.890 ;
        RECT 63.395 192.030 63.685 192.075 ;
        RECT 65.220 192.030 65.540 192.090 ;
        RECT 63.395 191.890 65.540 192.030 ;
        RECT 63.395 191.845 63.685 191.890 ;
        RECT 65.220 191.830 65.540 191.890 ;
        RECT 37.620 191.490 37.940 191.750 ;
        RECT 39.015 191.690 39.305 191.735 ;
        RECT 48.215 191.690 48.505 191.735 ;
        RECT 50.040 191.690 50.360 191.750 ;
        RECT 39.015 191.550 50.360 191.690 ;
        RECT 39.015 191.505 39.305 191.550 ;
        RECT 48.215 191.505 48.505 191.550 ;
        RECT 50.040 191.490 50.360 191.550 ;
        RECT 64.760 191.490 65.080 191.750 ;
        RECT 33.135 191.350 33.425 191.395 ;
        RECT 36.255 191.350 36.545 191.395 ;
        RECT 38.145 191.350 38.435 191.395 ;
        RECT 33.135 191.210 38.435 191.350 ;
        RECT 33.135 191.165 33.425 191.210 ;
        RECT 36.255 191.165 36.545 191.210 ;
        RECT 38.145 191.165 38.435 191.210 ;
        RECT 42.335 191.350 42.625 191.395 ;
        RECT 45.455 191.350 45.745 191.395 ;
        RECT 47.345 191.350 47.635 191.395 ;
        RECT 42.335 191.210 47.635 191.350 ;
        RECT 42.335 191.165 42.625 191.210 ;
        RECT 45.455 191.165 45.745 191.210 ;
        RECT 47.345 191.165 47.635 191.210 ;
        RECT 66.230 191.070 66.370 192.230 ;
        RECT 68.440 192.230 69.205 192.370 ;
        RECT 68.440 192.170 68.760 192.230 ;
        RECT 68.915 192.185 69.205 192.230 ;
        RECT 69.835 192.185 70.125 192.415 ;
        RECT 70.740 192.370 71.060 192.430 ;
        RECT 74.880 192.370 75.200 192.430 ;
        RECT 70.740 192.230 75.200 192.370 ;
        RECT 70.740 192.170 71.060 192.230 ;
        RECT 74.880 192.170 75.200 192.230 ;
        RECT 84.095 192.370 84.385 192.415 ;
        RECT 86.495 192.370 86.785 192.415 ;
        RECT 89.735 192.370 90.385 192.415 ;
        RECT 84.095 192.230 90.385 192.370 ;
        RECT 84.095 192.185 84.385 192.230 ;
        RECT 86.495 192.185 87.085 192.230 ;
        RECT 89.735 192.185 90.385 192.230 ;
        RECT 90.980 192.370 91.300 192.430 ;
        RECT 92.375 192.370 92.665 192.415 ;
        RECT 90.980 192.230 92.665 192.370 ;
        RECT 79.480 192.030 79.800 192.090 ;
        RECT 80.415 192.030 80.705 192.075 ;
        RECT 79.480 191.890 80.705 192.030 ;
        RECT 79.480 191.830 79.800 191.890 ;
        RECT 80.415 191.845 80.705 191.890 ;
        RECT 83.635 191.845 83.925 192.075 ;
        RECT 86.795 191.870 87.085 192.185 ;
        RECT 90.980 192.170 91.300 192.230 ;
        RECT 92.375 192.185 92.665 192.230 ;
        RECT 98.355 192.370 98.645 192.415 ;
        RECT 102.135 192.370 102.425 192.415 ;
        RECT 105.375 192.370 106.025 192.415 ;
        RECT 98.355 192.230 106.025 192.370 ;
        RECT 98.355 192.185 98.645 192.230 ;
        RECT 102.135 192.185 102.725 192.230 ;
        RECT 105.375 192.185 106.025 192.230 ;
        RECT 87.875 192.030 88.165 192.075 ;
        RECT 91.455 192.030 91.745 192.075 ;
        RECT 93.290 192.030 93.580 192.075 ;
        RECT 87.875 191.890 93.580 192.030 ;
        RECT 87.875 191.845 88.165 191.890 ;
        RECT 91.455 191.845 91.745 191.890 ;
        RECT 93.290 191.845 93.580 191.890 ;
        RECT 94.675 192.030 94.965 192.075 ;
        RECT 96.960 192.030 97.280 192.090 ;
        RECT 94.675 191.890 97.280 192.030 ;
        RECT 94.675 191.845 94.965 191.890 ;
        RECT 71.660 191.690 71.980 191.750 ;
        RECT 83.710 191.690 83.850 191.845 ;
        RECT 96.960 191.830 97.280 191.890 ;
        RECT 97.895 192.030 98.185 192.075 ;
        RECT 97.895 191.890 98.570 192.030 ;
        RECT 97.895 191.845 98.185 191.890 ;
        RECT 98.430 191.750 98.570 191.890 ;
        RECT 102.435 191.870 102.725 192.185 ;
        RECT 103.515 192.030 103.805 192.075 ;
        RECT 107.095 192.030 107.385 192.075 ;
        RECT 108.930 192.030 109.220 192.075 ;
        RECT 103.515 191.890 109.220 192.030 ;
        RECT 103.515 191.845 103.805 191.890 ;
        RECT 107.095 191.845 107.385 191.890 ;
        RECT 108.930 191.845 109.220 191.890 ;
        RECT 109.380 192.030 109.700 192.090 ;
        RECT 110.760 192.030 111.080 192.090 ;
        RECT 109.380 191.890 111.080 192.030 ;
        RECT 109.380 191.830 109.700 191.890 ;
        RECT 110.760 191.830 111.080 191.890 ;
        RECT 88.680 191.690 89.000 191.750 ;
        RECT 71.660 191.550 89.000 191.690 ;
        RECT 71.660 191.490 71.980 191.550 ;
        RECT 88.680 191.490 89.000 191.550 ;
        RECT 93.755 191.690 94.045 191.735 ;
        RECT 96.500 191.690 96.820 191.750 ;
        RECT 93.755 191.550 96.820 191.690 ;
        RECT 93.755 191.505 94.045 191.550 ;
        RECT 96.500 191.490 96.820 191.550 ;
        RECT 98.340 191.490 98.660 191.750 ;
        RECT 104.780 191.690 105.100 191.750 ;
        RECT 108.015 191.690 108.305 191.735 ;
        RECT 104.780 191.550 108.305 191.690 ;
        RECT 104.780 191.490 105.100 191.550 ;
        RECT 108.015 191.505 108.305 191.550 ;
        RECT 87.875 191.350 88.165 191.395 ;
        RECT 90.995 191.350 91.285 191.395 ;
        RECT 92.885 191.350 93.175 191.395 ;
        RECT 87.875 191.210 93.175 191.350 ;
        RECT 87.875 191.165 88.165 191.210 ;
        RECT 90.995 191.165 91.285 191.210 ;
        RECT 92.885 191.165 93.175 191.210 ;
        RECT 103.515 191.350 103.805 191.395 ;
        RECT 106.635 191.350 106.925 191.395 ;
        RECT 108.525 191.350 108.815 191.395 ;
        RECT 103.515 191.210 108.815 191.350 ;
        RECT 103.515 191.165 103.805 191.210 ;
        RECT 106.635 191.165 106.925 191.210 ;
        RECT 108.525 191.165 108.815 191.210 ;
        RECT 30.260 190.810 30.580 191.070 ;
        RECT 39.460 190.810 39.780 191.070 ;
        RECT 44.060 191.010 44.380 191.070 ;
        RECT 46.900 191.010 47.190 191.055 ;
        RECT 44.060 190.870 47.190 191.010 ;
        RECT 44.060 190.810 44.380 190.870 ;
        RECT 46.900 190.825 47.190 190.870 ;
        RECT 56.940 190.810 57.260 191.070 ;
        RECT 62.000 190.810 62.320 191.070 ;
        RECT 64.300 190.810 64.620 191.070 ;
        RECT 66.140 190.810 66.460 191.070 ;
        RECT 67.980 190.810 68.300 191.070 ;
        RECT 81.320 190.810 81.640 191.070 ;
        RECT 85.000 190.810 85.320 191.070 ;
        RECT 97.420 190.810 97.740 191.070 ;
        RECT 99.260 191.010 99.580 191.070 ;
        RECT 100.655 191.010 100.945 191.055 ;
        RECT 99.260 190.870 100.945 191.010 ;
        RECT 99.260 190.810 99.580 190.870 ;
        RECT 100.655 190.825 100.945 190.870 ;
        RECT 11.330 190.190 113.450 190.670 ;
        RECT 38.555 189.990 38.845 190.035 ;
        RECT 40.380 189.990 40.700 190.050 ;
        RECT 38.555 189.850 40.700 189.990 ;
        RECT 38.555 189.805 38.845 189.850 ;
        RECT 40.380 189.790 40.700 189.850 ;
        RECT 44.060 189.790 44.380 190.050 ;
        RECT 61.540 189.990 61.860 190.050 ;
        RECT 62.475 189.990 62.765 190.035 ;
        RECT 61.540 189.850 62.765 189.990 ;
        RECT 61.540 189.790 61.860 189.850 ;
        RECT 62.475 189.805 62.765 189.850 ;
        RECT 64.760 189.790 65.080 190.050 ;
        RECT 67.980 189.990 68.300 190.050 ;
        RECT 68.455 189.990 68.745 190.035 ;
        RECT 67.980 189.850 68.745 189.990 ;
        RECT 67.980 189.790 68.300 189.850 ;
        RECT 68.455 189.805 68.745 189.850 ;
        RECT 69.360 189.790 69.680 190.050 ;
        RECT 90.060 189.990 90.380 190.050 ;
        RECT 91.455 189.990 91.745 190.035 ;
        RECT 90.060 189.850 91.745 189.990 ;
        RECT 90.060 189.790 90.380 189.850 ;
        RECT 91.455 189.805 91.745 189.850 ;
        RECT 94.215 189.990 94.505 190.035 ;
        RECT 94.660 189.990 94.980 190.050 ;
        RECT 94.215 189.850 94.980 189.990 ;
        RECT 94.215 189.805 94.505 189.850 ;
        RECT 94.660 189.790 94.980 189.850 ;
        RECT 98.800 189.790 99.120 190.050 ;
        RECT 104.780 189.790 105.100 190.050 ;
        RECT 23.325 189.650 23.615 189.695 ;
        RECT 25.215 189.650 25.505 189.695 ;
        RECT 28.335 189.650 28.625 189.695 ;
        RECT 23.325 189.510 28.625 189.650 ;
        RECT 23.325 189.465 23.615 189.510 ;
        RECT 25.215 189.465 25.505 189.510 ;
        RECT 28.335 189.465 28.625 189.510 ;
        RECT 30.720 189.650 31.040 189.710 ;
        RECT 42.220 189.650 42.540 189.710 ;
        RECT 30.720 189.510 42.540 189.650 ;
        RECT 30.720 189.450 31.040 189.510 ;
        RECT 31.180 189.110 31.500 189.370 ;
        RECT 32.100 189.110 32.420 189.370 ;
        RECT 33.110 189.355 33.250 189.510 ;
        RECT 42.220 189.450 42.540 189.510 ;
        RECT 47.395 189.650 47.685 189.695 ;
        RECT 50.515 189.650 50.805 189.695 ;
        RECT 52.405 189.650 52.695 189.695 ;
        RECT 62.000 189.650 62.320 189.710 ;
        RECT 65.695 189.650 65.985 189.695 ;
        RECT 47.395 189.510 52.695 189.650 ;
        RECT 47.395 189.465 47.685 189.510 ;
        RECT 50.515 189.465 50.805 189.510 ;
        RECT 52.405 189.465 52.695 189.510 ;
        RECT 56.570 189.510 65.985 189.650 ;
        RECT 33.035 189.125 33.325 189.355 ;
        RECT 36.240 189.310 36.560 189.370 ;
        RECT 39.460 189.310 39.780 189.370 ;
        RECT 56.570 189.355 56.710 189.510 ;
        RECT 62.000 189.450 62.320 189.510 ;
        RECT 65.695 189.465 65.985 189.510 ;
        RECT 79.450 189.650 79.740 189.695 ;
        RECT 82.230 189.650 82.520 189.695 ;
        RECT 84.090 189.650 84.380 189.695 ;
        RECT 79.450 189.510 84.380 189.650 ;
        RECT 79.450 189.465 79.740 189.510 ;
        RECT 82.230 189.465 82.520 189.510 ;
        RECT 84.090 189.465 84.380 189.510 ;
        RECT 36.240 189.170 39.780 189.310 ;
        RECT 36.240 189.110 36.560 189.170 ;
        RECT 39.460 189.110 39.780 189.170 ;
        RECT 56.495 189.125 56.785 189.355 ;
        RECT 59.700 189.310 60.020 189.370 ;
        RECT 63.395 189.310 63.685 189.355 ;
        RECT 67.075 189.310 67.365 189.355 ;
        RECT 68.440 189.310 68.760 189.370 ;
        RECT 59.700 189.170 62.230 189.310 ;
        RECT 59.700 189.110 60.020 189.170 ;
        RECT 20.600 188.970 20.920 189.030 ;
        RECT 22.455 188.970 22.745 189.015 ;
        RECT 20.600 188.830 22.745 188.970 ;
        RECT 20.600 188.770 20.920 188.830 ;
        RECT 22.455 188.785 22.745 188.830 ;
        RECT 22.920 188.970 23.210 189.015 ;
        RECT 24.755 188.970 25.045 189.015 ;
        RECT 28.335 188.970 28.625 189.015 ;
        RECT 22.920 188.830 28.625 188.970 ;
        RECT 22.920 188.785 23.210 188.830 ;
        RECT 24.755 188.785 25.045 188.830 ;
        RECT 28.335 188.785 28.625 188.830 ;
        RECT 23.820 188.430 24.140 188.690 ;
        RECT 24.280 188.630 24.600 188.690 ;
        RECT 29.415 188.675 29.705 188.990 ;
        RECT 39.015 188.785 39.305 189.015 ;
        RECT 26.115 188.630 26.765 188.675 ;
        RECT 29.415 188.630 30.005 188.675 ;
        RECT 24.280 188.490 30.005 188.630 ;
        RECT 39.090 188.630 39.230 188.785 ;
        RECT 43.140 188.770 43.460 189.030 ;
        RECT 44.060 188.630 44.380 188.690 ;
        RECT 39.090 188.490 44.380 188.630 ;
        RECT 24.280 188.430 24.600 188.490 ;
        RECT 26.115 188.445 26.765 188.490 ;
        RECT 29.715 188.445 30.005 188.490 ;
        RECT 44.060 188.430 44.380 188.490 ;
        RECT 44.980 188.630 45.300 188.690 ;
        RECT 46.315 188.675 46.605 188.990 ;
        RECT 47.395 188.970 47.685 189.015 ;
        RECT 50.975 188.970 51.265 189.015 ;
        RECT 52.810 188.970 53.100 189.015 ;
        RECT 47.395 188.830 53.100 188.970 ;
        RECT 47.395 188.785 47.685 188.830 ;
        RECT 50.975 188.785 51.265 188.830 ;
        RECT 52.810 188.785 53.100 188.830 ;
        RECT 53.260 188.770 53.580 189.030 ;
        RECT 56.035 188.970 56.325 189.015 ;
        RECT 57.415 188.970 57.705 189.015 ;
        RECT 56.035 188.830 57.705 188.970 ;
        RECT 56.035 188.785 56.325 188.830 ;
        RECT 57.415 188.785 57.705 188.830 ;
        RECT 60.635 188.970 60.925 189.015 ;
        RECT 61.540 188.970 61.860 189.030 ;
        RECT 62.090 189.015 62.230 189.170 ;
        RECT 63.395 189.170 68.760 189.310 ;
        RECT 63.395 189.125 63.685 189.170 ;
        RECT 67.075 189.125 67.365 189.170 ;
        RECT 68.440 189.110 68.760 189.170 ;
        RECT 81.320 189.310 81.640 189.370 ;
        RECT 82.715 189.310 83.005 189.355 ;
        RECT 81.320 189.170 83.005 189.310 ;
        RECT 81.320 189.110 81.640 189.170 ;
        RECT 82.715 189.125 83.005 189.170 ;
        RECT 84.540 189.110 84.860 189.370 ;
        RECT 88.235 189.310 88.525 189.355 ;
        RECT 95.595 189.310 95.885 189.355 ;
        RECT 99.735 189.310 100.025 189.355 ;
        RECT 88.235 189.170 100.025 189.310 ;
        RECT 88.235 189.125 88.525 189.170 ;
        RECT 95.595 189.125 95.885 189.170 ;
        RECT 99.735 189.125 100.025 189.170 ;
        RECT 60.635 188.830 61.860 188.970 ;
        RECT 60.635 188.785 60.925 188.830 ;
        RECT 61.540 188.770 61.860 188.830 ;
        RECT 62.015 188.785 62.305 189.015 ;
        RECT 46.015 188.630 46.605 188.675 ;
        RECT 49.255 188.630 49.905 188.675 ;
        RECT 44.980 188.490 49.905 188.630 ;
        RECT 44.980 188.430 45.300 188.490 ;
        RECT 46.015 188.445 46.305 188.490 ;
        RECT 49.255 188.445 49.905 188.490 ;
        RECT 51.880 188.430 52.200 188.690 ;
        RECT 28.420 188.290 28.740 188.350 ;
        RECT 33.495 188.290 33.785 188.335 ;
        RECT 28.420 188.150 33.785 188.290 ;
        RECT 28.420 188.090 28.740 188.150 ;
        RECT 33.495 188.105 33.785 188.150 ;
        RECT 35.335 188.290 35.625 188.335 ;
        RECT 39.000 188.290 39.320 188.350 ;
        RECT 35.335 188.150 39.320 188.290 ;
        RECT 35.335 188.105 35.625 188.150 ;
        RECT 39.000 188.090 39.320 188.150 ;
        RECT 42.680 188.090 43.000 188.350 ;
        RECT 44.535 188.290 44.825 188.335 ;
        RECT 45.440 188.290 45.760 188.350 ;
        RECT 44.535 188.150 45.760 188.290 ;
        RECT 44.535 188.105 44.825 188.150 ;
        RECT 45.440 188.090 45.760 188.150 ;
        RECT 54.180 188.090 54.500 188.350 ;
        RECT 62.090 188.290 62.230 188.785 ;
        RECT 65.220 188.770 65.540 189.030 ;
        RECT 66.140 188.970 66.460 189.030 ;
        RECT 79.450 188.970 79.740 189.015 ;
        RECT 84.080 188.970 84.400 189.030 ;
        RECT 88.310 188.970 88.450 189.125 ;
        RECT 66.140 188.830 68.210 188.970 ;
        RECT 66.140 188.770 66.460 188.830 ;
        RECT 64.300 188.630 64.620 188.690 ;
        RECT 65.695 188.630 65.985 188.675 ;
        RECT 64.300 188.490 65.985 188.630 ;
        RECT 64.300 188.430 64.620 188.490 ;
        RECT 65.695 188.445 65.985 188.490 ;
        RECT 67.520 188.430 67.840 188.690 ;
        RECT 68.070 188.630 68.210 188.830 ;
        RECT 79.450 188.830 81.985 188.970 ;
        RECT 79.450 188.785 79.740 188.830 ;
        RECT 80.860 188.675 81.180 188.690 ;
        RECT 68.535 188.630 68.825 188.675 ;
        RECT 68.070 188.490 68.825 188.630 ;
        RECT 68.535 188.445 68.825 188.490 ;
        RECT 77.590 188.630 77.880 188.675 ;
        RECT 80.850 188.630 81.180 188.675 ;
        RECT 77.590 188.490 81.180 188.630 ;
        RECT 77.590 188.445 77.880 188.490 ;
        RECT 80.850 188.445 81.180 188.490 ;
        RECT 81.770 188.675 81.985 188.830 ;
        RECT 84.080 188.830 88.450 188.970 ;
        RECT 88.680 188.970 89.000 189.030 ;
        RECT 93.755 188.970 94.045 189.015 ;
        RECT 88.680 188.830 94.045 188.970 ;
        RECT 84.080 188.770 84.400 188.830 ;
        RECT 88.680 188.770 89.000 188.830 ;
        RECT 93.755 188.785 94.045 188.830 ;
        RECT 96.515 188.970 96.805 189.015 ;
        RECT 97.420 188.970 97.740 189.030 ;
        RECT 101.115 188.970 101.405 189.015 ;
        RECT 96.515 188.830 101.405 188.970 ;
        RECT 96.515 188.785 96.805 188.830 ;
        RECT 81.770 188.630 82.060 188.675 ;
        RECT 83.630 188.630 83.920 188.675 ;
        RECT 89.615 188.630 89.905 188.675 ;
        RECT 81.770 188.490 83.920 188.630 ;
        RECT 81.770 188.445 82.060 188.490 ;
        RECT 83.630 188.445 83.920 188.490 ;
        RECT 84.170 188.490 89.905 188.630 ;
        RECT 93.830 188.630 93.970 188.785 ;
        RECT 97.420 188.770 97.740 188.830 ;
        RECT 101.115 188.785 101.405 188.830 ;
        RECT 103.875 188.970 104.165 189.015 ;
        RECT 104.320 188.970 104.640 189.030 ;
        RECT 103.875 188.830 104.640 188.970 ;
        RECT 103.875 188.785 104.165 188.830 ;
        RECT 104.320 188.770 104.640 188.830 ;
        RECT 98.340 188.630 98.660 188.690 ;
        RECT 93.830 188.490 98.660 188.630 ;
        RECT 80.860 188.430 81.180 188.445 ;
        RECT 66.140 188.290 66.460 188.350 ;
        RECT 70.280 188.290 70.600 188.350 ;
        RECT 62.090 188.150 70.600 188.290 ;
        RECT 66.140 188.090 66.460 188.150 ;
        RECT 70.280 188.090 70.600 188.150 ;
        RECT 75.585 188.290 75.875 188.335 ;
        RECT 79.940 188.290 80.260 188.350 ;
        RECT 84.170 188.290 84.310 188.490 ;
        RECT 89.615 188.445 89.905 188.490 ;
        RECT 98.340 188.430 98.660 188.490 ;
        RECT 75.585 188.150 84.310 188.290 ;
        RECT 89.155 188.290 89.445 188.335 ;
        RECT 90.520 188.290 90.840 188.350 ;
        RECT 96.975 188.290 97.265 188.335 ;
        RECT 89.155 188.150 97.265 188.290 ;
        RECT 75.585 188.105 75.875 188.150 ;
        RECT 79.940 188.090 80.260 188.150 ;
        RECT 89.155 188.105 89.445 188.150 ;
        RECT 90.520 188.090 90.840 188.150 ;
        RECT 96.975 188.105 97.265 188.150 ;
        RECT 99.260 188.290 99.580 188.350 ;
        RECT 100.655 188.290 100.945 188.335 ;
        RECT 99.260 188.150 100.945 188.290 ;
        RECT 99.260 188.090 99.580 188.150 ;
        RECT 100.655 188.105 100.945 188.150 ;
        RECT 102.940 188.090 103.260 188.350 ;
        RECT 11.330 187.470 113.450 187.950 ;
        RECT 24.280 187.070 24.600 187.330 ;
        RECT 28.420 187.070 28.740 187.330 ;
        RECT 42.220 187.070 42.540 187.330 ;
        RECT 43.140 187.270 43.460 187.330 ;
        RECT 44.075 187.270 44.365 187.315 ;
        RECT 43.140 187.130 44.365 187.270 ;
        RECT 43.140 187.070 43.460 187.130 ;
        RECT 44.075 187.085 44.365 187.130 ;
        RECT 50.975 187.270 51.265 187.315 ;
        RECT 51.880 187.270 52.200 187.330 ;
        RECT 50.975 187.130 52.200 187.270 ;
        RECT 50.975 187.085 51.265 187.130 ;
        RECT 51.880 187.070 52.200 187.130 ;
        RECT 79.480 187.070 79.800 187.330 ;
        RECT 80.415 187.270 80.705 187.315 ;
        RECT 80.860 187.270 81.180 187.330 ;
        RECT 80.415 187.130 81.180 187.270 ;
        RECT 80.415 187.085 80.705 187.130 ;
        RECT 80.860 187.070 81.180 187.130 ;
        RECT 90.520 187.070 90.840 187.330 ;
        RECT 104.320 187.070 104.640 187.330 ;
        RECT 34.400 186.975 34.720 186.990 ;
        RECT 31.130 186.930 31.420 186.975 ;
        RECT 34.390 186.930 34.720 186.975 ;
        RECT 31.130 186.790 34.720 186.930 ;
        RECT 31.130 186.745 31.420 186.790 ;
        RECT 34.390 186.745 34.720 186.790 ;
        RECT 34.400 186.730 34.720 186.745 ;
        RECT 35.310 186.930 35.600 186.975 ;
        RECT 37.170 186.930 37.460 186.975 ;
        RECT 35.310 186.790 37.460 186.930 ;
        RECT 35.310 186.745 35.600 186.790 ;
        RECT 37.170 186.745 37.460 186.790 ;
        RECT 41.775 186.930 42.065 186.975 ;
        RECT 42.680 186.930 43.000 186.990 ;
        RECT 46.375 186.930 46.665 186.975 ;
        RECT 41.775 186.790 46.665 186.930 ;
        RECT 41.775 186.745 42.065 186.790 ;
        RECT 24.740 186.390 25.060 186.650 ;
        RECT 32.990 186.590 33.280 186.635 ;
        RECT 35.310 186.590 35.525 186.745 ;
        RECT 42.680 186.730 43.000 186.790 ;
        RECT 46.375 186.745 46.665 186.790 ;
        RECT 54.180 186.730 54.500 186.990 ;
        RECT 56.940 186.975 57.260 186.990 ;
        RECT 56.475 186.930 57.260 186.975 ;
        RECT 60.075 186.930 60.365 186.975 ;
        RECT 56.475 186.790 60.365 186.930 ;
        RECT 56.475 186.745 57.260 186.790 ;
        RECT 56.940 186.730 57.260 186.745 ;
        RECT 59.775 186.745 60.365 186.790 ;
        RECT 71.660 186.930 71.980 186.990 ;
        RECT 77.655 186.930 77.945 186.975 ;
        RECT 71.660 186.790 77.945 186.930 ;
        RECT 32.990 186.450 35.525 186.590 ;
        RECT 36.255 186.590 36.545 186.635 ;
        RECT 38.540 186.590 38.860 186.650 ;
        RECT 36.255 186.450 38.860 186.590 ;
        RECT 32.990 186.405 33.280 186.450 ;
        RECT 36.255 186.405 36.545 186.450 ;
        RECT 38.540 186.390 38.860 186.450 ;
        RECT 39.000 186.590 39.320 186.650 ;
        RECT 39.475 186.590 39.765 186.635 ;
        RECT 49.580 186.590 49.900 186.650 ;
        RECT 50.055 186.590 50.345 186.635 ;
        RECT 39.000 186.450 39.765 186.590 ;
        RECT 39.000 186.390 39.320 186.450 ;
        RECT 39.475 186.405 39.765 186.450 ;
        RECT 40.470 186.450 46.590 186.590 ;
        RECT 25.675 186.250 25.965 186.295 ;
        RECT 31.180 186.250 31.500 186.310 ;
        RECT 25.675 186.110 31.500 186.250 ;
        RECT 25.675 186.065 25.965 186.110 ;
        RECT 31.180 186.050 31.500 186.110 ;
        RECT 38.095 186.250 38.385 186.295 ;
        RECT 40.470 186.250 40.610 186.450 ;
        RECT 38.095 186.110 40.610 186.250 ;
        RECT 40.855 186.250 41.145 186.295 ;
        RECT 43.140 186.250 43.460 186.310 ;
        RECT 44.995 186.250 45.285 186.295 ;
        RECT 40.855 186.110 45.285 186.250 ;
        RECT 38.095 186.065 38.385 186.110 ;
        RECT 40.855 186.065 41.145 186.110 ;
        RECT 29.125 185.910 29.415 185.955 ;
        RECT 30.720 185.910 31.040 185.970 ;
        RECT 29.125 185.770 31.040 185.910 ;
        RECT 29.125 185.725 29.415 185.770 ;
        RECT 30.720 185.710 31.040 185.770 ;
        RECT 32.990 185.910 33.280 185.955 ;
        RECT 35.770 185.910 36.060 185.955 ;
        RECT 37.630 185.910 37.920 185.955 ;
        RECT 32.990 185.770 37.920 185.910 ;
        RECT 32.990 185.725 33.280 185.770 ;
        RECT 35.770 185.725 36.060 185.770 ;
        RECT 37.630 185.725 37.920 185.770 ;
        RECT 38.540 185.710 38.860 185.970 ;
        RECT 40.930 185.910 41.070 186.065 ;
        RECT 43.140 186.050 43.460 186.110 ;
        RECT 44.995 186.065 45.285 186.110 ;
        RECT 45.900 186.050 46.220 186.310 ;
        RECT 40.470 185.770 41.070 185.910 ;
        RECT 46.450 185.910 46.590 186.450 ;
        RECT 49.580 186.450 50.345 186.590 ;
        RECT 49.580 186.390 49.900 186.450 ;
        RECT 50.055 186.405 50.345 186.450 ;
        RECT 53.280 186.590 53.570 186.635 ;
        RECT 55.115 186.590 55.405 186.635 ;
        RECT 58.695 186.590 58.985 186.635 ;
        RECT 53.280 186.450 58.985 186.590 ;
        RECT 53.280 186.405 53.570 186.450 ;
        RECT 55.115 186.405 55.405 186.450 ;
        RECT 58.695 186.405 58.985 186.450 ;
        RECT 59.775 186.430 60.065 186.745 ;
        RECT 71.660 186.730 71.980 186.790 ;
        RECT 77.655 186.745 77.945 186.790 ;
        RECT 69.360 186.590 69.680 186.650 ;
        RECT 73.055 186.590 73.345 186.635 ;
        RECT 80.875 186.590 81.165 186.635 ;
        RECT 69.360 186.450 84.310 186.590 ;
        RECT 69.360 186.390 69.680 186.450 ;
        RECT 73.055 186.405 73.345 186.450 ;
        RECT 80.875 186.405 81.165 186.450 ;
        RECT 84.170 186.310 84.310 186.450 ;
        RECT 91.900 186.390 92.220 186.650 ;
        RECT 98.800 186.390 99.120 186.650 ;
        RECT 102.940 186.590 103.260 186.650 ;
        RECT 107.095 186.590 107.385 186.635 ;
        RECT 102.940 186.450 107.385 186.590 ;
        RECT 102.940 186.390 103.260 186.450 ;
        RECT 107.095 186.405 107.385 186.450 ;
        RECT 52.800 186.050 53.120 186.310 ;
        RECT 76.720 186.050 77.040 186.310 ;
        RECT 77.195 186.250 77.485 186.295 ;
        RECT 79.940 186.250 80.260 186.310 ;
        RECT 77.195 186.110 80.260 186.250 ;
        RECT 77.195 186.065 77.485 186.110 ;
        RECT 79.940 186.050 80.260 186.110 ;
        RECT 84.080 186.050 84.400 186.310 ;
        RECT 85.000 186.250 85.320 186.310 ;
        RECT 87.775 186.250 88.065 186.295 ;
        RECT 88.220 186.250 88.540 186.310 ;
        RECT 85.000 186.110 88.540 186.250 ;
        RECT 85.000 186.050 85.320 186.110 ;
        RECT 87.775 186.065 88.065 186.110 ;
        RECT 88.220 186.050 88.540 186.110 ;
        RECT 95.120 186.250 95.440 186.310 ;
        RECT 96.055 186.250 96.345 186.295 ;
        RECT 95.120 186.110 96.345 186.250 ;
        RECT 95.120 186.050 95.440 186.110 ;
        RECT 96.055 186.065 96.345 186.110 ;
        RECT 99.260 186.250 99.580 186.310 ;
        RECT 100.655 186.250 100.945 186.295 ;
        RECT 99.260 186.110 100.945 186.250 ;
        RECT 99.260 186.050 99.580 186.110 ;
        RECT 100.655 186.065 100.945 186.110 ;
        RECT 50.040 185.910 50.360 185.970 ;
        RECT 52.890 185.910 53.030 186.050 ;
        RECT 46.450 185.770 53.030 185.910 ;
        RECT 53.685 185.910 53.975 185.955 ;
        RECT 55.575 185.910 55.865 185.955 ;
        RECT 58.695 185.910 58.985 185.955 ;
        RECT 53.685 185.770 58.985 185.910 ;
        RECT 35.320 185.570 35.640 185.630 ;
        RECT 40.470 185.570 40.610 185.770 ;
        RECT 50.040 185.710 50.360 185.770 ;
        RECT 53.685 185.725 53.975 185.770 ;
        RECT 55.575 185.725 55.865 185.770 ;
        RECT 58.695 185.725 58.985 185.770 ;
        RECT 35.320 185.430 40.610 185.570 ;
        RECT 46.360 185.570 46.680 185.630 ;
        RECT 48.215 185.570 48.505 185.615 ;
        RECT 46.360 185.430 48.505 185.570 ;
        RECT 35.320 185.370 35.640 185.430 ;
        RECT 46.360 185.370 46.680 185.430 ;
        RECT 48.215 185.385 48.505 185.430 ;
        RECT 61.555 185.570 61.845 185.615 ;
        RECT 62.000 185.570 62.320 185.630 ;
        RECT 61.555 185.430 62.320 185.570 ;
        RECT 61.555 185.385 61.845 185.430 ;
        RECT 62.000 185.370 62.320 185.430 ;
        RECT 73.500 185.370 73.820 185.630 ;
        RECT 92.820 185.370 93.140 185.630 ;
        RECT 93.295 185.570 93.585 185.615 ;
        RECT 94.660 185.570 94.980 185.630 ;
        RECT 93.295 185.430 94.980 185.570 ;
        RECT 93.295 185.385 93.585 185.430 ;
        RECT 94.660 185.370 94.980 185.430 ;
        RECT 99.275 185.570 99.565 185.615 ;
        RECT 101.100 185.570 101.420 185.630 ;
        RECT 99.275 185.430 101.420 185.570 ;
        RECT 99.275 185.385 99.565 185.430 ;
        RECT 101.100 185.370 101.420 185.430 ;
        RECT 101.560 185.570 101.880 185.630 ;
        RECT 103.875 185.570 104.165 185.615 ;
        RECT 101.560 185.430 104.165 185.570 ;
        RECT 101.560 185.370 101.880 185.430 ;
        RECT 103.875 185.385 104.165 185.430 ;
        RECT 11.330 184.750 113.450 185.230 ;
        RECT 23.820 184.350 24.140 184.610 ;
        RECT 34.860 184.350 35.180 184.610 ;
        RECT 37.620 184.550 37.940 184.610 ;
        RECT 39.475 184.550 39.765 184.595 ;
        RECT 37.620 184.410 39.765 184.550 ;
        RECT 37.620 184.350 37.940 184.410 ;
        RECT 39.475 184.365 39.765 184.410 ;
        RECT 44.980 184.350 45.300 184.610 ;
        RECT 49.135 184.550 49.425 184.595 ;
        RECT 49.580 184.550 49.900 184.610 ;
        RECT 49.135 184.410 49.900 184.550 ;
        RECT 49.135 184.365 49.425 184.410 ;
        RECT 49.580 184.350 49.900 184.410 ;
        RECT 32.100 184.210 32.420 184.270 ;
        RECT 29.890 184.070 32.420 184.210 ;
        RECT 29.890 183.915 30.030 184.070 ;
        RECT 32.100 184.010 32.420 184.070 ;
        RECT 34.400 184.210 34.720 184.270 ;
        RECT 36.715 184.210 37.005 184.255 ;
        RECT 34.400 184.070 37.005 184.210 ;
        RECT 34.400 184.010 34.720 184.070 ;
        RECT 36.715 184.025 37.005 184.070 ;
        RECT 59.240 184.210 59.560 184.270 ;
        RECT 66.140 184.210 66.460 184.270 ;
        RECT 59.240 184.070 66.460 184.210 ;
        RECT 59.240 184.010 59.560 184.070 ;
        RECT 29.815 183.685 30.105 183.915 ;
        RECT 30.260 183.870 30.580 183.930 ;
        RECT 30.735 183.870 31.025 183.915 ;
        RECT 30.260 183.730 31.025 183.870 ;
        RECT 32.190 183.870 32.330 184.010 ;
        RECT 35.780 183.870 36.100 183.930 ;
        RECT 32.190 183.730 36.100 183.870 ;
        RECT 30.260 183.670 30.580 183.730 ;
        RECT 30.735 183.685 31.025 183.730 ;
        RECT 35.780 183.670 36.100 183.730 ;
        RECT 46.360 183.670 46.680 183.930 ;
        RECT 60.160 183.870 60.480 183.930 ;
        RECT 64.300 183.870 64.620 183.930 ;
        RECT 64.850 183.915 64.990 184.070 ;
        RECT 66.140 184.010 66.460 184.070 ;
        RECT 76.230 184.210 76.520 184.255 ;
        RECT 79.010 184.210 79.300 184.255 ;
        RECT 80.870 184.210 81.160 184.255 ;
        RECT 81.795 184.210 82.085 184.255 ;
        RECT 76.230 184.070 81.160 184.210 ;
        RECT 76.230 184.025 76.520 184.070 ;
        RECT 79.010 184.025 79.300 184.070 ;
        RECT 80.870 184.025 81.160 184.070 ;
        RECT 81.410 184.070 82.085 184.210 ;
        RECT 60.160 183.730 64.620 183.870 ;
        RECT 60.160 183.670 60.480 183.730 ;
        RECT 64.300 183.670 64.620 183.730 ;
        RECT 64.775 183.685 65.065 183.915 ;
        RECT 65.235 183.870 65.525 183.915 ;
        RECT 66.600 183.870 66.920 183.930 ;
        RECT 68.440 183.870 68.760 183.930 ;
        RECT 81.410 183.870 81.550 184.070 ;
        RECT 81.795 184.025 82.085 184.070 ;
        RECT 90.635 184.210 90.925 184.255 ;
        RECT 93.755 184.210 94.045 184.255 ;
        RECT 95.645 184.210 95.935 184.255 ;
        RECT 90.635 184.070 95.935 184.210 ;
        RECT 90.635 184.025 90.925 184.070 ;
        RECT 93.755 184.025 94.045 184.070 ;
        RECT 95.645 184.025 95.935 184.070 ;
        RECT 104.895 184.210 105.185 184.255 ;
        RECT 108.015 184.210 108.305 184.255 ;
        RECT 109.905 184.210 110.195 184.255 ;
        RECT 104.895 184.070 110.195 184.210 ;
        RECT 104.895 184.025 105.185 184.070 ;
        RECT 108.015 184.025 108.305 184.070 ;
        RECT 109.905 184.025 110.195 184.070 ;
        RECT 82.240 183.870 82.560 183.930 ;
        RECT 84.540 183.870 84.860 183.930 ;
        RECT 65.235 183.730 68.760 183.870 ;
        RECT 65.235 183.685 65.525 183.730 ;
        RECT 66.600 183.670 66.920 183.730 ;
        RECT 68.440 183.670 68.760 183.730 ;
        RECT 79.570 183.730 81.550 183.870 ;
        RECT 81.870 183.730 84.860 183.870 ;
        RECT 22.900 183.330 23.220 183.590 ;
        RECT 24.295 183.530 24.585 183.575 ;
        RECT 24.740 183.530 25.060 183.590 ;
        RECT 28.895 183.530 29.185 183.575 ;
        RECT 31.180 183.530 31.500 183.590 ;
        RECT 24.295 183.390 27.270 183.530 ;
        RECT 24.295 183.345 24.585 183.390 ;
        RECT 24.740 183.330 25.060 183.390 ;
        RECT 27.130 183.250 27.270 183.390 ;
        RECT 28.895 183.390 31.500 183.530 ;
        RECT 28.895 183.345 29.185 183.390 ;
        RECT 31.180 183.330 31.500 183.390 ;
        RECT 35.335 183.530 35.625 183.575 ;
        RECT 37.175 183.530 37.465 183.575 ;
        RECT 35.335 183.390 37.465 183.530 ;
        RECT 35.335 183.345 35.625 183.390 ;
        RECT 37.175 183.345 37.465 183.390 ;
        RECT 39.000 183.530 39.320 183.590 ;
        RECT 40.395 183.530 40.685 183.575 ;
        RECT 39.000 183.390 40.685 183.530 ;
        RECT 27.040 183.190 27.360 183.250 ;
        RECT 35.410 183.190 35.550 183.345 ;
        RECT 39.000 183.330 39.320 183.390 ;
        RECT 40.395 183.345 40.685 183.390 ;
        RECT 44.060 183.530 44.380 183.590 ;
        RECT 44.535 183.530 44.825 183.575 ;
        RECT 44.060 183.390 44.825 183.530 ;
        RECT 44.060 183.330 44.380 183.390 ;
        RECT 44.535 183.345 44.825 183.390 ;
        RECT 57.860 183.530 58.180 183.590 ;
        RECT 63.855 183.530 64.145 183.575 ;
        RECT 65.680 183.530 66.000 183.590 ;
        RECT 79.570 183.575 79.710 183.730 ;
        RECT 57.860 183.390 66.000 183.530 ;
        RECT 27.040 183.050 35.550 183.190 ;
        RECT 44.610 183.190 44.750 183.345 ;
        RECT 57.860 183.330 58.180 183.390 ;
        RECT 63.855 183.345 64.145 183.390 ;
        RECT 65.680 183.330 66.000 183.390 ;
        RECT 76.230 183.530 76.520 183.575 ;
        RECT 76.230 183.390 78.765 183.530 ;
        RECT 76.230 183.345 76.520 183.390 ;
        RECT 46.360 183.190 46.680 183.250 ;
        RECT 44.610 183.050 46.680 183.190 ;
        RECT 27.040 182.990 27.360 183.050 ;
        RECT 46.360 182.990 46.680 183.050 ;
        RECT 61.540 183.190 61.860 183.250 ;
        RECT 62.935 183.190 63.225 183.235 ;
        RECT 61.540 183.050 63.225 183.190 ;
        RECT 61.540 182.990 61.860 183.050 ;
        RECT 62.935 183.005 63.225 183.050 ;
        RECT 73.500 183.190 73.820 183.250 ;
        RECT 78.550 183.235 78.765 183.390 ;
        RECT 79.495 183.345 79.785 183.575 ;
        RECT 81.335 183.530 81.625 183.575 ;
        RECT 81.870 183.530 82.010 183.730 ;
        RECT 82.240 183.670 82.560 183.730 ;
        RECT 84.540 183.670 84.860 183.730 ;
        RECT 92.820 183.870 93.140 183.930 ;
        RECT 95.135 183.870 95.425 183.915 ;
        RECT 92.820 183.730 95.425 183.870 ;
        RECT 92.820 183.670 93.140 183.730 ;
        RECT 95.135 183.685 95.425 183.730 ;
        RECT 96.500 183.670 96.820 183.930 ;
        RECT 102.035 183.870 102.325 183.915 ;
        RECT 97.050 183.730 102.325 183.870 ;
        RECT 81.335 183.390 82.010 183.530 ;
        RECT 81.335 183.345 81.625 183.390 ;
        RECT 82.715 183.345 83.005 183.575 ;
        RECT 84.080 183.530 84.400 183.590 ;
        RECT 97.050 183.575 97.190 183.730 ;
        RECT 102.035 183.685 102.325 183.730 ;
        RECT 110.760 183.670 111.080 183.930 ;
        RECT 85.475 183.530 85.765 183.575 ;
        RECT 85.935 183.530 86.225 183.575 ;
        RECT 84.080 183.390 86.225 183.530 ;
        RECT 74.370 183.190 74.660 183.235 ;
        RECT 77.630 183.190 77.920 183.235 ;
        RECT 73.500 183.050 77.920 183.190 ;
        RECT 73.500 182.990 73.820 183.050 ;
        RECT 74.370 183.005 74.660 183.050 ;
        RECT 77.630 183.005 77.920 183.050 ;
        RECT 78.550 183.190 78.840 183.235 ;
        RECT 80.410 183.190 80.700 183.235 ;
        RECT 78.550 183.050 80.700 183.190 ;
        RECT 78.550 183.005 78.840 183.050 ;
        RECT 80.410 183.005 80.700 183.050 ;
        RECT 24.740 182.650 25.060 182.910 ;
        RECT 26.580 182.650 26.900 182.910 ;
        RECT 28.435 182.850 28.725 182.895 ;
        RECT 28.880 182.850 29.200 182.910 ;
        RECT 28.435 182.710 29.200 182.850 ;
        RECT 28.435 182.665 28.725 182.710 ;
        RECT 28.880 182.650 29.200 182.710 ;
        RECT 32.100 182.850 32.420 182.910 ;
        RECT 33.955 182.850 34.245 182.895 ;
        RECT 32.100 182.710 34.245 182.850 ;
        RECT 32.100 182.650 32.420 182.710 ;
        RECT 33.955 182.665 34.245 182.710 ;
        RECT 43.600 182.650 43.920 182.910 ;
        RECT 58.780 182.850 59.100 182.910 ;
        RECT 66.600 182.850 66.920 182.910 ;
        RECT 58.780 182.710 66.920 182.850 ;
        RECT 58.780 182.650 59.100 182.710 ;
        RECT 66.600 182.650 66.920 182.710 ;
        RECT 71.660 182.850 71.980 182.910 ;
        RECT 72.365 182.850 72.655 182.895 ;
        RECT 71.660 182.710 72.655 182.850 ;
        RECT 71.660 182.650 71.980 182.710 ;
        RECT 72.365 182.665 72.655 182.710 ;
        RECT 76.720 182.850 77.040 182.910 ;
        RECT 82.790 182.850 82.930 183.345 ;
        RECT 84.080 183.330 84.400 183.390 ;
        RECT 85.475 183.345 85.765 183.390 ;
        RECT 85.935 183.345 86.225 183.390 ;
        RECT 89.555 183.235 89.845 183.550 ;
        RECT 90.635 183.530 90.925 183.575 ;
        RECT 94.215 183.530 94.505 183.575 ;
        RECT 96.050 183.530 96.340 183.575 ;
        RECT 90.635 183.390 96.340 183.530 ;
        RECT 90.635 183.345 90.925 183.390 ;
        RECT 94.215 183.345 94.505 183.390 ;
        RECT 96.050 183.345 96.340 183.390 ;
        RECT 96.975 183.345 97.265 183.575 ;
        RECT 98.800 183.530 99.120 183.590 ;
        RECT 100.655 183.530 100.945 183.575 ;
        RECT 98.800 183.390 100.945 183.530 ;
        RECT 86.395 183.190 86.685 183.235 ;
        RECT 89.255 183.190 89.845 183.235 ;
        RECT 92.495 183.190 93.145 183.235 ;
        RECT 86.395 183.050 93.145 183.190 ;
        RECT 86.395 183.005 86.685 183.050 ;
        RECT 89.255 183.005 89.545 183.050 ;
        RECT 92.495 183.005 93.145 183.050 ;
        RECT 96.500 183.190 96.820 183.250 ;
        RECT 97.050 183.190 97.190 183.345 ;
        RECT 98.800 183.330 99.120 183.390 ;
        RECT 100.655 183.345 100.945 183.390 ;
        RECT 103.815 183.235 104.105 183.550 ;
        RECT 104.895 183.530 105.185 183.575 ;
        RECT 108.475 183.530 108.765 183.575 ;
        RECT 110.310 183.530 110.600 183.575 ;
        RECT 104.895 183.390 110.600 183.530 ;
        RECT 104.895 183.345 105.185 183.390 ;
        RECT 108.475 183.345 108.765 183.390 ;
        RECT 110.310 183.345 110.600 183.390 ;
        RECT 96.500 183.050 97.190 183.190 ;
        RECT 101.115 183.190 101.405 183.235 ;
        RECT 103.515 183.190 104.105 183.235 ;
        RECT 106.755 183.190 107.405 183.235 ;
        RECT 101.115 183.050 107.405 183.190 ;
        RECT 96.500 182.990 96.820 183.050 ;
        RECT 101.115 183.005 101.405 183.050 ;
        RECT 103.515 183.005 103.805 183.050 ;
        RECT 106.755 183.005 107.405 183.050 ;
        RECT 109.395 183.190 109.685 183.235 ;
        RECT 109.840 183.190 110.160 183.250 ;
        RECT 109.395 183.050 110.160 183.190 ;
        RECT 109.395 183.005 109.685 183.050 ;
        RECT 109.840 182.990 110.160 183.050 ;
        RECT 76.720 182.710 82.930 182.850 ;
        RECT 76.720 182.650 77.040 182.710 ;
        RECT 85.000 182.650 85.320 182.910 ;
        RECT 87.760 182.650 88.080 182.910 ;
        RECT 100.180 182.650 100.500 182.910 ;
        RECT 11.330 182.030 113.450 182.510 ;
        RECT 22.455 181.830 22.745 181.875 ;
        RECT 22.900 181.830 23.220 181.890 ;
        RECT 22.455 181.690 23.220 181.830 ;
        RECT 22.455 181.645 22.745 181.690 ;
        RECT 22.900 181.630 23.220 181.690 ;
        RECT 32.100 181.830 32.420 181.890 ;
        RECT 36.715 181.830 37.005 181.875 ;
        RECT 32.100 181.690 37.005 181.830 ;
        RECT 32.100 181.630 32.420 181.690 ;
        RECT 36.715 181.645 37.005 181.690 ;
        RECT 39.000 181.630 39.320 181.890 ;
        RECT 60.160 181.830 60.480 181.890 ;
        RECT 58.410 181.690 60.480 181.830 ;
        RECT 26.580 181.490 26.900 181.550 ;
        RECT 30.720 181.490 31.040 181.550 ;
        RECT 19.770 181.350 26.900 181.490 ;
        RECT 19.770 181.195 19.910 181.350 ;
        RECT 26.580 181.290 26.900 181.350 ;
        RECT 28.970 181.350 31.040 181.490 ;
        RECT 28.970 181.195 29.110 181.350 ;
        RECT 30.720 181.290 31.040 181.350 ;
        RECT 34.875 181.490 35.165 181.535 ;
        RECT 37.175 181.490 37.465 181.535 ;
        RECT 34.875 181.350 37.465 181.490 ;
        RECT 34.875 181.305 35.165 181.350 ;
        RECT 37.175 181.305 37.465 181.350 ;
        RECT 40.955 181.490 41.245 181.535 ;
        RECT 43.600 181.490 43.920 181.550 ;
        RECT 44.195 181.490 44.845 181.535 ;
        RECT 40.955 181.350 44.845 181.490 ;
        RECT 40.955 181.305 41.545 181.350 ;
        RECT 19.695 180.965 19.985 181.195 ;
        RECT 27.975 181.150 28.265 181.195 ;
        RECT 27.975 181.010 28.650 181.150 ;
        RECT 27.975 180.965 28.265 181.010 ;
        RECT 24.755 180.810 25.045 180.855 ;
        RECT 25.200 180.810 25.520 180.870 ;
        RECT 24.755 180.670 25.520 180.810 ;
        RECT 24.755 180.625 25.045 180.670 ;
        RECT 25.200 180.610 25.520 180.670 ;
        RECT 28.510 180.470 28.650 181.010 ;
        RECT 28.895 180.965 29.185 181.195 ;
        RECT 29.340 180.950 29.660 181.210 ;
        RECT 30.045 181.150 30.335 181.195 ;
        RECT 32.115 181.150 32.405 181.195 ;
        RECT 30.045 181.010 31.870 181.150 ;
        RECT 30.045 180.965 30.335 181.010 ;
        RECT 31.730 180.810 31.870 181.010 ;
        RECT 32.115 181.010 39.690 181.150 ;
        RECT 32.115 180.965 32.405 181.010 ;
        RECT 33.940 180.810 34.260 180.870 ;
        RECT 31.730 180.670 34.260 180.810 ;
        RECT 33.940 180.610 34.260 180.670 ;
        RECT 35.780 180.610 36.100 180.870 ;
        RECT 38.080 180.810 38.400 180.870 ;
        RECT 39.550 180.855 39.690 181.010 ;
        RECT 41.255 180.990 41.545 181.305 ;
        RECT 43.600 181.290 43.920 181.350 ;
        RECT 44.195 181.305 44.845 181.350 ;
        RECT 58.410 181.195 58.550 181.690 ;
        RECT 60.160 181.630 60.480 181.690 ;
        RECT 60.620 181.830 60.940 181.890 ;
        RECT 64.760 181.830 65.080 181.890 ;
        RECT 66.155 181.830 66.445 181.875 ;
        RECT 60.620 181.690 63.150 181.830 ;
        RECT 60.620 181.630 60.940 181.690 ;
        RECT 63.010 181.535 63.150 181.690 ;
        RECT 64.760 181.690 66.445 181.830 ;
        RECT 64.760 181.630 65.080 181.690 ;
        RECT 66.155 181.645 66.445 181.690 ;
        RECT 66.600 181.630 66.920 181.890 ;
        RECT 73.975 181.830 74.265 181.875 ;
        RECT 76.720 181.830 77.040 181.890 ;
        RECT 73.975 181.690 77.040 181.830 ;
        RECT 73.975 181.645 74.265 181.690 ;
        RECT 76.720 181.630 77.040 181.690 ;
        RECT 79.035 181.645 79.325 181.875 ;
        RECT 90.995 181.830 91.285 181.875 ;
        RECT 91.900 181.830 92.220 181.890 ;
        RECT 90.995 181.690 92.220 181.830 ;
        RECT 90.995 181.645 91.285 181.690 ;
        RECT 58.870 181.350 61.310 181.490 ;
        RECT 58.870 181.210 59.010 181.350 ;
        RECT 42.335 181.150 42.625 181.195 ;
        RECT 45.915 181.150 46.205 181.195 ;
        RECT 47.750 181.150 48.040 181.195 ;
        RECT 42.335 181.010 48.040 181.150 ;
        RECT 42.335 180.965 42.625 181.010 ;
        RECT 45.915 180.965 46.205 181.010 ;
        RECT 47.750 180.965 48.040 181.010 ;
        RECT 58.335 180.965 58.625 181.195 ;
        RECT 58.780 180.950 59.100 181.210 ;
        RECT 59.240 180.950 59.560 181.210 ;
        RECT 60.160 181.150 60.480 181.210 ;
        RECT 61.170 181.195 61.310 181.350 ;
        RECT 62.935 181.305 63.225 181.535 ;
        RECT 63.855 181.490 64.145 181.535 ;
        RECT 65.680 181.490 66.000 181.550 ;
        RECT 63.855 181.350 66.000 181.490 ;
        RECT 63.855 181.305 64.145 181.350 ;
        RECT 60.635 181.150 60.925 181.195 ;
        RECT 60.160 181.010 60.925 181.150 ;
        RECT 60.160 180.950 60.480 181.010 ;
        RECT 60.635 180.965 60.925 181.010 ;
        RECT 61.095 180.965 61.385 181.195 ;
        RECT 61.555 181.150 61.845 181.195 ;
        RECT 63.930 181.150 64.070 181.305 ;
        RECT 65.680 181.290 66.000 181.350 ;
        RECT 76.260 181.490 76.580 181.550 ;
        RECT 79.110 181.490 79.250 181.645 ;
        RECT 91.900 181.630 92.220 181.690 ;
        RECT 76.260 181.350 79.250 181.490 ;
        RECT 82.815 181.490 83.105 181.535 ;
        RECT 85.000 181.490 85.320 181.550 ;
        RECT 86.055 181.490 86.705 181.535 ;
        RECT 82.815 181.350 86.705 181.490 ;
        RECT 76.260 181.290 76.580 181.350 ;
        RECT 82.815 181.305 83.405 181.350 ;
        RECT 61.555 181.010 64.070 181.150 ;
        RECT 61.555 180.965 61.845 181.010 ;
        RECT 69.360 180.950 69.680 181.210 ;
        RECT 72.135 181.150 72.425 181.195 ;
        RECT 73.040 181.150 73.360 181.210 ;
        RECT 76.735 181.150 77.025 181.195 ;
        RECT 72.135 181.010 77.025 181.150 ;
        RECT 72.135 180.965 72.425 181.010 ;
        RECT 73.040 180.950 73.360 181.010 ;
        RECT 76.735 180.965 77.025 181.010 ;
        RECT 77.195 181.150 77.485 181.195 ;
        RECT 79.480 181.150 79.800 181.210 ;
        RECT 77.195 181.010 81.550 181.150 ;
        RECT 77.195 180.965 77.485 181.010 ;
        RECT 79.480 180.950 79.800 181.010 ;
        RECT 36.330 180.670 38.400 180.810 ;
        RECT 29.800 180.470 30.120 180.530 ;
        RECT 28.510 180.330 30.120 180.470 ;
        RECT 29.800 180.270 30.120 180.330 ;
        RECT 27.515 180.130 27.805 180.175 ;
        RECT 28.880 180.130 29.200 180.190 ;
        RECT 27.515 179.990 29.200 180.130 ;
        RECT 27.515 179.945 27.805 179.990 ;
        RECT 28.880 179.930 29.200 179.990 ;
        RECT 31.195 180.130 31.485 180.175 ;
        RECT 36.330 180.130 36.470 180.670 ;
        RECT 38.080 180.610 38.400 180.670 ;
        RECT 39.475 180.810 39.765 180.855 ;
        RECT 41.760 180.810 42.080 180.870 ;
        RECT 39.475 180.670 42.080 180.810 ;
        RECT 39.475 180.625 39.765 180.670 ;
        RECT 41.760 180.610 42.080 180.670 ;
        RECT 48.215 180.810 48.505 180.855 ;
        RECT 50.040 180.810 50.360 180.870 ;
        RECT 48.215 180.670 50.360 180.810 ;
        RECT 48.215 180.625 48.505 180.670 ;
        RECT 50.040 180.610 50.360 180.670 ;
        RECT 57.860 180.610 58.180 180.870 ;
        RECT 62.015 180.625 62.305 180.855 ;
        RECT 67.060 180.810 67.380 180.870 ;
        RECT 67.535 180.810 67.825 180.855 ;
        RECT 67.060 180.670 67.825 180.810 ;
        RECT 42.335 180.470 42.625 180.515 ;
        RECT 45.455 180.470 45.745 180.515 ;
        RECT 47.345 180.470 47.635 180.515 ;
        RECT 42.335 180.330 47.635 180.470 ;
        RECT 62.090 180.470 62.230 180.625 ;
        RECT 67.060 180.610 67.380 180.670 ;
        RECT 67.535 180.625 67.825 180.670 ;
        RECT 68.915 180.810 69.205 180.855 ;
        RECT 70.740 180.810 71.060 180.870 ;
        RECT 68.915 180.670 71.060 180.810 ;
        RECT 68.915 180.625 69.205 180.670 ;
        RECT 70.740 180.610 71.060 180.670 ;
        RECT 71.200 180.610 71.520 180.870 ;
        RECT 71.660 180.610 71.980 180.870 ;
        RECT 75.815 180.810 76.105 180.855 ;
        RECT 77.640 180.810 77.960 180.870 ;
        RECT 81.410 180.855 81.550 181.010 ;
        RECT 83.115 180.990 83.405 181.305 ;
        RECT 85.000 181.290 85.320 181.350 ;
        RECT 86.055 181.305 86.705 181.350 ;
        RECT 92.835 181.490 93.125 181.535 ;
        RECT 94.660 181.490 94.980 181.550 ;
        RECT 97.435 181.490 97.725 181.535 ;
        RECT 92.835 181.350 97.725 181.490 ;
        RECT 92.835 181.305 93.125 181.350 ;
        RECT 94.660 181.290 94.980 181.350 ;
        RECT 97.435 181.305 97.725 181.350 ;
        RECT 97.895 181.490 98.185 181.535 ;
        RECT 100.180 181.490 100.500 181.550 ;
        RECT 97.895 181.350 100.500 181.490 ;
        RECT 97.895 181.305 98.185 181.350 ;
        RECT 100.180 181.290 100.500 181.350 ;
        RECT 101.100 181.490 101.420 181.550 ;
        RECT 102.135 181.490 102.425 181.535 ;
        RECT 105.375 181.490 106.025 181.535 ;
        RECT 101.100 181.350 106.025 181.490 ;
        RECT 101.100 181.290 101.420 181.350 ;
        RECT 102.135 181.305 102.725 181.350 ;
        RECT 105.375 181.305 106.025 181.350 ;
        RECT 84.195 181.150 84.485 181.195 ;
        RECT 87.775 181.150 88.065 181.195 ;
        RECT 89.610 181.150 89.900 181.195 ;
        RECT 84.195 181.010 89.900 181.150 ;
        RECT 84.195 180.965 84.485 181.010 ;
        RECT 87.775 180.965 88.065 181.010 ;
        RECT 89.610 180.965 89.900 181.010 ;
        RECT 102.435 180.990 102.725 181.305 ;
        RECT 103.515 181.150 103.805 181.195 ;
        RECT 107.095 181.150 107.385 181.195 ;
        RECT 108.930 181.150 109.220 181.195 ;
        RECT 103.515 181.010 109.220 181.150 ;
        RECT 103.515 180.965 103.805 181.010 ;
        RECT 107.095 180.965 107.385 181.010 ;
        RECT 108.930 180.965 109.220 181.010 ;
        RECT 109.395 181.150 109.685 181.195 ;
        RECT 110.760 181.150 111.080 181.210 ;
        RECT 109.395 181.010 111.080 181.150 ;
        RECT 109.395 180.965 109.685 181.010 ;
        RECT 110.760 180.950 111.080 181.010 ;
        RECT 75.815 180.670 77.960 180.810 ;
        RECT 75.815 180.625 76.105 180.670 ;
        RECT 62.460 180.470 62.780 180.530 ;
        RECT 62.090 180.330 62.780 180.470 ;
        RECT 42.335 180.285 42.625 180.330 ;
        RECT 45.455 180.285 45.745 180.330 ;
        RECT 47.345 180.285 47.635 180.330 ;
        RECT 62.460 180.270 62.780 180.330 ;
        RECT 63.855 180.470 64.145 180.515 ;
        RECT 66.140 180.470 66.460 180.530 ;
        RECT 63.855 180.330 66.460 180.470 ;
        RECT 71.290 180.470 71.430 180.610 ;
        RECT 75.890 180.470 76.030 180.625 ;
        RECT 77.640 180.610 77.960 180.670 ;
        RECT 81.335 180.625 81.625 180.855 ;
        RECT 82.240 180.810 82.560 180.870 ;
        RECT 90.075 180.810 90.365 180.855 ;
        RECT 82.240 180.670 90.365 180.810 ;
        RECT 82.240 180.610 82.560 180.670 ;
        RECT 90.075 180.625 90.365 180.670 ;
        RECT 90.980 180.810 91.300 180.870 ;
        RECT 93.295 180.810 93.585 180.855 ;
        RECT 90.980 180.670 93.585 180.810 ;
        RECT 90.980 180.610 91.300 180.670 ;
        RECT 93.295 180.625 93.585 180.670 ;
        RECT 93.740 180.810 94.060 180.870 ;
        RECT 96.515 180.810 96.805 180.855 ;
        RECT 100.655 180.810 100.945 180.855 ;
        RECT 93.740 180.670 96.805 180.810 ;
        RECT 93.740 180.610 94.060 180.670 ;
        RECT 96.515 180.625 96.805 180.670 ;
        RECT 97.510 180.670 100.945 180.810 ;
        RECT 71.290 180.330 76.030 180.470 ;
        RECT 77.730 180.470 77.870 180.610 ;
        RECT 83.620 180.470 83.940 180.530 ;
        RECT 77.730 180.330 83.940 180.470 ;
        RECT 63.855 180.285 64.145 180.330 ;
        RECT 66.140 180.270 66.460 180.330 ;
        RECT 83.620 180.270 83.940 180.330 ;
        RECT 84.195 180.470 84.485 180.515 ;
        RECT 87.315 180.470 87.605 180.515 ;
        RECT 89.205 180.470 89.495 180.515 ;
        RECT 84.195 180.330 89.495 180.470 ;
        RECT 84.195 180.285 84.485 180.330 ;
        RECT 87.315 180.285 87.605 180.330 ;
        RECT 89.205 180.285 89.495 180.330 ;
        RECT 95.120 180.470 95.440 180.530 ;
        RECT 97.510 180.470 97.650 180.670 ;
        RECT 100.655 180.625 100.945 180.670 ;
        RECT 95.120 180.330 97.650 180.470 ;
        RECT 103.515 180.470 103.805 180.515 ;
        RECT 106.635 180.470 106.925 180.515 ;
        RECT 108.525 180.470 108.815 180.515 ;
        RECT 103.515 180.330 108.815 180.470 ;
        RECT 95.120 180.270 95.440 180.330 ;
        RECT 103.515 180.285 103.805 180.330 ;
        RECT 106.635 180.285 106.925 180.330 ;
        RECT 108.525 180.285 108.815 180.330 ;
        RECT 31.195 179.990 36.470 180.130 ;
        RECT 46.820 180.175 47.140 180.190 ;
        RECT 31.195 179.945 31.485 179.990 ;
        RECT 46.820 179.945 47.190 180.175 ;
        RECT 56.955 180.130 57.245 180.175 ;
        RECT 58.780 180.130 59.100 180.190 ;
        RECT 56.955 179.990 59.100 180.130 ;
        RECT 56.955 179.945 57.245 179.990 ;
        RECT 46.820 179.930 47.140 179.945 ;
        RECT 58.780 179.930 59.100 179.990 ;
        RECT 88.790 180.130 89.080 180.175 ;
        RECT 91.440 180.130 91.760 180.190 ;
        RECT 88.790 179.990 91.760 180.130 ;
        RECT 88.790 179.945 89.080 179.990 ;
        RECT 91.440 179.930 91.760 179.990 ;
        RECT 99.735 180.130 100.025 180.175 ;
        RECT 104.320 180.130 104.640 180.190 ;
        RECT 99.735 179.990 104.640 180.130 ;
        RECT 99.735 179.945 100.025 179.990 ;
        RECT 104.320 179.930 104.640 179.990 ;
        RECT 105.240 180.130 105.560 180.190 ;
        RECT 108.080 180.130 108.370 180.175 ;
        RECT 105.240 179.990 108.370 180.130 ;
        RECT 105.240 179.930 105.560 179.990 ;
        RECT 108.080 179.945 108.370 179.990 ;
        RECT 11.330 179.310 113.450 179.790 ;
        RECT 31.180 179.110 31.500 179.170 ;
        RECT 40.380 179.110 40.700 179.170 ;
        RECT 31.180 178.970 40.700 179.110 ;
        RECT 31.180 178.910 31.500 178.970 ;
        RECT 40.380 178.910 40.700 178.970 ;
        RECT 46.820 178.910 47.140 179.170 ;
        RECT 66.140 179.110 66.460 179.170 ;
        RECT 64.850 178.970 66.460 179.110 ;
        RECT 21.485 178.770 21.775 178.815 ;
        RECT 23.375 178.770 23.665 178.815 ;
        RECT 26.495 178.770 26.785 178.815 ;
        RECT 21.485 178.630 26.785 178.770 ;
        RECT 21.485 178.585 21.775 178.630 ;
        RECT 23.375 178.585 23.665 178.630 ;
        RECT 26.495 178.585 26.785 178.630 ;
        RECT 29.340 178.770 29.660 178.830 ;
        RECT 30.720 178.770 31.040 178.830 ;
        RECT 33.940 178.770 34.260 178.830 ;
        RECT 51.420 178.770 51.740 178.830 ;
        RECT 62.000 178.770 62.320 178.830 ;
        RECT 63.395 178.770 63.685 178.815 ;
        RECT 29.340 178.630 33.710 178.770 ;
        RECT 29.340 178.570 29.660 178.630 ;
        RECT 30.720 178.570 31.040 178.630 ;
        RECT 20.600 178.230 20.920 178.490 ;
        RECT 30.260 178.430 30.580 178.490 ;
        RECT 33.570 178.430 33.710 178.630 ;
        RECT 33.940 178.630 51.740 178.770 ;
        RECT 33.940 178.570 34.260 178.630 ;
        RECT 51.420 178.570 51.740 178.630 ;
        RECT 56.800 178.630 61.770 178.770 ;
        RECT 56.800 178.430 56.940 178.630 ;
        RECT 30.260 178.290 33.250 178.430 ;
        RECT 30.260 178.230 30.580 178.290 ;
        RECT 33.110 178.135 33.250 178.290 ;
        RECT 33.570 178.290 56.940 178.430 ;
        RECT 33.570 178.135 33.710 178.290 ;
        RECT 58.320 178.230 58.640 178.490 ;
        RECT 61.630 178.430 61.770 178.630 ;
        RECT 62.000 178.630 63.685 178.770 ;
        RECT 62.000 178.570 62.320 178.630 ;
        RECT 63.395 178.585 63.685 178.630 ;
        RECT 61.630 178.290 64.070 178.430 ;
        RECT 21.080 178.090 21.370 178.135 ;
        RECT 22.915 178.090 23.205 178.135 ;
        RECT 26.495 178.090 26.785 178.135 ;
        RECT 21.080 177.950 26.785 178.090 ;
        RECT 21.080 177.905 21.370 177.950 ;
        RECT 22.915 177.905 23.205 177.950 ;
        RECT 26.495 177.905 26.785 177.950 ;
        RECT 21.980 177.550 22.300 177.810 ;
        RECT 24.740 177.795 25.060 177.810 ;
        RECT 24.275 177.750 25.060 177.795 ;
        RECT 27.575 177.795 27.865 178.110 ;
        RECT 32.115 177.905 32.405 178.135 ;
        RECT 33.035 177.905 33.325 178.135 ;
        RECT 33.495 177.905 33.785 178.135 ;
        RECT 27.575 177.750 28.165 177.795 ;
        RECT 24.275 177.610 28.165 177.750 ;
        RECT 32.190 177.750 32.330 177.905 ;
        RECT 33.940 177.890 34.260 178.150 ;
        RECT 37.160 178.090 37.480 178.150 ;
        RECT 40.855 178.090 41.145 178.135 ;
        RECT 37.160 177.950 41.145 178.090 ;
        RECT 37.160 177.890 37.480 177.950 ;
        RECT 40.855 177.905 41.145 177.950 ;
        RECT 41.315 177.905 41.605 178.135 ;
        RECT 38.540 177.750 38.860 177.810 ;
        RECT 32.190 177.610 38.860 177.750 ;
        RECT 24.275 177.565 25.060 177.610 ;
        RECT 27.875 177.565 28.165 177.610 ;
        RECT 24.740 177.550 25.060 177.565 ;
        RECT 38.540 177.550 38.860 177.610 ;
        RECT 39.000 177.750 39.320 177.810 ;
        RECT 41.390 177.750 41.530 177.905 ;
        RECT 41.760 177.890 42.080 178.150 ;
        RECT 42.680 177.890 43.000 178.150 ;
        RECT 43.615 178.090 43.905 178.135 ;
        RECT 44.980 178.090 45.300 178.150 ;
        RECT 43.615 177.950 45.300 178.090 ;
        RECT 43.615 177.905 43.905 177.950 ;
        RECT 44.980 177.890 45.300 177.950 ;
        RECT 46.375 178.090 46.665 178.135 ;
        RECT 47.755 178.090 48.045 178.135 ;
        RECT 46.375 177.950 48.045 178.090 ;
        RECT 46.375 177.905 46.665 177.950 ;
        RECT 47.755 177.905 48.045 177.950 ;
        RECT 49.580 178.090 49.900 178.150 ;
        RECT 50.975 178.090 51.265 178.135 ;
        RECT 49.580 177.950 51.265 178.090 ;
        RECT 49.580 177.890 49.900 177.950 ;
        RECT 50.975 177.905 51.265 177.950 ;
        RECT 56.940 178.090 57.260 178.150 ;
        RECT 57.415 178.090 57.705 178.135 ;
        RECT 56.940 177.950 57.705 178.090 ;
        RECT 56.940 177.890 57.260 177.950 ;
        RECT 57.415 177.905 57.705 177.950 ;
        RECT 62.015 178.090 62.305 178.135 ;
        RECT 62.460 178.090 62.780 178.150 ;
        RECT 62.015 177.950 62.780 178.090 ;
        RECT 63.930 178.090 64.070 178.290 ;
        RECT 64.300 178.230 64.620 178.490 ;
        RECT 64.850 178.475 64.990 178.970 ;
        RECT 66.140 178.910 66.460 178.970 ;
        RECT 68.915 179.110 69.205 179.155 ;
        RECT 71.200 179.110 71.520 179.170 ;
        RECT 68.915 178.970 71.520 179.110 ;
        RECT 68.915 178.925 69.205 178.970 ;
        RECT 71.200 178.910 71.520 178.970 ;
        RECT 73.040 178.910 73.360 179.170 ;
        RECT 91.440 178.910 91.760 179.170 ;
        RECT 105.240 178.910 105.560 179.170 ;
        RECT 107.555 179.110 107.845 179.155 ;
        RECT 109.840 179.110 110.160 179.170 ;
        RECT 107.555 178.970 110.160 179.110 ;
        RECT 107.555 178.925 107.845 178.970 ;
        RECT 109.840 178.910 110.160 178.970 ;
        RECT 66.600 178.770 66.920 178.830 ;
        RECT 65.310 178.630 66.920 178.770 ;
        RECT 65.310 178.475 65.450 178.630 ;
        RECT 66.600 178.570 66.920 178.630 ;
        RECT 76.375 178.770 76.665 178.815 ;
        RECT 79.495 178.770 79.785 178.815 ;
        RECT 81.385 178.770 81.675 178.815 ;
        RECT 93.740 178.770 94.060 178.830 ;
        RECT 76.375 178.630 81.675 178.770 ;
        RECT 76.375 178.585 76.665 178.630 ;
        RECT 79.495 178.585 79.785 178.630 ;
        RECT 81.385 178.585 81.675 178.630 ;
        RECT 86.010 178.630 94.060 178.770 ;
        RECT 64.775 178.245 65.065 178.475 ;
        RECT 65.235 178.245 65.525 178.475 ;
        RECT 65.680 178.230 66.000 178.490 ;
        RECT 67.980 178.430 68.300 178.490 ;
        RECT 66.230 178.290 68.300 178.430 ;
        RECT 66.230 178.090 66.370 178.290 ;
        RECT 67.980 178.230 68.300 178.290 ;
        RECT 73.515 178.245 73.805 178.475 ;
        RECT 63.930 177.950 66.370 178.090 ;
        RECT 66.600 178.090 66.920 178.150 ;
        RECT 69.835 178.090 70.125 178.135 ;
        RECT 73.590 178.090 73.730 178.245 ;
        RECT 82.240 178.230 82.560 178.490 ;
        RECT 83.620 178.430 83.940 178.490 ;
        RECT 86.010 178.475 86.150 178.630 ;
        RECT 93.740 178.570 94.060 178.630 ;
        RECT 85.935 178.430 86.225 178.475 ;
        RECT 83.620 178.290 86.225 178.430 ;
        RECT 83.620 178.230 83.940 178.290 ;
        RECT 85.935 178.245 86.225 178.290 ;
        RECT 87.760 178.430 88.080 178.490 ;
        RECT 90.520 178.430 90.840 178.490 ;
        RECT 87.760 178.290 90.840 178.430 ;
        RECT 93.830 178.430 93.970 178.570 ;
        RECT 100.655 178.430 100.945 178.475 ;
        RECT 93.830 178.290 100.945 178.430 ;
        RECT 87.760 178.230 88.080 178.290 ;
        RECT 90.520 178.230 90.840 178.290 ;
        RECT 100.655 178.245 100.945 178.290 ;
        RECT 66.600 177.950 73.730 178.090 ;
        RECT 62.015 177.905 62.305 177.950 ;
        RECT 62.460 177.890 62.780 177.950 ;
        RECT 66.600 177.890 66.920 177.950 ;
        RECT 69.835 177.905 70.125 177.950 ;
        RECT 39.000 177.610 41.530 177.750 ;
        RECT 43.140 177.750 43.460 177.810 ;
        RECT 52.355 177.750 52.645 177.795 ;
        RECT 43.140 177.610 52.645 177.750 ;
        RECT 39.000 177.550 39.320 177.610 ;
        RECT 43.140 177.550 43.460 177.610 ;
        RECT 52.355 177.565 52.645 177.610 ;
        RECT 54.195 177.750 54.485 177.795 ;
        RECT 67.520 177.750 67.840 177.810 ;
        RECT 54.195 177.610 67.840 177.750 ;
        RECT 54.195 177.565 54.485 177.610 ;
        RECT 67.520 177.550 67.840 177.610 ;
        RECT 70.740 177.750 71.060 177.810 ;
        RECT 75.295 177.795 75.585 178.110 ;
        RECT 76.375 178.090 76.665 178.135 ;
        RECT 79.955 178.090 80.245 178.135 ;
        RECT 81.790 178.090 82.080 178.135 ;
        RECT 85.475 178.090 85.765 178.135 ;
        RECT 76.375 177.950 82.080 178.090 ;
        RECT 76.375 177.905 76.665 177.950 ;
        RECT 79.955 177.905 80.245 177.950 ;
        RECT 81.790 177.905 82.080 177.950 ;
        RECT 82.330 177.950 85.765 178.090 ;
        RECT 74.995 177.750 75.585 177.795 ;
        RECT 78.235 177.750 78.885 177.795 ;
        RECT 70.740 177.610 78.885 177.750 ;
        RECT 70.740 177.550 71.060 177.610 ;
        RECT 74.995 177.565 75.285 177.610 ;
        RECT 78.235 177.565 78.885 177.610 ;
        RECT 80.860 177.550 81.180 177.810 ;
        RECT 82.330 177.750 82.470 177.950 ;
        RECT 85.475 177.905 85.765 177.950 ;
        RECT 87.300 178.090 87.620 178.150 ;
        RECT 92.375 178.090 92.665 178.135 ;
        RECT 87.300 177.950 92.665 178.090 ;
        RECT 87.300 177.890 87.620 177.950 ;
        RECT 92.375 177.905 92.665 177.950 ;
        RECT 94.200 177.890 94.520 178.150 ;
        RECT 94.675 177.905 94.965 178.135 ;
        RECT 81.410 177.610 82.470 177.750 ;
        RECT 85.015 177.750 85.305 177.795 ;
        RECT 90.980 177.750 91.300 177.810 ;
        RECT 85.015 177.610 91.300 177.750 ;
        RECT 94.750 177.750 94.890 177.905 ;
        RECT 95.120 177.890 95.440 178.150 ;
        RECT 96.040 177.890 96.360 178.150 ;
        RECT 100.180 178.090 100.500 178.150 ;
        RECT 101.115 178.090 101.405 178.135 ;
        RECT 100.180 177.950 101.405 178.090 ;
        RECT 100.180 177.890 100.500 177.950 ;
        RECT 101.115 177.905 101.405 177.950 ;
        RECT 101.560 177.890 101.880 178.150 ;
        RECT 104.320 177.890 104.640 178.150 ;
        RECT 106.635 177.905 106.925 178.135 ;
        RECT 97.420 177.750 97.740 177.810 ;
        RECT 106.710 177.750 106.850 177.905 ;
        RECT 94.750 177.610 97.740 177.750 ;
        RECT 25.200 177.410 25.520 177.470 ;
        RECT 29.340 177.410 29.660 177.470 ;
        RECT 25.200 177.270 29.660 177.410 ;
        RECT 25.200 177.210 25.520 177.270 ;
        RECT 29.340 177.210 29.660 177.270 ;
        RECT 30.260 177.410 30.580 177.470 ;
        RECT 33.940 177.410 34.260 177.470 ;
        RECT 30.260 177.270 34.260 177.410 ;
        RECT 30.260 177.210 30.580 177.270 ;
        RECT 33.940 177.210 34.260 177.270 ;
        RECT 35.320 177.210 35.640 177.470 ;
        RECT 39.460 177.210 39.780 177.470 ;
        RECT 51.895 177.410 52.185 177.455 ;
        RECT 56.480 177.410 56.800 177.470 ;
        RECT 51.895 177.270 56.800 177.410 ;
        RECT 51.895 177.225 52.185 177.270 ;
        RECT 56.480 177.210 56.800 177.270 ;
        RECT 62.475 177.410 62.765 177.455 ;
        RECT 64.760 177.410 65.080 177.470 ;
        RECT 62.475 177.270 65.080 177.410 ;
        RECT 62.475 177.225 62.765 177.270 ;
        RECT 64.760 177.210 65.080 177.270 ;
        RECT 79.480 177.410 79.800 177.470 ;
        RECT 81.410 177.410 81.550 177.610 ;
        RECT 85.015 177.565 85.305 177.610 ;
        RECT 90.980 177.550 91.300 177.610 ;
        RECT 97.420 177.550 97.740 177.610 ;
        RECT 105.100 177.610 106.850 177.750 ;
        RECT 79.480 177.270 81.550 177.410 ;
        RECT 79.480 177.210 79.800 177.270 ;
        RECT 83.160 177.210 83.480 177.470 ;
        RECT 92.835 177.410 93.125 177.455 ;
        RECT 95.120 177.410 95.440 177.470 ;
        RECT 92.835 177.270 95.440 177.410 ;
        RECT 92.835 177.225 93.125 177.270 ;
        RECT 95.120 177.210 95.440 177.270 ;
        RECT 103.415 177.410 103.705 177.455 ;
        RECT 105.100 177.410 105.240 177.610 ;
        RECT 103.415 177.270 105.240 177.410 ;
        RECT 103.415 177.225 103.705 177.270 ;
        RECT 11.330 176.590 113.450 177.070 ;
        RECT 21.980 176.390 22.300 176.450 ;
        RECT 23.835 176.390 24.125 176.435 ;
        RECT 21.980 176.250 24.125 176.390 ;
        RECT 21.980 176.190 22.300 176.250 ;
        RECT 23.835 176.205 24.125 176.250 ;
        RECT 28.880 176.190 29.200 176.450 ;
        RECT 32.100 176.390 32.420 176.450 ;
        RECT 32.575 176.390 32.865 176.435 ;
        RECT 32.100 176.250 32.865 176.390 ;
        RECT 32.100 176.190 32.420 176.250 ;
        RECT 32.575 176.205 32.865 176.250 ;
        RECT 41.760 176.390 42.080 176.450 ;
        RECT 44.075 176.390 44.365 176.435 ;
        RECT 41.760 176.250 44.365 176.390 ;
        RECT 41.760 176.190 42.080 176.250 ;
        RECT 44.075 176.205 44.365 176.250 ;
        RECT 44.980 176.390 45.300 176.450 ;
        RECT 46.375 176.390 46.665 176.435 ;
        RECT 49.135 176.390 49.425 176.435 ;
        RECT 44.980 176.250 46.665 176.390 ;
        RECT 44.980 176.190 45.300 176.250 ;
        RECT 46.375 176.205 46.665 176.250 ;
        RECT 46.910 176.250 49.425 176.390 ;
        RECT 38.540 176.050 38.860 176.110 ;
        RECT 46.910 176.050 47.050 176.250 ;
        RECT 49.135 176.205 49.425 176.250 ;
        RECT 51.420 176.390 51.740 176.450 ;
        RECT 59.715 176.390 60.005 176.435 ;
        RECT 80.415 176.390 80.705 176.435 ;
        RECT 80.860 176.390 81.180 176.450 ;
        RECT 51.420 176.250 80.170 176.390 ;
        RECT 51.420 176.190 51.740 176.250 ;
        RECT 59.715 176.205 60.005 176.250 ;
        RECT 35.410 175.910 38.860 176.050 ;
        RECT 24.755 175.525 25.045 175.755 ;
        RECT 25.215 175.710 25.505 175.755 ;
        RECT 26.580 175.710 26.900 175.770 ;
        RECT 25.215 175.570 26.900 175.710 ;
        RECT 25.215 175.525 25.505 175.570 ;
        RECT 24.830 175.370 24.970 175.525 ;
        RECT 26.580 175.510 26.900 175.570 ;
        RECT 28.420 175.710 28.740 175.770 ;
        RECT 35.410 175.755 35.550 175.910 ;
        RECT 38.540 175.850 38.860 175.910 ;
        RECT 39.550 175.910 47.050 176.050 ;
        RECT 47.755 176.050 48.045 176.095 ;
        RECT 50.615 176.050 50.905 176.095 ;
        RECT 53.855 176.050 54.505 176.095 ;
        RECT 47.755 175.910 54.505 176.050 ;
        RECT 32.115 175.710 32.405 175.755 ;
        RECT 28.420 175.570 32.405 175.710 ;
        RECT 28.420 175.510 28.740 175.570 ;
        RECT 32.115 175.525 32.405 175.570 ;
        RECT 35.335 175.525 35.625 175.755 ;
        RECT 36.240 175.510 36.560 175.770 ;
        RECT 36.715 175.525 37.005 175.755 ;
        RECT 29.815 175.370 30.105 175.415 ;
        RECT 31.655 175.370 31.945 175.415 ;
        RECT 35.780 175.370 36.100 175.430 ;
        RECT 24.830 175.230 26.810 175.370 ;
        RECT 26.670 175.075 26.810 175.230 ;
        RECT 29.815 175.230 36.100 175.370 ;
        RECT 36.790 175.370 36.930 175.525 ;
        RECT 37.160 175.510 37.480 175.770 ;
        RECT 39.550 175.755 39.690 175.910 ;
        RECT 44.150 175.770 44.290 175.910 ;
        RECT 47.755 175.865 48.045 175.910 ;
        RECT 50.615 175.865 51.205 175.910 ;
        RECT 53.855 175.865 54.505 175.910 ;
        RECT 39.475 175.525 39.765 175.755 ;
        RECT 44.060 175.510 44.380 175.770 ;
        RECT 44.535 175.525 44.825 175.755 ;
        RECT 46.820 175.710 47.140 175.770 ;
        RECT 47.295 175.710 47.585 175.755 ;
        RECT 46.820 175.570 47.585 175.710 ;
        RECT 39.000 175.370 39.320 175.430 ;
        RECT 36.790 175.230 39.320 175.370 ;
        RECT 29.815 175.185 30.105 175.230 ;
        RECT 31.655 175.185 31.945 175.230 ;
        RECT 35.780 175.170 36.100 175.230 ;
        RECT 39.000 175.170 39.320 175.230 ;
        RECT 43.140 175.170 43.460 175.430 ;
        RECT 26.595 174.845 26.885 175.075 ;
        RECT 44.610 175.030 44.750 175.525 ;
        RECT 46.820 175.510 47.140 175.570 ;
        RECT 47.295 175.525 47.585 175.570 ;
        RECT 50.915 175.550 51.205 175.865 ;
        RECT 56.480 175.850 56.800 176.110 ;
        RECT 64.760 176.050 65.080 176.110 ;
        RECT 66.615 176.050 66.905 176.095 ;
        RECT 67.520 176.050 67.840 176.110 ;
        RECT 58.870 175.910 62.690 176.050 ;
        RECT 58.870 175.770 59.010 175.910 ;
        RECT 51.995 175.710 52.285 175.755 ;
        RECT 55.575 175.710 55.865 175.755 ;
        RECT 57.410 175.710 57.700 175.755 ;
        RECT 51.995 175.570 57.700 175.710 ;
        RECT 51.995 175.525 52.285 175.570 ;
        RECT 55.575 175.525 55.865 175.570 ;
        RECT 57.410 175.525 57.700 175.570 ;
        RECT 58.780 175.510 59.100 175.770 ;
        RECT 62.000 175.510 62.320 175.770 ;
        RECT 62.550 175.755 62.690 175.910 ;
        RECT 64.760 175.910 66.370 176.050 ;
        RECT 64.760 175.850 65.080 175.910 ;
        RECT 62.475 175.710 62.765 175.755 ;
        RECT 64.315 175.710 64.605 175.755 ;
        RECT 62.475 175.570 64.605 175.710 ;
        RECT 62.475 175.525 62.765 175.570 ;
        RECT 64.315 175.525 64.605 175.570 ;
        RECT 65.220 175.710 65.540 175.770 ;
        RECT 66.230 175.755 66.370 175.910 ;
        RECT 66.615 175.910 67.840 176.050 ;
        RECT 80.030 176.050 80.170 176.250 ;
        RECT 80.415 176.250 81.180 176.390 ;
        RECT 80.415 176.205 80.705 176.250 ;
        RECT 80.860 176.190 81.180 176.250 ;
        RECT 84.095 176.390 84.385 176.435 ;
        RECT 87.300 176.390 87.620 176.450 ;
        RECT 84.095 176.250 87.620 176.390 ;
        RECT 84.095 176.205 84.385 176.250 ;
        RECT 87.300 176.190 87.620 176.250 ;
        RECT 91.440 176.390 91.760 176.450 ;
        RECT 91.440 176.250 95.350 176.390 ;
        RECT 91.440 176.190 91.760 176.250 ;
        RECT 86.380 176.050 86.700 176.110 ;
        RECT 87.775 176.050 88.065 176.095 ;
        RECT 80.030 175.910 84.770 176.050 ;
        RECT 66.615 175.865 66.905 175.910 ;
        RECT 67.520 175.850 67.840 175.910 ;
        RECT 65.695 175.710 65.985 175.755 ;
        RECT 65.220 175.570 65.985 175.710 ;
        RECT 65.220 175.510 65.540 175.570 ;
        RECT 65.695 175.525 65.985 175.570 ;
        RECT 66.155 175.525 66.445 175.755 ;
        RECT 67.075 175.525 67.365 175.755 ;
        RECT 70.740 175.710 71.060 175.770 ;
        RECT 71.675 175.710 71.965 175.755 ;
        RECT 70.740 175.570 71.965 175.710 ;
        RECT 50.040 175.370 50.360 175.430 ;
        RECT 57.860 175.370 58.180 175.430 ;
        RECT 50.040 175.230 58.180 175.370 ;
        RECT 62.090 175.370 62.230 175.510 ;
        RECT 64.775 175.370 65.065 175.415 ;
        RECT 67.150 175.370 67.290 175.525 ;
        RECT 70.740 175.510 71.060 175.570 ;
        RECT 71.675 175.525 71.965 175.570 ;
        RECT 72.120 175.510 72.440 175.770 ;
        RECT 72.595 175.525 72.885 175.755 ;
        RECT 73.040 175.710 73.360 175.770 ;
        RECT 73.515 175.710 73.805 175.755 ;
        RECT 73.040 175.570 73.805 175.710 ;
        RECT 62.090 175.230 67.290 175.370 ;
        RECT 72.670 175.370 72.810 175.525 ;
        RECT 73.040 175.510 73.360 175.570 ;
        RECT 73.515 175.525 73.805 175.570 ;
        RECT 76.260 175.510 76.580 175.770 ;
        RECT 79.035 175.710 79.325 175.755 ;
        RECT 79.495 175.710 79.785 175.755 ;
        RECT 79.035 175.570 79.785 175.710 ;
        RECT 79.035 175.525 79.325 175.570 ;
        RECT 79.495 175.525 79.785 175.570 ;
        RECT 81.335 175.710 81.625 175.755 ;
        RECT 83.160 175.710 83.480 175.770 ;
        RECT 81.335 175.570 83.480 175.710 ;
        RECT 84.630 175.710 84.770 175.910 ;
        RECT 86.380 175.910 88.065 176.050 ;
        RECT 86.380 175.850 86.700 175.910 ;
        RECT 87.775 175.865 88.065 175.910 ;
        RECT 88.220 176.050 88.540 176.110 ;
        RECT 88.220 175.910 94.890 176.050 ;
        RECT 88.220 175.850 88.540 175.910 ;
        RECT 89.600 175.710 89.920 175.770 ;
        RECT 84.630 175.570 89.920 175.710 ;
        RECT 81.335 175.525 81.625 175.570 ;
        RECT 83.160 175.510 83.480 175.570 ;
        RECT 89.600 175.510 89.920 175.570 ;
        RECT 90.075 175.525 90.365 175.755 ;
        RECT 79.940 175.370 80.260 175.430 ;
        RECT 72.670 175.230 80.260 175.370 ;
        RECT 50.040 175.170 50.360 175.230 ;
        RECT 57.860 175.170 58.180 175.230 ;
        RECT 64.775 175.185 65.065 175.230 ;
        RECT 79.940 175.170 80.260 175.230 ;
        RECT 85.015 175.370 85.305 175.415 ;
        RECT 85.920 175.370 86.240 175.430 ;
        RECT 90.150 175.370 90.290 175.525 ;
        RECT 90.520 175.510 90.840 175.770 ;
        RECT 91.440 175.510 91.760 175.770 ;
        RECT 93.280 175.725 93.600 175.770 ;
        RECT 94.750 175.755 94.890 175.910 ;
        RECT 93.755 175.725 94.045 175.755 ;
        RECT 93.280 175.585 94.045 175.725 ;
        RECT 93.280 175.510 93.600 175.585 ;
        RECT 93.755 175.525 94.045 175.585 ;
        RECT 94.215 175.525 94.505 175.755 ;
        RECT 94.675 175.525 94.965 175.755 ;
        RECT 95.210 175.710 95.350 176.250 ;
        RECT 95.595 175.710 95.885 175.755 ;
        RECT 96.040 175.710 96.360 175.770 ;
        RECT 95.210 175.570 96.360 175.710 ;
        RECT 95.595 175.525 95.885 175.570 ;
        RECT 92.820 175.370 93.140 175.430 ;
        RECT 94.290 175.370 94.430 175.525 ;
        RECT 96.040 175.510 96.360 175.570 ;
        RECT 96.960 175.510 97.280 175.770 ;
        RECT 97.420 175.510 97.740 175.770 ;
        RECT 97.895 175.525 98.185 175.755 ;
        RECT 99.720 175.710 100.040 175.770 ;
        RECT 107.095 175.710 107.385 175.755 ;
        RECT 99.720 175.570 107.385 175.710 ;
        RECT 97.510 175.370 97.650 175.510 ;
        RECT 85.015 175.230 86.240 175.370 ;
        RECT 85.015 175.185 85.305 175.230 ;
        RECT 85.920 175.170 86.240 175.230 ;
        RECT 89.690 175.230 97.650 175.370 ;
        RECT 43.690 174.890 44.750 175.030 ;
        RECT 51.995 175.030 52.285 175.075 ;
        RECT 55.115 175.030 55.405 175.075 ;
        RECT 57.005 175.030 57.295 175.075 ;
        RECT 51.995 174.890 57.295 175.030 ;
        RECT 43.690 174.750 43.830 174.890 ;
        RECT 51.995 174.845 52.285 174.890 ;
        RECT 55.115 174.845 55.405 174.890 ;
        RECT 57.005 174.845 57.295 174.890 ;
        RECT 67.980 175.030 68.300 175.090 ;
        RECT 89.140 175.030 89.460 175.090 ;
        RECT 89.690 175.030 89.830 175.230 ;
        RECT 92.820 175.170 93.140 175.230 ;
        RECT 67.980 174.890 89.830 175.030 ;
        RECT 93.280 175.030 93.600 175.090 ;
        RECT 94.200 175.030 94.520 175.090 ;
        RECT 97.970 175.030 98.110 175.525 ;
        RECT 99.720 175.510 100.040 175.570 ;
        RECT 107.095 175.525 107.385 175.570 ;
        RECT 93.280 174.890 98.110 175.030 ;
        RECT 67.980 174.830 68.300 174.890 ;
        RECT 89.140 174.830 89.460 174.890 ;
        RECT 93.280 174.830 93.600 174.890 ;
        RECT 94.200 174.830 94.520 174.890 ;
        RECT 25.660 174.490 25.980 174.750 ;
        RECT 34.415 174.690 34.705 174.735 ;
        RECT 35.320 174.690 35.640 174.750 ;
        RECT 34.415 174.550 35.640 174.690 ;
        RECT 34.415 174.505 34.705 174.550 ;
        RECT 35.320 174.490 35.640 174.550 ;
        RECT 38.555 174.690 38.845 174.735 ;
        RECT 39.920 174.690 40.240 174.750 ;
        RECT 38.555 174.550 40.240 174.690 ;
        RECT 38.555 174.505 38.845 174.550 ;
        RECT 39.920 174.490 40.240 174.550 ;
        RECT 42.235 174.690 42.525 174.735 ;
        RECT 43.600 174.690 43.920 174.750 ;
        RECT 42.235 174.550 43.920 174.690 ;
        RECT 42.235 174.505 42.525 174.550 ;
        RECT 43.600 174.490 43.920 174.550 ;
        RECT 61.095 174.690 61.385 174.735 ;
        RECT 62.000 174.690 62.320 174.750 ;
        RECT 61.095 174.550 62.320 174.690 ;
        RECT 61.095 174.505 61.385 174.550 ;
        RECT 62.000 174.490 62.320 174.550 ;
        RECT 63.380 174.690 63.700 174.750 ;
        RECT 67.520 174.690 67.840 174.750 ;
        RECT 63.380 174.550 67.840 174.690 ;
        RECT 63.380 174.490 63.700 174.550 ;
        RECT 67.520 174.490 67.840 174.550 ;
        RECT 70.280 174.490 70.600 174.750 ;
        RECT 86.840 174.690 87.160 174.750 ;
        RECT 88.235 174.690 88.525 174.735 ;
        RECT 86.840 174.550 88.525 174.690 ;
        RECT 86.840 174.490 87.160 174.550 ;
        RECT 88.235 174.505 88.525 174.550 ;
        RECT 91.900 174.690 92.220 174.750 ;
        RECT 92.375 174.690 92.665 174.735 ;
        RECT 91.900 174.550 92.665 174.690 ;
        RECT 91.900 174.490 92.220 174.550 ;
        RECT 92.375 174.505 92.665 174.550 ;
        RECT 94.660 174.690 94.980 174.750 ;
        RECT 99.275 174.690 99.565 174.735 ;
        RECT 94.660 174.550 99.565 174.690 ;
        RECT 94.660 174.490 94.980 174.550 ;
        RECT 99.275 174.505 99.565 174.550 ;
        RECT 108.015 174.690 108.305 174.735 ;
        RECT 109.840 174.690 110.160 174.750 ;
        RECT 108.015 174.550 110.160 174.690 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 108.015 174.505 108.305 174.550 ;
        RECT 109.840 174.490 110.160 174.550 ;
        RECT 11.330 173.870 113.450 174.350 ;
        RECT 45.915 173.670 46.205 173.715 ;
        RECT 49.580 173.670 49.900 173.730 ;
        RECT 63.380 173.670 63.700 173.730 ;
        RECT 45.915 173.530 49.900 173.670 ;
        RECT 45.915 173.485 46.205 173.530 ;
        RECT 49.580 173.470 49.900 173.530 ;
        RECT 50.130 173.530 63.700 173.670 ;
        RECT 25.675 173.330 25.965 173.375 ;
        RECT 28.420 173.330 28.740 173.390 ;
        RECT 25.675 173.190 28.740 173.330 ;
        RECT 25.675 173.145 25.965 173.190 ;
        RECT 28.420 173.130 28.740 173.190 ;
        RECT 28.995 173.330 29.285 173.375 ;
        RECT 32.115 173.330 32.405 173.375 ;
        RECT 34.005 173.330 34.295 173.375 ;
        RECT 28.995 173.190 34.295 173.330 ;
        RECT 28.995 173.145 29.285 173.190 ;
        RECT 32.115 173.145 32.405 173.190 ;
        RECT 34.005 173.145 34.295 173.190 ;
        RECT 36.255 173.145 36.545 173.375 ;
        RECT 37.160 173.330 37.480 173.390 ;
        RECT 41.300 173.330 41.620 173.390 ;
        RECT 46.360 173.330 46.680 173.390 ;
        RECT 50.130 173.330 50.270 173.530 ;
        RECT 63.380 173.470 63.700 173.530 ;
        RECT 86.380 173.470 86.700 173.730 ;
        RECT 89.600 173.670 89.920 173.730 ;
        RECT 93.280 173.670 93.600 173.730 ;
        RECT 89.600 173.530 93.600 173.670 ;
        RECT 89.600 173.470 89.920 173.530 ;
        RECT 93.280 173.470 93.600 173.530 ;
        RECT 99.720 173.470 100.040 173.730 ;
        RECT 37.160 173.190 50.270 173.330 ;
        RECT 53.375 173.330 53.665 173.375 ;
        RECT 56.495 173.330 56.785 173.375 ;
        RECT 58.385 173.330 58.675 173.375 ;
        RECT 53.375 173.190 58.675 173.330 ;
        RECT 33.495 172.990 33.785 173.035 ;
        RECT 36.330 172.990 36.470 173.145 ;
        RECT 37.160 173.130 37.480 173.190 ;
        RECT 33.495 172.850 36.470 172.990 ;
        RECT 39.000 172.990 39.320 173.050 ;
        RECT 39.000 172.850 40.150 172.990 ;
        RECT 33.495 172.805 33.785 172.850 ;
        RECT 39.000 172.790 39.320 172.850 ;
        RECT 22.915 172.465 23.205 172.695 ;
        RECT 22.990 171.970 23.130 172.465 ;
        RECT 25.660 172.310 25.980 172.370 ;
        RECT 27.915 172.355 28.205 172.670 ;
        RECT 28.995 172.650 29.285 172.695 ;
        RECT 32.575 172.650 32.865 172.695 ;
        RECT 34.410 172.650 34.700 172.695 ;
        RECT 28.995 172.510 34.700 172.650 ;
        RECT 28.995 172.465 29.285 172.510 ;
        RECT 32.575 172.465 32.865 172.510 ;
        RECT 34.410 172.465 34.700 172.510 ;
        RECT 34.860 172.450 35.180 172.710 ;
        RECT 35.320 172.650 35.640 172.710 ;
        RECT 37.175 172.650 37.465 172.695 ;
        RECT 35.320 172.510 37.465 172.650 ;
        RECT 35.320 172.450 35.640 172.510 ;
        RECT 37.175 172.465 37.465 172.510 ;
        RECT 38.540 172.450 38.860 172.710 ;
        RECT 40.010 172.695 40.150 172.850 ;
        RECT 40.470 172.695 40.610 173.190 ;
        RECT 41.300 173.130 41.620 173.190 ;
        RECT 46.360 173.130 46.680 173.190 ;
        RECT 53.375 173.145 53.665 173.190 ;
        RECT 56.495 173.145 56.785 173.190 ;
        RECT 58.385 173.145 58.675 173.190 ;
        RECT 80.975 173.330 81.265 173.375 ;
        RECT 84.095 173.330 84.385 173.375 ;
        RECT 85.985 173.330 86.275 173.375 ;
        RECT 80.975 173.190 86.275 173.330 ;
        RECT 86.470 173.330 86.610 173.470 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 105.355 173.330 105.645 173.375 ;
        RECT 108.475 173.330 108.765 173.375 ;
        RECT 110.365 173.330 110.655 173.375 ;
        RECT 86.470 173.190 98.110 173.330 ;
        RECT 80.975 173.145 81.265 173.190 ;
        RECT 84.095 173.145 84.385 173.190 ;
        RECT 85.985 173.145 86.275 173.190 ;
        RECT 43.140 172.790 43.460 173.050 ;
        RECT 43.600 172.790 43.920 173.050 ;
        RECT 46.835 172.990 47.125 173.035 ;
        RECT 44.150 172.850 47.125 172.990 ;
        RECT 39.475 172.465 39.765 172.695 ;
        RECT 39.935 172.465 40.225 172.695 ;
        RECT 40.395 172.465 40.685 172.695 ;
        RECT 43.230 172.650 43.370 172.790 ;
        RECT 44.150 172.650 44.290 172.850 ;
        RECT 46.835 172.805 47.125 172.850 ;
        RECT 47.280 172.990 47.600 173.050 ;
        RECT 54.640 172.990 54.960 173.050 ;
        RECT 47.280 172.850 54.960 172.990 ;
        RECT 47.280 172.790 47.600 172.850 ;
        RECT 54.640 172.790 54.960 172.850 ;
        RECT 56.020 172.990 56.340 173.050 ;
        RECT 57.875 172.990 58.165 173.035 ;
        RECT 56.020 172.850 58.165 172.990 ;
        RECT 56.020 172.790 56.340 172.850 ;
        RECT 57.875 172.805 58.165 172.850 ;
        RECT 62.000 172.990 62.320 173.050 ;
        RECT 72.120 172.990 72.440 173.050 ;
        RECT 78.115 172.990 78.405 173.035 ;
        RECT 85.460 172.990 85.780 173.050 ;
        RECT 96.500 172.990 96.820 173.050 ;
        RECT 62.000 172.850 72.440 172.990 ;
        RECT 62.000 172.790 62.320 172.850 ;
        RECT 43.230 172.510 44.290 172.650 ;
        RECT 27.615 172.310 28.205 172.355 ;
        RECT 30.855 172.310 31.505 172.355 ;
        RECT 25.660 172.170 31.505 172.310 ;
        RECT 39.550 172.310 39.690 172.465 ;
        RECT 45.900 172.450 46.220 172.710 ;
        RECT 45.990 172.310 46.130 172.450 ;
        RECT 48.215 172.310 48.505 172.355 ;
        RECT 39.550 172.170 48.505 172.310 ;
        RECT 25.660 172.110 25.980 172.170 ;
        RECT 27.615 172.125 27.905 172.170 ;
        RECT 30.855 172.125 31.505 172.170 ;
        RECT 48.215 172.125 48.505 172.170 ;
        RECT 48.660 172.310 48.980 172.370 ;
        RECT 52.295 172.355 52.585 172.670 ;
        RECT 53.375 172.650 53.665 172.695 ;
        RECT 56.955 172.650 57.245 172.695 ;
        RECT 58.790 172.650 59.080 172.695 ;
        RECT 53.375 172.510 59.080 172.650 ;
        RECT 53.375 172.465 53.665 172.510 ;
        RECT 56.955 172.465 57.245 172.510 ;
        RECT 58.790 172.465 59.080 172.510 ;
        RECT 59.255 172.465 59.545 172.695 ;
        RECT 51.995 172.310 52.585 172.355 ;
        RECT 54.180 172.310 54.500 172.370 ;
        RECT 55.235 172.310 55.885 172.355 ;
        RECT 48.660 172.170 51.190 172.310 ;
        RECT 48.660 172.110 48.980 172.170 ;
        RECT 26.135 171.970 26.425 172.015 ;
        RECT 32.100 171.970 32.420 172.030 ;
        RECT 22.990 171.830 32.420 171.970 ;
        RECT 26.135 171.785 26.425 171.830 ;
        RECT 32.100 171.770 32.420 171.830 ;
        RECT 41.760 171.770 42.080 172.030 ;
        RECT 44.075 171.970 44.365 172.015 ;
        RECT 45.900 171.970 46.220 172.030 ;
        RECT 47.755 171.970 48.045 172.015 ;
        RECT 44.075 171.830 48.045 171.970 ;
        RECT 44.075 171.785 44.365 171.830 ;
        RECT 45.900 171.770 46.220 171.830 ;
        RECT 47.755 171.785 48.045 171.830 ;
        RECT 50.040 171.770 50.360 172.030 ;
        RECT 50.500 171.770 50.820 172.030 ;
        RECT 51.050 171.970 51.190 172.170 ;
        RECT 51.995 172.170 55.885 172.310 ;
        RECT 51.995 172.125 52.285 172.170 ;
        RECT 54.180 172.110 54.500 172.170 ;
        RECT 55.235 172.125 55.885 172.170 ;
        RECT 57.860 172.310 58.180 172.370 ;
        RECT 59.330 172.310 59.470 172.465 ;
        RECT 64.760 172.450 65.080 172.710 ;
        RECT 65.695 172.465 65.985 172.695 ;
        RECT 65.770 172.310 65.910 172.465 ;
        RECT 66.600 172.450 66.920 172.710 ;
        RECT 67.150 172.695 67.290 172.850 ;
        RECT 67.075 172.465 67.365 172.695 ;
        RECT 67.520 172.650 67.840 172.710 ;
        RECT 70.740 172.650 71.060 172.710 ;
        RECT 71.290 172.695 71.430 172.850 ;
        RECT 72.120 172.790 72.440 172.850 ;
        RECT 73.590 172.850 76.490 172.990 ;
        RECT 67.520 172.510 71.060 172.650 ;
        RECT 67.520 172.450 67.840 172.510 ;
        RECT 70.740 172.450 71.060 172.510 ;
        RECT 71.215 172.465 71.505 172.695 ;
        RECT 71.660 172.450 71.980 172.710 ;
        RECT 73.590 172.695 73.730 172.850 ;
        RECT 72.595 172.465 72.885 172.695 ;
        RECT 73.515 172.465 73.805 172.695 ;
        RECT 72.670 172.310 72.810 172.465 ;
        RECT 74.880 172.450 75.200 172.710 ;
        RECT 76.350 172.695 76.490 172.850 ;
        RECT 78.115 172.850 85.780 172.990 ;
        RECT 78.115 172.805 78.405 172.850 ;
        RECT 85.460 172.790 85.780 172.850 ;
        RECT 87.850 172.850 90.290 172.990 ;
        RECT 76.275 172.650 76.565 172.695 ;
        RECT 77.640 172.650 77.960 172.710 ;
        RECT 76.275 172.510 77.960 172.650 ;
        RECT 76.275 172.465 76.565 172.510 ;
        RECT 77.640 172.450 77.960 172.510 ;
        RECT 73.040 172.310 73.360 172.370 ;
        RECT 79.895 172.355 80.185 172.670 ;
        RECT 80.975 172.650 81.265 172.695 ;
        RECT 84.555 172.650 84.845 172.695 ;
        RECT 86.390 172.650 86.680 172.695 ;
        RECT 80.975 172.510 86.680 172.650 ;
        RECT 80.975 172.465 81.265 172.510 ;
        RECT 84.555 172.465 84.845 172.510 ;
        RECT 86.390 172.465 86.680 172.510 ;
        RECT 86.855 172.465 87.145 172.695 ;
        RECT 87.300 172.650 87.620 172.710 ;
        RECT 87.850 172.695 87.990 172.850 ;
        RECT 87.775 172.650 88.065 172.695 ;
        RECT 87.300 172.510 88.065 172.650 ;
        RECT 57.860 172.170 59.470 172.310 ;
        RECT 63.930 172.170 73.360 172.310 ;
        RECT 57.860 172.110 58.180 172.170 ;
        RECT 63.930 172.015 64.070 172.170 ;
        RECT 73.040 172.110 73.360 172.170 ;
        RECT 73.975 172.310 74.265 172.355 ;
        RECT 79.595 172.310 80.185 172.355 ;
        RECT 82.835 172.310 83.485 172.355 ;
        RECT 73.975 172.170 83.485 172.310 ;
        RECT 73.975 172.125 74.265 172.170 ;
        RECT 79.595 172.125 79.885 172.170 ;
        RECT 82.835 172.125 83.485 172.170 ;
        RECT 85.460 172.110 85.780 172.370 ;
        RECT 86.930 172.310 87.070 172.465 ;
        RECT 87.300 172.450 87.620 172.510 ;
        RECT 87.775 172.465 88.065 172.510 ;
        RECT 88.695 172.465 88.985 172.695 ;
        RECT 86.470 172.170 87.070 172.310 ;
        RECT 88.770 172.310 88.910 172.465 ;
        RECT 89.140 172.450 89.460 172.710 ;
        RECT 89.600 172.450 89.920 172.710 ;
        RECT 90.150 172.650 90.290 172.850 ;
        RECT 92.450 172.850 96.820 172.990 ;
        RECT 91.440 172.650 91.760 172.710 ;
        RECT 92.450 172.695 92.590 172.850 ;
        RECT 96.500 172.790 96.820 172.850 ;
        RECT 96.975 172.990 97.265 173.035 ;
        RECT 97.420 172.990 97.740 173.050 ;
        RECT 96.975 172.850 97.740 172.990 ;
        RECT 96.975 172.805 97.265 172.850 ;
        RECT 97.420 172.790 97.740 172.850 ;
        RECT 90.150 172.510 91.760 172.650 ;
        RECT 91.440 172.450 91.760 172.510 ;
        RECT 92.375 172.465 92.665 172.695 ;
        RECT 92.820 172.450 93.140 172.710 ;
        RECT 93.280 172.450 93.600 172.710 ;
        RECT 97.970 172.695 98.110 173.190 ;
        RECT 105.355 173.190 110.655 173.330 ;
        RECT 105.355 173.145 105.645 173.190 ;
        RECT 108.475 173.145 108.765 173.190 ;
        RECT 110.365 173.145 110.655 173.190 ;
        RECT 109.840 172.790 110.160 173.050 ;
        RECT 97.895 172.465 98.185 172.695 ;
        RECT 101.100 172.450 101.420 172.710 ;
        RECT 99.260 172.310 99.580 172.370 ;
        RECT 104.275 172.355 104.565 172.670 ;
        RECT 105.355 172.650 105.645 172.695 ;
        RECT 108.935 172.650 109.225 172.695 ;
        RECT 110.770 172.650 111.060 172.695 ;
        RECT 105.355 172.510 111.060 172.650 ;
        RECT 105.355 172.465 105.645 172.510 ;
        RECT 108.935 172.465 109.225 172.510 ;
        RECT 110.770 172.465 111.060 172.510 ;
        RECT 111.235 172.650 111.525 172.695 ;
        RECT 111.680 172.650 112.000 172.710 ;
        RECT 111.235 172.510 112.000 172.650 ;
        RECT 111.235 172.465 111.525 172.510 ;
        RECT 111.680 172.450 112.000 172.510 ;
        RECT 88.770 172.170 99.580 172.310 ;
        RECT 63.855 171.970 64.145 172.015 ;
        RECT 51.050 171.830 64.145 171.970 ;
        RECT 63.855 171.785 64.145 171.830 ;
        RECT 68.900 171.770 69.220 172.030 ;
        RECT 69.360 171.770 69.680 172.030 ;
        RECT 82.240 171.970 82.560 172.030 ;
        RECT 86.470 171.970 86.610 172.170 ;
        RECT 99.260 172.110 99.580 172.170 ;
        RECT 101.575 172.310 101.865 172.355 ;
        RECT 103.975 172.310 104.565 172.355 ;
        RECT 107.215 172.310 107.865 172.355 ;
        RECT 101.575 172.170 107.865 172.310 ;
        RECT 101.575 172.125 101.865 172.170 ;
        RECT 103.975 172.125 104.265 172.170 ;
        RECT 107.215 172.125 107.865 172.170 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 82.240 171.830 86.610 171.970 ;
        RECT 82.240 171.770 82.560 171.830 ;
        RECT 90.980 171.770 91.300 172.030 ;
        RECT 94.675 171.970 94.965 172.015 ;
        RECT 96.040 171.970 96.360 172.030 ;
        RECT 94.675 171.830 96.360 171.970 ;
        RECT 94.675 171.785 94.965 171.830 ;
        RECT 96.040 171.770 96.360 171.830 ;
        RECT 97.420 171.770 97.740 172.030 ;
        RECT 100.640 171.970 100.960 172.030 ;
        RECT 102.495 171.970 102.785 172.015 ;
        RECT 100.640 171.830 102.785 171.970 ;
        RECT 100.640 171.770 100.960 171.830 ;
        RECT 102.495 171.785 102.785 171.830 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 11.330 171.150 113.450 171.630 ;
        RECT 30.720 170.950 31.040 171.010 ;
        RECT 31.640 170.950 31.960 171.010 ;
        RECT 30.720 170.810 31.960 170.950 ;
        RECT 30.720 170.750 31.040 170.810 ;
        RECT 31.640 170.750 31.960 170.810 ;
        RECT 32.100 170.950 32.420 171.010 ;
        RECT 38.540 170.950 38.860 171.010 ;
        RECT 42.680 170.950 43.000 171.010 ;
        RECT 48.660 170.950 48.980 171.010 ;
        RECT 32.100 170.810 32.790 170.950 ;
        RECT 32.100 170.750 32.420 170.810 ;
        RECT 30.260 170.610 30.580 170.670 ;
        RECT 28.050 170.470 31.870 170.610 ;
        RECT 24.755 170.270 25.045 170.315 ;
        RECT 26.580 170.270 26.900 170.330 ;
        RECT 28.050 170.315 28.190 170.470 ;
        RECT 30.260 170.410 30.580 170.470 ;
        RECT 24.755 170.130 26.900 170.270 ;
        RECT 24.755 170.085 25.045 170.130 ;
        RECT 26.580 170.070 26.900 170.130 ;
        RECT 27.975 170.085 28.265 170.315 ;
        RECT 28.435 170.085 28.725 170.315 ;
        RECT 24.295 169.930 24.585 169.975 ;
        RECT 28.510 169.930 28.650 170.085 ;
        RECT 28.880 170.070 29.200 170.330 ;
        RECT 29.800 170.270 30.120 170.330 ;
        RECT 31.730 170.315 31.870 170.470 ;
        RECT 29.800 170.130 31.410 170.270 ;
        RECT 29.800 170.070 30.120 170.130 ;
        RECT 30.720 169.930 31.040 169.990 ;
        RECT 24.295 169.790 28.190 169.930 ;
        RECT 28.510 169.790 31.040 169.930 ;
        RECT 31.270 169.930 31.410 170.130 ;
        RECT 31.655 170.085 31.945 170.315 ;
        RECT 32.100 170.070 32.420 170.330 ;
        RECT 32.650 170.315 32.790 170.810 ;
        RECT 38.540 170.810 48.980 170.950 ;
        RECT 38.540 170.750 38.860 170.810 ;
        RECT 42.680 170.750 43.000 170.810 ;
        RECT 41.300 170.610 41.620 170.670 ;
        RECT 39.090 170.470 42.910 170.610 ;
        RECT 39.090 170.315 39.230 170.470 ;
        RECT 41.300 170.410 41.620 170.470 ;
        RECT 32.575 170.085 32.865 170.315 ;
        RECT 33.495 170.085 33.785 170.315 ;
        RECT 39.015 170.085 39.305 170.315 ;
        RECT 33.570 169.930 33.710 170.085 ;
        RECT 39.460 170.070 39.780 170.330 ;
        RECT 39.935 170.260 40.225 170.315 ;
        RECT 40.380 170.260 40.700 170.330 ;
        RECT 39.935 170.120 40.700 170.260 ;
        RECT 39.935 170.085 40.225 170.120 ;
        RECT 40.380 170.070 40.700 170.120 ;
        RECT 40.855 170.270 41.145 170.315 ;
        RECT 42.220 170.270 42.540 170.330 ;
        RECT 42.770 170.315 42.910 170.470 ;
        RECT 40.855 170.130 42.540 170.270 ;
        RECT 40.855 170.085 41.145 170.130 ;
        RECT 42.220 170.070 42.540 170.130 ;
        RECT 42.695 170.085 42.985 170.315 ;
        RECT 43.155 170.085 43.445 170.315 ;
        RECT 43.615 170.270 43.905 170.315 ;
        RECT 44.060 170.270 44.380 170.330 ;
        RECT 43.615 170.130 44.380 170.270 ;
        RECT 43.615 170.085 43.905 170.130 ;
        RECT 38.080 169.930 38.400 169.990 ;
        RECT 31.270 169.790 38.400 169.930 ;
        RECT 39.550 169.930 39.690 170.070 ;
        RECT 43.230 169.930 43.370 170.085 ;
        RECT 44.060 170.070 44.380 170.130 ;
        RECT 44.535 170.270 44.825 170.315 ;
        RECT 45.070 170.270 45.210 170.810 ;
        RECT 48.660 170.750 48.980 170.810 ;
        RECT 54.180 170.750 54.500 171.010 ;
        RECT 56.020 170.750 56.340 171.010 ;
        RECT 62.920 170.950 63.240 171.010 ;
        RECT 74.880 170.950 75.200 171.010 ;
        RECT 62.920 170.810 75.200 170.950 ;
        RECT 62.920 170.750 63.240 170.810 ;
        RECT 74.880 170.750 75.200 170.810 ;
        RECT 82.240 170.750 82.560 171.010 ;
        RECT 101.100 170.950 101.420 171.010 ;
        RECT 106.620 170.950 106.940 171.010 ;
        RECT 86.930 170.810 93.970 170.950 ;
        RECT 50.500 170.610 50.820 170.670 ;
        RECT 47.370 170.470 50.820 170.610 ;
        RECT 44.535 170.130 45.210 170.270 ;
        RECT 44.535 170.085 44.825 170.130 ;
        RECT 46.360 170.070 46.680 170.330 ;
        RECT 47.370 170.315 47.510 170.470 ;
        RECT 50.500 170.410 50.820 170.470 ;
        RECT 52.355 170.610 52.645 170.655 ;
        RECT 61.080 170.610 61.400 170.670 ;
        RECT 63.380 170.610 63.700 170.670 ;
        RECT 79.480 170.610 79.800 170.670 ;
        RECT 52.355 170.470 55.330 170.610 ;
        RECT 52.355 170.425 52.645 170.470 ;
        RECT 46.835 170.085 47.125 170.315 ;
        RECT 47.295 170.085 47.585 170.315 ;
        RECT 48.215 170.270 48.505 170.315 ;
        RECT 48.660 170.270 48.980 170.330 ;
        RECT 48.215 170.130 48.980 170.270 ;
        RECT 48.215 170.085 48.505 170.130 ;
        RECT 46.910 169.930 47.050 170.085 ;
        RECT 48.660 170.070 48.980 170.130 ;
        RECT 49.595 170.270 49.885 170.315 ;
        RECT 50.040 170.270 50.360 170.330 ;
        RECT 49.595 170.130 50.360 170.270 ;
        RECT 49.595 170.085 49.885 170.130 ;
        RECT 50.040 170.070 50.360 170.130 ;
        RECT 54.640 170.070 54.960 170.330 ;
        RECT 55.190 170.315 55.330 170.470 ;
        RECT 61.080 170.470 63.700 170.610 ;
        RECT 61.080 170.410 61.400 170.470 ;
        RECT 63.380 170.410 63.700 170.470 ;
        RECT 72.670 170.470 79.800 170.610 ;
        RECT 55.115 170.085 55.405 170.315 ;
        RECT 60.160 170.270 60.480 170.330 ;
        RECT 64.315 170.270 64.605 170.315 ;
        RECT 64.760 170.270 65.080 170.330 ;
        RECT 65.680 170.270 66.000 170.330 ;
        RECT 60.160 170.130 66.000 170.270 ;
        RECT 60.160 170.070 60.480 170.130 ;
        RECT 64.315 170.085 64.605 170.130 ;
        RECT 64.760 170.070 65.080 170.130 ;
        RECT 65.680 170.070 66.000 170.130 ;
        RECT 70.740 170.270 71.060 170.330 ;
        RECT 71.675 170.270 71.965 170.315 ;
        RECT 70.740 170.130 71.965 170.270 ;
        RECT 70.740 170.070 71.060 170.130 ;
        RECT 71.675 170.085 71.965 170.130 ;
        RECT 72.120 170.070 72.440 170.330 ;
        RECT 72.670 170.315 72.810 170.470 ;
        RECT 79.480 170.410 79.800 170.470 ;
        RECT 72.595 170.085 72.885 170.315 ;
        RECT 73.040 170.270 73.360 170.330 ;
        RECT 73.515 170.270 73.805 170.315 ;
        RECT 73.040 170.130 73.805 170.270 ;
        RECT 73.040 170.070 73.360 170.130 ;
        RECT 73.515 170.085 73.805 170.130 ;
        RECT 75.800 170.070 76.120 170.330 ;
        RECT 77.640 170.270 77.960 170.330 ;
        RECT 84.080 170.270 84.400 170.330 ;
        RECT 86.930 170.315 87.070 170.810 ;
        RECT 87.315 170.610 87.605 170.655 ;
        RECT 89.715 170.610 90.005 170.655 ;
        RECT 92.955 170.610 93.605 170.655 ;
        RECT 87.315 170.470 93.605 170.610 ;
        RECT 93.830 170.610 93.970 170.810 ;
        RECT 101.100 170.810 106.940 170.950 ;
        RECT 101.100 170.750 101.420 170.810 ;
        RECT 101.650 170.610 101.790 170.810 ;
        RECT 106.620 170.750 106.940 170.810 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 107.080 170.655 107.400 170.670 ;
        RECT 93.830 170.470 101.790 170.610 ;
        RECT 87.315 170.425 87.605 170.470 ;
        RECT 89.715 170.425 90.305 170.470 ;
        RECT 92.955 170.425 93.605 170.470 ;
        RECT 86.855 170.270 87.145 170.315 ;
        RECT 77.640 170.130 87.145 170.270 ;
        RECT 77.640 170.070 77.960 170.130 ;
        RECT 84.080 170.070 84.400 170.130 ;
        RECT 86.855 170.085 87.145 170.130 ;
        RECT 90.015 170.110 90.305 170.425 ;
        RECT 91.095 170.270 91.385 170.315 ;
        RECT 94.675 170.270 94.965 170.315 ;
        RECT 96.510 170.270 96.800 170.315 ;
        RECT 91.095 170.130 96.800 170.270 ;
        RECT 91.095 170.085 91.385 170.130 ;
        RECT 94.675 170.085 94.965 170.130 ;
        RECT 96.510 170.085 96.800 170.130 ;
        RECT 97.880 170.270 98.200 170.330 ;
        RECT 101.650 170.315 101.790 170.470 ;
        RECT 103.975 170.610 104.265 170.655 ;
        RECT 107.080 170.610 107.865 170.655 ;
        RECT 103.975 170.470 107.865 170.610 ;
        RECT 103.975 170.425 104.565 170.470 ;
        RECT 98.355 170.270 98.645 170.315 ;
        RECT 97.880 170.130 98.645 170.270 ;
        RECT 97.880 170.070 98.200 170.130 ;
        RECT 98.355 170.085 98.645 170.130 ;
        RECT 101.575 170.085 101.865 170.315 ;
        RECT 104.275 170.110 104.565 170.425 ;
        RECT 107.080 170.425 107.865 170.470 ;
        RECT 107.080 170.410 107.400 170.425 ;
        RECT 109.840 170.410 110.160 170.670 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 105.355 170.270 105.645 170.315 ;
        RECT 108.935 170.270 109.225 170.315 ;
        RECT 110.770 170.270 111.060 170.315 ;
        RECT 105.355 170.130 111.060 170.270 ;
        RECT 105.355 170.085 105.645 170.130 ;
        RECT 108.935 170.085 109.225 170.130 ;
        RECT 110.770 170.085 111.060 170.130 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 62.000 169.930 62.320 169.990 ;
        RECT 39.550 169.790 62.320 169.930 ;
        RECT 24.295 169.745 24.585 169.790 ;
        RECT 26.120 169.250 26.440 169.310 ;
        RECT 26.595 169.250 26.885 169.295 ;
        RECT 26.120 169.110 26.885 169.250 ;
        RECT 28.050 169.250 28.190 169.790 ;
        RECT 30.720 169.730 31.040 169.790 ;
        RECT 38.080 169.730 38.400 169.790 ;
        RECT 62.000 169.730 62.320 169.790 ;
        RECT 95.595 169.930 95.885 169.975 ;
        RECT 96.960 169.930 97.280 169.990 ;
        RECT 111.235 169.930 111.525 169.975 ;
        RECT 111.680 169.930 112.000 169.990 ;
        RECT 95.595 169.790 96.730 169.930 ;
        RECT 95.595 169.745 95.885 169.790 ;
        RECT 63.395 169.590 63.685 169.635 ;
        RECT 87.300 169.590 87.620 169.650 ;
        RECT 40.470 169.450 87.620 169.590 ;
        RECT 29.800 169.250 30.120 169.310 ;
        RECT 28.050 169.110 30.120 169.250 ;
        RECT 26.120 169.050 26.440 169.110 ;
        RECT 26.595 169.065 26.885 169.110 ;
        RECT 29.800 169.050 30.120 169.110 ;
        RECT 30.275 169.250 30.565 169.295 ;
        RECT 30.720 169.250 31.040 169.310 ;
        RECT 30.275 169.110 31.040 169.250 ;
        RECT 30.275 169.065 30.565 169.110 ;
        RECT 30.720 169.050 31.040 169.110 ;
        RECT 31.640 169.250 31.960 169.310 ;
        RECT 37.635 169.250 37.925 169.295 ;
        RECT 31.640 169.110 37.925 169.250 ;
        RECT 31.640 169.050 31.960 169.110 ;
        RECT 37.635 169.065 37.925 169.110 ;
        RECT 38.080 169.250 38.400 169.310 ;
        RECT 40.470 169.250 40.610 169.450 ;
        RECT 63.395 169.405 63.685 169.450 ;
        RECT 87.300 169.390 87.620 169.450 ;
        RECT 91.095 169.590 91.385 169.635 ;
        RECT 94.215 169.590 94.505 169.635 ;
        RECT 96.105 169.590 96.395 169.635 ;
        RECT 91.095 169.450 96.395 169.590 ;
        RECT 96.590 169.590 96.730 169.790 ;
        RECT 96.960 169.790 112.000 169.930 ;
        RECT 96.960 169.730 97.280 169.790 ;
        RECT 111.235 169.745 111.525 169.790 ;
        RECT 111.680 169.730 112.000 169.790 ;
        RECT 97.435 169.590 97.725 169.635 ;
        RECT 96.590 169.450 97.725 169.590 ;
        RECT 91.095 169.405 91.385 169.450 ;
        RECT 94.215 169.405 94.505 169.450 ;
        RECT 96.105 169.405 96.395 169.450 ;
        RECT 97.435 169.405 97.725 169.450 ;
        RECT 105.355 169.590 105.645 169.635 ;
        RECT 108.475 169.590 108.765 169.635 ;
        RECT 110.365 169.590 110.655 169.635 ;
        RECT 105.355 169.450 110.655 169.590 ;
        RECT 105.355 169.405 105.645 169.450 ;
        RECT 108.475 169.405 108.765 169.450 ;
        RECT 110.365 169.405 110.655 169.450 ;
        RECT 38.080 169.110 40.610 169.250 ;
        RECT 38.080 169.050 38.400 169.110 ;
        RECT 41.300 169.050 41.620 169.310 ;
        RECT 44.980 169.050 45.300 169.310 ;
        RECT 55.560 169.250 55.880 169.310 ;
        RECT 56.480 169.250 56.800 169.310 ;
        RECT 62.920 169.250 63.240 169.310 ;
        RECT 55.560 169.110 63.240 169.250 ;
        RECT 55.560 169.050 55.880 169.110 ;
        RECT 56.480 169.050 56.800 169.110 ;
        RECT 62.920 169.050 63.240 169.110 ;
        RECT 65.220 169.250 65.540 169.310 ;
        RECT 70.295 169.250 70.585 169.295 ;
        RECT 65.220 169.110 70.585 169.250 ;
        RECT 65.220 169.050 65.540 169.110 ;
        RECT 70.295 169.065 70.585 169.110 ;
        RECT 88.220 169.050 88.540 169.310 ;
        RECT 101.100 169.050 101.420 169.310 ;
        RECT 102.020 169.250 102.340 169.310 ;
        RECT 102.495 169.250 102.785 169.295 ;
        RECT 102.020 169.110 102.785 169.250 ;
        RECT 102.020 169.050 102.340 169.110 ;
        RECT 102.495 169.065 102.785 169.110 ;
        RECT 11.330 168.430 113.450 168.910 ;
        RECT 24.370 168.090 41.070 168.230 ;
        RECT 18.780 167.890 19.070 167.935 ;
        RECT 20.640 167.890 20.930 167.935 ;
        RECT 23.420 167.890 23.710 167.935 ;
        RECT 18.780 167.750 23.710 167.890 ;
        RECT 18.780 167.705 19.070 167.750 ;
        RECT 20.640 167.705 20.930 167.750 ;
        RECT 23.420 167.705 23.710 167.750 ;
        RECT 24.370 167.550 24.510 168.090 ;
        RECT 17.010 167.410 24.510 167.550 ;
        RECT 25.200 167.550 25.520 167.610 ;
        RECT 27.285 167.550 27.575 167.595 ;
        RECT 36.240 167.550 36.560 167.610 ;
        RECT 25.200 167.410 27.575 167.550 ;
        RECT 13.255 167.210 13.545 167.255 ;
        RECT 13.700 167.210 14.020 167.270 ;
        RECT 13.255 167.070 14.020 167.210 ;
        RECT 13.255 167.025 13.545 167.070 ;
        RECT 13.700 167.010 14.020 167.070 ;
        RECT 14.160 167.210 14.480 167.270 ;
        RECT 17.010 167.255 17.150 167.410 ;
        RECT 25.200 167.350 25.520 167.410 ;
        RECT 27.285 167.365 27.575 167.410 ;
        RECT 33.570 167.410 36.560 167.550 ;
        RECT 40.930 167.550 41.070 168.090 ;
        RECT 45.900 168.030 46.220 168.290 ;
        RECT 60.710 168.090 76.490 168.230 ;
        RECT 43.140 167.890 43.460 167.950 ;
        RECT 44.060 167.890 44.380 167.950 ;
        RECT 60.175 167.890 60.465 167.935 ;
        RECT 43.140 167.750 60.465 167.890 ;
        RECT 43.140 167.690 43.460 167.750 ;
        RECT 44.060 167.690 44.380 167.750 ;
        RECT 60.175 167.705 60.465 167.750 ;
        RECT 46.360 167.550 46.680 167.610 ;
        RECT 49.135 167.550 49.425 167.595 ;
        RECT 50.500 167.550 50.820 167.610 ;
        RECT 40.930 167.410 48.430 167.550 ;
        RECT 14.635 167.210 14.925 167.255 ;
        RECT 16.935 167.210 17.225 167.255 ;
        RECT 14.160 167.070 17.225 167.210 ;
        RECT 14.160 167.010 14.480 167.070 ;
        RECT 14.635 167.025 14.925 167.070 ;
        RECT 16.935 167.025 17.225 167.070 ;
        RECT 18.315 167.210 18.605 167.255 ;
        RECT 19.680 167.210 20.000 167.270 ;
        RECT 18.315 167.070 20.000 167.210 ;
        RECT 18.315 167.025 18.605 167.070 ;
        RECT 19.680 167.010 20.000 167.070 ;
        RECT 20.140 167.010 20.460 167.270 ;
        RECT 33.570 167.255 33.710 167.410 ;
        RECT 36.240 167.350 36.560 167.410 ;
        RECT 46.360 167.350 46.680 167.410 ;
        RECT 23.420 167.210 23.710 167.255 ;
        RECT 21.175 167.070 23.710 167.210 ;
        RECT 15.080 166.670 15.400 166.930 ;
        RECT 21.175 166.915 21.390 167.070 ;
        RECT 23.420 167.025 23.710 167.070 ;
        RECT 33.495 167.025 33.785 167.255 ;
        RECT 33.955 167.025 34.245 167.255 ;
        RECT 34.415 167.025 34.705 167.255 ;
        RECT 35.395 167.210 35.685 167.255 ;
        RECT 38.080 167.210 38.400 167.270 ;
        RECT 35.395 167.070 38.400 167.210 ;
        RECT 35.395 167.025 35.685 167.070 ;
        RECT 19.240 166.870 19.530 166.915 ;
        RECT 21.100 166.870 21.390 166.915 ;
        RECT 22.020 166.870 22.310 166.915 ;
        RECT 25.280 166.870 25.570 166.915 ;
        RECT 19.240 166.730 21.390 166.870 ;
        RECT 19.240 166.685 19.530 166.730 ;
        RECT 21.100 166.685 21.390 166.730 ;
        RECT 21.610 166.730 25.570 166.870 ;
        RECT 14.175 166.530 14.465 166.575 ;
        RECT 14.620 166.530 14.940 166.590 ;
        RECT 14.175 166.390 14.940 166.530 ;
        RECT 14.175 166.345 14.465 166.390 ;
        RECT 14.620 166.330 14.940 166.390 ;
        RECT 17.395 166.530 17.685 166.575 ;
        RECT 21.610 166.530 21.750 166.730 ;
        RECT 22.020 166.685 22.310 166.730 ;
        RECT 25.280 166.685 25.570 166.730 ;
        RECT 27.040 166.870 27.360 166.930 ;
        RECT 31.180 166.870 31.500 166.930 ;
        RECT 32.115 166.870 32.405 166.915 ;
        RECT 27.040 166.730 30.950 166.870 ;
        RECT 27.040 166.670 27.360 166.730 ;
        RECT 17.395 166.390 21.750 166.530 ;
        RECT 30.810 166.530 30.950 166.730 ;
        RECT 31.180 166.730 32.405 166.870 ;
        RECT 31.180 166.670 31.500 166.730 ;
        RECT 32.115 166.685 32.405 166.730 ;
        RECT 32.560 166.870 32.880 166.930 ;
        RECT 34.030 166.870 34.170 167.025 ;
        RECT 32.560 166.730 34.170 166.870 ;
        RECT 32.560 166.670 32.880 166.730 ;
        RECT 34.490 166.530 34.630 167.025 ;
        RECT 38.080 167.010 38.400 167.070 ;
        RECT 38.555 167.210 38.845 167.255 ;
        RECT 48.290 167.210 48.430 167.410 ;
        RECT 49.135 167.410 50.820 167.550 ;
        RECT 49.135 167.365 49.425 167.410 ;
        RECT 50.500 167.350 50.820 167.410 ;
        RECT 50.960 167.550 51.280 167.610 ;
        RECT 55.575 167.550 55.865 167.595 ;
        RECT 60.710 167.550 60.850 168.090 ;
        RECT 70.295 167.705 70.585 167.935 ;
        RECT 71.220 167.890 71.510 167.935 ;
        RECT 73.080 167.890 73.370 167.935 ;
        RECT 75.860 167.890 76.150 167.935 ;
        RECT 71.220 167.750 76.150 167.890 ;
        RECT 76.350 167.890 76.490 168.090 ;
        RECT 85.460 168.030 85.780 168.290 ;
        RECT 86.010 168.090 105.930 168.230 ;
        RECT 86.010 167.890 86.150 168.090 ;
        RECT 76.350 167.750 86.150 167.890 ;
        RECT 100.295 167.890 100.585 167.935 ;
        RECT 103.415 167.890 103.705 167.935 ;
        RECT 105.305 167.890 105.595 167.935 ;
        RECT 100.295 167.750 105.595 167.890 ;
        RECT 105.790 167.890 105.930 168.090 ;
        RECT 107.080 168.030 107.400 168.290 ;
        RECT 109.840 168.030 110.160 168.290 ;
        RECT 107.540 167.890 107.860 167.950 ;
        RECT 108.015 167.890 108.305 167.935 ;
        RECT 105.790 167.750 108.305 167.890 ;
        RECT 71.220 167.705 71.510 167.750 ;
        RECT 73.080 167.705 73.370 167.750 ;
        RECT 75.860 167.705 76.150 167.750 ;
        RECT 100.295 167.705 100.585 167.750 ;
        RECT 103.415 167.705 103.705 167.750 ;
        RECT 105.305 167.705 105.595 167.750 ;
        RECT 50.960 167.410 55.865 167.550 ;
        RECT 50.960 167.350 51.280 167.410 ;
        RECT 55.575 167.365 55.865 167.410 ;
        RECT 59.330 167.410 60.850 167.550 ;
        RECT 52.815 167.210 53.105 167.255 ;
        RECT 38.555 167.070 47.970 167.210 ;
        RECT 48.290 167.070 53.105 167.210 ;
        RECT 38.555 167.025 38.845 167.070 ;
        RECT 36.715 166.870 37.005 166.915 ;
        RECT 39.000 166.870 39.320 166.930 ;
        RECT 36.715 166.730 39.320 166.870 ;
        RECT 36.715 166.685 37.005 166.730 ;
        RECT 39.000 166.670 39.320 166.730 ;
        RECT 44.075 166.685 44.365 166.915 ;
        RECT 47.830 166.870 47.970 167.070 ;
        RECT 52.815 167.025 53.105 167.070 ;
        RECT 54.195 167.210 54.485 167.255 ;
        RECT 55.100 167.210 55.420 167.270 ;
        RECT 57.010 167.210 57.300 167.255 ;
        RECT 59.330 167.210 59.470 167.410 ;
        RECT 63.380 167.350 63.700 167.610 ;
        RECT 64.300 167.350 64.620 167.610 ;
        RECT 70.370 167.550 70.510 167.705 ;
        RECT 107.540 167.690 107.860 167.750 ;
        RECT 108.015 167.705 108.305 167.750 ;
        RECT 72.595 167.550 72.885 167.595 ;
        RECT 78.560 167.550 78.880 167.610 ;
        RECT 82.240 167.550 82.560 167.610 ;
        RECT 70.370 167.410 72.885 167.550 ;
        RECT 72.595 167.365 72.885 167.410 ;
        RECT 73.130 167.410 82.560 167.550 ;
        RECT 54.195 167.195 56.710 167.210 ;
        RECT 57.010 167.195 59.470 167.210 ;
        RECT 54.195 167.070 59.470 167.195 ;
        RECT 60.160 167.210 60.480 167.270 ;
        RECT 61.095 167.210 61.385 167.255 ;
        RECT 60.160 167.070 61.385 167.210 ;
        RECT 54.195 167.025 54.485 167.070 ;
        RECT 55.100 167.010 55.420 167.070 ;
        RECT 56.570 167.055 57.300 167.070 ;
        RECT 57.010 167.025 57.300 167.055 ;
        RECT 60.160 167.010 60.480 167.070 ;
        RECT 61.095 167.025 61.385 167.070 ;
        RECT 61.540 167.210 61.860 167.270 ;
        RECT 62.935 167.210 63.225 167.255 ;
        RECT 61.540 167.070 63.225 167.210 ;
        RECT 61.540 167.010 61.860 167.070 ;
        RECT 62.935 167.025 63.225 167.070 ;
        RECT 64.775 167.210 65.065 167.255 ;
        RECT 65.680 167.210 66.000 167.270 ;
        RECT 64.775 167.070 66.000 167.210 ;
        RECT 64.775 167.025 65.065 167.070 ;
        RECT 65.680 167.010 66.000 167.070 ;
        RECT 69.375 167.210 69.665 167.255 ;
        RECT 69.820 167.210 70.140 167.270 ;
        RECT 69.375 167.070 70.140 167.210 ;
        RECT 69.375 167.025 69.665 167.070 ;
        RECT 69.820 167.010 70.140 167.070 ;
        RECT 70.755 167.210 71.045 167.255 ;
        RECT 73.130 167.210 73.270 167.410 ;
        RECT 78.560 167.350 78.880 167.410 ;
        RECT 82.240 167.350 82.560 167.410 ;
        RECT 96.515 167.550 96.805 167.595 ;
        RECT 96.960 167.550 97.280 167.610 ;
        RECT 96.515 167.410 97.280 167.550 ;
        RECT 96.515 167.365 96.805 167.410 ;
        RECT 96.960 167.350 97.280 167.410 ;
        RECT 106.175 167.550 106.465 167.595 ;
        RECT 111.680 167.550 112.000 167.610 ;
        RECT 106.175 167.410 112.000 167.550 ;
        RECT 106.175 167.365 106.465 167.410 ;
        RECT 111.680 167.350 112.000 167.410 ;
        RECT 75.860 167.210 76.150 167.255 ;
        RECT 70.755 167.070 73.270 167.210 ;
        RECT 73.615 167.070 76.150 167.210 ;
        RECT 82.330 167.210 82.470 167.350 ;
        RECT 85.015 167.210 85.305 167.255 ;
        RECT 82.330 167.070 85.305 167.210 ;
        RECT 70.755 167.025 71.045 167.070 ;
        RECT 62.000 166.870 62.320 166.930 ;
        RECT 73.615 166.915 73.830 167.070 ;
        RECT 75.860 167.025 76.150 167.070 ;
        RECT 85.015 167.025 85.305 167.070 ;
        RECT 86.395 167.025 86.685 167.255 ;
        RECT 65.235 166.870 65.525 166.915 ;
        RECT 47.830 166.730 65.525 166.870 ;
        RECT 30.810 166.390 34.630 166.530 ;
        RECT 34.860 166.530 35.180 166.590 ;
        RECT 44.150 166.530 44.290 166.685 ;
        RECT 62.000 166.670 62.320 166.730 ;
        RECT 65.235 166.685 65.525 166.730 ;
        RECT 71.680 166.870 71.970 166.915 ;
        RECT 73.540 166.870 73.830 166.915 ;
        RECT 71.680 166.730 73.830 166.870 ;
        RECT 71.680 166.685 71.970 166.730 ;
        RECT 73.540 166.685 73.830 166.730 ;
        RECT 74.460 166.870 74.750 166.915 ;
        RECT 76.720 166.870 77.040 166.930 ;
        RECT 77.720 166.870 78.010 166.915 ;
        RECT 74.460 166.730 78.010 166.870 ;
        RECT 74.460 166.685 74.750 166.730 ;
        RECT 76.720 166.670 77.040 166.730 ;
        RECT 77.720 166.685 78.010 166.730 ;
        RECT 84.080 166.870 84.400 166.930 ;
        RECT 86.470 166.870 86.610 167.025 ;
        RECT 87.760 167.010 88.080 167.270 ;
        RECT 99.215 166.915 99.505 167.230 ;
        RECT 100.295 167.210 100.585 167.255 ;
        RECT 103.875 167.210 104.165 167.255 ;
        RECT 105.710 167.210 106.000 167.255 ;
        RECT 100.295 167.070 106.000 167.210 ;
        RECT 100.295 167.025 100.585 167.070 ;
        RECT 103.875 167.025 104.165 167.070 ;
        RECT 105.710 167.025 106.000 167.070 ;
        RECT 106.620 167.010 106.940 167.270 ;
        RECT 110.760 167.010 111.080 167.270 ;
        RECT 84.080 166.730 86.610 166.870 ;
        RECT 98.915 166.870 99.505 166.915 ;
        RECT 101.100 166.870 101.420 166.930 ;
        RECT 102.155 166.870 102.805 166.915 ;
        RECT 98.915 166.730 102.805 166.870 ;
        RECT 84.080 166.670 84.400 166.730 ;
        RECT 98.915 166.685 99.205 166.730 ;
        RECT 101.100 166.670 101.420 166.730 ;
        RECT 102.155 166.685 102.805 166.730 ;
        RECT 104.780 166.670 105.100 166.930 ;
        RECT 108.935 166.870 109.225 166.915 ;
        RECT 113.520 166.870 113.840 166.930 ;
        RECT 108.935 166.730 113.840 166.870 ;
        RECT 108.935 166.685 109.225 166.730 ;
        RECT 113.520 166.670 113.840 166.730 ;
        RECT 47.280 166.530 47.600 166.590 ;
        RECT 79.940 166.575 80.260 166.590 ;
        RECT 34.860 166.390 47.600 166.530 ;
        RECT 17.395 166.345 17.685 166.390 ;
        RECT 34.860 166.330 35.180 166.390 ;
        RECT 47.280 166.330 47.600 166.390 ;
        RECT 79.725 166.345 80.260 166.575 ;
        RECT 79.940 166.330 80.260 166.345 ;
        RECT 95.580 166.530 95.900 166.590 ;
        RECT 97.435 166.530 97.725 166.575 ;
        RECT 95.580 166.390 97.725 166.530 ;
        RECT 95.580 166.330 95.900 166.390 ;
        RECT 97.435 166.345 97.725 166.390 ;
        RECT 11.330 165.710 113.450 166.190 ;
        RECT 15.080 165.510 15.400 165.570 ;
        RECT 21.765 165.510 22.055 165.555 ;
        RECT 24.280 165.510 24.600 165.570 ;
        RECT 27.040 165.510 27.360 165.570 ;
        RECT 15.080 165.370 16.230 165.510 ;
        RECT 15.080 165.310 15.400 165.370 ;
        RECT 13.720 165.170 14.010 165.215 ;
        RECT 15.580 165.170 15.870 165.215 ;
        RECT 13.720 165.030 15.870 165.170 ;
        RECT 16.090 165.170 16.230 165.370 ;
        RECT 21.765 165.370 27.360 165.510 ;
        RECT 21.765 165.325 22.055 165.370 ;
        RECT 24.280 165.310 24.600 165.370 ;
        RECT 27.040 165.310 27.360 165.370 ;
        RECT 34.860 165.510 35.180 165.570 ;
        RECT 35.795 165.510 36.085 165.555 ;
        RECT 34.860 165.370 36.085 165.510 ;
        RECT 34.860 165.310 35.180 165.370 ;
        RECT 35.795 165.325 36.085 165.370 ;
        RECT 38.555 165.510 38.845 165.555 ;
        RECT 41.760 165.510 42.080 165.570 ;
        RECT 75.800 165.510 76.120 165.570 ;
        RECT 38.555 165.370 42.080 165.510 ;
        RECT 38.555 165.325 38.845 165.370 ;
        RECT 41.760 165.310 42.080 165.370 ;
        RECT 70.830 165.370 76.120 165.510 ;
        RECT 16.500 165.170 16.790 165.215 ;
        RECT 19.760 165.170 20.050 165.215 ;
        RECT 16.090 165.030 20.050 165.170 ;
        RECT 13.720 164.985 14.010 165.030 ;
        RECT 15.580 164.985 15.870 165.030 ;
        RECT 16.500 164.985 16.790 165.030 ;
        RECT 19.760 164.985 20.050 165.030 ;
        RECT 35.320 165.170 35.640 165.230 ;
        RECT 40.035 165.170 40.325 165.215 ;
        RECT 43.275 165.170 43.925 165.215 ;
        RECT 55.100 165.170 55.420 165.230 ;
        RECT 35.320 165.030 43.925 165.170 ;
        RECT 14.620 164.630 14.940 164.890 ;
        RECT 15.655 164.830 15.870 164.985 ;
        RECT 35.320 164.970 35.640 165.030 ;
        RECT 40.035 164.985 40.625 165.030 ;
        RECT 43.275 164.985 43.925 165.030 ;
        RECT 52.890 165.030 55.420 165.170 ;
        RECT 17.900 164.830 18.190 164.875 ;
        RECT 15.655 164.690 18.190 164.830 ;
        RECT 17.900 164.645 18.190 164.690 ;
        RECT 24.740 164.630 25.060 164.890 ;
        RECT 25.200 164.830 25.520 164.890 ;
        RECT 27.055 164.830 27.345 164.875 ;
        RECT 25.200 164.690 27.345 164.830 ;
        RECT 25.200 164.630 25.520 164.690 ;
        RECT 27.055 164.645 27.345 164.690 ;
        RECT 29.340 164.630 29.660 164.890 ;
        RECT 40.335 164.670 40.625 164.985 ;
        RECT 41.415 164.830 41.705 164.875 ;
        RECT 44.995 164.830 45.285 164.875 ;
        RECT 46.830 164.830 47.120 164.875 ;
        RECT 41.415 164.690 47.120 164.830 ;
        RECT 41.415 164.645 41.705 164.690 ;
        RECT 44.995 164.645 45.285 164.690 ;
        RECT 46.830 164.645 47.120 164.690 ;
        RECT 47.280 164.830 47.600 164.890 ;
        RECT 49.580 164.830 49.900 164.890 ;
        RECT 52.890 164.875 53.030 165.030 ;
        RECT 55.100 164.970 55.420 165.030 ;
        RECT 62.000 165.170 62.320 165.230 ;
        RECT 62.475 165.170 62.765 165.215 ;
        RECT 62.000 165.030 62.765 165.170 ;
        RECT 62.000 164.970 62.320 165.030 ;
        RECT 62.475 164.985 62.765 165.030 ;
        RECT 67.010 165.170 67.300 165.215 ;
        RECT 70.270 165.170 70.560 165.215 ;
        RECT 70.830 165.170 70.970 165.370 ;
        RECT 75.800 165.310 76.120 165.370 ;
        RECT 104.780 165.510 105.100 165.570 ;
        RECT 108.475 165.510 108.765 165.555 ;
        RECT 104.780 165.370 108.765 165.510 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 104.780 165.310 105.100 165.370 ;
        RECT 108.475 165.325 108.765 165.370 ;
        RECT 82.700 165.215 83.020 165.230 ;
        RECT 67.010 165.030 70.970 165.170 ;
        RECT 71.190 165.170 71.480 165.215 ;
        RECT 73.050 165.170 73.340 165.215 ;
        RECT 71.190 165.030 73.340 165.170 ;
        RECT 67.010 164.985 67.300 165.030 ;
        RECT 70.270 164.985 70.560 165.030 ;
        RECT 71.190 164.985 71.480 165.030 ;
        RECT 73.050 164.985 73.340 165.030 ;
        RECT 76.740 165.170 77.030 165.215 ;
        RECT 78.600 165.170 78.890 165.215 ;
        RECT 76.740 165.030 78.890 165.170 ;
        RECT 76.740 164.985 77.030 165.030 ;
        RECT 78.600 164.985 78.890 165.030 ;
        RECT 79.520 165.170 79.810 165.215 ;
        RECT 82.700 165.170 83.070 165.215 ;
        RECT 96.960 165.170 97.280 165.230 ;
        RECT 79.520 165.030 83.070 165.170 ;
        RECT 79.520 164.985 79.810 165.030 ;
        RECT 82.700 164.985 83.070 165.030 ;
        RECT 96.130 165.030 97.280 165.170 ;
        RECT 47.280 164.690 49.900 164.830 ;
        RECT 47.280 164.630 47.600 164.690 ;
        RECT 49.580 164.630 49.900 164.690 ;
        RECT 52.815 164.645 53.105 164.875 ;
        RECT 68.870 164.830 69.160 164.875 ;
        RECT 71.190 164.830 71.405 164.985 ;
        RECT 68.870 164.690 71.405 164.830 ;
        RECT 68.870 164.645 69.160 164.690 ;
        RECT 77.640 164.630 77.960 164.890 ;
        RECT 78.675 164.830 78.890 164.985 ;
        RECT 82.700 164.970 83.020 164.985 ;
        RECT 96.130 164.875 96.270 165.030 ;
        RECT 96.960 164.970 97.280 165.030 ;
        RECT 102.020 165.170 102.340 165.230 ;
        RECT 102.495 165.170 102.785 165.215 ;
        RECT 102.020 165.030 102.785 165.170 ;
        RECT 102.020 164.970 102.340 165.030 ;
        RECT 102.495 164.985 102.785 165.030 ;
        RECT 80.920 164.830 81.210 164.875 ;
        RECT 78.675 164.690 81.210 164.830 ;
        RECT 80.920 164.645 81.210 164.690 ;
        RECT 96.055 164.645 96.345 164.875 ;
        RECT 108.015 164.830 108.305 164.875 ;
        RECT 109.395 164.830 109.685 164.875 ;
        RECT 108.015 164.690 109.685 164.830 ;
        RECT 108.015 164.645 108.305 164.690 ;
        RECT 109.395 164.645 109.685 164.690 ;
        RECT 12.780 164.490 13.100 164.550 ;
        RECT 19.680 164.490 20.000 164.550 ;
        RECT 12.780 164.350 20.000 164.490 ;
        RECT 12.780 164.290 13.100 164.350 ;
        RECT 19.680 164.290 20.000 164.350 ;
        RECT 27.500 164.290 27.820 164.550 ;
        RECT 28.435 164.490 28.725 164.535 ;
        RECT 39.000 164.490 39.320 164.550 ;
        RECT 28.435 164.350 39.320 164.490 ;
        RECT 28.435 164.305 28.725 164.350 ;
        RECT 13.260 164.150 13.550 164.195 ;
        RECT 15.120 164.150 15.410 164.195 ;
        RECT 17.900 164.150 18.190 164.195 ;
        RECT 13.260 164.010 18.190 164.150 ;
        RECT 13.260 163.965 13.550 164.010 ;
        RECT 15.120 163.965 15.410 164.010 ;
        RECT 17.900 163.965 18.190 164.010 ;
        RECT 20.140 164.150 20.460 164.210 ;
        RECT 23.835 164.150 24.125 164.195 ;
        RECT 20.140 164.010 24.125 164.150 ;
        RECT 20.140 163.950 20.460 164.010 ;
        RECT 23.835 163.965 24.125 164.010 ;
        RECT 25.660 164.150 25.980 164.210 ;
        RECT 28.510 164.150 28.650 164.305 ;
        RECT 39.000 164.290 39.320 164.350 ;
        RECT 45.900 164.290 46.220 164.550 ;
        RECT 51.895 164.490 52.185 164.535 ;
        RECT 54.640 164.490 54.960 164.550 ;
        RECT 56.480 164.490 56.800 164.550 ;
        RECT 51.895 164.350 56.800 164.490 ;
        RECT 51.895 164.305 52.185 164.350 ;
        RECT 54.640 164.290 54.960 164.350 ;
        RECT 56.480 164.290 56.800 164.350 ;
        RECT 70.740 164.490 71.060 164.550 ;
        RECT 72.135 164.490 72.425 164.535 ;
        RECT 70.740 164.350 72.425 164.490 ;
        RECT 70.740 164.290 71.060 164.350 ;
        RECT 72.135 164.305 72.425 164.350 ;
        RECT 73.975 164.490 74.265 164.535 ;
        RECT 75.815 164.490 76.105 164.535 ;
        RECT 78.560 164.490 78.880 164.550 ;
        RECT 73.975 164.350 78.880 164.490 ;
        RECT 73.975 164.305 74.265 164.350 ;
        RECT 75.815 164.305 76.105 164.350 ;
        RECT 78.560 164.290 78.880 164.350 ;
        RECT 95.580 164.490 95.900 164.550 ;
        RECT 96.975 164.490 97.265 164.535 ;
        RECT 95.580 164.350 97.265 164.490 ;
        RECT 95.580 164.290 95.900 164.350 ;
        RECT 96.975 164.305 97.265 164.350 ;
        RECT 98.340 164.490 98.660 164.550 ;
        RECT 101.115 164.490 101.405 164.535 ;
        RECT 101.560 164.490 101.880 164.550 ;
        RECT 98.340 164.350 101.880 164.490 ;
        RECT 98.340 164.290 98.660 164.350 ;
        RECT 101.115 164.305 101.405 164.350 ;
        RECT 101.560 164.290 101.880 164.350 ;
        RECT 102.035 164.305 102.325 164.535 ;
        RECT 104.795 164.305 105.085 164.535 ;
        RECT 84.540 164.195 84.860 164.210 ;
        RECT 25.660 164.010 28.650 164.150 ;
        RECT 41.415 164.150 41.705 164.195 ;
        RECT 44.535 164.150 44.825 164.195 ;
        RECT 46.425 164.150 46.715 164.195 ;
        RECT 41.415 164.010 46.715 164.150 ;
        RECT 25.660 163.950 25.980 164.010 ;
        RECT 41.415 163.965 41.705 164.010 ;
        RECT 44.535 163.965 44.825 164.010 ;
        RECT 46.425 163.965 46.715 164.010 ;
        RECT 63.855 164.150 64.145 164.195 ;
        RECT 68.870 164.150 69.160 164.195 ;
        RECT 71.650 164.150 71.940 164.195 ;
        RECT 73.510 164.150 73.800 164.195 ;
        RECT 63.855 164.010 68.670 164.150 ;
        RECT 63.855 163.965 64.145 164.010 ;
        RECT 23.360 163.810 23.680 163.870 ;
        RECT 25.215 163.810 25.505 163.855 ;
        RECT 23.360 163.670 25.505 163.810 ;
        RECT 23.360 163.610 23.680 163.670 ;
        RECT 25.215 163.625 25.505 163.670 ;
        RECT 54.655 163.810 54.945 163.855 ;
        RECT 55.100 163.810 55.420 163.870 ;
        RECT 54.655 163.670 55.420 163.810 ;
        RECT 54.655 163.625 54.945 163.670 ;
        RECT 55.100 163.610 55.420 163.670 ;
        RECT 65.005 163.810 65.295 163.855 ;
        RECT 67.520 163.810 67.840 163.870 ;
        RECT 65.005 163.670 67.840 163.810 ;
        RECT 68.530 163.810 68.670 164.010 ;
        RECT 68.870 164.010 73.800 164.150 ;
        RECT 68.870 163.965 69.160 164.010 ;
        RECT 71.650 163.965 71.940 164.010 ;
        RECT 73.510 163.965 73.800 164.010 ;
        RECT 76.280 164.150 76.570 164.195 ;
        RECT 78.140 164.150 78.430 164.195 ;
        RECT 80.920 164.150 81.210 164.195 ;
        RECT 76.280 164.010 81.210 164.150 ;
        RECT 76.280 163.965 76.570 164.010 ;
        RECT 78.140 163.965 78.430 164.010 ;
        RECT 80.920 163.965 81.210 164.010 ;
        RECT 84.540 163.965 85.075 164.195 ;
        RECT 102.110 164.150 102.250 164.305 ;
        RECT 99.810 164.010 102.250 164.150 ;
        RECT 104.335 164.150 104.625 164.195 ;
        RECT 104.870 164.150 105.010 164.305 ;
        RECT 104.335 164.010 105.010 164.150 ;
        RECT 84.540 163.950 84.860 163.965 ;
        RECT 99.810 163.870 99.950 164.010 ;
        RECT 104.335 163.965 104.625 164.010 ;
        RECT 74.420 163.810 74.740 163.870 ;
        RECT 68.530 163.670 74.740 163.810 ;
        RECT 65.005 163.625 65.295 163.670 ;
        RECT 67.520 163.610 67.840 163.670 ;
        RECT 74.420 163.610 74.740 163.670 ;
        RECT 77.640 163.810 77.960 163.870 ;
        RECT 91.440 163.810 91.760 163.870 ;
        RECT 77.640 163.670 91.760 163.810 ;
        RECT 77.640 163.610 77.960 163.670 ;
        RECT 91.440 163.610 91.760 163.670 ;
        RECT 99.720 163.610 100.040 163.870 ;
        RECT 11.330 162.990 113.450 163.470 ;
        RECT 13.700 162.790 14.020 162.850 ;
        RECT 17.395 162.790 17.685 162.835 ;
        RECT 13.700 162.650 17.685 162.790 ;
        RECT 13.700 162.590 14.020 162.650 ;
        RECT 17.395 162.605 17.685 162.650 ;
        RECT 22.455 162.790 22.745 162.835 ;
        RECT 24.740 162.790 25.060 162.850 ;
        RECT 22.455 162.650 25.060 162.790 ;
        RECT 22.455 162.605 22.745 162.650 ;
        RECT 24.740 162.590 25.060 162.650 ;
        RECT 36.240 162.790 36.560 162.850 ;
        RECT 64.775 162.790 65.065 162.835 ;
        RECT 67.980 162.790 68.300 162.850 ;
        RECT 36.240 162.650 68.300 162.790 ;
        RECT 36.240 162.590 36.560 162.650 ;
        RECT 64.775 162.605 65.065 162.650 ;
        RECT 67.980 162.590 68.300 162.650 ;
        RECT 70.740 162.590 71.060 162.850 ;
        RECT 75.800 162.590 76.120 162.850 ;
        RECT 76.720 162.790 77.040 162.850 ;
        RECT 77.195 162.790 77.485 162.835 ;
        RECT 76.720 162.650 77.485 162.790 ;
        RECT 76.720 162.590 77.040 162.650 ;
        RECT 77.195 162.605 77.485 162.650 ;
        RECT 82.715 162.790 83.005 162.835 ;
        RECT 84.080 162.790 84.400 162.850 ;
        RECT 82.715 162.650 84.400 162.790 ;
        RECT 82.715 162.605 83.005 162.650 ;
        RECT 84.080 162.590 84.400 162.650 ;
        RECT 84.630 162.650 87.530 162.790 ;
        RECT 27.465 162.450 27.755 162.495 ;
        RECT 29.355 162.450 29.645 162.495 ;
        RECT 32.475 162.450 32.765 162.495 ;
        RECT 27.465 162.310 32.765 162.450 ;
        RECT 27.465 162.265 27.755 162.310 ;
        RECT 29.355 162.265 29.645 162.310 ;
        RECT 32.475 162.265 32.765 162.310 ;
        RECT 35.335 162.450 35.625 162.495 ;
        RECT 35.780 162.450 36.100 162.510 ;
        RECT 39.460 162.450 39.780 162.510 ;
        RECT 35.335 162.310 39.780 162.450 ;
        RECT 35.335 162.265 35.625 162.310 ;
        RECT 35.780 162.250 36.100 162.310 ;
        RECT 39.460 162.250 39.780 162.310 ;
        RECT 39.935 162.265 40.225 162.495 ;
        RECT 43.255 162.450 43.545 162.495 ;
        RECT 46.375 162.450 46.665 162.495 ;
        RECT 48.265 162.450 48.555 162.495 ;
        RECT 69.820 162.450 70.140 162.510 ;
        RECT 71.215 162.450 71.505 162.495 ;
        RECT 43.255 162.310 48.555 162.450 ;
        RECT 43.255 162.265 43.545 162.310 ;
        RECT 46.375 162.265 46.665 162.310 ;
        RECT 48.265 162.265 48.555 162.310 ;
        RECT 48.750 162.310 50.730 162.450 ;
        RECT 20.140 162.110 20.460 162.170 ;
        RECT 20.615 162.110 20.905 162.155 ;
        RECT 25.660 162.110 25.980 162.170 ;
        RECT 20.140 161.970 25.980 162.110 ;
        RECT 20.140 161.910 20.460 161.970 ;
        RECT 20.615 161.925 20.905 161.970 ;
        RECT 25.660 161.910 25.980 161.970 ;
        RECT 27.960 162.110 28.280 162.170 ;
        RECT 37.175 162.110 37.465 162.155 ;
        RECT 39.000 162.110 39.320 162.170 ;
        RECT 27.960 161.970 34.170 162.110 ;
        RECT 27.960 161.910 28.280 161.970 ;
        RECT 13.715 161.770 14.005 161.815 ;
        RECT 14.160 161.770 14.480 161.830 ;
        RECT 13.715 161.630 14.480 161.770 ;
        RECT 13.715 161.585 14.005 161.630 ;
        RECT 14.160 161.570 14.480 161.630 ;
        RECT 16.475 161.770 16.765 161.815 ;
        RECT 19.220 161.770 19.540 161.830 ;
        RECT 16.475 161.630 19.540 161.770 ;
        RECT 16.475 161.585 16.765 161.630 ;
        RECT 19.220 161.570 19.540 161.630 ;
        RECT 19.695 161.770 19.985 161.815 ;
        RECT 24.280 161.770 24.600 161.830 ;
        RECT 19.695 161.630 24.600 161.770 ;
        RECT 19.695 161.585 19.985 161.630 ;
        RECT 24.280 161.570 24.600 161.630 ;
        RECT 24.755 161.770 25.045 161.815 ;
        RECT 25.200 161.770 25.520 161.830 ;
        RECT 24.755 161.630 25.520 161.770 ;
        RECT 24.755 161.585 25.045 161.630 ;
        RECT 25.200 161.570 25.520 161.630 ;
        RECT 26.595 161.585 26.885 161.815 ;
        RECT 27.060 161.770 27.350 161.815 ;
        RECT 28.895 161.770 29.185 161.815 ;
        RECT 32.475 161.770 32.765 161.815 ;
        RECT 27.060 161.630 32.765 161.770 ;
        RECT 27.060 161.585 27.350 161.630 ;
        RECT 28.895 161.585 29.185 161.630 ;
        RECT 32.475 161.585 32.765 161.630 ;
        RECT 19.310 161.430 19.450 161.570 ;
        RECT 22.440 161.430 22.760 161.490 ;
        RECT 26.670 161.430 26.810 161.585 ;
        RECT 30.260 161.475 30.580 161.490 ;
        RECT 33.555 161.475 33.845 161.790 ;
        RECT 34.030 161.770 34.170 161.970 ;
        RECT 37.175 161.970 39.320 162.110 ;
        RECT 40.010 162.110 40.150 162.265 ;
        RECT 48.750 162.110 48.890 162.310 ;
        RECT 40.010 161.970 48.890 162.110 ;
        RECT 49.135 162.110 49.425 162.155 ;
        RECT 49.580 162.110 49.900 162.170 ;
        RECT 49.135 161.970 49.900 162.110 ;
        RECT 37.175 161.925 37.465 161.970 ;
        RECT 39.000 161.910 39.320 161.970 ;
        RECT 49.135 161.925 49.425 161.970 ;
        RECT 49.580 161.910 49.900 161.970 ;
        RECT 38.095 161.770 38.385 161.815 ;
        RECT 34.030 161.630 38.385 161.770 ;
        RECT 38.095 161.585 38.385 161.630 ;
        RECT 19.310 161.290 26.810 161.430 ;
        RECT 22.440 161.230 22.760 161.290 ;
        RECT 27.975 161.245 28.265 161.475 ;
        RECT 30.255 161.430 30.905 161.475 ;
        RECT 33.555 161.430 34.145 161.475 ;
        RECT 30.255 161.290 34.145 161.430 ;
        RECT 30.255 161.245 30.905 161.290 ;
        RECT 33.855 161.245 34.145 161.290 ;
        RECT 34.860 161.430 35.180 161.490 ;
        RECT 42.175 161.475 42.465 161.790 ;
        RECT 43.255 161.770 43.545 161.815 ;
        RECT 46.835 161.770 47.125 161.815 ;
        RECT 48.670 161.770 48.960 161.815 ;
        RECT 43.255 161.630 48.960 161.770 ;
        RECT 43.255 161.585 43.545 161.630 ;
        RECT 46.835 161.585 47.125 161.630 ;
        RECT 48.670 161.585 48.960 161.630 ;
        RECT 41.875 161.430 42.465 161.475 ;
        RECT 45.115 161.430 45.765 161.475 ;
        RECT 34.860 161.290 45.765 161.430 ;
        RECT 13.255 161.090 13.545 161.135 ;
        RECT 16.920 161.090 17.240 161.150 ;
        RECT 13.255 160.950 17.240 161.090 ;
        RECT 13.255 160.905 13.545 160.950 ;
        RECT 16.920 160.890 17.240 160.950 ;
        RECT 19.235 161.090 19.525 161.135 ;
        RECT 19.680 161.090 20.000 161.150 ;
        RECT 19.235 160.950 20.000 161.090 ;
        RECT 19.235 160.905 19.525 160.950 ;
        RECT 19.680 160.890 20.000 160.950 ;
        RECT 24.280 161.090 24.600 161.150 ;
        RECT 28.050 161.090 28.190 161.245 ;
        RECT 30.260 161.230 30.580 161.245 ;
        RECT 34.860 161.230 35.180 161.290 ;
        RECT 41.875 161.245 42.165 161.290 ;
        RECT 45.115 161.245 45.765 161.290 ;
        RECT 47.755 161.245 48.045 161.475 ;
        RECT 49.670 161.430 49.810 161.910 ;
        RECT 50.590 161.815 50.730 162.310 ;
        RECT 69.820 162.310 71.505 162.450 ;
        RECT 69.820 162.250 70.140 162.310 ;
        RECT 71.215 162.265 71.505 162.310 ;
        RECT 61.540 162.110 61.860 162.170 ;
        RECT 74.420 162.110 74.740 162.170 ;
        RECT 79.955 162.110 80.245 162.155 ;
        RECT 81.780 162.110 82.100 162.170 ;
        RECT 84.095 162.110 84.385 162.155 ;
        RECT 84.630 162.110 84.770 162.650 ;
        RECT 86.855 162.265 87.145 162.495 ;
        RECT 87.390 162.450 87.530 162.650 ;
        RECT 91.440 162.590 91.760 162.850 ;
        RECT 97.420 162.790 97.740 162.850 ;
        RECT 108.475 162.790 108.765 162.835 ;
        RECT 110.760 162.790 111.080 162.850 ;
        RECT 97.420 162.650 100.410 162.790 ;
        RECT 97.420 162.590 97.740 162.650 ;
        RECT 96.515 162.450 96.805 162.495 ;
        RECT 97.880 162.450 98.200 162.510 ;
        RECT 87.390 162.310 93.970 162.450 ;
        RECT 59.330 161.970 64.070 162.110 ;
        RECT 50.515 161.585 50.805 161.815 ;
        RECT 55.100 161.770 55.420 161.830 ;
        RECT 59.330 161.815 59.470 161.970 ;
        RECT 61.540 161.910 61.860 161.970 ;
        RECT 56.495 161.770 56.785 161.815 ;
        RECT 55.100 161.630 56.785 161.770 ;
        RECT 55.100 161.570 55.420 161.630 ;
        RECT 56.495 161.585 56.785 161.630 ;
        RECT 59.255 161.585 59.545 161.815 ;
        RECT 61.080 161.770 61.400 161.830 ;
        RECT 63.930 161.815 64.070 161.970 ;
        RECT 74.420 161.970 84.770 162.110 ;
        RECT 74.420 161.910 74.740 161.970 ;
        RECT 79.955 161.925 80.245 161.970 ;
        RECT 81.780 161.910 82.100 161.970 ;
        RECT 84.095 161.925 84.385 161.970 ;
        RECT 62.015 161.770 62.305 161.815 ;
        RECT 61.080 161.630 62.305 161.770 ;
        RECT 61.080 161.570 61.400 161.630 ;
        RECT 62.015 161.585 62.305 161.630 ;
        RECT 63.855 161.585 64.145 161.815 ;
        RECT 69.820 161.570 70.140 161.830 ;
        RECT 76.275 161.770 76.565 161.815 ;
        RECT 77.655 161.770 77.945 161.815 ;
        RECT 79.020 161.770 79.340 161.830 ;
        RECT 76.275 161.630 79.340 161.770 ;
        RECT 76.275 161.585 76.565 161.630 ;
        RECT 77.655 161.585 77.945 161.630 ;
        RECT 79.020 161.570 79.340 161.630 ;
        RECT 80.415 161.770 80.705 161.815 ;
        RECT 86.380 161.770 86.700 161.830 ;
        RECT 80.415 161.630 86.700 161.770 ;
        RECT 86.930 161.770 87.070 162.265 ;
        RECT 88.220 162.110 88.540 162.170 ;
        RECT 90.520 162.110 90.840 162.170 ;
        RECT 93.830 162.155 93.970 162.310 ;
        RECT 96.515 162.310 98.200 162.450 ;
        RECT 96.515 162.265 96.805 162.310 ;
        RECT 97.880 162.250 98.200 162.310 ;
        RECT 88.220 161.970 90.840 162.110 ;
        RECT 88.220 161.910 88.540 161.970 ;
        RECT 90.520 161.910 90.840 161.970 ;
        RECT 93.755 162.110 94.045 162.155 ;
        RECT 98.340 162.110 98.660 162.170 ;
        RECT 93.755 161.970 98.660 162.110 ;
        RECT 93.755 161.925 94.045 161.970 ;
        RECT 98.340 161.910 98.660 161.970 ;
        RECT 92.375 161.770 92.665 161.815 ;
        RECT 86.930 161.630 92.665 161.770 ;
        RECT 80.415 161.585 80.705 161.630 ;
        RECT 86.380 161.570 86.700 161.630 ;
        RECT 92.375 161.585 92.665 161.630 ;
        RECT 94.675 161.770 94.965 161.815 ;
        RECT 99.720 161.770 100.040 161.830 ;
        RECT 94.675 161.630 100.040 161.770 ;
        RECT 100.270 161.770 100.410 162.650 ;
        RECT 108.475 162.650 111.080 162.790 ;
        RECT 108.475 162.605 108.765 162.650 ;
        RECT 110.760 162.590 111.080 162.650 ;
        RECT 102.480 162.450 102.800 162.510 ;
        RECT 100.730 162.310 102.800 162.450 ;
        RECT 100.730 162.170 100.870 162.310 ;
        RECT 102.480 162.250 102.800 162.310 ;
        RECT 104.795 162.450 105.085 162.495 ;
        RECT 104.795 162.310 105.470 162.450 ;
        RECT 104.795 162.265 105.085 162.310 ;
        RECT 100.640 161.910 100.960 162.170 ;
        RECT 101.560 161.910 101.880 162.170 ;
        RECT 105.330 162.155 105.470 162.310 ;
        RECT 105.255 161.925 105.545 162.155 ;
        RECT 102.955 161.770 103.245 161.815 ;
        RECT 100.270 161.630 103.245 161.770 ;
        RECT 94.675 161.585 94.965 161.630 ;
        RECT 99.720 161.570 100.040 161.630 ;
        RECT 102.955 161.585 103.245 161.630 ;
        RECT 107.080 161.770 107.400 161.830 ;
        RECT 108.935 161.770 109.225 161.815 ;
        RECT 107.080 161.630 109.225 161.770 ;
        RECT 107.080 161.570 107.400 161.630 ;
        RECT 108.935 161.585 109.225 161.630 ;
        RECT 57.860 161.430 58.180 161.490 ;
        RECT 49.670 161.290 58.180 161.430 ;
        RECT 24.280 160.950 28.190 161.090 ;
        RECT 24.280 160.890 24.600 160.950 ;
        RECT 37.620 160.890 37.940 161.150 ;
        RECT 40.380 160.890 40.700 161.150 ;
        RECT 47.830 161.090 47.970 161.245 ;
        RECT 57.860 161.230 58.180 161.290 ;
        RECT 85.015 161.430 85.305 161.475 ;
        RECT 87.775 161.430 88.065 161.475 ;
        RECT 94.215 161.430 94.505 161.475 ;
        RECT 85.015 161.290 94.505 161.430 ;
        RECT 85.015 161.245 85.305 161.290 ;
        RECT 87.775 161.245 88.065 161.290 ;
        RECT 94.215 161.245 94.505 161.290 ;
        RECT 105.700 161.430 106.020 161.490 ;
        RECT 110.315 161.430 110.605 161.475 ;
        RECT 105.700 161.290 110.605 161.430 ;
        RECT 105.700 161.230 106.020 161.290 ;
        RECT 110.315 161.245 110.605 161.290 ;
        RECT 49.595 161.090 49.885 161.135 ;
        RECT 47.830 160.950 49.885 161.090 ;
        RECT 49.595 160.905 49.885 160.950 ;
        RECT 56.955 161.090 57.245 161.135 ;
        RECT 57.400 161.090 57.720 161.150 ;
        RECT 56.955 160.950 57.720 161.090 ;
        RECT 56.955 160.905 57.245 160.950 ;
        RECT 57.400 160.890 57.720 160.950 ;
        RECT 58.320 160.890 58.640 161.150 ;
        RECT 59.700 161.090 60.020 161.150 ;
        RECT 60.175 161.090 60.465 161.135 ;
        RECT 59.700 160.950 60.465 161.090 ;
        RECT 59.700 160.890 60.020 160.950 ;
        RECT 60.175 160.905 60.465 160.950 ;
        RECT 62.935 161.090 63.225 161.135 ;
        RECT 64.760 161.090 65.080 161.150 ;
        RECT 62.935 160.950 65.080 161.090 ;
        RECT 62.935 160.905 63.225 160.950 ;
        RECT 64.760 160.890 65.080 160.950 ;
        RECT 67.520 161.090 67.840 161.150 ;
        RECT 73.055 161.090 73.345 161.135 ;
        RECT 67.520 160.950 73.345 161.090 ;
        RECT 67.520 160.890 67.840 160.950 ;
        RECT 73.055 160.905 73.345 160.950 ;
        RECT 73.500 161.090 73.820 161.150 ;
        RECT 79.940 161.090 80.260 161.150 ;
        RECT 80.875 161.090 81.165 161.135 ;
        RECT 73.500 160.950 81.165 161.090 ;
        RECT 73.500 160.890 73.820 160.950 ;
        RECT 79.940 160.890 80.260 160.950 ;
        RECT 80.875 160.905 81.165 160.950 ;
        RECT 84.540 160.890 84.860 161.150 ;
        RECT 102.020 161.090 102.340 161.150 ;
        RECT 102.495 161.090 102.785 161.135 ;
        RECT 102.020 160.950 102.785 161.090 ;
        RECT 102.020 160.890 102.340 160.950 ;
        RECT 102.495 160.905 102.785 160.950 ;
        RECT 11.330 160.270 113.450 160.750 ;
        RECT 24.280 159.870 24.600 160.130 ;
        RECT 24.755 160.070 25.045 160.115 ;
        RECT 27.500 160.070 27.820 160.130 ;
        RECT 50.960 160.070 51.280 160.130 ;
        RECT 24.755 159.930 27.820 160.070 ;
        RECT 24.755 159.885 25.045 159.930 ;
        RECT 27.500 159.870 27.820 159.930 ;
        RECT 32.190 159.930 51.280 160.070 ;
        RECT 16.920 159.775 17.240 159.790 ;
        RECT 14.180 159.730 14.470 159.775 ;
        RECT 16.040 159.730 16.330 159.775 ;
        RECT 14.180 159.590 16.330 159.730 ;
        RECT 14.180 159.545 14.470 159.590 ;
        RECT 16.040 159.545 16.330 159.590 ;
        RECT 12.780 159.390 13.100 159.450 ;
        RECT 13.255 159.390 13.545 159.435 ;
        RECT 12.780 159.250 13.545 159.390 ;
        RECT 16.115 159.390 16.330 159.545 ;
        RECT 16.920 159.730 17.250 159.775 ;
        RECT 20.220 159.730 20.510 159.775 ;
        RECT 16.920 159.590 20.510 159.730 ;
        RECT 16.920 159.545 17.250 159.590 ;
        RECT 20.220 159.545 20.510 159.590 ;
        RECT 25.200 159.730 25.520 159.790 ;
        RECT 25.200 159.590 29.570 159.730 ;
        RECT 16.920 159.530 17.240 159.545 ;
        RECT 25.200 159.530 25.520 159.590 ;
        RECT 18.360 159.390 18.650 159.435 ;
        RECT 16.115 159.250 18.650 159.390 ;
        RECT 12.780 159.190 13.100 159.250 ;
        RECT 13.255 159.205 13.545 159.250 ;
        RECT 18.360 159.205 18.650 159.250 ;
        RECT 23.360 159.190 23.680 159.450 ;
        RECT 28.420 159.190 28.740 159.450 ;
        RECT 29.430 159.435 29.570 159.590 ;
        RECT 29.355 159.205 29.645 159.435 ;
        RECT 29.800 159.190 30.120 159.450 ;
        RECT 30.260 159.190 30.580 159.450 ;
        RECT 32.190 159.435 32.330 159.930 ;
        RECT 50.960 159.870 51.280 159.930 ;
        RECT 53.720 159.870 54.040 160.130 ;
        RECT 67.520 159.870 67.840 160.130 ;
        RECT 69.820 159.870 70.140 160.130 ;
        RECT 73.975 159.885 74.265 160.115 ;
        RECT 107.080 160.070 107.400 160.130 ;
        RECT 91.530 159.930 96.270 160.070 ;
        RECT 32.575 159.730 32.865 159.775 ;
        RECT 34.860 159.730 35.180 159.790 ;
        RECT 32.575 159.590 35.180 159.730 ;
        RECT 32.575 159.545 32.865 159.590 ;
        RECT 34.860 159.530 35.180 159.590 ;
        RECT 36.715 159.730 37.005 159.775 ;
        RECT 37.620 159.730 37.940 159.790 ;
        RECT 42.695 159.730 42.985 159.775 ;
        RECT 36.715 159.590 42.985 159.730 ;
        RECT 36.715 159.545 37.005 159.590 ;
        RECT 37.620 159.530 37.940 159.590 ;
        RECT 42.695 159.545 42.985 159.590 ;
        RECT 46.375 159.730 46.665 159.775 ;
        RECT 52.340 159.730 52.660 159.790 ;
        RECT 46.375 159.590 52.660 159.730 ;
        RECT 53.810 159.730 53.950 159.870 ;
        RECT 57.400 159.775 57.720 159.790 ;
        RECT 57.350 159.730 57.720 159.775 ;
        RECT 60.610 159.730 60.900 159.775 ;
        RECT 53.810 159.590 54.870 159.730 ;
        RECT 46.375 159.545 46.665 159.590 ;
        RECT 52.340 159.530 52.660 159.590 ;
        RECT 32.115 159.390 32.405 159.435 ;
        RECT 33.020 159.390 33.340 159.450 ;
        RECT 32.115 159.250 33.340 159.390 ;
        RECT 32.115 159.205 32.405 159.250 ;
        RECT 33.020 159.190 33.340 159.250 ;
        RECT 33.955 159.390 34.245 159.435 ;
        RECT 38.080 159.390 38.400 159.450 ;
        RECT 40.380 159.390 40.700 159.450 ;
        RECT 33.955 159.250 40.700 159.390 ;
        RECT 33.955 159.205 34.245 159.250 ;
        RECT 38.080 159.190 38.400 159.250 ;
        RECT 40.380 159.190 40.700 159.250 ;
        RECT 41.760 159.390 42.080 159.450 ;
        RECT 43.155 159.390 43.445 159.435 ;
        RECT 41.760 159.250 43.445 159.390 ;
        RECT 41.760 159.190 42.080 159.250 ;
        RECT 43.155 159.205 43.445 159.250 ;
        RECT 45.440 159.190 45.760 159.450 ;
        RECT 46.820 159.190 47.140 159.450 ;
        RECT 47.295 159.205 47.585 159.435 ;
        RECT 50.055 159.390 50.345 159.435 ;
        RECT 50.055 159.250 52.570 159.390 ;
        RECT 50.055 159.205 50.345 159.250 ;
        RECT 15.080 158.850 15.400 159.110 ;
        RECT 27.975 159.050 28.265 159.095 ;
        RECT 35.780 159.050 36.100 159.110 ;
        RECT 27.975 158.910 36.100 159.050 ;
        RECT 27.975 158.865 28.265 158.910 ;
        RECT 35.780 158.850 36.100 158.910 ;
        RECT 37.635 158.865 37.925 159.095 ;
        RECT 39.000 159.050 39.320 159.110 ;
        RECT 43.600 159.050 43.920 159.110 ;
        RECT 39.000 158.910 43.920 159.050 ;
        RECT 13.720 158.710 14.010 158.755 ;
        RECT 15.580 158.710 15.870 158.755 ;
        RECT 18.360 158.710 18.650 158.755 ;
        RECT 13.720 158.570 18.650 158.710 ;
        RECT 13.720 158.525 14.010 158.570 ;
        RECT 15.580 158.525 15.870 158.570 ;
        RECT 18.360 158.525 18.650 158.570 ;
        RECT 32.100 158.710 32.420 158.770 ;
        RECT 34.860 158.710 35.180 158.770 ;
        RECT 32.100 158.570 35.180 158.710 ;
        RECT 37.710 158.710 37.850 158.865 ;
        RECT 39.000 158.850 39.320 158.910 ;
        RECT 43.600 158.850 43.920 158.910 ;
        RECT 44.520 159.050 44.840 159.110 ;
        RECT 47.370 159.050 47.510 159.205 ;
        RECT 51.435 159.050 51.725 159.095 ;
        RECT 44.520 158.910 51.725 159.050 ;
        RECT 44.520 158.850 44.840 158.910 ;
        RECT 51.435 158.865 51.725 158.910 ;
        RECT 40.855 158.710 41.145 158.755 ;
        RECT 37.710 158.570 41.145 158.710 ;
        RECT 52.430 158.710 52.570 159.250 ;
        RECT 52.800 159.190 53.120 159.450 ;
        RECT 53.260 159.190 53.580 159.450 ;
        RECT 53.735 159.390 54.025 159.435 ;
        RECT 54.180 159.390 54.500 159.450 ;
        RECT 54.730 159.435 54.870 159.590 ;
        RECT 57.350 159.590 60.900 159.730 ;
        RECT 57.350 159.545 57.720 159.590 ;
        RECT 60.610 159.545 60.900 159.590 ;
        RECT 61.530 159.730 61.820 159.775 ;
        RECT 63.390 159.730 63.680 159.775 ;
        RECT 61.530 159.590 63.680 159.730 ;
        RECT 61.530 159.545 61.820 159.590 ;
        RECT 63.390 159.545 63.680 159.590 ;
        RECT 67.995 159.730 68.285 159.775 ;
        RECT 68.440 159.730 68.760 159.790 ;
        RECT 71.675 159.730 71.965 159.775 ;
        RECT 67.995 159.590 71.965 159.730 ;
        RECT 67.995 159.545 68.285 159.590 ;
        RECT 57.400 159.530 57.720 159.545 ;
        RECT 53.735 159.250 54.500 159.390 ;
        RECT 53.735 159.205 54.025 159.250 ;
        RECT 54.180 159.190 54.500 159.250 ;
        RECT 54.655 159.205 54.945 159.435 ;
        RECT 59.210 159.390 59.500 159.435 ;
        RECT 61.530 159.390 61.745 159.545 ;
        RECT 68.440 159.530 68.760 159.590 ;
        RECT 71.675 159.545 71.965 159.590 ;
        RECT 72.120 159.530 72.440 159.790 ;
        RECT 74.050 159.730 74.190 159.885 ;
        RECT 79.430 159.730 79.720 159.775 ;
        RECT 79.940 159.730 80.260 159.790 ;
        RECT 82.690 159.730 82.980 159.775 ;
        RECT 74.050 159.590 75.570 159.730 ;
        RECT 75.430 159.435 75.570 159.590 ;
        RECT 79.430 159.590 82.980 159.730 ;
        RECT 79.430 159.545 79.720 159.590 ;
        RECT 79.940 159.530 80.260 159.590 ;
        RECT 82.690 159.545 82.980 159.590 ;
        RECT 83.610 159.730 83.900 159.775 ;
        RECT 85.470 159.730 85.760 159.775 ;
        RECT 83.610 159.590 85.760 159.730 ;
        RECT 83.610 159.545 83.900 159.590 ;
        RECT 85.470 159.545 85.760 159.590 ;
        RECT 85.920 159.730 86.240 159.790 ;
        RECT 91.530 159.730 91.670 159.930 ;
        RECT 95.580 159.730 95.900 159.790 ;
        RECT 85.920 159.590 91.670 159.730 ;
        RECT 91.990 159.590 95.900 159.730 ;
        RECT 96.130 159.730 96.270 159.930 ;
        RECT 105.100 159.930 107.400 160.070 ;
        RECT 96.130 159.590 97.190 159.730 ;
        RECT 59.210 159.250 61.745 159.390 ;
        RECT 64.315 159.390 64.605 159.435 ;
        RECT 64.315 159.250 75.110 159.390 ;
        RECT 59.210 159.205 59.500 159.250 ;
        RECT 64.315 159.205 64.605 159.250 ;
        RECT 54.270 159.050 54.410 159.190 ;
        RECT 55.345 159.050 55.635 159.095 ;
        RECT 54.270 158.910 55.635 159.050 ;
        RECT 55.345 158.865 55.635 158.910 ;
        RECT 62.460 158.850 62.780 159.110 ;
        RECT 67.075 159.050 67.365 159.095 ;
        RECT 71.215 159.050 71.505 159.095 ;
        RECT 74.420 159.050 74.740 159.110 ;
        RECT 67.075 158.910 74.740 159.050 ;
        RECT 74.970 159.050 75.110 159.250 ;
        RECT 75.355 159.205 75.645 159.435 ;
        RECT 81.290 159.390 81.580 159.435 ;
        RECT 83.610 159.390 83.825 159.545 ;
        RECT 85.920 159.530 86.240 159.590 ;
        RECT 81.290 159.250 83.825 159.390 ;
        RECT 84.555 159.390 84.845 159.435 ;
        RECT 85.000 159.390 85.320 159.450 ;
        RECT 84.555 159.250 85.320 159.390 ;
        RECT 81.290 159.205 81.580 159.250 ;
        RECT 84.555 159.205 84.845 159.250 ;
        RECT 85.000 159.190 85.320 159.250 ;
        RECT 88.680 159.190 89.000 159.450 ;
        RECT 90.060 159.390 90.380 159.450 ;
        RECT 91.990 159.435 92.130 159.590 ;
        RECT 95.580 159.530 95.900 159.590 ;
        RECT 90.995 159.390 91.285 159.435 ;
        RECT 90.060 159.250 91.285 159.390 ;
        RECT 90.060 159.190 90.380 159.250 ;
        RECT 90.995 159.205 91.285 159.250 ;
        RECT 91.915 159.205 92.205 159.435 ;
        RECT 82.240 159.050 82.560 159.110 ;
        RECT 86.395 159.050 86.685 159.095 ;
        RECT 74.970 158.910 86.685 159.050 ;
        RECT 67.075 158.865 67.365 158.910 ;
        RECT 71.215 158.865 71.505 158.910 ;
        RECT 74.420 158.850 74.740 158.910 ;
        RECT 82.240 158.850 82.560 158.910 ;
        RECT 86.395 158.865 86.685 158.910 ;
        RECT 54.640 158.710 54.960 158.770 ;
        RECT 52.430 158.570 54.960 158.710 ;
        RECT 32.100 158.510 32.420 158.570 ;
        RECT 34.860 158.510 35.180 158.570 ;
        RECT 40.855 158.525 41.145 158.570 ;
        RECT 54.640 158.510 54.960 158.570 ;
        RECT 59.210 158.710 59.500 158.755 ;
        RECT 61.990 158.710 62.280 158.755 ;
        RECT 63.850 158.710 64.140 158.755 ;
        RECT 59.210 158.570 64.140 158.710 ;
        RECT 59.210 158.525 59.500 158.570 ;
        RECT 61.990 158.525 62.280 158.570 ;
        RECT 63.850 158.525 64.140 158.570 ;
        RECT 72.120 158.710 72.440 158.770 ;
        RECT 77.425 158.710 77.715 158.755 ;
        RECT 80.400 158.710 80.720 158.770 ;
        RECT 72.120 158.570 80.720 158.710 ;
        RECT 72.120 158.510 72.440 158.570 ;
        RECT 77.425 158.525 77.715 158.570 ;
        RECT 80.400 158.510 80.720 158.570 ;
        RECT 81.290 158.710 81.580 158.755 ;
        RECT 84.070 158.710 84.360 158.755 ;
        RECT 85.930 158.710 86.220 158.755 ;
        RECT 81.290 158.570 86.220 158.710 ;
        RECT 91.070 158.710 91.210 159.205 ;
        RECT 92.360 159.190 92.680 159.450 ;
        RECT 92.820 159.190 93.140 159.450 ;
        RECT 93.370 159.250 95.810 159.390 ;
        RECT 93.370 158.710 93.510 159.250 ;
        RECT 94.660 159.050 94.980 159.110 ;
        RECT 91.070 158.570 93.510 158.710 ;
        RECT 93.830 158.910 94.980 159.050 ;
        RECT 95.670 159.050 95.810 159.250 ;
        RECT 96.040 159.190 96.360 159.450 ;
        RECT 96.500 159.190 96.820 159.450 ;
        RECT 97.050 159.435 97.190 159.590 ;
        RECT 96.975 159.205 97.265 159.435 ;
        RECT 97.895 159.205 98.185 159.435 ;
        RECT 103.415 159.390 103.705 159.435 ;
        RECT 105.100 159.390 105.240 159.930 ;
        RECT 107.080 159.870 107.400 159.930 ;
        RECT 103.415 159.250 105.240 159.390 ;
        RECT 103.415 159.205 103.705 159.250 ;
        RECT 97.970 159.050 98.110 159.205 ;
        RECT 102.940 159.050 103.260 159.110 ;
        RECT 95.670 158.910 103.260 159.050 ;
        RECT 81.290 158.525 81.580 158.570 ;
        RECT 84.070 158.525 84.360 158.570 ;
        RECT 85.930 158.525 86.220 158.570 ;
        RECT 19.680 158.370 20.000 158.430 ;
        RECT 22.225 158.370 22.515 158.415 ;
        RECT 19.680 158.230 22.515 158.370 ;
        RECT 19.680 158.170 20.000 158.230 ;
        RECT 22.225 158.185 22.515 158.230 ;
        RECT 31.655 158.370 31.945 158.415 ;
        RECT 37.160 158.370 37.480 158.430 ;
        RECT 31.655 158.230 37.480 158.370 ;
        RECT 31.655 158.185 31.945 158.230 ;
        RECT 37.160 158.170 37.480 158.230 ;
        RECT 40.395 158.370 40.685 158.415 ;
        RECT 43.600 158.370 43.920 158.430 ;
        RECT 40.395 158.230 43.920 158.370 ;
        RECT 40.395 158.185 40.685 158.230 ;
        RECT 43.600 158.170 43.920 158.230 ;
        RECT 48.215 158.370 48.505 158.415 ;
        RECT 49.580 158.370 49.900 158.430 ;
        RECT 48.215 158.230 49.900 158.370 ;
        RECT 48.215 158.185 48.505 158.230 ;
        RECT 49.580 158.170 49.900 158.230 ;
        RECT 50.500 158.170 50.820 158.430 ;
        RECT 64.300 158.370 64.620 158.430 ;
        RECT 65.680 158.370 66.000 158.430 ;
        RECT 66.600 158.370 66.920 158.430 ;
        RECT 64.300 158.230 66.920 158.370 ;
        RECT 64.300 158.170 64.620 158.230 ;
        RECT 65.680 158.170 66.000 158.230 ;
        RECT 66.600 158.170 66.920 158.230 ;
        RECT 76.275 158.370 76.565 158.415 ;
        RECT 76.720 158.370 77.040 158.430 ;
        RECT 76.275 158.230 77.040 158.370 ;
        RECT 76.275 158.185 76.565 158.230 ;
        RECT 76.720 158.170 77.040 158.230 ;
        RECT 82.700 158.370 83.020 158.430 ;
        RECT 88.235 158.370 88.525 158.415 ;
        RECT 82.700 158.230 88.525 158.370 ;
        RECT 82.700 158.170 83.020 158.230 ;
        RECT 88.235 158.185 88.525 158.230 ;
        RECT 91.440 158.370 91.760 158.430 ;
        RECT 93.830 158.370 93.970 158.910 ;
        RECT 94.660 158.850 94.980 158.910 ;
        RECT 102.940 158.850 103.260 158.910 ;
        RECT 104.320 158.850 104.640 159.110 ;
        RECT 94.215 158.710 94.505 158.755 ;
        RECT 99.260 158.710 99.580 158.770 ;
        RECT 94.215 158.570 99.580 158.710 ;
        RECT 94.215 158.525 94.505 158.570 ;
        RECT 99.260 158.510 99.580 158.570 ;
        RECT 91.440 158.230 93.970 158.370 ;
        RECT 91.440 158.170 91.760 158.230 ;
        RECT 94.660 158.170 94.980 158.430 ;
        RECT 11.330 157.550 113.450 158.030 ;
        RECT 14.635 157.350 14.925 157.395 ;
        RECT 15.080 157.350 15.400 157.410 ;
        RECT 14.635 157.210 15.400 157.350 ;
        RECT 14.635 157.165 14.925 157.210 ;
        RECT 15.080 157.150 15.400 157.210 ;
        RECT 22.440 157.350 22.760 157.410 ;
        RECT 27.040 157.350 27.360 157.410 ;
        RECT 22.440 157.210 27.360 157.350 ;
        RECT 22.440 157.150 22.760 157.210 ;
        RECT 27.040 157.150 27.360 157.210 ;
        RECT 31.655 157.350 31.945 157.395 ;
        RECT 32.100 157.350 32.420 157.410 ;
        RECT 36.255 157.350 36.545 157.395 ;
        RECT 31.655 157.210 32.420 157.350 ;
        RECT 31.655 157.165 31.945 157.210 ;
        RECT 32.100 157.150 32.420 157.210 ;
        RECT 32.650 157.210 36.545 157.350 ;
        RECT 19.680 157.010 20.000 157.070 ;
        RECT 18.390 156.870 20.000 157.010 ;
        RECT 18.390 156.730 18.530 156.870 ;
        RECT 19.680 156.810 20.000 156.870 ;
        RECT 22.900 157.010 23.220 157.070 ;
        RECT 32.650 157.010 32.790 157.210 ;
        RECT 36.255 157.165 36.545 157.210 ;
        RECT 37.635 157.165 37.925 157.395 ;
        RECT 39.460 157.350 39.780 157.410 ;
        RECT 44.995 157.350 45.285 157.395 ;
        RECT 45.440 157.350 45.760 157.410 ;
        RECT 39.460 157.210 41.990 157.350 ;
        RECT 22.900 156.870 32.790 157.010 ;
        RECT 22.900 156.810 23.220 156.870 ;
        RECT 18.300 156.470 18.620 156.730 ;
        RECT 19.235 156.670 19.525 156.715 ;
        RECT 20.140 156.670 20.460 156.730 ;
        RECT 19.235 156.530 20.460 156.670 ;
        RECT 19.235 156.485 19.525 156.530 ;
        RECT 20.140 156.470 20.460 156.530 ;
        RECT 29.340 156.670 29.660 156.730 ;
        RECT 29.340 156.530 32.330 156.670 ;
        RECT 29.340 156.470 29.660 156.530 ;
        RECT 15.555 156.330 15.845 156.375 ;
        RECT 15.555 156.190 16.230 156.330 ;
        RECT 15.555 156.145 15.845 156.190 ;
        RECT 16.090 155.695 16.230 156.190 ;
        RECT 28.880 156.130 29.200 156.390 ;
        RECT 30.275 156.145 30.565 156.375 ;
        RECT 30.735 156.330 31.025 156.375 ;
        RECT 31.180 156.330 31.500 156.390 ;
        RECT 30.735 156.190 31.500 156.330 ;
        RECT 30.735 156.145 31.025 156.190 ;
        RECT 24.740 155.990 25.060 156.050 ;
        RECT 26.580 155.990 26.900 156.050 ;
        RECT 30.350 155.990 30.490 156.145 ;
        RECT 31.180 156.130 31.500 156.190 ;
        RECT 31.640 156.130 31.960 156.390 ;
        RECT 32.190 156.330 32.330 156.530 ;
        RECT 32.560 156.470 32.880 156.730 ;
        RECT 37.710 156.670 37.850 157.165 ;
        RECT 39.460 157.150 39.780 157.210 ;
        RECT 36.790 156.530 37.850 156.670 ;
        RECT 38.095 156.670 38.385 156.715 ;
        RECT 38.540 156.670 38.860 156.730 ;
        RECT 38.095 156.530 38.860 156.670 ;
        RECT 36.790 156.330 36.930 156.530 ;
        RECT 38.095 156.485 38.385 156.530 ;
        RECT 38.540 156.470 38.860 156.530 ;
        RECT 39.000 156.470 39.320 156.730 ;
        RECT 32.190 156.190 36.930 156.330 ;
        RECT 37.160 156.130 37.480 156.390 ;
        RECT 39.460 156.330 39.780 156.390 ;
        RECT 40.395 156.330 40.685 156.375 ;
        RECT 39.460 156.190 40.685 156.330 ;
        RECT 39.460 156.130 39.780 156.190 ;
        RECT 40.395 156.145 40.685 156.190 ;
        RECT 40.840 156.130 41.160 156.390 ;
        RECT 41.315 156.330 41.605 156.375 ;
        RECT 41.850 156.330 41.990 157.210 ;
        RECT 44.995 157.210 45.760 157.350 ;
        RECT 44.995 157.165 45.285 157.210 ;
        RECT 45.440 157.150 45.760 157.210 ;
        RECT 53.720 157.350 54.040 157.410 ;
        RECT 61.095 157.350 61.385 157.395 ;
        RECT 62.460 157.350 62.780 157.410 ;
        RECT 74.420 157.350 74.740 157.410 ;
        RECT 53.720 157.210 59.470 157.350 ;
        RECT 53.720 157.150 54.040 157.210 ;
        RECT 44.535 157.010 44.825 157.055 ;
        RECT 45.900 157.010 46.220 157.070 ;
        RECT 44.535 156.870 46.220 157.010 ;
        RECT 44.535 156.825 44.825 156.870 ;
        RECT 45.900 156.810 46.220 156.870 ;
        RECT 49.580 157.010 49.900 157.070 ;
        RECT 54.150 157.010 54.440 157.055 ;
        RECT 56.930 157.010 57.220 157.055 ;
        RECT 58.790 157.010 59.080 157.055 ;
        RECT 49.580 156.870 51.190 157.010 ;
        RECT 49.580 156.810 49.900 156.870 ;
        RECT 50.285 156.485 50.575 156.715 ;
        RECT 51.050 156.670 51.190 156.870 ;
        RECT 54.150 156.870 59.080 157.010 ;
        RECT 59.330 157.010 59.470 157.210 ;
        RECT 61.095 157.210 62.780 157.350 ;
        RECT 61.095 157.165 61.385 157.210 ;
        RECT 62.460 157.150 62.780 157.210 ;
        RECT 64.390 157.210 74.740 157.350 ;
        RECT 64.390 157.055 64.530 157.210 ;
        RECT 74.420 157.150 74.740 157.210 ;
        RECT 79.940 157.150 80.260 157.410 ;
        RECT 85.000 157.150 85.320 157.410 ;
        RECT 88.680 157.350 89.000 157.410 ;
        RECT 88.680 157.210 104.550 157.350 ;
        RECT 88.680 157.150 89.000 157.210 ;
        RECT 64.315 157.010 64.605 157.055 ;
        RECT 59.330 156.870 64.605 157.010 ;
        RECT 54.150 156.825 54.440 156.870 ;
        RECT 56.930 156.825 57.220 156.870 ;
        RECT 58.790 156.825 59.080 156.870 ;
        RECT 64.315 156.825 64.605 156.870 ;
        RECT 67.520 156.810 67.840 157.070 ;
        RECT 68.900 156.810 69.220 157.070 ;
        RECT 73.470 157.010 73.760 157.055 ;
        RECT 76.250 157.010 76.540 157.055 ;
        RECT 78.110 157.010 78.400 157.055 ;
        RECT 82.240 157.010 82.560 157.070 ;
        RECT 73.470 156.870 78.400 157.010 ;
        RECT 73.470 156.825 73.760 156.870 ;
        RECT 76.250 156.825 76.540 156.870 ;
        RECT 78.110 156.825 78.400 156.870 ;
        RECT 78.650 156.870 82.560 157.010 ;
        RECT 57.415 156.670 57.705 156.715 ;
        RECT 51.050 156.530 57.705 156.670 ;
        RECT 57.415 156.485 57.705 156.530 ;
        RECT 64.760 156.670 65.080 156.730 ;
        RECT 67.610 156.670 67.750 156.810 ;
        RECT 64.760 156.530 66.370 156.670 ;
        RECT 41.315 156.190 41.990 156.330 ;
        RECT 41.315 156.145 41.605 156.190 ;
        RECT 42.235 156.145 42.525 156.375 ;
        RECT 37.620 155.990 37.940 156.050 ;
        RECT 24.740 155.850 30.030 155.990 ;
        RECT 30.350 155.850 37.940 155.990 ;
        RECT 24.740 155.790 25.060 155.850 ;
        RECT 26.580 155.790 26.900 155.850 ;
        RECT 16.015 155.465 16.305 155.695 ;
        RECT 17.840 155.450 18.160 155.710 ;
        RECT 24.280 155.650 24.600 155.710 ;
        RECT 29.355 155.650 29.645 155.695 ;
        RECT 24.280 155.510 29.645 155.650 ;
        RECT 29.890 155.650 30.030 155.850 ;
        RECT 37.620 155.790 37.940 155.850 ;
        RECT 38.555 155.990 38.845 156.035 ;
        RECT 41.760 155.990 42.080 156.050 ;
        RECT 42.310 155.990 42.450 156.145 ;
        RECT 43.600 156.130 43.920 156.390 ;
        RECT 47.740 156.330 48.060 156.390 ;
        RECT 50.360 156.330 50.500 156.485 ;
        RECT 64.760 156.470 65.080 156.530 ;
        RECT 47.740 156.190 50.500 156.330 ;
        RECT 54.150 156.330 54.440 156.375 ;
        RECT 57.860 156.330 58.180 156.390 ;
        RECT 59.255 156.330 59.545 156.375 ;
        RECT 54.150 156.190 56.685 156.330 ;
        RECT 47.740 156.130 48.060 156.190 ;
        RECT 54.150 156.145 54.440 156.190 ;
        RECT 50.500 155.990 50.820 156.050 ;
        RECT 56.470 156.035 56.685 156.190 ;
        RECT 57.860 156.190 59.545 156.330 ;
        RECT 57.860 156.130 58.180 156.190 ;
        RECT 59.255 156.145 59.545 156.190 ;
        RECT 60.160 156.130 60.480 156.390 ;
        RECT 64.300 156.330 64.620 156.390 ;
        RECT 65.235 156.330 65.525 156.375 ;
        RECT 64.300 156.190 65.525 156.330 ;
        RECT 64.300 156.130 64.620 156.190 ;
        RECT 65.235 156.145 65.525 156.190 ;
        RECT 65.695 156.145 65.985 156.375 ;
        RECT 52.290 155.990 52.580 156.035 ;
        RECT 55.550 155.990 55.840 156.035 ;
        RECT 38.555 155.850 41.070 155.990 ;
        RECT 38.555 155.805 38.845 155.850 ;
        RECT 40.930 155.710 41.070 155.850 ;
        RECT 41.760 155.850 50.270 155.990 ;
        RECT 41.760 155.790 42.080 155.850 ;
        RECT 31.640 155.650 31.960 155.710 ;
        RECT 33.020 155.650 33.340 155.710 ;
        RECT 29.890 155.510 33.340 155.650 ;
        RECT 24.280 155.450 24.600 155.510 ;
        RECT 29.355 155.465 29.645 155.510 ;
        RECT 31.640 155.450 31.960 155.510 ;
        RECT 33.020 155.450 33.340 155.510 ;
        RECT 35.335 155.650 35.625 155.695 ;
        RECT 35.780 155.650 36.100 155.710 ;
        RECT 35.335 155.510 36.100 155.650 ;
        RECT 35.335 155.465 35.625 155.510 ;
        RECT 35.780 155.450 36.100 155.510 ;
        RECT 40.840 155.450 41.160 155.710 ;
        RECT 42.220 155.650 42.540 155.710 ;
        RECT 43.600 155.650 43.920 155.710 ;
        RECT 42.220 155.510 43.920 155.650 ;
        RECT 50.130 155.650 50.270 155.850 ;
        RECT 50.500 155.850 55.840 155.990 ;
        RECT 50.500 155.790 50.820 155.850 ;
        RECT 52.290 155.805 52.580 155.850 ;
        RECT 55.550 155.805 55.840 155.850 ;
        RECT 56.470 155.990 56.760 156.035 ;
        RECT 58.330 155.990 58.620 156.035 ;
        RECT 56.470 155.850 58.620 155.990 ;
        RECT 56.470 155.805 56.760 155.850 ;
        RECT 58.330 155.805 58.620 155.850 ;
        RECT 65.770 155.650 65.910 156.145 ;
        RECT 66.230 155.990 66.370 156.530 ;
        RECT 66.690 156.530 67.750 156.670 ;
        RECT 68.440 156.670 68.760 156.730 ;
        RECT 69.605 156.670 69.895 156.715 ;
        RECT 68.440 156.530 69.895 156.670 ;
        RECT 66.690 156.375 66.830 156.530 ;
        RECT 68.440 156.470 68.760 156.530 ;
        RECT 69.605 156.485 69.895 156.530 ;
        RECT 76.720 156.470 77.040 156.730 ;
        RECT 78.650 156.715 78.790 156.870 ;
        RECT 82.240 156.810 82.560 156.870 ;
        RECT 84.555 156.825 84.845 157.055 ;
        RECT 78.575 156.485 78.865 156.715 ;
        RECT 81.780 156.470 82.100 156.730 ;
        RECT 66.615 156.145 66.905 156.375 ;
        RECT 67.075 156.145 67.365 156.375 ;
        RECT 67.150 155.990 67.290 156.145 ;
        RECT 67.520 156.130 67.840 156.390 ;
        RECT 73.470 156.330 73.760 156.375 ;
        RECT 73.470 156.190 76.005 156.330 ;
        RECT 73.470 156.145 73.760 156.190 ;
        RECT 66.230 155.850 67.290 155.990 ;
        RECT 71.610 155.990 71.900 156.035 ;
        RECT 73.960 155.990 74.280 156.050 ;
        RECT 75.790 156.035 76.005 156.190 ;
        RECT 79.480 156.130 79.800 156.390 ;
        RECT 80.400 156.330 80.720 156.390 ;
        RECT 82.255 156.330 82.545 156.375 ;
        RECT 80.400 156.190 82.545 156.330 ;
        RECT 84.630 156.330 84.770 156.825 ;
        RECT 85.935 156.330 86.225 156.375 ;
        RECT 84.630 156.190 86.225 156.330 ;
        RECT 80.400 156.130 80.720 156.190 ;
        RECT 82.255 156.145 82.545 156.190 ;
        RECT 85.935 156.145 86.225 156.190 ;
        RECT 74.870 155.990 75.160 156.035 ;
        RECT 71.610 155.850 75.160 155.990 ;
        RECT 71.610 155.805 71.900 155.850 ;
        RECT 73.960 155.790 74.280 155.850 ;
        RECT 74.870 155.805 75.160 155.850 ;
        RECT 75.790 155.990 76.080 156.035 ;
        RECT 77.650 155.990 77.940 156.035 ;
        RECT 75.790 155.850 77.940 155.990 ;
        RECT 79.570 155.990 79.710 156.130 ;
        RECT 84.080 155.990 84.400 156.050 ;
        RECT 88.770 155.990 88.910 157.150 ;
        RECT 96.500 157.010 96.820 157.070 ;
        RECT 96.500 156.870 102.250 157.010 ;
        RECT 96.500 156.810 96.820 156.870 ;
        RECT 90.520 156.670 90.840 156.730 ;
        RECT 90.520 156.530 92.130 156.670 ;
        RECT 90.520 156.470 90.840 156.530 ;
        RECT 91.990 156.375 92.130 156.530 ;
        RECT 96.130 156.530 101.790 156.670 ;
        RECT 96.130 156.390 96.270 156.530 ;
        RECT 90.995 156.145 91.285 156.375 ;
        RECT 91.915 156.145 92.205 156.375 ;
        RECT 79.570 155.850 88.910 155.990 ;
        RECT 90.520 155.990 90.840 156.050 ;
        RECT 91.070 155.990 91.210 156.145 ;
        RECT 92.360 156.130 92.680 156.390 ;
        RECT 92.820 156.330 93.140 156.390 ;
        RECT 96.040 156.330 96.360 156.390 ;
        RECT 92.820 156.190 96.360 156.330 ;
        RECT 92.820 156.130 93.140 156.190 ;
        RECT 96.040 156.130 96.360 156.190 ;
        RECT 97.880 156.130 98.200 156.390 ;
        RECT 98.355 156.145 98.645 156.375 ;
        RECT 92.450 155.990 92.590 156.130 ;
        RECT 90.520 155.850 91.210 155.990 ;
        RECT 91.990 155.850 92.590 155.990 ;
        RECT 97.420 155.990 97.740 156.050 ;
        RECT 98.430 155.990 98.570 156.145 ;
        RECT 98.800 156.130 99.120 156.390 ;
        RECT 99.735 156.330 100.025 156.375 ;
        RECT 100.640 156.330 100.960 156.390 ;
        RECT 101.650 156.375 101.790 156.530 ;
        RECT 102.110 156.375 102.250 156.870 ;
        RECT 99.735 156.190 100.960 156.330 ;
        RECT 99.735 156.145 100.025 156.190 ;
        RECT 100.640 156.130 100.960 156.190 ;
        RECT 101.575 156.145 101.865 156.375 ;
        RECT 102.035 156.145 102.325 156.375 ;
        RECT 102.480 156.130 102.800 156.390 ;
        RECT 102.940 156.330 103.260 156.390 ;
        RECT 104.410 156.375 104.550 157.210 ;
        RECT 103.415 156.330 103.705 156.375 ;
        RECT 102.940 156.190 103.705 156.330 ;
        RECT 102.940 156.130 103.260 156.190 ;
        RECT 103.415 156.145 103.705 156.190 ;
        RECT 104.335 156.330 104.625 156.375 ;
        RECT 105.700 156.330 106.020 156.390 ;
        RECT 107.080 156.330 107.400 156.390 ;
        RECT 104.335 156.190 107.400 156.330 ;
        RECT 104.335 156.145 104.625 156.190 ;
        RECT 105.700 156.130 106.020 156.190 ;
        RECT 107.080 156.130 107.400 156.190 ;
        RECT 107.555 156.145 107.845 156.375 ;
        RECT 97.420 155.850 98.570 155.990 ;
        RECT 103.860 155.990 104.180 156.050 ;
        RECT 107.630 155.990 107.770 156.145 ;
        RECT 103.860 155.850 107.770 155.990 ;
        RECT 75.790 155.805 76.080 155.850 ;
        RECT 77.650 155.805 77.940 155.850 ;
        RECT 84.080 155.790 84.400 155.850 ;
        RECT 90.520 155.790 90.840 155.850 ;
        RECT 67.520 155.650 67.840 155.710 ;
        RECT 50.130 155.510 67.840 155.650 ;
        RECT 42.220 155.450 42.540 155.510 ;
        RECT 43.600 155.450 43.920 155.510 ;
        RECT 67.520 155.450 67.840 155.510 ;
        RECT 82.715 155.650 83.005 155.695 ;
        RECT 84.540 155.650 84.860 155.710 ;
        RECT 87.300 155.650 87.620 155.710 ;
        RECT 82.715 155.510 87.620 155.650 ;
        RECT 82.715 155.465 83.005 155.510 ;
        RECT 84.540 155.450 84.860 155.510 ;
        RECT 87.300 155.450 87.620 155.510 ;
        RECT 87.760 155.650 88.080 155.710 ;
        RECT 91.990 155.650 92.130 155.850 ;
        RECT 97.420 155.790 97.740 155.850 ;
        RECT 103.860 155.790 104.180 155.850 ;
        RECT 87.760 155.510 92.130 155.650 ;
        RECT 94.215 155.650 94.505 155.695 ;
        RECT 95.580 155.650 95.900 155.710 ;
        RECT 94.215 155.510 95.900 155.650 ;
        RECT 87.760 155.450 88.080 155.510 ;
        RECT 94.215 155.465 94.505 155.510 ;
        RECT 95.580 155.450 95.900 155.510 ;
        RECT 96.500 155.450 96.820 155.710 ;
        RECT 100.180 155.450 100.500 155.710 ;
        RECT 104.780 155.450 105.100 155.710 ;
        RECT 106.160 155.450 106.480 155.710 ;
        RECT 108.460 155.450 108.780 155.710 ;
        RECT 11.330 154.830 113.450 155.310 ;
        RECT 16.935 154.445 17.225 154.675 ;
        RECT 17.840 154.630 18.160 154.690 ;
        RECT 19.235 154.630 19.525 154.675 ;
        RECT 21.520 154.630 21.840 154.690 ;
        RECT 32.575 154.630 32.865 154.675 ;
        RECT 35.320 154.630 35.640 154.690 ;
        RECT 38.540 154.630 38.860 154.690 ;
        RECT 17.840 154.490 29.570 154.630 ;
        RECT 14.160 153.750 14.480 154.010 ;
        RECT 16.475 153.950 16.765 153.995 ;
        RECT 17.010 153.950 17.150 154.445 ;
        RECT 17.840 154.430 18.160 154.490 ;
        RECT 19.235 154.445 19.525 154.490 ;
        RECT 21.520 154.430 21.840 154.490 ;
        RECT 18.300 154.290 18.620 154.350 ;
        RECT 18.300 154.150 27.270 154.290 ;
        RECT 18.300 154.090 18.620 154.150 ;
        RECT 16.475 153.810 17.150 153.950 ;
        RECT 18.775 153.950 19.065 153.995 ;
        RECT 21.060 153.950 21.380 154.010 ;
        RECT 18.775 153.810 21.380 153.950 ;
        RECT 16.475 153.765 16.765 153.810 ;
        RECT 18.775 153.765 19.065 153.810 ;
        RECT 21.060 153.750 21.380 153.810 ;
        RECT 24.295 153.950 24.585 153.995 ;
        RECT 24.740 153.950 25.060 154.010 ;
        RECT 27.130 153.995 27.270 154.150 ;
        RECT 24.295 153.810 25.060 153.950 ;
        RECT 24.295 153.765 24.585 153.810 ;
        RECT 24.740 153.750 25.060 153.810 ;
        RECT 26.135 153.765 26.425 153.995 ;
        RECT 26.595 153.765 26.885 153.995 ;
        RECT 27.055 153.765 27.345 153.995 ;
        RECT 27.975 153.950 28.265 153.995 ;
        RECT 28.420 153.950 28.740 154.010 ;
        RECT 29.430 153.995 29.570 154.490 ;
        RECT 32.575 154.490 35.640 154.630 ;
        RECT 32.575 154.445 32.865 154.490 ;
        RECT 35.320 154.430 35.640 154.490 ;
        RECT 36.100 154.490 38.860 154.630 ;
        RECT 36.100 154.290 36.240 154.490 ;
        RECT 38.540 154.430 38.860 154.490 ;
        RECT 40.840 154.430 41.160 154.690 ;
        RECT 52.800 154.630 53.120 154.690 ;
        RECT 54.640 154.630 54.960 154.690 ;
        RECT 42.310 154.490 54.960 154.630 ;
        RECT 39.460 154.290 39.780 154.350 ;
        RECT 34.950 154.150 36.240 154.290 ;
        RECT 36.790 154.150 39.780 154.290 ;
        RECT 34.950 154.010 35.090 154.150 ;
        RECT 27.975 153.810 28.740 153.950 ;
        RECT 27.975 153.765 28.265 153.810 ;
        RECT 20.140 153.410 20.460 153.670 ;
        RECT 26.210 153.270 26.350 153.765 ;
        RECT 26.670 153.610 26.810 153.765 ;
        RECT 28.420 153.750 28.740 153.810 ;
        RECT 29.355 153.765 29.645 153.995 ;
        RECT 29.800 153.750 30.120 154.010 ;
        RECT 30.260 153.950 30.580 154.010 ;
        RECT 31.180 153.950 31.500 154.010 ;
        RECT 30.260 153.810 31.500 153.950 ;
        RECT 30.260 153.750 30.580 153.810 ;
        RECT 31.180 153.750 31.500 153.810 ;
        RECT 31.640 153.950 31.960 154.010 ;
        RECT 32.115 153.950 32.405 153.995 ;
        RECT 31.640 153.810 32.405 153.950 ;
        RECT 31.640 153.750 31.960 153.810 ;
        RECT 32.115 153.765 32.405 153.810 ;
        RECT 33.495 153.950 33.785 153.995 ;
        RECT 33.940 153.950 34.260 154.010 ;
        RECT 33.495 153.810 34.260 153.950 ;
        RECT 33.495 153.765 33.785 153.810 ;
        RECT 33.940 153.750 34.260 153.810 ;
        RECT 34.415 153.765 34.705 153.995 ;
        RECT 29.890 153.610 30.030 153.750 ;
        RECT 34.490 153.610 34.630 153.765 ;
        RECT 34.860 153.750 35.180 154.010 ;
        RECT 35.335 153.950 35.625 153.995 ;
        RECT 36.240 153.950 36.560 154.010 ;
        RECT 36.790 153.950 36.930 154.150 ;
        RECT 35.335 153.810 36.930 153.950 ;
        RECT 35.335 153.765 35.625 153.810 ;
        RECT 36.240 153.750 36.560 153.810 ;
        RECT 37.175 153.765 37.465 153.995 ;
        RECT 37.250 153.610 37.390 153.765 ;
        RECT 38.080 153.750 38.400 154.010 ;
        RECT 38.540 153.750 38.860 154.010 ;
        RECT 39.090 153.995 39.230 154.150 ;
        RECT 39.460 154.090 39.780 154.150 ;
        RECT 39.015 153.765 39.305 153.995 ;
        RECT 40.380 153.950 40.700 154.010 ;
        RECT 42.310 153.995 42.450 154.490 ;
        RECT 52.800 154.430 53.120 154.490 ;
        RECT 54.640 154.430 54.960 154.490 ;
        RECT 55.560 154.430 55.880 154.690 ;
        RECT 64.760 154.430 65.080 154.690 ;
        RECT 67.520 154.630 67.840 154.690 ;
        RECT 71.660 154.630 71.980 154.690 ;
        RECT 67.520 154.490 71.980 154.630 ;
        RECT 67.520 154.430 67.840 154.490 ;
        RECT 71.660 154.430 71.980 154.490 ;
        RECT 73.515 154.630 73.805 154.675 ;
        RECT 73.960 154.630 74.280 154.690 ;
        RECT 100.180 154.630 100.500 154.690 ;
        RECT 73.515 154.490 74.280 154.630 ;
        RECT 73.515 154.445 73.805 154.490 ;
        RECT 73.960 154.430 74.280 154.490 ;
        RECT 91.070 154.490 100.500 154.630 ;
        RECT 47.740 154.290 48.060 154.350 ;
        RECT 50.975 154.290 51.265 154.335 ;
        RECT 43.690 154.150 51.265 154.290 ;
        RECT 40.380 153.810 41.990 153.950 ;
        RECT 40.380 153.750 40.700 153.810 ;
        RECT 40.840 153.610 41.160 153.670 ;
        RECT 26.670 153.470 30.030 153.610 ;
        RECT 30.350 153.470 34.630 153.610 ;
        RECT 36.100 153.470 41.160 153.610 ;
        RECT 41.850 153.610 41.990 153.810 ;
        RECT 42.235 153.765 42.525 153.995 ;
        RECT 42.695 153.765 42.985 153.995 ;
        RECT 43.260 153.950 43.550 153.995 ;
        RECT 43.690 153.950 43.830 154.150 ;
        RECT 47.740 154.090 48.060 154.150 ;
        RECT 50.975 154.105 51.265 154.150 ;
        RECT 64.850 154.290 64.990 154.430 ;
        RECT 72.120 154.290 72.440 154.350 ;
        RECT 64.850 154.150 65.975 154.290 ;
        RECT 43.260 153.810 43.830 153.950 ;
        RECT 43.260 153.765 43.550 153.810 ;
        RECT 42.770 153.610 42.910 153.765 ;
        RECT 44.060 153.750 44.380 154.010 ;
        RECT 53.260 153.950 53.580 154.010 ;
        RECT 44.610 153.810 53.580 153.950 ;
        RECT 44.610 153.610 44.750 153.810 ;
        RECT 53.260 153.750 53.580 153.810 ;
        RECT 62.000 153.750 62.320 154.010 ;
        RECT 41.850 153.470 42.450 153.610 ;
        RECT 42.770 153.470 44.750 153.610 ;
        RECT 44.995 153.610 45.285 153.655 ;
        RECT 45.900 153.610 46.220 153.670 ;
        RECT 44.995 153.470 46.220 153.610 ;
        RECT 28.420 153.270 28.740 153.330 ;
        RECT 30.350 153.270 30.490 153.470 ;
        RECT 26.210 153.130 26.810 153.270 ;
        RECT 14.620 152.730 14.940 152.990 ;
        RECT 15.540 152.730 15.860 152.990 ;
        RECT 23.820 152.730 24.140 152.990 ;
        RECT 24.755 152.930 25.045 152.975 ;
        RECT 25.200 152.930 25.520 152.990 ;
        RECT 24.755 152.790 25.520 152.930 ;
        RECT 26.670 152.930 26.810 153.130 ;
        RECT 28.420 153.130 30.490 153.270 ;
        RECT 32.560 153.270 32.880 153.330 ;
        RECT 33.940 153.270 34.260 153.330 ;
        RECT 36.100 153.270 36.240 153.470 ;
        RECT 40.840 153.410 41.160 153.470 ;
        RECT 32.560 153.130 36.240 153.270 ;
        RECT 40.930 153.270 41.070 153.410 ;
        RECT 41.760 153.270 42.080 153.330 ;
        RECT 40.930 153.130 42.080 153.270 ;
        RECT 42.310 153.270 42.450 153.470 ;
        RECT 44.995 153.425 45.285 153.470 ;
        RECT 45.900 153.410 46.220 153.470 ;
        RECT 47.755 153.610 48.045 153.655 ;
        RECT 51.435 153.610 51.725 153.655 ;
        RECT 51.880 153.610 52.200 153.670 ;
        RECT 47.755 153.470 52.200 153.610 ;
        RECT 47.755 153.425 48.045 153.470 ;
        RECT 51.435 153.425 51.725 153.470 ;
        RECT 51.880 153.410 52.200 153.470 ;
        RECT 52.340 153.610 52.660 153.670 ;
        RECT 56.480 153.610 56.800 153.670 ;
        RECT 52.340 153.470 56.800 153.610 ;
        RECT 52.340 153.410 52.660 153.470 ;
        RECT 56.480 153.410 56.800 153.470 ;
        RECT 64.850 153.270 64.990 154.150 ;
        RECT 65.835 153.995 65.975 154.150 ;
        RECT 66.230 154.150 72.440 154.290 ;
        RECT 66.230 153.995 66.370 154.150 ;
        RECT 72.120 154.090 72.440 154.150 ;
        RECT 74.420 154.290 74.740 154.350 ;
        RECT 74.420 154.150 88.450 154.290 ;
        RECT 74.420 154.090 74.740 154.150 ;
        RECT 65.135 153.950 65.425 153.995 ;
        RECT 65.135 153.765 65.450 153.950 ;
        RECT 65.695 153.765 65.985 153.995 ;
        RECT 66.155 153.765 66.445 153.995 ;
        RECT 67.075 153.950 67.365 153.995 ;
        RECT 67.520 153.950 67.840 154.010 ;
        RECT 67.075 153.810 67.840 153.950 ;
        RECT 67.075 153.765 67.365 153.810 ;
        RECT 42.310 153.130 64.990 153.270 ;
        RECT 65.310 153.270 65.450 153.765 ;
        RECT 65.835 153.610 65.975 153.765 ;
        RECT 67.520 153.750 67.840 153.810 ;
        RECT 68.440 153.750 68.760 154.010 ;
        RECT 69.820 153.995 70.140 154.010 ;
        RECT 68.915 153.765 69.205 153.995 ;
        RECT 69.605 153.765 70.140 153.995 ;
        RECT 73.975 153.950 74.265 153.995 ;
        RECT 79.480 153.950 79.800 154.010 ;
        RECT 73.975 153.810 79.800 153.950 ;
        RECT 86.395 153.940 86.685 153.995 ;
        RECT 73.975 153.765 74.265 153.810 ;
        RECT 68.990 153.610 69.130 153.765 ;
        RECT 69.820 153.750 70.140 153.765 ;
        RECT 79.480 153.750 79.800 153.810 ;
        RECT 86.370 153.765 86.685 153.940 ;
        RECT 86.855 153.765 87.145 153.995 ;
        RECT 65.835 153.470 69.130 153.610 ;
        RECT 65.310 153.130 65.910 153.270 ;
        RECT 28.420 153.070 28.740 153.130 ;
        RECT 32.560 153.070 32.880 153.130 ;
        RECT 33.940 153.070 34.260 153.130 ;
        RECT 41.760 153.070 42.080 153.130 ;
        RECT 29.800 152.930 30.120 152.990 ;
        RECT 26.670 152.790 30.120 152.930 ;
        RECT 24.755 152.745 25.045 152.790 ;
        RECT 25.200 152.730 25.520 152.790 ;
        RECT 29.800 152.730 30.120 152.790 ;
        RECT 30.260 152.930 30.580 152.990 ;
        RECT 31.655 152.930 31.945 152.975 ;
        RECT 30.260 152.790 31.945 152.930 ;
        RECT 30.260 152.730 30.580 152.790 ;
        RECT 31.655 152.745 31.945 152.790 ;
        RECT 36.715 152.930 37.005 152.975 ;
        RECT 37.160 152.930 37.480 152.990 ;
        RECT 36.715 152.790 37.480 152.930 ;
        RECT 36.715 152.745 37.005 152.790 ;
        RECT 37.160 152.730 37.480 152.790 ;
        RECT 40.395 152.930 40.685 152.975 ;
        RECT 42.680 152.930 43.000 152.990 ;
        RECT 40.395 152.790 43.000 152.930 ;
        RECT 40.395 152.745 40.685 152.790 ;
        RECT 42.680 152.730 43.000 152.790 ;
        RECT 49.135 152.930 49.425 152.975 ;
        RECT 49.580 152.930 49.900 152.990 ;
        RECT 49.135 152.790 49.900 152.930 ;
        RECT 49.135 152.745 49.425 152.790 ;
        RECT 49.580 152.730 49.900 152.790 ;
        RECT 63.855 152.930 64.145 152.975 ;
        RECT 64.760 152.930 65.080 152.990 ;
        RECT 63.855 152.790 65.080 152.930 ;
        RECT 65.770 152.930 65.910 153.130 ;
        RECT 67.980 152.930 68.300 152.990 ;
        RECT 65.770 152.790 68.300 152.930 ;
        RECT 68.990 152.930 69.130 153.470 ;
        RECT 86.370 153.270 86.510 153.765 ;
        RECT 86.930 153.610 87.070 153.765 ;
        RECT 87.300 153.750 87.620 154.010 ;
        RECT 88.310 153.995 88.450 154.150 ;
        RECT 91.070 153.995 91.210 154.490 ;
        RECT 100.180 154.430 100.500 154.490 ;
        RECT 92.375 154.290 92.665 154.335 ;
        RECT 96.500 154.290 96.820 154.350 ;
        RECT 92.375 154.150 96.820 154.290 ;
        RECT 92.375 154.105 92.665 154.150 ;
        RECT 96.500 154.090 96.820 154.150 ;
        RECT 103.975 154.290 104.265 154.335 ;
        RECT 104.780 154.290 105.100 154.350 ;
        RECT 107.215 154.290 107.865 154.335 ;
        RECT 103.975 154.150 107.865 154.290 ;
        RECT 103.975 154.105 104.565 154.150 ;
        RECT 88.235 153.765 88.525 153.995 ;
        RECT 90.995 153.765 91.285 153.995 ;
        RECT 87.760 153.610 88.080 153.670 ;
        RECT 86.930 153.470 88.080 153.610 ;
        RECT 88.310 153.610 88.450 153.765 ;
        RECT 91.440 153.750 91.760 154.010 ;
        RECT 92.835 153.765 93.125 153.995 ;
        RECT 90.520 153.610 90.840 153.670 ;
        RECT 92.910 153.610 93.050 153.765 ;
        RECT 93.740 153.750 94.060 154.010 ;
        RECT 94.200 153.750 94.520 154.010 ;
        RECT 94.675 153.950 94.965 153.995 ;
        RECT 96.040 153.950 96.360 154.010 ;
        RECT 94.675 153.810 96.360 153.950 ;
        RECT 94.675 153.765 94.965 153.810 ;
        RECT 94.750 153.610 94.890 153.765 ;
        RECT 96.040 153.750 96.360 153.810 ;
        RECT 104.275 153.790 104.565 154.105 ;
        RECT 104.780 154.090 105.100 154.150 ;
        RECT 107.215 154.105 107.865 154.150 ;
        RECT 108.460 154.290 108.780 154.350 ;
        RECT 109.855 154.290 110.145 154.335 ;
        RECT 108.460 154.150 110.145 154.290 ;
        RECT 108.460 154.090 108.780 154.150 ;
        RECT 109.855 154.105 110.145 154.150 ;
        RECT 105.355 153.950 105.645 153.995 ;
        RECT 108.935 153.950 109.225 153.995 ;
        RECT 110.770 153.950 111.060 153.995 ;
        RECT 105.355 153.810 111.060 153.950 ;
        RECT 105.355 153.765 105.645 153.810 ;
        RECT 108.935 153.765 109.225 153.810 ;
        RECT 110.770 153.765 111.060 153.810 ;
        RECT 88.310 153.470 93.050 153.610 ;
        RECT 94.290 153.470 94.890 153.610 ;
        RECT 96.975 153.610 97.265 153.655 ;
        RECT 98.800 153.610 99.120 153.670 ;
        RECT 102.495 153.610 102.785 153.655 ;
        RECT 96.975 153.470 102.785 153.610 ;
        RECT 87.760 153.410 88.080 153.470 ;
        RECT 90.520 153.410 90.840 153.470 ;
        RECT 94.290 153.270 94.430 153.470 ;
        RECT 96.975 153.425 97.265 153.470 ;
        RECT 98.800 153.410 99.120 153.470 ;
        RECT 102.495 153.425 102.785 153.470 ;
        RECT 111.235 153.610 111.525 153.655 ;
        RECT 111.680 153.610 112.000 153.670 ;
        RECT 111.235 153.470 112.000 153.610 ;
        RECT 111.235 153.425 111.525 153.470 ;
        RECT 111.680 153.410 112.000 153.470 ;
        RECT 102.020 153.270 102.340 153.330 ;
        RECT 70.370 153.130 94.430 153.270 ;
        RECT 95.670 153.130 102.340 153.270 ;
        RECT 70.370 152.990 70.510 153.130 ;
        RECT 69.360 152.930 69.680 152.990 ;
        RECT 68.990 152.790 69.680 152.930 ;
        RECT 63.855 152.745 64.145 152.790 ;
        RECT 64.760 152.730 65.080 152.790 ;
        RECT 67.980 152.730 68.300 152.790 ;
        RECT 69.360 152.730 69.680 152.790 ;
        RECT 70.280 152.730 70.600 152.990 ;
        RECT 70.740 152.730 71.060 152.990 ;
        RECT 85.015 152.930 85.305 152.975 ;
        RECT 85.920 152.930 86.240 152.990 ;
        RECT 85.015 152.790 86.240 152.930 ;
        RECT 85.015 152.745 85.305 152.790 ;
        RECT 85.920 152.730 86.240 152.790 ;
        RECT 89.140 152.930 89.460 152.990 ;
        RECT 90.075 152.930 90.365 152.975 ;
        RECT 89.140 152.790 90.365 152.930 ;
        RECT 89.140 152.730 89.460 152.790 ;
        RECT 90.075 152.745 90.365 152.790 ;
        RECT 92.360 152.730 92.680 152.990 ;
        RECT 93.740 152.930 94.060 152.990 ;
        RECT 95.670 152.930 95.810 153.130 ;
        RECT 102.020 153.070 102.340 153.130 ;
        RECT 105.355 153.270 105.645 153.315 ;
        RECT 108.475 153.270 108.765 153.315 ;
        RECT 110.365 153.270 110.655 153.315 ;
        RECT 105.355 153.130 110.655 153.270 ;
        RECT 105.355 153.085 105.645 153.130 ;
        RECT 108.475 153.085 108.765 153.130 ;
        RECT 110.365 153.085 110.655 153.130 ;
        RECT 93.740 152.790 95.810 152.930 ;
        RECT 93.740 152.730 94.060 152.790 ;
        RECT 96.040 152.730 96.360 152.990 ;
        RECT 99.720 152.730 100.040 152.990 ;
        RECT 11.330 152.110 113.450 152.590 ;
        RECT 21.520 151.955 21.840 151.970 ;
        RECT 21.520 151.725 22.055 151.955 ;
        RECT 27.040 151.910 27.360 151.970 ;
        RECT 31.640 151.910 31.960 151.970 ;
        RECT 27.040 151.770 31.960 151.910 ;
        RECT 21.520 151.710 21.840 151.725 ;
        RECT 27.040 151.710 27.360 151.770 ;
        RECT 31.640 151.710 31.960 151.770 ;
        RECT 34.860 151.910 35.180 151.970 ;
        RECT 42.220 151.910 42.540 151.970 ;
        RECT 43.600 151.910 43.920 151.970 ;
        RECT 34.860 151.770 40.150 151.910 ;
        RECT 34.860 151.710 35.180 151.770 ;
        RECT 13.260 151.570 13.550 151.615 ;
        RECT 15.120 151.570 15.410 151.615 ;
        RECT 17.900 151.570 18.190 151.615 ;
        RECT 13.260 151.430 18.190 151.570 ;
        RECT 13.260 151.385 13.550 151.430 ;
        RECT 15.120 151.385 15.410 151.430 ;
        RECT 17.900 151.385 18.190 151.430 ;
        RECT 25.775 151.570 26.065 151.615 ;
        RECT 28.895 151.570 29.185 151.615 ;
        RECT 30.785 151.570 31.075 151.615 ;
        RECT 33.020 151.570 33.340 151.630 ;
        RECT 25.775 151.430 31.075 151.570 ;
        RECT 25.775 151.385 26.065 151.430 ;
        RECT 28.895 151.385 29.185 151.430 ;
        RECT 30.785 151.385 31.075 151.430 ;
        RECT 31.270 151.430 32.330 151.570 ;
        RECT 14.635 151.230 14.925 151.275 ;
        RECT 15.540 151.230 15.860 151.290 ;
        RECT 14.635 151.090 15.860 151.230 ;
        RECT 14.635 151.045 14.925 151.090 ;
        RECT 15.540 151.030 15.860 151.090 ;
        RECT 21.060 151.230 21.380 151.290 ;
        RECT 31.270 151.230 31.410 151.430 ;
        RECT 21.060 151.090 31.410 151.230 ;
        RECT 21.060 151.030 21.380 151.090 ;
        RECT 31.640 151.030 31.960 151.290 ;
        RECT 32.190 151.230 32.330 151.430 ;
        RECT 33.020 151.430 37.390 151.570 ;
        RECT 33.020 151.370 33.340 151.430 ;
        RECT 32.190 151.090 33.250 151.230 ;
        RECT 12.795 150.890 13.085 150.935 ;
        RECT 13.240 150.890 13.560 150.950 ;
        RECT 17.900 150.890 18.190 150.935 ;
        RECT 12.795 150.750 13.560 150.890 ;
        RECT 12.795 150.705 13.085 150.750 ;
        RECT 13.240 150.690 13.560 150.750 ;
        RECT 15.655 150.750 18.190 150.890 ;
        RECT 15.655 150.595 15.870 150.750 ;
        RECT 17.900 150.705 18.190 150.750 ;
        RECT 13.720 150.550 14.010 150.595 ;
        RECT 15.580 150.550 15.870 150.595 ;
        RECT 16.500 150.550 16.790 150.595 ;
        RECT 19.760 150.550 20.050 150.595 ;
        RECT 13.720 150.410 15.870 150.550 ;
        RECT 13.720 150.365 14.010 150.410 ;
        RECT 15.580 150.365 15.870 150.410 ;
        RECT 16.090 150.410 20.050 150.550 ;
        RECT 14.620 150.210 14.940 150.270 ;
        RECT 16.090 150.210 16.230 150.410 ;
        RECT 16.500 150.365 16.790 150.410 ;
        RECT 19.760 150.365 20.050 150.410 ;
        RECT 23.820 150.550 24.140 150.610 ;
        RECT 24.695 150.595 24.985 150.910 ;
        RECT 25.775 150.890 26.065 150.935 ;
        RECT 29.355 150.890 29.645 150.935 ;
        RECT 31.190 150.890 31.480 150.935 ;
        RECT 25.775 150.750 31.480 150.890 ;
        RECT 25.775 150.705 26.065 150.750 ;
        RECT 29.355 150.705 29.645 150.750 ;
        RECT 31.190 150.705 31.480 150.750 ;
        RECT 32.115 150.890 32.405 150.935 ;
        RECT 32.560 150.890 32.880 150.950 ;
        RECT 33.110 150.935 33.250 151.090 ;
        RECT 32.115 150.750 32.880 150.890 ;
        RECT 32.115 150.705 32.405 150.750 ;
        RECT 32.560 150.690 32.880 150.750 ;
        RECT 33.035 150.705 33.325 150.935 ;
        RECT 33.480 150.690 33.800 150.950 ;
        RECT 33.940 150.690 34.260 150.950 ;
        RECT 37.250 150.935 37.390 151.430 ;
        RECT 40.010 151.275 40.150 151.770 ;
        RECT 42.220 151.770 43.920 151.910 ;
        RECT 42.220 151.710 42.540 151.770 ;
        RECT 43.600 151.710 43.920 151.770 ;
        RECT 44.060 151.910 44.380 151.970 ;
        RECT 53.260 151.910 53.580 151.970 ;
        RECT 44.060 151.770 53.580 151.910 ;
        RECT 44.060 151.710 44.380 151.770 ;
        RECT 53.260 151.710 53.580 151.770 ;
        RECT 54.640 151.910 54.960 151.970 ;
        RECT 59.715 151.910 60.005 151.955 ;
        RECT 60.160 151.910 60.480 151.970 ;
        RECT 67.075 151.910 67.365 151.955 ;
        RECT 67.980 151.910 68.300 151.970 ;
        RECT 91.440 151.910 91.760 151.970 ;
        RECT 92.375 151.910 92.665 151.955 ;
        RECT 97.420 151.910 97.740 151.970 ;
        RECT 54.640 151.770 59.470 151.910 ;
        RECT 54.640 151.710 54.960 151.770 ;
        RECT 47.855 151.570 48.145 151.615 ;
        RECT 50.975 151.570 51.265 151.615 ;
        RECT 52.865 151.570 53.155 151.615 ;
        RECT 57.860 151.570 58.180 151.630 ;
        RECT 47.855 151.430 53.155 151.570 ;
        RECT 47.855 151.385 48.145 151.430 ;
        RECT 50.975 151.385 51.265 151.430 ;
        RECT 52.865 151.385 53.155 151.430 ;
        RECT 53.810 151.430 58.180 151.570 ;
        RECT 59.330 151.570 59.470 151.770 ;
        RECT 59.715 151.770 60.480 151.910 ;
        RECT 59.715 151.725 60.005 151.770 ;
        RECT 60.160 151.710 60.480 151.770 ;
        RECT 66.690 151.770 67.750 151.910 ;
        RECT 66.690 151.570 66.830 151.770 ;
        RECT 67.075 151.725 67.365 151.770 ;
        RECT 59.330 151.430 66.830 151.570 ;
        RECT 67.610 151.570 67.750 151.770 ;
        RECT 67.980 151.770 91.210 151.910 ;
        RECT 67.980 151.710 68.300 151.770 ;
        RECT 72.580 151.570 72.900 151.630 ;
        RECT 67.610 151.430 72.900 151.570 ;
        RECT 91.070 151.570 91.210 151.770 ;
        RECT 91.440 151.770 92.665 151.910 ;
        RECT 91.440 151.710 91.760 151.770 ;
        RECT 92.375 151.725 92.665 151.770 ;
        RECT 93.830 151.770 97.740 151.910 ;
        RECT 93.830 151.570 93.970 151.770 ;
        RECT 97.420 151.710 97.740 151.770 ;
        RECT 97.895 151.910 98.185 151.955 ;
        RECT 98.340 151.910 98.660 151.970 ;
        RECT 105.700 151.910 106.020 151.970 ;
        RECT 97.895 151.770 98.660 151.910 ;
        RECT 97.895 151.725 98.185 151.770 ;
        RECT 98.340 151.710 98.660 151.770 ;
        RECT 99.810 151.770 106.020 151.910 ;
        RECT 91.070 151.430 93.970 151.570 ;
        RECT 39.935 151.045 40.225 151.275 ;
        RECT 40.855 151.230 41.145 151.275 ;
        RECT 43.140 151.230 43.460 151.290 ;
        RECT 53.810 151.275 53.950 151.430 ;
        RECT 57.860 151.370 58.180 151.430 ;
        RECT 72.580 151.370 72.900 151.430 ;
        RECT 40.855 151.090 43.460 151.230 ;
        RECT 40.855 151.045 41.145 151.090 ;
        RECT 43.140 151.030 43.460 151.090 ;
        RECT 53.735 151.045 54.025 151.275 ;
        RECT 56.480 151.230 56.800 151.290 ;
        RECT 56.955 151.230 57.245 151.275 ;
        RECT 62.475 151.230 62.765 151.275 ;
        RECT 67.060 151.230 67.380 151.290 ;
        RECT 56.480 151.090 62.765 151.230 ;
        RECT 56.480 151.030 56.800 151.090 ;
        RECT 56.955 151.045 57.245 151.090 ;
        RECT 62.475 151.045 62.765 151.090 ;
        RECT 66.230 151.090 67.380 151.230 ;
        RECT 37.175 150.705 37.465 150.935 ;
        RECT 38.540 150.890 38.860 150.950 ;
        RECT 40.380 150.890 40.700 150.950 ;
        RECT 38.540 150.750 40.700 150.890 ;
        RECT 38.540 150.690 38.860 150.750 ;
        RECT 40.380 150.690 40.700 150.750 ;
        RECT 24.395 150.550 24.985 150.595 ;
        RECT 27.635 150.550 28.285 150.595 ;
        RECT 30.275 150.550 30.565 150.595 ;
        RECT 23.820 150.410 28.285 150.550 ;
        RECT 23.820 150.350 24.140 150.410 ;
        RECT 24.395 150.365 24.685 150.410 ;
        RECT 27.635 150.365 28.285 150.410 ;
        RECT 29.430 150.410 30.565 150.550 ;
        RECT 29.430 150.270 29.570 150.410 ;
        RECT 30.275 150.365 30.565 150.410 ;
        RECT 35.780 150.550 36.100 150.610 ;
        RECT 46.775 150.595 47.065 150.910 ;
        RECT 47.855 150.890 48.145 150.935 ;
        RECT 51.435 150.890 51.725 150.935 ;
        RECT 53.270 150.890 53.560 150.935 ;
        RECT 47.855 150.750 53.560 150.890 ;
        RECT 47.855 150.705 48.145 150.750 ;
        RECT 51.435 150.705 51.725 150.750 ;
        RECT 53.270 150.705 53.560 150.750 ;
        RECT 54.180 150.890 54.500 150.950 ;
        RECT 66.230 150.935 66.370 151.090 ;
        RECT 67.060 151.030 67.380 151.090 ;
        RECT 69.360 151.230 69.680 151.290 ;
        RECT 73.500 151.230 73.820 151.290 ;
        RECT 69.360 151.090 70.510 151.230 ;
        RECT 69.360 151.030 69.680 151.090 ;
        RECT 57.415 150.890 57.705 150.935 ;
        RECT 54.180 150.750 57.705 150.890 ;
        RECT 54.180 150.690 54.500 150.750 ;
        RECT 57.415 150.705 57.705 150.750 ;
        RECT 66.155 150.705 66.445 150.935 ;
        RECT 67.995 150.875 68.285 150.935 ;
        RECT 67.610 150.735 68.285 150.875 ;
        RECT 39.475 150.550 39.765 150.595 ;
        RECT 35.780 150.410 39.765 150.550 ;
        RECT 35.780 150.350 36.100 150.410 ;
        RECT 39.475 150.365 39.765 150.410 ;
        RECT 46.475 150.550 47.065 150.595 ;
        RECT 47.280 150.550 47.600 150.610 ;
        RECT 49.715 150.550 50.365 150.595 ;
        RECT 46.475 150.410 50.365 150.550 ;
        RECT 46.475 150.365 46.765 150.410 ;
        RECT 47.280 150.350 47.600 150.410 ;
        RECT 49.715 150.365 50.365 150.410 ;
        RECT 52.355 150.365 52.645 150.595 ;
        RECT 53.720 150.550 54.040 150.610 ;
        RECT 63.855 150.550 64.145 150.595 ;
        RECT 67.060 150.550 67.380 150.610 ;
        RECT 53.720 150.410 58.550 150.550 ;
        RECT 14.620 150.070 16.230 150.210 ;
        RECT 22.440 150.210 22.760 150.270 ;
        RECT 22.915 150.210 23.205 150.255 ;
        RECT 28.420 150.210 28.740 150.270 ;
        RECT 22.440 150.070 28.740 150.210 ;
        RECT 14.620 150.010 14.940 150.070 ;
        RECT 22.440 150.010 22.760 150.070 ;
        RECT 22.915 150.025 23.205 150.070 ;
        RECT 28.420 150.010 28.740 150.070 ;
        RECT 29.340 150.010 29.660 150.270 ;
        RECT 35.320 150.010 35.640 150.270 ;
        RECT 36.240 150.210 36.560 150.270 ;
        RECT 36.715 150.210 37.005 150.255 ;
        RECT 36.240 150.070 37.005 150.210 ;
        RECT 36.240 150.010 36.560 150.070 ;
        RECT 36.715 150.025 37.005 150.070 ;
        RECT 37.635 150.210 37.925 150.255 ;
        RECT 38.080 150.210 38.400 150.270 ;
        RECT 37.635 150.070 38.400 150.210 ;
        RECT 37.635 150.025 37.925 150.070 ;
        RECT 38.080 150.010 38.400 150.070 ;
        RECT 44.995 150.210 45.285 150.255 ;
        RECT 45.900 150.210 46.220 150.270 ;
        RECT 44.995 150.070 46.220 150.210 ;
        RECT 44.995 150.025 45.285 150.070 ;
        RECT 45.900 150.010 46.220 150.070 ;
        RECT 51.420 150.210 51.740 150.270 ;
        RECT 52.430 150.210 52.570 150.365 ;
        RECT 53.720 150.350 54.040 150.410 ;
        RECT 51.420 150.070 52.570 150.210 ;
        RECT 57.400 150.210 57.720 150.270 ;
        RECT 57.875 150.210 58.165 150.255 ;
        RECT 57.400 150.070 58.165 150.210 ;
        RECT 58.410 150.210 58.550 150.410 ;
        RECT 63.855 150.410 67.380 150.550 ;
        RECT 67.610 150.550 67.750 150.735 ;
        RECT 67.995 150.705 68.285 150.735 ;
        RECT 68.440 150.890 68.760 150.950 ;
        RECT 69.820 150.890 70.140 150.950 ;
        RECT 70.370 150.935 70.510 151.090 ;
        RECT 70.830 151.090 73.820 151.230 ;
        RECT 70.830 150.935 70.970 151.090 ;
        RECT 73.500 151.030 73.820 151.090 ;
        RECT 91.900 151.230 92.220 151.290 ;
        RECT 92.375 151.230 92.665 151.275 ;
        RECT 91.900 151.090 92.665 151.230 ;
        RECT 93.830 151.230 93.970 151.430 ;
        RECT 94.215 151.570 94.505 151.615 ;
        RECT 99.810 151.570 99.950 151.770 ;
        RECT 105.700 151.710 106.020 151.770 ;
        RECT 94.215 151.430 99.950 151.570 ;
        RECT 102.035 151.570 102.325 151.615 ;
        RECT 103.860 151.570 104.180 151.630 ;
        RECT 102.035 151.430 104.180 151.570 ;
        RECT 94.215 151.385 94.505 151.430 ;
        RECT 102.035 151.385 102.325 151.430 ;
        RECT 103.860 151.370 104.180 151.430 ;
        RECT 106.590 151.570 106.880 151.615 ;
        RECT 109.370 151.570 109.660 151.615 ;
        RECT 111.230 151.570 111.520 151.615 ;
        RECT 106.590 151.430 111.520 151.570 ;
        RECT 106.590 151.385 106.880 151.430 ;
        RECT 109.370 151.385 109.660 151.430 ;
        RECT 111.230 151.385 111.520 151.430 ;
        RECT 98.800 151.230 99.120 151.290 ;
        RECT 93.830 151.090 96.270 151.230 ;
        RECT 91.900 151.030 92.220 151.090 ;
        RECT 92.375 151.045 92.665 151.090 ;
        RECT 68.440 150.750 70.140 150.890 ;
        RECT 68.440 150.690 68.760 150.750 ;
        RECT 69.820 150.690 70.140 150.750 ;
        RECT 70.295 150.705 70.585 150.935 ;
        RECT 70.755 150.705 71.045 150.935 ;
        RECT 71.660 150.690 71.980 150.950 ;
        RECT 72.120 150.690 72.440 150.950 ;
        RECT 84.080 150.690 84.400 150.950 ;
        RECT 85.475 150.705 85.765 150.935 ;
        RECT 93.295 150.890 93.585 150.935 ;
        RECT 94.200 150.890 94.520 150.950 ;
        RECT 93.295 150.750 94.520 150.890 ;
        RECT 93.295 150.705 93.585 150.750 ;
        RECT 67.610 150.410 70.050 150.550 ;
        RECT 63.855 150.365 64.145 150.410 ;
        RECT 67.060 150.350 67.380 150.410 ;
        RECT 69.910 150.270 70.050 150.410 ;
        RECT 65.235 150.210 65.525 150.255 ;
        RECT 67.980 150.210 68.300 150.270 ;
        RECT 58.410 150.070 68.300 150.210 ;
        RECT 51.420 150.010 51.740 150.070 ;
        RECT 57.400 150.010 57.720 150.070 ;
        RECT 57.875 150.025 58.165 150.070 ;
        RECT 65.235 150.025 65.525 150.070 ;
        RECT 67.980 150.010 68.300 150.070 ;
        RECT 68.440 150.010 68.760 150.270 ;
        RECT 69.820 150.010 70.140 150.270 ;
        RECT 71.750 150.210 71.890 150.690 ;
        RECT 79.940 150.550 80.260 150.610 ;
        RECT 85.550 150.550 85.690 150.705 ;
        RECT 94.200 150.690 94.520 150.750 ;
        RECT 94.675 150.705 94.965 150.935 ;
        RECT 79.940 150.410 85.690 150.550 ;
        RECT 79.940 150.350 80.260 150.410 ;
        RECT 91.900 150.350 92.220 150.610 ;
        RECT 94.750 150.550 94.890 150.705 ;
        RECT 94.290 150.410 94.890 150.550 ;
        RECT 73.055 150.210 73.345 150.255 ;
        RECT 71.750 150.070 73.345 150.210 ;
        RECT 73.055 150.025 73.345 150.070 ;
        RECT 83.635 150.210 83.925 150.255 ;
        RECT 84.080 150.210 84.400 150.270 ;
        RECT 83.635 150.070 84.400 150.210 ;
        RECT 83.635 150.025 83.925 150.070 ;
        RECT 84.080 150.010 84.400 150.070 ;
        RECT 86.380 150.010 86.700 150.270 ;
        RECT 89.600 150.210 89.920 150.270 ;
        RECT 94.290 150.210 94.430 150.410 ;
        RECT 89.600 150.070 94.430 150.210 ;
        RECT 94.660 150.210 94.980 150.270 ;
        RECT 95.210 150.210 95.350 151.090 ;
        RECT 96.130 150.935 96.270 151.090 ;
        RECT 96.590 151.090 99.120 151.230 ;
        RECT 96.590 150.935 96.730 151.090 ;
        RECT 98.800 151.030 99.120 151.090 ;
        RECT 99.275 151.230 99.565 151.275 ;
        RECT 99.275 151.090 100.870 151.230 ;
        RECT 99.275 151.045 99.565 151.090 ;
        RECT 95.595 150.705 95.885 150.935 ;
        RECT 96.055 150.705 96.345 150.935 ;
        RECT 96.515 150.705 96.805 150.935 ;
        RECT 97.420 150.890 97.740 150.950 ;
        RECT 100.195 150.890 100.485 150.935 ;
        RECT 97.420 150.750 100.485 150.890 ;
        RECT 100.730 150.890 100.870 151.090 ;
        RECT 111.680 151.030 112.000 151.290 ;
        RECT 102.020 150.890 102.340 150.950 ;
        RECT 100.730 150.750 102.340 150.890 ;
        RECT 95.670 150.550 95.810 150.705 ;
        RECT 97.420 150.690 97.740 150.750 ;
        RECT 100.195 150.705 100.485 150.750 ;
        RECT 102.020 150.690 102.340 150.750 ;
        RECT 106.590 150.890 106.880 150.935 ;
        RECT 106.590 150.750 109.125 150.890 ;
        RECT 106.590 150.705 106.880 150.750 ;
        RECT 102.725 150.550 103.015 150.595 ;
        RECT 103.860 150.550 104.180 150.610 ;
        RECT 95.670 150.410 104.180 150.550 ;
        RECT 102.725 150.365 103.015 150.410 ;
        RECT 103.860 150.350 104.180 150.410 ;
        RECT 104.730 150.550 105.020 150.595 ;
        RECT 106.160 150.550 106.480 150.610 ;
        RECT 108.910 150.595 109.125 150.750 ;
        RECT 109.840 150.690 110.160 150.950 ;
        RECT 107.990 150.550 108.280 150.595 ;
        RECT 104.730 150.410 108.280 150.550 ;
        RECT 104.730 150.365 105.020 150.410 ;
        RECT 106.160 150.350 106.480 150.410 ;
        RECT 107.990 150.365 108.280 150.410 ;
        RECT 108.910 150.550 109.200 150.595 ;
        RECT 110.770 150.550 111.060 150.595 ;
        RECT 108.910 150.410 111.060 150.550 ;
        RECT 108.910 150.365 109.200 150.410 ;
        RECT 110.770 150.365 111.060 150.410 ;
        RECT 98.800 150.210 99.120 150.270 ;
        RECT 94.660 150.070 99.120 150.210 ;
        RECT 89.600 150.010 89.920 150.070 ;
        RECT 94.660 150.010 94.980 150.070 ;
        RECT 98.800 150.010 99.120 150.070 ;
        RECT 99.735 150.210 100.025 150.255 ;
        RECT 100.180 150.210 100.500 150.270 ;
        RECT 99.735 150.070 100.500 150.210 ;
        RECT 99.735 150.025 100.025 150.070 ;
        RECT 100.180 150.010 100.500 150.070 ;
        RECT 11.330 149.390 113.450 149.870 ;
        RECT 14.620 149.190 14.940 149.250 ;
        RECT 21.060 149.190 21.380 149.250 ;
        RECT 22.225 149.190 22.515 149.235 ;
        RECT 14.620 149.050 16.690 149.190 ;
        RECT 14.620 148.990 14.940 149.050 ;
        RECT 14.180 148.850 14.470 148.895 ;
        RECT 16.040 148.850 16.330 148.895 ;
        RECT 14.180 148.710 16.330 148.850 ;
        RECT 16.550 148.850 16.690 149.050 ;
        RECT 21.060 149.050 22.515 149.190 ;
        RECT 21.060 148.990 21.380 149.050 ;
        RECT 22.225 149.005 22.515 149.050 ;
        RECT 28.420 148.990 28.740 149.250 ;
        RECT 28.895 149.190 29.185 149.235 ;
        RECT 31.180 149.190 31.500 149.250 ;
        RECT 33.940 149.190 34.260 149.250 ;
        RECT 47.280 149.190 47.600 149.250 ;
        RECT 47.755 149.190 48.045 149.235 ;
        RECT 28.895 149.050 34.260 149.190 ;
        RECT 28.895 149.005 29.185 149.050 ;
        RECT 31.180 148.990 31.500 149.050 ;
        RECT 33.940 148.990 34.260 149.050 ;
        RECT 34.490 149.050 39.230 149.190 ;
        RECT 16.960 148.850 17.250 148.895 ;
        RECT 20.220 148.850 20.510 148.895 ;
        RECT 16.550 148.710 20.510 148.850 ;
        RECT 14.180 148.665 14.470 148.710 ;
        RECT 16.040 148.665 16.330 148.710 ;
        RECT 16.960 148.665 17.250 148.710 ;
        RECT 20.220 148.665 20.510 148.710 ;
        RECT 26.595 148.850 26.885 148.895 ;
        RECT 34.490 148.850 34.630 149.050 ;
        RECT 26.595 148.710 34.630 148.850 ;
        RECT 34.855 148.850 35.505 148.895 ;
        RECT 36.240 148.850 36.560 148.910 ;
        RECT 38.455 148.850 38.745 148.895 ;
        RECT 34.855 148.710 38.745 148.850 ;
        RECT 39.090 148.850 39.230 149.050 ;
        RECT 47.280 149.050 48.045 149.190 ;
        RECT 47.280 148.990 47.600 149.050 ;
        RECT 47.755 149.005 48.045 149.050 ;
        RECT 51.420 148.990 51.740 149.250 ;
        RECT 53.260 149.190 53.580 149.250 ;
        RECT 54.180 149.190 54.500 149.250 ;
        RECT 67.060 149.190 67.380 149.250 ;
        RECT 67.995 149.190 68.285 149.235 ;
        RECT 53.260 149.050 55.330 149.190 ;
        RECT 53.260 148.990 53.580 149.050 ;
        RECT 54.180 148.990 54.500 149.050 ;
        RECT 51.895 148.850 52.185 148.895 ;
        RECT 54.640 148.850 54.960 148.910 ;
        RECT 39.090 148.710 52.185 148.850 ;
        RECT 26.595 148.665 26.885 148.710 ;
        RECT 34.855 148.665 35.505 148.710 ;
        RECT 13.240 148.310 13.560 148.570 ;
        RECT 16.115 148.510 16.330 148.665 ;
        RECT 36.240 148.650 36.560 148.710 ;
        RECT 38.155 148.665 38.745 148.710 ;
        RECT 51.895 148.665 52.185 148.710 ;
        RECT 53.350 148.710 54.960 148.850 ;
        RECT 18.360 148.510 18.650 148.555 ;
        RECT 16.115 148.370 18.650 148.510 ;
        RECT 18.360 148.325 18.650 148.370 ;
        RECT 25.200 148.310 25.520 148.570 ;
        RECT 27.040 148.510 27.360 148.570 ;
        RECT 31.195 148.510 31.485 148.555 ;
        RECT 27.040 148.370 31.485 148.510 ;
        RECT 27.040 148.310 27.360 148.370 ;
        RECT 31.195 148.325 31.485 148.370 ;
        RECT 31.660 148.510 31.950 148.555 ;
        RECT 33.495 148.510 33.785 148.555 ;
        RECT 37.075 148.510 37.365 148.555 ;
        RECT 31.660 148.370 37.365 148.510 ;
        RECT 31.660 148.325 31.950 148.370 ;
        RECT 33.495 148.325 33.785 148.370 ;
        RECT 37.075 148.325 37.365 148.370 ;
        RECT 38.155 148.350 38.445 148.665 ;
        RECT 40.855 148.510 41.145 148.555 ;
        RECT 41.300 148.510 41.620 148.570 ;
        RECT 40.855 148.370 41.620 148.510 ;
        RECT 40.855 148.325 41.145 148.370 ;
        RECT 41.300 148.310 41.620 148.370 ;
        RECT 41.760 148.310 42.080 148.570 ;
        RECT 42.235 148.325 42.525 148.555 ;
        RECT 42.695 148.325 42.985 148.555 ;
        RECT 46.820 148.510 47.140 148.570 ;
        RECT 47.295 148.510 47.585 148.555 ;
        RECT 46.820 148.370 47.585 148.510 ;
        RECT 15.080 147.970 15.400 148.230 ;
        RECT 26.120 147.970 26.440 148.230 ;
        RECT 27.515 147.985 27.805 148.215 ;
        RECT 13.720 147.830 14.010 147.875 ;
        RECT 15.580 147.830 15.870 147.875 ;
        RECT 18.360 147.830 18.650 147.875 ;
        RECT 13.720 147.690 18.650 147.830 ;
        RECT 13.720 147.645 14.010 147.690 ;
        RECT 15.580 147.645 15.870 147.690 ;
        RECT 18.360 147.645 18.650 147.690 ;
        RECT 20.140 147.830 20.460 147.890 ;
        RECT 27.590 147.830 27.730 147.985 ;
        RECT 32.560 147.970 32.880 148.230 ;
        RECT 39.460 147.970 39.780 148.230 ;
        RECT 40.380 148.170 40.700 148.230 ;
        RECT 42.310 148.170 42.450 148.325 ;
        RECT 40.380 148.030 42.450 148.170 ;
        RECT 40.380 147.970 40.700 148.030 ;
        RECT 20.140 147.690 27.730 147.830 ;
        RECT 32.065 147.830 32.355 147.875 ;
        RECT 33.955 147.830 34.245 147.875 ;
        RECT 37.075 147.830 37.365 147.875 ;
        RECT 32.065 147.690 37.365 147.830 ;
        RECT 39.550 147.830 39.690 147.970 ;
        RECT 40.840 147.830 41.160 147.890 ;
        RECT 42.770 147.830 42.910 148.325 ;
        RECT 46.820 148.310 47.140 148.370 ;
        RECT 47.295 148.325 47.585 148.370 ;
        RECT 49.580 148.510 49.900 148.570 ;
        RECT 50.515 148.510 50.805 148.555 ;
        RECT 49.580 148.370 50.805 148.510 ;
        RECT 49.580 148.310 49.900 148.370 ;
        RECT 50.515 148.325 50.805 148.370 ;
        RECT 52.340 148.510 52.660 148.570 ;
        RECT 53.350 148.555 53.490 148.710 ;
        RECT 54.640 148.650 54.960 148.710 ;
        RECT 53.275 148.510 53.565 148.555 ;
        RECT 52.340 148.370 53.565 148.510 ;
        RECT 52.340 148.310 52.660 148.370 ;
        RECT 53.275 148.325 53.565 148.370 ;
        RECT 53.720 148.310 54.040 148.570 ;
        RECT 55.190 148.555 55.330 149.050 ;
        RECT 67.060 149.050 69.590 149.190 ;
        RECT 67.060 148.990 67.380 149.050 ;
        RECT 67.995 149.005 68.285 149.050 ;
        RECT 58.730 148.850 59.020 148.895 ;
        RECT 60.160 148.850 60.480 148.910 ;
        RECT 61.990 148.850 62.280 148.895 ;
        RECT 58.730 148.710 62.280 148.850 ;
        RECT 58.730 148.665 59.020 148.710 ;
        RECT 60.160 148.650 60.480 148.710 ;
        RECT 61.990 148.665 62.280 148.710 ;
        RECT 62.910 148.850 63.200 148.895 ;
        RECT 64.770 148.850 65.060 148.895 ;
        RECT 62.910 148.710 65.060 148.850 ;
        RECT 62.910 148.665 63.200 148.710 ;
        RECT 64.770 148.665 65.060 148.710 ;
        RECT 65.680 148.850 66.000 148.910 ;
        RECT 69.450 148.895 69.590 149.050 ;
        RECT 79.940 148.990 80.260 149.250 ;
        RECT 80.415 149.190 80.705 149.235 ;
        RECT 80.415 149.050 89.370 149.190 ;
        RECT 80.415 149.005 80.705 149.050 ;
        RECT 65.680 148.710 67.750 148.850 ;
        RECT 54.195 148.325 54.485 148.555 ;
        RECT 55.115 148.325 55.405 148.555 ;
        RECT 60.590 148.510 60.880 148.555 ;
        RECT 62.910 148.510 63.125 148.665 ;
        RECT 65.680 148.650 66.000 148.710 ;
        RECT 60.590 148.370 63.125 148.510 ;
        RECT 60.590 148.325 60.880 148.370 ;
        RECT 54.270 148.170 54.410 148.325 ;
        RECT 66.140 148.310 66.460 148.570 ;
        RECT 66.600 148.310 66.920 148.570 ;
        RECT 67.610 148.230 67.750 148.710 ;
        RECT 69.375 148.665 69.665 148.895 ;
        RECT 81.895 148.850 82.185 148.895 ;
        RECT 84.080 148.850 84.400 148.910 ;
        RECT 85.135 148.850 85.785 148.895 ;
        RECT 81.895 148.710 85.785 148.850 ;
        RECT 81.895 148.665 82.485 148.710 ;
        RECT 67.980 148.510 68.300 148.570 ;
        RECT 72.120 148.510 72.440 148.570 ;
        RECT 67.980 148.370 72.440 148.510 ;
        RECT 67.980 148.310 68.300 148.370 ;
        RECT 72.120 148.310 72.440 148.370 ;
        RECT 76.720 148.510 77.040 148.570 ;
        RECT 78.115 148.510 78.405 148.555 ;
        RECT 76.720 148.370 78.405 148.510 ;
        RECT 76.720 148.310 77.040 148.370 ;
        RECT 78.115 148.325 78.405 148.370 ;
        RECT 82.195 148.350 82.485 148.665 ;
        RECT 84.080 148.650 84.400 148.710 ;
        RECT 85.135 148.665 85.785 148.710 ;
        RECT 86.380 148.850 86.700 148.910 ;
        RECT 87.775 148.850 88.065 148.895 ;
        RECT 86.380 148.710 88.065 148.850 ;
        RECT 86.380 148.650 86.700 148.710 ;
        RECT 87.775 148.665 88.065 148.710 ;
        RECT 83.275 148.510 83.565 148.555 ;
        RECT 86.855 148.510 87.145 148.555 ;
        RECT 88.690 148.510 88.980 148.555 ;
        RECT 83.275 148.370 88.980 148.510 ;
        RECT 89.230 148.510 89.370 149.050 ;
        RECT 94.660 148.990 94.980 149.250 ;
        RECT 96.040 149.190 96.360 149.250 ;
        RECT 96.040 149.050 99.030 149.190 ;
        RECT 96.040 148.990 96.360 149.050 ;
        RECT 91.900 148.850 92.220 148.910 ;
        RECT 93.755 148.850 94.045 148.895 ;
        RECT 91.900 148.710 94.045 148.850 ;
        RECT 94.750 148.850 94.890 148.990 ;
        RECT 97.435 148.850 97.725 148.895 ;
        RECT 98.340 148.850 98.660 148.910 ;
        RECT 94.750 148.710 95.810 148.850 ;
        RECT 91.900 148.650 92.220 148.710 ;
        RECT 93.755 148.665 94.045 148.710 ;
        RECT 89.615 148.510 89.905 148.555 ;
        RECT 89.230 148.370 89.905 148.510 ;
        RECT 83.275 148.325 83.565 148.370 ;
        RECT 86.855 148.325 87.145 148.370 ;
        RECT 88.690 148.325 88.980 148.370 ;
        RECT 89.615 148.325 89.905 148.370 ;
        RECT 90.520 148.510 90.840 148.570 ;
        RECT 95.670 148.555 95.810 148.710 ;
        RECT 97.435 148.710 98.660 148.850 ;
        RECT 97.435 148.665 97.725 148.710 ;
        RECT 98.340 148.650 98.660 148.710 ;
        RECT 95.035 148.510 95.325 148.555 ;
        RECT 90.520 148.370 95.325 148.510 ;
        RECT 56.725 148.170 57.015 148.215 ;
        RECT 57.400 148.170 57.720 148.230 ;
        RECT 54.270 148.030 57.720 148.170 ;
        RECT 56.725 147.985 57.015 148.030 ;
        RECT 57.400 147.970 57.720 148.030 ;
        RECT 62.000 148.170 62.320 148.230 ;
        RECT 63.855 148.170 64.145 148.215 ;
        RECT 62.000 148.030 64.145 148.170 ;
        RECT 62.000 147.970 62.320 148.030 ;
        RECT 63.855 147.985 64.145 148.030 ;
        RECT 65.695 147.985 65.985 148.215 ;
        RECT 39.550 147.690 42.910 147.830 ;
        RECT 60.590 147.830 60.880 147.875 ;
        RECT 63.370 147.830 63.660 147.875 ;
        RECT 65.230 147.830 65.520 147.875 ;
        RECT 60.590 147.690 65.520 147.830 ;
        RECT 65.770 147.830 65.910 147.985 ;
        RECT 67.520 147.970 67.840 148.230 ;
        RECT 70.755 148.170 71.045 148.215 ;
        RECT 75.800 148.170 76.120 148.230 ;
        RECT 77.195 148.170 77.485 148.215 ;
        RECT 70.755 148.030 77.485 148.170 ;
        RECT 70.755 147.985 71.045 148.030 ;
        RECT 75.800 147.970 76.120 148.030 ;
        RECT 77.195 147.985 77.485 148.030 ;
        RECT 77.655 148.170 77.945 148.215 ;
        RECT 77.655 148.030 88.910 148.170 ;
        RECT 77.655 147.985 77.945 148.030 ;
        RECT 82.240 147.830 82.560 147.890 ;
        RECT 65.770 147.690 82.560 147.830 ;
        RECT 20.140 147.630 20.460 147.690 ;
        RECT 32.065 147.645 32.355 147.690 ;
        RECT 33.955 147.645 34.245 147.690 ;
        RECT 37.075 147.645 37.365 147.690 ;
        RECT 40.840 147.630 41.160 147.690 ;
        RECT 60.590 147.645 60.880 147.690 ;
        RECT 63.370 147.645 63.660 147.690 ;
        RECT 65.230 147.645 65.520 147.690 ;
        RECT 82.240 147.630 82.560 147.690 ;
        RECT 83.275 147.830 83.565 147.875 ;
        RECT 86.395 147.830 86.685 147.875 ;
        RECT 88.285 147.830 88.575 147.875 ;
        RECT 83.275 147.690 88.575 147.830 ;
        RECT 83.275 147.645 83.565 147.690 ;
        RECT 86.395 147.645 86.685 147.690 ;
        RECT 88.285 147.645 88.575 147.690 ;
        RECT 23.820 147.490 24.140 147.550 ;
        RECT 24.295 147.490 24.585 147.535 ;
        RECT 23.820 147.350 24.585 147.490 ;
        RECT 23.820 147.290 24.140 147.350 ;
        RECT 24.295 147.305 24.585 147.350 ;
        RECT 26.120 147.290 26.440 147.550 ;
        RECT 27.500 147.490 27.820 147.550 ;
        RECT 30.735 147.490 31.025 147.535 ;
        RECT 27.500 147.350 31.025 147.490 ;
        RECT 27.500 147.290 27.820 147.350 ;
        RECT 30.735 147.305 31.025 147.350 ;
        RECT 39.000 147.490 39.320 147.550 ;
        RECT 39.935 147.490 40.225 147.535 ;
        RECT 39.000 147.350 40.225 147.490 ;
        RECT 39.000 147.290 39.320 147.350 ;
        RECT 39.935 147.305 40.225 147.350 ;
        RECT 44.060 147.290 44.380 147.550 ;
        RECT 88.770 147.490 88.910 148.030 ;
        RECT 89.155 147.985 89.445 148.215 ;
        RECT 89.690 148.170 89.830 148.325 ;
        RECT 90.520 148.310 90.840 148.370 ;
        RECT 95.035 148.325 95.325 148.370 ;
        RECT 95.595 148.325 95.885 148.555 ;
        RECT 96.160 148.525 96.450 148.570 ;
        RECT 98.890 148.555 99.030 149.050 ;
        RECT 103.860 148.990 104.180 149.250 ;
        RECT 108.935 149.190 109.225 149.235 ;
        RECT 109.840 149.190 110.160 149.250 ;
        RECT 108.935 149.050 110.160 149.190 ;
        RECT 108.935 149.005 109.225 149.050 ;
        RECT 109.840 148.990 110.160 149.050 ;
        RECT 100.180 148.850 100.500 148.910 ;
        RECT 104.335 148.850 104.625 148.895 ;
        RECT 100.180 148.710 104.625 148.850 ;
        RECT 100.180 148.650 100.500 148.710 ;
        RECT 104.335 148.665 104.625 148.710 ;
        RECT 96.160 148.385 96.730 148.525 ;
        RECT 96.160 148.340 96.450 148.385 ;
        RECT 96.590 148.170 96.730 148.385 ;
        RECT 96.975 148.510 97.265 148.555 ;
        RECT 96.975 148.370 98.570 148.510 ;
        RECT 96.975 148.325 97.265 148.370 ;
        RECT 89.690 148.030 96.730 148.170 ;
        RECT 89.230 147.830 89.370 147.985 ;
        RECT 97.880 147.970 98.200 148.230 ;
        RECT 98.430 148.170 98.570 148.370 ;
        RECT 98.815 148.325 99.105 148.555 ;
        RECT 108.015 148.510 108.305 148.555 ;
        RECT 106.250 148.370 108.305 148.510 ;
        RECT 100.180 148.170 100.500 148.230 ;
        RECT 98.430 148.030 100.500 148.170 ;
        RECT 100.180 147.970 100.500 148.030 ;
        RECT 102.020 148.170 102.340 148.230 ;
        RECT 102.955 148.170 103.245 148.215 ;
        RECT 102.020 148.030 103.245 148.170 ;
        RECT 102.020 147.970 102.340 148.030 ;
        RECT 102.955 147.985 103.245 148.030 ;
        RECT 98.340 147.830 98.660 147.890 ;
        RECT 106.250 147.875 106.390 148.370 ;
        RECT 108.015 148.325 108.305 148.370 ;
        RECT 89.230 147.690 98.660 147.830 ;
        RECT 98.340 147.630 98.660 147.690 ;
        RECT 106.175 147.645 106.465 147.875 ;
        RECT 92.835 147.490 93.125 147.535 ;
        RECT 97.420 147.490 97.740 147.550 ;
        RECT 88.770 147.350 97.740 147.490 ;
        RECT 92.835 147.305 93.125 147.350 ;
        RECT 97.420 147.290 97.740 147.350 ;
        RECT 97.880 147.290 98.200 147.550 ;
        RECT 99.720 147.290 100.040 147.550 ;
        RECT 11.330 146.670 113.450 147.150 ;
        RECT 14.175 146.470 14.465 146.515 ;
        RECT 14.620 146.470 14.940 146.530 ;
        RECT 14.175 146.330 14.940 146.470 ;
        RECT 14.175 146.285 14.465 146.330 ;
        RECT 14.620 146.270 14.940 146.330 ;
        RECT 15.080 146.270 15.400 146.530 ;
        RECT 22.440 146.470 22.760 146.530 ;
        RECT 19.770 146.330 22.760 146.470 ;
        RECT 16.935 145.790 17.225 145.835 ;
        RECT 19.770 145.790 19.910 146.330 ;
        RECT 22.440 146.270 22.760 146.330 ;
        RECT 29.340 146.470 29.660 146.530 ;
        RECT 34.415 146.470 34.705 146.515 ;
        RECT 29.340 146.330 34.705 146.470 ;
        RECT 29.340 146.270 29.660 146.330 ;
        RECT 34.415 146.285 34.705 146.330 ;
        RECT 65.235 146.470 65.525 146.515 ;
        RECT 91.900 146.470 92.220 146.530 ;
        RECT 92.375 146.470 92.665 146.515 ;
        RECT 100.180 146.470 100.500 146.530 ;
        RECT 65.235 146.330 66.830 146.470 ;
        RECT 65.235 146.285 65.525 146.330 ;
        RECT 20.140 146.130 20.460 146.190 ;
        RECT 20.140 145.990 23.130 146.130 ;
        RECT 20.140 145.930 20.460 145.990 ;
        RECT 16.935 145.650 19.910 145.790 ;
        RECT 21.060 145.790 21.380 145.850 ;
        RECT 22.990 145.835 23.130 145.990 ;
        RECT 56.110 145.990 61.310 146.130 ;
        RECT 22.455 145.790 22.745 145.835 ;
        RECT 21.060 145.650 22.745 145.790 ;
        RECT 16.935 145.605 17.225 145.650 ;
        RECT 21.060 145.590 21.380 145.650 ;
        RECT 22.455 145.605 22.745 145.650 ;
        RECT 22.915 145.605 23.205 145.835 ;
        RECT 27.500 145.590 27.820 145.850 ;
        RECT 30.735 145.790 31.025 145.835 ;
        RECT 31.180 145.790 31.500 145.850 ;
        RECT 30.735 145.650 31.500 145.790 ;
        RECT 30.735 145.605 31.025 145.650 ;
        RECT 31.180 145.590 31.500 145.650 ;
        RECT 33.955 145.790 34.245 145.835 ;
        RECT 39.000 145.790 39.320 145.850 ;
        RECT 44.520 145.790 44.840 145.850 ;
        RECT 55.560 145.790 55.880 145.850 ;
        RECT 56.110 145.790 56.250 145.990 ;
        RECT 33.955 145.650 39.690 145.790 ;
        RECT 33.955 145.605 34.245 145.650 ;
        RECT 39.000 145.590 39.320 145.650 ;
        RECT 13.715 145.450 14.005 145.495 ;
        RECT 14.160 145.450 14.480 145.510 ;
        RECT 13.715 145.310 14.480 145.450 ;
        RECT 13.715 145.265 14.005 145.310 ;
        RECT 14.160 145.250 14.480 145.310 ;
        RECT 16.015 145.265 16.305 145.495 ;
        RECT 19.695 145.450 19.985 145.495 ;
        RECT 21.995 145.450 22.285 145.495 ;
        RECT 19.695 145.310 22.285 145.450 ;
        RECT 19.695 145.265 19.985 145.310 ;
        RECT 21.995 145.265 22.285 145.310 ;
        RECT 30.275 145.450 30.565 145.495 ;
        RECT 35.335 145.450 35.625 145.495 ;
        RECT 30.275 145.310 35.625 145.450 ;
        RECT 30.275 145.265 30.565 145.310 ;
        RECT 35.335 145.265 35.625 145.310 ;
        RECT 16.090 145.110 16.230 145.265 ;
        RECT 38.080 145.250 38.400 145.510 ;
        RECT 39.550 145.495 39.690 145.650 ;
        RECT 44.520 145.650 54.870 145.790 ;
        RECT 44.520 145.590 44.840 145.650 ;
        RECT 38.555 145.265 38.845 145.495 ;
        RECT 39.475 145.265 39.765 145.495 ;
        RECT 38.630 145.110 38.770 145.265 ;
        RECT 39.920 145.250 40.240 145.510 ;
        RECT 40.395 145.450 40.685 145.495 ;
        RECT 40.840 145.450 41.160 145.510 ;
        RECT 40.395 145.310 41.160 145.450 ;
        RECT 40.395 145.265 40.685 145.310 ;
        RECT 40.840 145.250 41.160 145.310 ;
        RECT 52.340 145.250 52.660 145.510 ;
        RECT 52.800 145.250 53.120 145.510 ;
        RECT 53.275 145.265 53.565 145.495 ;
        RECT 41.300 145.110 41.620 145.170 ;
        RECT 16.090 144.970 20.370 145.110 ;
        RECT 38.630 144.970 41.620 145.110 ;
        RECT 53.350 145.110 53.490 145.265 ;
        RECT 54.180 145.250 54.500 145.510 ;
        RECT 54.730 145.450 54.870 145.650 ;
        RECT 55.560 145.650 56.250 145.790 ;
        RECT 55.560 145.590 55.880 145.650 ;
        RECT 56.480 145.590 56.800 145.850 ;
        RECT 57.400 145.590 57.720 145.850 ;
        RECT 60.160 145.790 60.480 145.850 ;
        RECT 60.635 145.790 60.925 145.835 ;
        RECT 60.160 145.650 60.925 145.790 ;
        RECT 60.160 145.590 60.480 145.650 ;
        RECT 60.635 145.605 60.925 145.650 ;
        RECT 61.170 145.495 61.310 145.990 ;
        RECT 66.140 145.930 66.460 146.190 ;
        RECT 66.230 145.790 66.370 145.930 ;
        RECT 63.930 145.650 66.370 145.790 ;
        RECT 61.095 145.450 61.385 145.495 ;
        RECT 61.540 145.450 61.860 145.510 ;
        RECT 63.930 145.495 64.070 145.650 ;
        RECT 54.730 145.310 60.850 145.450 ;
        RECT 57.860 145.110 58.180 145.170 ;
        RECT 53.350 144.970 58.375 145.110 ;
        RECT 20.230 144.815 20.370 144.970 ;
        RECT 41.300 144.910 41.620 144.970 ;
        RECT 57.860 144.910 58.180 144.970 ;
        RECT 20.155 144.585 20.445 144.815 ;
        RECT 32.560 144.770 32.880 144.830 ;
        RECT 37.175 144.770 37.465 144.815 ;
        RECT 32.560 144.630 37.465 144.770 ;
        RECT 32.560 144.570 32.880 144.630 ;
        RECT 37.175 144.585 37.465 144.630 ;
        RECT 41.760 144.570 42.080 144.830 ;
        RECT 50.960 144.570 51.280 144.830 ;
        RECT 59.700 144.570 60.020 144.830 ;
        RECT 60.710 144.770 60.850 145.310 ;
        RECT 61.095 145.310 61.860 145.450 ;
        RECT 61.095 145.265 61.385 145.310 ;
        RECT 61.540 145.250 61.860 145.310 ;
        RECT 63.855 145.265 64.145 145.495 ;
        RECT 64.315 145.265 64.605 145.495 ;
        RECT 64.390 145.110 64.530 145.265 ;
        RECT 66.140 145.250 66.460 145.510 ;
        RECT 66.690 145.450 66.830 146.330 ;
        RECT 91.900 146.330 92.665 146.470 ;
        RECT 91.900 146.270 92.220 146.330 ;
        RECT 92.375 146.285 92.665 146.330 ;
        RECT 97.050 146.330 100.500 146.470 ;
        RECT 67.075 146.130 67.365 146.175 ;
        RECT 78.070 146.130 78.360 146.175 ;
        RECT 80.850 146.130 81.140 146.175 ;
        RECT 82.710 146.130 83.000 146.175 ;
        RECT 67.075 145.990 70.740 146.130 ;
        RECT 67.075 145.945 67.365 145.990 ;
        RECT 70.600 145.790 70.740 145.990 ;
        RECT 78.070 145.990 83.000 146.130 ;
        RECT 78.070 145.945 78.360 145.990 ;
        RECT 80.850 145.945 81.140 145.990 ;
        RECT 82.710 145.945 83.000 145.990 ;
        RECT 72.120 145.790 72.440 145.850 ;
        RECT 70.600 145.650 72.440 145.790 ;
        RECT 72.120 145.590 72.440 145.650 ;
        RECT 82.240 145.790 82.560 145.850 ;
        RECT 83.175 145.790 83.465 145.835 ;
        RECT 84.080 145.790 84.400 145.850 ;
        RECT 82.240 145.650 84.400 145.790 ;
        RECT 82.240 145.590 82.560 145.650 ;
        RECT 83.175 145.605 83.465 145.650 ;
        RECT 84.080 145.590 84.400 145.650 ;
        RECT 93.295 145.790 93.585 145.835 ;
        RECT 95.120 145.790 95.440 145.850 ;
        RECT 93.295 145.650 95.440 145.790 ;
        RECT 93.295 145.605 93.585 145.650 ;
        RECT 95.120 145.590 95.440 145.650 ;
        RECT 72.580 145.450 72.900 145.510 ;
        RECT 66.690 145.310 72.900 145.450 ;
        RECT 72.580 145.250 72.900 145.310 ;
        RECT 73.500 145.250 73.820 145.510 ;
        RECT 74.205 145.450 74.495 145.495 ;
        RECT 76.720 145.450 77.040 145.510 ;
        RECT 74.205 145.310 77.040 145.450 ;
        RECT 74.205 145.265 74.495 145.310 ;
        RECT 76.720 145.250 77.040 145.310 ;
        RECT 78.070 145.450 78.360 145.495 ;
        RECT 78.070 145.310 80.605 145.450 ;
        RECT 78.070 145.265 78.360 145.310 ;
        RECT 67.980 145.110 68.300 145.170 ;
        RECT 80.390 145.155 80.605 145.310 ;
        RECT 81.320 145.250 81.640 145.510 ;
        RECT 92.375 145.450 92.665 145.495 ;
        RECT 96.500 145.450 96.820 145.510 ;
        RECT 97.050 145.495 97.190 146.330 ;
        RECT 100.180 146.270 100.500 146.330 ;
        RECT 98.800 145.930 99.120 146.190 ;
        RECT 102.020 146.130 102.340 146.190 ;
        RECT 102.020 145.990 103.170 146.130 ;
        RECT 102.020 145.930 102.340 145.990 ;
        RECT 98.890 145.790 99.030 145.930 ;
        RECT 103.030 145.835 103.170 145.990 ;
        RECT 98.430 145.650 99.030 145.790 ;
        RECT 98.430 145.495 98.570 145.650 ;
        RECT 102.955 145.605 103.245 145.835 ;
        RECT 92.375 145.310 96.820 145.450 ;
        RECT 92.375 145.265 92.665 145.310 ;
        RECT 96.500 145.250 96.820 145.310 ;
        RECT 96.975 145.265 97.265 145.495 ;
        RECT 97.790 145.450 98.080 145.495 ;
        RECT 97.510 145.310 98.080 145.450 ;
        RECT 64.390 144.970 68.300 145.110 ;
        RECT 67.980 144.910 68.300 144.970 ;
        RECT 73.055 145.110 73.345 145.155 ;
        RECT 76.210 145.110 76.500 145.155 ;
        RECT 79.470 145.110 79.760 145.155 ;
        RECT 73.055 144.970 79.760 145.110 ;
        RECT 73.055 144.925 73.345 144.970 ;
        RECT 76.210 144.925 76.500 144.970 ;
        RECT 79.470 144.925 79.760 144.970 ;
        RECT 80.390 145.110 80.680 145.155 ;
        RECT 82.250 145.110 82.540 145.155 ;
        RECT 80.390 144.970 82.540 145.110 ;
        RECT 80.390 144.925 80.680 144.970 ;
        RECT 82.250 144.925 82.540 144.970 ;
        RECT 93.755 145.110 94.045 145.155 ;
        RECT 94.660 145.110 94.980 145.170 ;
        RECT 97.050 145.110 97.190 145.265 ;
        RECT 93.755 144.970 94.980 145.110 ;
        RECT 93.755 144.925 94.045 144.970 ;
        RECT 94.660 144.910 94.980 144.970 ;
        RECT 96.590 144.970 97.190 145.110 ;
        RECT 96.590 144.830 96.730 144.970 ;
        RECT 62.935 144.770 63.225 144.815 ;
        RECT 71.660 144.770 71.980 144.830 ;
        RECT 60.710 144.630 71.980 144.770 ;
        RECT 62.935 144.585 63.225 144.630 ;
        RECT 71.660 144.570 71.980 144.630 ;
        RECT 91.455 144.770 91.745 144.815 ;
        RECT 96.040 144.770 96.360 144.830 ;
        RECT 91.455 144.630 96.360 144.770 ;
        RECT 91.455 144.585 91.745 144.630 ;
        RECT 96.040 144.570 96.360 144.630 ;
        RECT 96.500 144.570 96.820 144.830 ;
        RECT 97.510 144.770 97.650 145.310 ;
        RECT 97.790 145.265 98.080 145.310 ;
        RECT 98.370 145.265 98.660 145.495 ;
        RECT 98.915 145.450 99.205 145.495 ;
        RECT 101.100 145.450 101.420 145.510 ;
        RECT 98.915 145.310 101.420 145.450 ;
        RECT 98.915 145.265 99.205 145.310 ;
        RECT 101.100 145.250 101.420 145.310 ;
        RECT 103.860 145.450 104.180 145.510 ;
        RECT 104.335 145.450 104.625 145.495 ;
        RECT 103.860 145.310 104.625 145.450 ;
        RECT 103.860 145.250 104.180 145.310 ;
        RECT 104.335 145.265 104.625 145.310 ;
        RECT 105.700 145.450 106.020 145.510 ;
        RECT 107.080 145.450 107.400 145.510 ;
        RECT 107.555 145.450 107.845 145.495 ;
        RECT 105.700 145.310 107.845 145.450 ;
        RECT 105.700 145.250 106.020 145.310 ;
        RECT 107.080 145.250 107.400 145.310 ;
        RECT 107.555 145.265 107.845 145.310 ;
        RECT 108.015 145.265 108.305 145.495 ;
        RECT 108.090 145.110 108.230 145.265 ;
        RECT 98.890 144.970 103.170 145.110 ;
        RECT 98.890 144.770 99.030 144.970 ;
        RECT 103.030 144.830 103.170 144.970 ;
        RECT 106.250 144.970 108.230 145.110 ;
        RECT 97.510 144.630 99.030 144.770 ;
        RECT 100.180 144.570 100.500 144.830 ;
        RECT 102.940 144.770 103.260 144.830 ;
        RECT 106.250 144.815 106.390 144.970 ;
        RECT 103.875 144.770 104.165 144.815 ;
        RECT 102.940 144.630 104.165 144.770 ;
        RECT 102.940 144.570 103.260 144.630 ;
        RECT 103.875 144.585 104.165 144.630 ;
        RECT 106.175 144.585 106.465 144.815 ;
        RECT 107.080 144.570 107.400 144.830 ;
        RECT 108.935 144.770 109.225 144.815 ;
        RECT 109.840 144.770 110.160 144.830 ;
        RECT 108.935 144.630 110.160 144.770 ;
        RECT 108.935 144.585 109.225 144.630 ;
        RECT 109.840 144.570 110.160 144.630 ;
        RECT 11.330 143.950 113.450 144.430 ;
        RECT 51.895 143.750 52.185 143.795 ;
        RECT 52.340 143.750 52.660 143.810 ;
        RECT 51.895 143.610 52.660 143.750 ;
        RECT 51.895 143.565 52.185 143.610 ;
        RECT 52.340 143.550 52.660 143.610 ;
        RECT 54.195 143.565 54.485 143.795 ;
        RECT 54.640 143.750 54.960 143.810 ;
        RECT 62.000 143.750 62.320 143.810 ;
        RECT 62.475 143.750 62.765 143.795 ;
        RECT 54.640 143.610 56.940 143.750 ;
        RECT 31.655 143.410 31.945 143.455 ;
        RECT 50.960 143.410 51.280 143.470 ;
        RECT 31.655 143.270 51.280 143.410 ;
        RECT 31.655 143.225 31.945 143.270 ;
        RECT 50.960 143.210 51.280 143.270 ;
        RECT 30.260 142.870 30.580 143.130 ;
        RECT 30.720 142.870 31.040 143.130 ;
        RECT 44.520 143.070 44.840 143.130 ;
        RECT 44.995 143.070 45.285 143.115 ;
        RECT 44.520 142.930 45.285 143.070 ;
        RECT 44.520 142.870 44.840 142.930 ;
        RECT 44.995 142.885 45.285 142.930 ;
        RECT 45.440 142.870 45.760 143.130 ;
        RECT 45.900 142.870 46.220 143.130 ;
        RECT 46.835 143.070 47.125 143.115 ;
        RECT 50.040 143.070 50.360 143.130 ;
        RECT 46.835 142.930 50.360 143.070 ;
        RECT 46.835 142.885 47.125 142.930 ;
        RECT 50.040 142.870 50.360 142.930 ;
        RECT 51.880 143.070 52.200 143.130 ;
        RECT 52.355 143.070 52.645 143.115 ;
        RECT 51.880 142.930 52.645 143.070 ;
        RECT 54.270 143.070 54.410 143.565 ;
        RECT 54.640 143.550 54.960 143.610 ;
        RECT 56.800 143.410 56.940 143.610 ;
        RECT 62.000 143.610 62.765 143.750 ;
        RECT 62.000 143.550 62.320 143.610 ;
        RECT 62.475 143.565 62.765 143.610 ;
        RECT 76.720 143.550 77.040 143.810 ;
        RECT 79.035 143.565 79.325 143.795 ;
        RECT 80.415 143.750 80.705 143.795 ;
        RECT 81.320 143.750 81.640 143.810 ;
        RECT 90.520 143.750 90.840 143.810 ;
        RECT 80.415 143.610 81.640 143.750 ;
        RECT 80.415 143.565 80.705 143.610 ;
        RECT 69.835 143.410 70.125 143.455 ;
        RECT 70.295 143.410 70.585 143.455 ;
        RECT 76.810 143.410 76.950 143.550 ;
        RECT 56.800 143.270 69.590 143.410 ;
        RECT 55.115 143.070 55.405 143.115 ;
        RECT 54.270 142.930 55.405 143.070 ;
        RECT 51.880 142.870 52.200 142.930 ;
        RECT 52.355 142.885 52.645 142.930 ;
        RECT 55.115 142.885 55.405 142.930 ;
        RECT 59.700 143.070 60.020 143.130 ;
        RECT 61.555 143.070 61.845 143.115 ;
        RECT 59.700 142.930 61.845 143.070 ;
        RECT 59.700 142.870 60.020 142.930 ;
        RECT 61.555 142.885 61.845 142.930 ;
        RECT 68.440 142.870 68.760 143.130 ;
        RECT 69.450 143.070 69.590 143.270 ;
        RECT 69.835 143.270 70.585 143.410 ;
        RECT 69.835 143.225 70.125 143.270 ;
        RECT 70.295 143.225 70.585 143.270 ;
        RECT 72.670 143.270 76.950 143.410 ;
        RECT 69.450 142.930 71.430 143.070 ;
        RECT 51.435 142.730 51.725 142.775 ;
        RECT 53.720 142.730 54.040 142.790 ;
        RECT 56.480 142.730 56.800 142.790 ;
        RECT 51.435 142.590 56.800 142.730 ;
        RECT 51.435 142.545 51.725 142.590 ;
        RECT 53.720 142.530 54.040 142.590 ;
        RECT 56.480 142.530 56.800 142.590 ;
        RECT 67.060 142.730 67.380 142.790 ;
        RECT 68.915 142.730 69.205 142.775 ;
        RECT 67.060 142.590 69.205 142.730 ;
        RECT 71.290 142.730 71.430 142.930 ;
        RECT 71.660 142.870 71.980 143.130 ;
        RECT 72.120 142.870 72.440 143.130 ;
        RECT 72.670 143.115 72.810 143.270 ;
        RECT 72.595 142.885 72.885 143.115 ;
        RECT 73.040 143.070 73.360 143.130 ;
        RECT 73.515 143.070 73.805 143.115 ;
        RECT 73.040 142.930 73.805 143.070 ;
        RECT 73.040 142.870 73.360 142.930 ;
        RECT 73.515 142.885 73.805 142.930 ;
        RECT 76.720 143.070 77.040 143.130 ;
        RECT 77.195 143.070 77.485 143.115 ;
        RECT 76.720 142.930 77.485 143.070 ;
        RECT 79.110 143.070 79.250 143.565 ;
        RECT 81.320 143.550 81.640 143.610 ;
        RECT 89.230 143.610 90.840 143.750 ;
        RECT 87.315 143.410 87.605 143.455 ;
        RECT 87.775 143.410 88.065 143.455 ;
        RECT 87.315 143.270 88.065 143.410 ;
        RECT 87.315 143.225 87.605 143.270 ;
        RECT 87.775 143.225 88.065 143.270 ;
        RECT 79.495 143.070 79.785 143.115 ;
        RECT 79.110 142.930 79.785 143.070 ;
        RECT 76.720 142.870 77.040 142.930 ;
        RECT 77.195 142.885 77.485 142.930 ;
        RECT 79.495 142.885 79.785 142.930 ;
        RECT 85.920 142.870 86.240 143.130 ;
        RECT 89.230 143.115 89.370 143.610 ;
        RECT 90.520 143.550 90.840 143.610 ;
        RECT 93.755 143.750 94.045 143.795 ;
        RECT 94.660 143.750 94.980 143.810 ;
        RECT 93.755 143.610 94.980 143.750 ;
        RECT 93.755 143.565 94.045 143.610 ;
        RECT 94.660 143.550 94.980 143.610 ;
        RECT 95.580 143.750 95.900 143.810 ;
        RECT 97.435 143.750 97.725 143.795 ;
        RECT 95.580 143.610 97.725 143.750 ;
        RECT 95.580 143.550 95.900 143.610 ;
        RECT 97.435 143.565 97.725 143.610 ;
        RECT 98.800 143.410 99.120 143.470 ;
        RECT 89.690 143.270 99.120 143.410 ;
        RECT 89.690 143.115 89.830 143.270 ;
        RECT 89.155 142.885 89.445 143.115 ;
        RECT 89.615 142.885 89.905 143.115 ;
        RECT 90.060 142.870 90.380 143.130 ;
        RECT 95.670 143.115 95.810 143.270 ;
        RECT 98.800 143.210 99.120 143.270 ;
        RECT 99.260 143.210 99.580 143.470 ;
        RECT 99.735 143.410 100.025 143.455 ;
        RECT 100.180 143.410 100.500 143.470 ;
        RECT 102.940 143.455 103.260 143.470 ;
        RECT 99.735 143.270 100.500 143.410 ;
        RECT 99.735 143.225 100.025 143.270 ;
        RECT 100.180 143.210 100.500 143.270 ;
        RECT 102.725 143.225 103.260 143.455 ;
        RECT 104.730 143.410 105.020 143.455 ;
        RECT 107.080 143.410 107.400 143.470 ;
        RECT 107.990 143.410 108.280 143.455 ;
        RECT 104.730 143.270 108.280 143.410 ;
        RECT 104.730 143.225 105.020 143.270 ;
        RECT 102.940 143.210 103.260 143.225 ;
        RECT 107.080 143.210 107.400 143.270 ;
        RECT 107.990 143.225 108.280 143.270 ;
        RECT 108.910 143.410 109.200 143.455 ;
        RECT 110.770 143.410 111.060 143.455 ;
        RECT 108.910 143.270 111.060 143.410 ;
        RECT 108.910 143.225 109.200 143.270 ;
        RECT 110.770 143.225 111.060 143.270 ;
        RECT 90.995 143.070 91.285 143.115 ;
        RECT 90.610 142.930 91.285 143.070 ;
        RECT 71.290 142.590 75.570 142.730 ;
        RECT 67.060 142.530 67.380 142.590 ;
        RECT 68.915 142.545 69.205 142.590 ;
        RECT 67.535 142.390 67.825 142.435 ;
        RECT 73.500 142.390 73.820 142.450 ;
        RECT 67.535 142.250 73.820 142.390 ;
        RECT 75.430 142.390 75.570 142.590 ;
        RECT 75.800 142.530 76.120 142.790 ;
        RECT 86.840 142.530 87.160 142.790 ;
        RECT 89.600 142.390 89.920 142.450 ;
        RECT 90.610 142.390 90.750 142.930 ;
        RECT 90.995 142.885 91.285 142.930 ;
        RECT 95.135 142.885 95.425 143.115 ;
        RECT 95.595 142.885 95.885 143.115 ;
        RECT 96.055 142.885 96.345 143.115 ;
        RECT 96.500 143.070 96.820 143.130 ;
        RECT 96.975 143.070 97.265 143.115 ;
        RECT 96.500 142.930 97.265 143.070 ;
        RECT 95.210 142.730 95.350 142.885 ;
        RECT 91.070 142.590 95.350 142.730 ;
        RECT 96.130 142.730 96.270 142.885 ;
        RECT 96.500 142.870 96.820 142.930 ;
        RECT 96.975 142.885 97.265 142.930 ;
        RECT 98.355 143.070 98.645 143.115 ;
        RECT 99.350 143.070 99.490 143.210 ;
        RECT 98.355 142.930 99.490 143.070 ;
        RECT 101.115 143.070 101.405 143.115 ;
        RECT 105.700 143.070 106.020 143.130 ;
        RECT 101.115 142.930 106.020 143.070 ;
        RECT 98.355 142.885 98.645 142.930 ;
        RECT 101.115 142.885 101.405 142.930 ;
        RECT 105.700 142.870 106.020 142.930 ;
        RECT 106.590 143.070 106.880 143.115 ;
        RECT 108.910 143.070 109.125 143.225 ;
        RECT 106.590 142.930 109.125 143.070 ;
        RECT 106.590 142.885 106.880 142.930 ;
        RECT 109.840 142.870 110.160 143.130 ;
        RECT 98.800 142.730 99.120 142.790 ;
        RECT 96.130 142.590 99.120 142.730 ;
        RECT 91.070 142.450 91.210 142.590 ;
        RECT 98.800 142.530 99.120 142.590 ;
        RECT 99.275 142.545 99.565 142.775 ;
        RECT 75.430 142.250 90.750 142.390 ;
        RECT 67.535 142.205 67.825 142.250 ;
        RECT 73.500 142.190 73.820 142.250 ;
        RECT 89.600 142.190 89.920 142.250 ;
        RECT 27.960 142.050 28.280 142.110 ;
        RECT 29.355 142.050 29.645 142.095 ;
        RECT 27.960 141.910 29.645 142.050 ;
        RECT 27.960 141.850 28.280 141.910 ;
        RECT 29.355 141.865 29.645 141.910 ;
        RECT 30.260 141.850 30.580 142.110 ;
        RECT 38.540 142.050 38.860 142.110 ;
        RECT 43.615 142.050 43.905 142.095 ;
        RECT 38.540 141.910 43.905 142.050 ;
        RECT 38.540 141.850 38.860 141.910 ;
        RECT 43.615 141.865 43.905 141.910 ;
        RECT 56.035 142.050 56.325 142.095 ;
        RECT 56.480 142.050 56.800 142.110 ;
        RECT 56.035 141.910 56.800 142.050 ;
        RECT 56.035 141.865 56.325 141.910 ;
        RECT 56.480 141.850 56.800 141.910 ;
        RECT 69.820 141.850 70.140 142.110 ;
        RECT 85.015 142.050 85.305 142.095 ;
        RECT 85.460 142.050 85.780 142.110 ;
        RECT 85.015 141.910 85.780 142.050 ;
        RECT 85.015 141.865 85.305 141.910 ;
        RECT 85.460 141.850 85.780 141.910 ;
        RECT 86.840 141.850 87.160 142.110 ;
        RECT 90.610 142.050 90.750 142.250 ;
        RECT 90.980 142.190 91.300 142.450 ;
        RECT 94.660 142.390 94.980 142.450 ;
        RECT 96.040 142.390 96.360 142.450 ;
        RECT 94.660 142.250 96.360 142.390 ;
        RECT 94.660 142.190 94.980 142.250 ;
        RECT 96.040 142.190 96.360 142.250 ;
        RECT 96.960 142.390 97.280 142.450 ;
        RECT 99.350 142.390 99.490 142.545 ;
        RECT 111.680 142.530 112.000 142.790 ;
        RECT 96.960 142.250 99.490 142.390 ;
        RECT 106.590 142.390 106.880 142.435 ;
        RECT 109.370 142.390 109.660 142.435 ;
        RECT 111.230 142.390 111.520 142.435 ;
        RECT 106.590 142.250 111.520 142.390 ;
        RECT 96.960 142.190 97.280 142.250 ;
        RECT 106.590 142.205 106.880 142.250 ;
        RECT 109.370 142.205 109.660 142.250 ;
        RECT 111.230 142.205 111.520 142.250 ;
        RECT 96.500 142.050 96.820 142.110 ;
        RECT 90.610 141.910 96.820 142.050 ;
        RECT 96.500 141.850 96.820 141.910 ;
        RECT 97.420 142.050 97.740 142.110 ;
        RECT 98.355 142.050 98.645 142.095 ;
        RECT 97.420 141.910 98.645 142.050 ;
        RECT 97.420 141.850 97.740 141.910 ;
        RECT 98.355 141.865 98.645 141.910 ;
        RECT 101.560 141.850 101.880 142.110 ;
        RECT 11.330 141.230 113.450 141.710 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 26.120 140.830 26.440 141.090 ;
        RECT 30.260 140.830 30.580 141.090 ;
        RECT 35.780 141.030 36.100 141.090 ;
        RECT 38.555 141.030 38.845 141.075 ;
        RECT 35.780 140.890 38.845 141.030 ;
        RECT 35.780 140.830 36.100 140.890 ;
        RECT 38.555 140.845 38.845 140.890 ;
        RECT 39.920 141.030 40.240 141.090 ;
        RECT 41.315 141.030 41.605 141.075 ;
        RECT 57.400 141.030 57.720 141.090 ;
        RECT 39.920 140.890 41.605 141.030 ;
        RECT 39.920 140.830 40.240 140.890 ;
        RECT 41.315 140.845 41.605 140.890 ;
        RECT 50.130 140.890 57.720 141.030 ;
        RECT 25.200 140.690 25.520 140.750 ;
        RECT 17.930 140.550 25.520 140.690 ;
        RECT 17.930 140.055 18.070 140.550 ;
        RECT 25.200 140.490 25.520 140.550 ;
        RECT 40.855 140.690 41.145 140.735 ;
        RECT 43.615 140.690 43.905 140.735 ;
        RECT 50.130 140.690 50.270 140.890 ;
        RECT 57.400 140.830 57.720 140.890 ;
        RECT 40.855 140.550 43.370 140.690 ;
        RECT 40.855 140.505 41.145 140.550 ;
        RECT 21.520 140.350 21.840 140.410 ;
        RECT 21.995 140.350 22.285 140.395 ;
        RECT 27.975 140.350 28.265 140.395 ;
        RECT 21.520 140.210 22.285 140.350 ;
        RECT 21.520 140.150 21.840 140.210 ;
        RECT 21.995 140.165 22.285 140.210 ;
        RECT 22.990 140.210 28.265 140.350 ;
        RECT 17.855 139.825 18.145 140.055 ;
        RECT 21.060 140.010 21.380 140.070 ;
        RECT 22.990 140.010 23.130 140.210 ;
        RECT 27.975 140.165 28.265 140.210 ;
        RECT 39.460 140.150 39.780 140.410 ;
        RECT 42.220 140.150 42.540 140.410 ;
        RECT 43.230 140.350 43.370 140.550 ;
        RECT 43.615 140.550 50.270 140.690 ;
        RECT 53.230 140.690 53.520 140.735 ;
        RECT 56.010 140.690 56.300 140.735 ;
        RECT 57.870 140.690 58.160 140.735 ;
        RECT 53.230 140.550 58.160 140.690 ;
        RECT 43.615 140.505 43.905 140.550 ;
        RECT 53.230 140.505 53.520 140.550 ;
        RECT 56.010 140.505 56.300 140.550 ;
        RECT 57.870 140.505 58.160 140.550 ;
        RECT 71.660 140.490 71.980 140.750 ;
        RECT 98.800 140.690 99.120 140.750 ;
        RECT 100.885 140.690 101.175 140.735 ;
        RECT 102.480 140.690 102.800 140.750 ;
        RECT 97.970 140.550 102.800 140.690 ;
        RECT 43.230 140.210 56.250 140.350 ;
        RECT 21.060 139.870 23.130 140.010 ;
        RECT 24.295 140.010 24.585 140.055 ;
        RECT 25.200 140.010 25.520 140.070 ;
        RECT 24.295 139.870 25.520 140.010 ;
        RECT 21.060 139.810 21.380 139.870 ;
        RECT 24.295 139.825 24.585 139.870 ;
        RECT 25.200 139.810 25.520 139.870 ;
        RECT 27.055 139.825 27.345 140.055 ;
        RECT 21.535 139.670 21.825 139.715 ;
        RECT 22.440 139.670 22.760 139.730 ;
        RECT 21.535 139.530 22.760 139.670 ;
        RECT 27.130 139.670 27.270 139.825 ;
        RECT 28.420 139.810 28.740 140.070 ;
        RECT 29.355 140.010 29.645 140.055 ;
        RECT 31.180 140.010 31.500 140.070 ;
        RECT 29.355 139.870 31.500 140.010 ;
        RECT 29.355 139.825 29.645 139.870 ;
        RECT 29.430 139.670 29.570 139.825 ;
        RECT 31.180 139.810 31.500 139.870 ;
        RECT 38.540 139.810 38.860 140.070 ;
        RECT 39.000 140.010 39.320 140.070 ;
        RECT 39.935 140.010 40.225 140.055 ;
        RECT 39.000 139.870 40.225 140.010 ;
        RECT 39.000 139.810 39.320 139.870 ;
        RECT 39.935 139.825 40.225 139.870 ;
        RECT 42.680 139.810 43.000 140.070 ;
        RECT 44.520 140.010 44.840 140.070 ;
        RECT 46.360 140.010 46.680 140.070 ;
        RECT 46.835 140.010 47.125 140.055 ;
        RECT 44.520 139.870 47.125 140.010 ;
        RECT 44.520 139.810 44.840 139.870 ;
        RECT 46.360 139.810 46.680 139.870 ;
        RECT 46.835 139.825 47.125 139.870 ;
        RECT 47.295 139.825 47.585 140.055 ;
        RECT 47.755 139.825 48.045 140.055 ;
        RECT 48.675 140.010 48.965 140.055 ;
        RECT 50.040 140.010 50.360 140.070 ;
        RECT 48.675 139.870 50.360 140.010 ;
        RECT 48.675 139.825 48.965 139.870 ;
        RECT 27.130 139.530 29.570 139.670 ;
        RECT 41.315 139.670 41.605 139.715 ;
        RECT 45.455 139.670 45.745 139.715 ;
        RECT 41.315 139.530 45.745 139.670 ;
        RECT 21.535 139.485 21.825 139.530 ;
        RECT 22.440 139.470 22.760 139.530 ;
        RECT 41.315 139.485 41.605 139.530 ;
        RECT 45.455 139.485 45.745 139.530 ;
        RECT 45.900 139.670 46.220 139.730 ;
        RECT 47.370 139.670 47.510 139.825 ;
        RECT 45.900 139.530 47.510 139.670 ;
        RECT 45.900 139.470 46.220 139.530 ;
        RECT 17.395 139.330 17.685 139.375 ;
        RECT 17.840 139.330 18.160 139.390 ;
        RECT 17.395 139.190 18.160 139.330 ;
        RECT 17.395 139.145 17.685 139.190 ;
        RECT 17.840 139.130 18.160 139.190 ;
        RECT 19.235 139.330 19.525 139.375 ;
        RECT 21.980 139.330 22.300 139.390 ;
        RECT 19.235 139.190 22.300 139.330 ;
        RECT 19.235 139.145 19.525 139.190 ;
        RECT 21.980 139.130 22.300 139.190 ;
        RECT 24.740 139.130 25.060 139.390 ;
        RECT 47.830 139.330 47.970 139.825 ;
        RECT 50.040 139.810 50.360 139.870 ;
        RECT 53.230 140.010 53.520 140.055 ;
        RECT 56.110 140.010 56.250 140.210 ;
        RECT 56.480 140.150 56.800 140.410 ;
        RECT 71.750 140.350 71.890 140.490 ;
        RECT 70.830 140.210 71.890 140.350 ;
        RECT 74.420 140.350 74.740 140.410 ;
        RECT 75.800 140.350 76.120 140.410 ;
        RECT 74.420 140.210 76.120 140.350 ;
        RECT 58.335 140.010 58.625 140.055 ;
        RECT 61.080 140.010 61.400 140.070 ;
        RECT 70.830 140.055 70.970 140.210 ;
        RECT 74.420 140.150 74.740 140.210 ;
        RECT 75.800 140.150 76.120 140.210 ;
        RECT 76.260 140.150 76.580 140.410 ;
        RECT 77.180 140.350 77.500 140.410 ;
        RECT 94.215 140.350 94.505 140.395 ;
        RECT 96.040 140.350 96.360 140.410 ;
        RECT 77.180 140.210 81.090 140.350 ;
        RECT 77.180 140.150 77.500 140.210 ;
        RECT 53.230 139.870 55.765 140.010 ;
        RECT 56.110 139.870 58.090 140.010 ;
        RECT 53.230 139.825 53.520 139.870 ;
        RECT 51.370 139.670 51.660 139.715 ;
        RECT 51.880 139.670 52.200 139.730 ;
        RECT 55.550 139.715 55.765 139.870 ;
        RECT 54.630 139.670 54.920 139.715 ;
        RECT 51.370 139.530 54.920 139.670 ;
        RECT 51.370 139.485 51.660 139.530 ;
        RECT 51.880 139.470 52.200 139.530 ;
        RECT 54.630 139.485 54.920 139.530 ;
        RECT 55.550 139.670 55.840 139.715 ;
        RECT 57.410 139.670 57.700 139.715 ;
        RECT 55.550 139.530 57.700 139.670 ;
        RECT 57.950 139.670 58.090 139.870 ;
        RECT 58.335 139.870 61.400 140.010 ;
        RECT 58.335 139.825 58.625 139.870 ;
        RECT 61.080 139.810 61.400 139.870 ;
        RECT 70.755 139.825 71.045 140.055 ;
        RECT 71.215 139.825 71.505 140.055 ;
        RECT 71.675 139.825 71.965 140.055 ;
        RECT 72.595 140.010 72.885 140.055 ;
        RECT 73.040 140.010 73.360 140.070 ;
        RECT 80.950 140.055 81.090 140.210 ;
        RECT 94.215 140.210 96.360 140.350 ;
        RECT 94.215 140.165 94.505 140.210 ;
        RECT 96.040 140.150 96.360 140.210 ;
        RECT 79.495 140.010 79.785 140.055 ;
        RECT 72.595 139.870 73.360 140.010 ;
        RECT 72.595 139.825 72.885 139.870 ;
        RECT 60.160 139.670 60.480 139.730 ;
        RECT 57.950 139.530 60.480 139.670 ;
        RECT 55.550 139.485 55.840 139.530 ;
        RECT 57.410 139.485 57.700 139.530 ;
        RECT 60.160 139.470 60.480 139.530 ;
        RECT 49.365 139.330 49.655 139.375 ;
        RECT 52.340 139.330 52.660 139.390 ;
        RECT 47.830 139.190 52.660 139.330 ;
        RECT 49.365 139.145 49.655 139.190 ;
        RECT 52.340 139.130 52.660 139.190 ;
        RECT 69.375 139.330 69.665 139.375 ;
        RECT 70.280 139.330 70.600 139.390 ;
        RECT 69.375 139.190 70.600 139.330 ;
        RECT 71.290 139.330 71.430 139.825 ;
        RECT 71.750 139.670 71.890 139.825 ;
        RECT 73.040 139.810 73.360 139.870 ;
        RECT 78.650 139.870 79.785 140.010 ;
        RECT 76.260 139.670 76.580 139.730 ;
        RECT 71.750 139.530 76.580 139.670 ;
        RECT 76.260 139.470 76.580 139.530 ;
        RECT 71.660 139.330 71.980 139.390 ;
        RECT 71.290 139.190 71.980 139.330 ;
        RECT 69.375 139.145 69.665 139.190 ;
        RECT 70.280 139.130 70.600 139.190 ;
        RECT 71.660 139.130 71.980 139.190 ;
        RECT 74.880 139.330 75.200 139.390 ;
        RECT 78.650 139.375 78.790 139.870 ;
        RECT 79.495 139.825 79.785 139.870 ;
        RECT 80.875 139.825 81.165 140.055 ;
        RECT 90.060 140.010 90.380 140.070 ;
        RECT 94.675 140.010 94.965 140.055 ;
        RECT 90.060 139.870 94.965 140.010 ;
        RECT 90.060 139.810 90.380 139.870 ;
        RECT 94.675 139.825 94.965 139.870 ;
        RECT 95.135 140.010 95.425 140.055 ;
        RECT 97.970 140.010 98.110 140.550 ;
        RECT 98.800 140.490 99.120 140.550 ;
        RECT 100.885 140.505 101.175 140.550 ;
        RECT 102.480 140.490 102.800 140.550 ;
        RECT 104.750 140.690 105.040 140.735 ;
        RECT 107.530 140.690 107.820 140.735 ;
        RECT 109.390 140.690 109.680 140.735 ;
        RECT 104.750 140.550 109.680 140.690 ;
        RECT 104.750 140.505 105.040 140.550 ;
        RECT 107.530 140.505 107.820 140.550 ;
        RECT 109.390 140.505 109.680 140.550 ;
        RECT 98.340 140.350 98.660 140.410 ;
        RECT 98.340 140.210 107.770 140.350 ;
        RECT 98.340 140.150 98.660 140.210 ;
        RECT 95.135 139.870 98.110 140.010 ;
        RECT 104.750 140.010 105.040 140.055 ;
        RECT 107.630 140.010 107.770 140.210 ;
        RECT 108.000 140.150 108.320 140.410 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 109.855 140.010 110.145 140.055 ;
        RECT 111.680 140.010 112.000 140.070 ;
        RECT 104.750 139.870 107.285 140.010 ;
        RECT 107.630 139.870 112.000 140.010 ;
        RECT 95.135 139.825 95.425 139.870 ;
        RECT 104.750 139.825 105.040 139.870 ;
        RECT 101.560 139.670 101.880 139.730 ;
        RECT 107.070 139.715 107.285 139.870 ;
        RECT 109.855 139.825 110.145 139.870 ;
        RECT 111.680 139.810 112.000 139.870 ;
        RECT 102.890 139.670 103.180 139.715 ;
        RECT 106.150 139.670 106.440 139.715 ;
        RECT 101.560 139.530 106.440 139.670 ;
        RECT 101.560 139.470 101.880 139.530 ;
        RECT 102.890 139.485 103.180 139.530 ;
        RECT 106.150 139.485 106.440 139.530 ;
        RECT 107.070 139.670 107.360 139.715 ;
        RECT 108.930 139.670 109.220 139.715 ;
        RECT 107.070 139.530 109.220 139.670 ;
        RECT 107.070 139.485 107.360 139.530 ;
        RECT 108.930 139.485 109.220 139.530 ;
        RECT 76.735 139.330 77.025 139.375 ;
        RECT 74.880 139.190 77.025 139.330 ;
        RECT 74.880 139.130 75.200 139.190 ;
        RECT 76.735 139.145 77.025 139.190 ;
        RECT 78.575 139.145 78.865 139.375 ;
        RECT 80.400 139.130 80.720 139.390 ;
        RECT 81.795 139.330 82.085 139.375 ;
        RECT 82.240 139.330 82.560 139.390 ;
        RECT 81.795 139.190 82.560 139.330 ;
        RECT 81.795 139.145 82.085 139.190 ;
        RECT 82.240 139.130 82.560 139.190 ;
        RECT 96.960 139.130 97.280 139.390 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 11.330 138.510 113.450 138.990 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 13.485 138.310 13.775 138.355 ;
        RECT 21.060 138.310 21.380 138.370 ;
        RECT 13.485 138.170 21.380 138.310 ;
        RECT 13.485 138.125 13.775 138.170 ;
        RECT 21.060 138.110 21.380 138.170 ;
        RECT 22.440 138.310 22.760 138.370 ;
        RECT 23.605 138.310 23.895 138.355 ;
        RECT 28.420 138.310 28.740 138.370 ;
        RECT 22.440 138.170 28.740 138.310 ;
        RECT 22.440 138.110 22.760 138.170 ;
        RECT 23.605 138.125 23.895 138.170 ;
        RECT 28.420 138.110 28.740 138.170 ;
        RECT 32.100 138.310 32.420 138.370 ;
        RECT 33.035 138.310 33.325 138.355 ;
        RECT 32.100 138.170 33.325 138.310 ;
        RECT 32.100 138.110 32.420 138.170 ;
        RECT 33.035 138.125 33.325 138.170 ;
        RECT 46.820 138.110 47.140 138.370 ;
        RECT 51.880 138.110 52.200 138.370 ;
        RECT 52.340 138.310 52.660 138.370 ;
        RECT 54.655 138.310 54.945 138.355 ;
        RECT 52.340 138.170 54.945 138.310 ;
        RECT 52.340 138.110 52.660 138.170 ;
        RECT 54.655 138.125 54.945 138.170 ;
        RECT 75.125 138.310 75.415 138.355 ;
        RECT 76.260 138.310 76.580 138.370 ;
        RECT 75.125 138.170 76.580 138.310 ;
        RECT 75.125 138.125 75.415 138.170 ;
        RECT 76.260 138.110 76.580 138.170 ;
        RECT 86.855 138.310 87.145 138.355 ;
        RECT 89.385 138.310 89.675 138.355 ;
        RECT 90.060 138.310 90.380 138.370 ;
        RECT 96.040 138.310 96.360 138.370 ;
        RECT 102.020 138.310 102.340 138.370 ;
        RECT 86.855 138.170 90.380 138.310 ;
        RECT 86.855 138.125 87.145 138.170 ;
        RECT 89.385 138.125 89.675 138.170 ;
        RECT 90.060 138.110 90.380 138.170 ;
        RECT 91.070 138.170 102.340 138.310 ;
        RECT 15.490 137.970 15.780 138.015 ;
        RECT 17.840 137.970 18.160 138.030 ;
        RECT 18.750 137.970 19.040 138.015 ;
        RECT 15.490 137.830 19.040 137.970 ;
        RECT 15.490 137.785 15.780 137.830 ;
        RECT 17.840 137.770 18.160 137.830 ;
        RECT 18.750 137.785 19.040 137.830 ;
        RECT 19.670 137.970 19.960 138.015 ;
        RECT 21.530 137.970 21.820 138.015 ;
        RECT 19.670 137.830 21.820 137.970 ;
        RECT 19.670 137.785 19.960 137.830 ;
        RECT 21.530 137.785 21.820 137.830 ;
        RECT 24.740 137.970 25.060 138.030 ;
        RECT 25.610 137.970 25.900 138.015 ;
        RECT 28.870 137.970 29.160 138.015 ;
        RECT 24.740 137.830 29.160 137.970 ;
        RECT 17.350 137.630 17.640 137.675 ;
        RECT 19.670 137.630 19.885 137.785 ;
        RECT 24.740 137.770 25.060 137.830 ;
        RECT 25.610 137.785 25.900 137.830 ;
        RECT 28.870 137.785 29.160 137.830 ;
        RECT 29.790 137.970 30.080 138.015 ;
        RECT 31.650 137.970 31.940 138.015 ;
        RECT 46.910 137.970 47.050 138.110 ;
        RECT 59.700 137.970 60.020 138.030 ;
        RECT 60.620 137.970 60.940 138.030 ;
        RECT 63.855 137.970 64.145 138.015 ;
        RECT 29.790 137.830 31.940 137.970 ;
        RECT 29.790 137.785 30.080 137.830 ;
        RECT 31.650 137.785 31.940 137.830 ;
        RECT 34.030 137.830 38.310 137.970 ;
        RECT 46.910 137.830 51.650 137.970 ;
        RECT 17.350 137.490 19.885 137.630 ;
        RECT 27.470 137.630 27.760 137.675 ;
        RECT 29.790 137.630 30.005 137.785 ;
        RECT 27.470 137.490 30.005 137.630 ;
        RECT 17.350 137.445 17.640 137.490 ;
        RECT 27.470 137.445 27.760 137.490 ;
        RECT 30.720 137.430 31.040 137.690 ;
        RECT 31.180 137.630 31.500 137.690 ;
        RECT 34.030 137.675 34.170 137.830 ;
        RECT 33.955 137.630 34.245 137.675 ;
        RECT 31.180 137.490 34.245 137.630 ;
        RECT 31.180 137.430 31.500 137.490 ;
        RECT 33.955 137.445 34.245 137.490 ;
        RECT 35.320 137.630 35.640 137.690 ;
        RECT 37.175 137.630 37.465 137.675 ;
        RECT 35.320 137.490 37.465 137.630 ;
        RECT 35.320 137.430 35.640 137.490 ;
        RECT 37.175 137.445 37.465 137.490 ;
        RECT 37.620 137.430 37.940 137.690 ;
        RECT 20.600 137.090 20.920 137.350 ;
        RECT 22.455 137.290 22.745 137.335 ;
        RECT 24.740 137.290 25.060 137.350 ;
        RECT 32.575 137.290 32.865 137.335 ;
        RECT 22.455 137.150 32.865 137.290 ;
        RECT 22.455 137.105 22.745 137.150 ;
        RECT 24.740 137.090 25.060 137.150 ;
        RECT 32.575 137.105 32.865 137.150 ;
        RECT 34.875 137.105 35.165 137.335 ;
        RECT 17.350 136.950 17.640 136.995 ;
        RECT 20.130 136.950 20.420 136.995 ;
        RECT 21.990 136.950 22.280 136.995 ;
        RECT 17.350 136.810 22.280 136.950 ;
        RECT 17.350 136.765 17.640 136.810 ;
        RECT 20.130 136.765 20.420 136.810 ;
        RECT 21.990 136.765 22.280 136.810 ;
        RECT 27.470 136.950 27.760 136.995 ;
        RECT 30.250 136.950 30.540 136.995 ;
        RECT 32.110 136.950 32.400 136.995 ;
        RECT 27.470 136.810 32.400 136.950 ;
        RECT 27.470 136.765 27.760 136.810 ;
        RECT 30.250 136.765 30.540 136.810 ;
        RECT 32.110 136.765 32.400 136.810 ;
        RECT 19.680 136.610 20.000 136.670 ;
        RECT 34.950 136.610 35.090 137.105 ;
        RECT 36.240 136.750 36.560 137.010 ;
        RECT 38.170 136.950 38.310 137.830 ;
        RECT 38.540 137.430 38.860 137.690 ;
        RECT 46.360 137.430 46.680 137.690 ;
        RECT 46.835 137.445 47.125 137.675 ;
        RECT 47.295 137.445 47.585 137.675 ;
        RECT 48.215 137.630 48.505 137.675 ;
        RECT 50.040 137.630 50.360 137.690 ;
        RECT 51.510 137.675 51.650 137.830 ;
        RECT 51.970 137.830 60.390 137.970 ;
        RECT 48.215 137.490 50.360 137.630 ;
        RECT 48.215 137.445 48.505 137.490 ;
        RECT 45.440 137.290 45.760 137.350 ;
        RECT 46.910 137.290 47.050 137.445 ;
        RECT 45.440 137.150 47.050 137.290 ;
        RECT 47.370 137.290 47.510 137.445 ;
        RECT 50.040 137.430 50.360 137.490 ;
        RECT 51.435 137.445 51.725 137.675 ;
        RECT 49.580 137.290 49.900 137.350 ;
        RECT 47.370 137.150 49.900 137.290 ;
        RECT 45.440 137.090 45.760 137.150 ;
        RECT 49.580 137.090 49.900 137.150 ;
        RECT 51.970 136.950 52.110 137.830 ;
        RECT 59.700 137.770 60.020 137.830 ;
        RECT 57.875 137.630 58.165 137.675 ;
        RECT 56.570 137.490 58.165 137.630 ;
        RECT 60.250 137.630 60.390 137.830 ;
        RECT 60.620 137.830 64.145 137.970 ;
        RECT 60.620 137.770 60.940 137.830 ;
        RECT 63.855 137.785 64.145 137.830 ;
        RECT 70.280 137.770 70.600 138.030 ;
        RECT 73.515 137.970 73.805 138.015 ;
        RECT 77.130 137.970 77.420 138.015 ;
        RECT 80.390 137.970 80.680 138.015 ;
        RECT 73.515 137.830 80.680 137.970 ;
        RECT 73.515 137.785 73.805 137.830 ;
        RECT 77.130 137.785 77.420 137.830 ;
        RECT 80.390 137.785 80.680 137.830 ;
        RECT 81.310 137.970 81.600 138.015 ;
        RECT 83.170 137.970 83.460 138.015 ;
        RECT 91.070 137.970 91.210 138.170 ;
        RECT 96.040 138.110 96.360 138.170 ;
        RECT 81.310 137.830 83.460 137.970 ;
        RECT 81.310 137.785 81.600 137.830 ;
        RECT 83.170 137.785 83.460 137.830 ;
        RECT 85.550 137.830 91.210 137.970 ;
        RECT 91.390 137.970 91.680 138.015 ;
        RECT 93.740 137.970 94.060 138.030 ;
        RECT 94.650 137.970 94.940 138.015 ;
        RECT 91.390 137.830 94.940 137.970 ;
        RECT 62.935 137.630 63.225 137.675 ;
        RECT 60.250 137.490 63.225 137.630 ;
        RECT 53.720 137.090 54.040 137.350 ;
        RECT 54.180 137.090 54.500 137.350 ;
        RECT 56.570 136.995 56.710 137.490 ;
        RECT 57.875 137.445 58.165 137.490 ;
        RECT 62.935 137.445 63.225 137.490 ;
        RECT 68.900 137.430 69.220 137.690 ;
        RECT 69.360 137.430 69.680 137.690 ;
        RECT 73.960 137.630 74.280 137.690 ;
        RECT 75.800 137.630 76.120 137.690 ;
        RECT 73.960 137.490 76.120 137.630 ;
        RECT 73.960 137.430 74.280 137.490 ;
        RECT 75.800 137.430 76.120 137.490 ;
        RECT 78.990 137.630 79.280 137.675 ;
        RECT 81.310 137.630 81.525 137.785 ;
        RECT 78.990 137.490 81.525 137.630 ;
        RECT 78.990 137.445 79.280 137.490 ;
        RECT 84.080 137.430 84.400 137.690 ;
        RECT 80.400 137.290 80.720 137.350 ;
        RECT 85.550 137.335 85.690 137.830 ;
        RECT 91.390 137.785 91.680 137.830 ;
        RECT 93.740 137.770 94.060 137.830 ;
        RECT 94.650 137.785 94.940 137.830 ;
        RECT 95.570 137.970 95.860 138.015 ;
        RECT 97.430 137.970 97.720 138.015 ;
        RECT 95.570 137.830 97.720 137.970 ;
        RECT 95.570 137.785 95.860 137.830 ;
        RECT 97.430 137.785 97.720 137.830 ;
        RECT 93.250 137.630 93.540 137.675 ;
        RECT 95.570 137.630 95.785 137.785 ;
        RECT 93.250 137.490 95.785 137.630 ;
        RECT 93.250 137.445 93.540 137.490 ;
        RECT 98.340 137.430 98.660 137.690 ;
        RECT 82.255 137.290 82.545 137.335 ;
        RECT 85.475 137.290 85.765 137.335 ;
        RECT 80.400 137.150 82.545 137.290 ;
        RECT 80.400 137.090 80.720 137.150 ;
        RECT 82.255 137.105 82.545 137.150 ;
        RECT 85.090 137.150 85.765 137.290 ;
        RECT 38.170 136.810 52.110 136.950 ;
        RECT 56.495 136.765 56.785 136.995 ;
        RECT 78.990 136.950 79.280 136.995 ;
        RECT 81.770 136.950 82.060 136.995 ;
        RECT 83.630 136.950 83.920 136.995 ;
        RECT 78.990 136.810 83.920 136.950 ;
        RECT 78.990 136.765 79.280 136.810 ;
        RECT 81.770 136.765 82.060 136.810 ;
        RECT 83.630 136.765 83.920 136.810 ;
        RECT 19.680 136.470 35.090 136.610 ;
        RECT 35.320 136.610 35.640 136.670 ;
        RECT 37.175 136.610 37.465 136.655 ;
        RECT 35.320 136.470 37.465 136.610 ;
        RECT 19.680 136.410 20.000 136.470 ;
        RECT 35.320 136.410 35.640 136.470 ;
        RECT 37.175 136.425 37.465 136.470 ;
        RECT 40.380 136.610 40.700 136.670 ;
        RECT 44.995 136.610 45.285 136.655 ;
        RECT 40.380 136.470 45.285 136.610 ;
        RECT 40.380 136.410 40.700 136.470 ;
        RECT 44.995 136.425 45.285 136.470 ;
        RECT 58.795 136.610 59.085 136.655 ;
        RECT 59.240 136.610 59.560 136.670 ;
        RECT 58.795 136.470 59.560 136.610 ;
        RECT 58.795 136.425 59.085 136.470 ;
        RECT 59.240 136.410 59.560 136.470 ;
        RECT 67.995 136.610 68.285 136.655 ;
        RECT 68.440 136.610 68.760 136.670 ;
        RECT 67.995 136.470 68.760 136.610 ;
        RECT 67.995 136.425 68.285 136.470 ;
        RECT 68.440 136.410 68.760 136.470 ;
        RECT 69.820 136.410 70.140 136.670 ;
        RECT 74.420 136.610 74.740 136.670 ;
        RECT 85.090 136.610 85.230 137.150 ;
        RECT 85.475 137.105 85.765 137.150 ;
        RECT 85.920 137.290 86.240 137.350 ;
        RECT 86.395 137.290 86.685 137.335 ;
        RECT 85.920 137.150 86.685 137.290 ;
        RECT 85.920 137.090 86.240 137.150 ;
        RECT 86.395 137.105 86.685 137.150 ;
        RECT 96.500 137.090 96.820 137.350 ;
        RECT 101.650 137.335 101.790 138.170 ;
        RECT 102.020 138.110 102.340 138.170 ;
        RECT 102.480 138.110 102.800 138.370 ;
        RECT 102.940 138.110 103.260 138.370 ;
        RECT 104.795 138.125 105.085 138.355 ;
        RECT 107.095 138.310 107.385 138.355 ;
        RECT 108.000 138.310 108.320 138.370 ;
        RECT 107.095 138.170 108.320 138.310 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 107.095 138.125 107.385 138.170 ;
        RECT 104.870 137.630 105.010 138.125 ;
        RECT 108.000 138.110 108.320 138.170 ;
        RECT 106.175 137.630 106.465 137.675 ;
        RECT 104.870 137.490 106.465 137.630 ;
        RECT 106.175 137.445 106.465 137.490 ;
        RECT 101.575 137.105 101.865 137.335 ;
        RECT 93.250 136.950 93.540 136.995 ;
        RECT 96.030 136.950 96.320 136.995 ;
        RECT 97.890 136.950 98.180 136.995 ;
        RECT 93.250 136.810 98.180 136.950 ;
        RECT 93.250 136.765 93.540 136.810 ;
        RECT 96.030 136.765 96.320 136.810 ;
        RECT 97.890 136.765 98.180 136.810 ;
        RECT 74.420 136.470 85.230 136.610 ;
        RECT 88.695 136.610 88.985 136.655 ;
        RECT 90.060 136.610 90.380 136.670 ;
        RECT 88.695 136.470 90.380 136.610 ;
        RECT 74.420 136.410 74.740 136.470 ;
        RECT 88.695 136.425 88.985 136.470 ;
        RECT 90.060 136.410 90.380 136.470 ;
        RECT 11.330 135.790 113.450 136.270 ;
        RECT 20.600 135.590 20.920 135.650 ;
        RECT 21.075 135.590 21.365 135.635 ;
        RECT 20.600 135.450 21.365 135.590 ;
        RECT 20.600 135.390 20.920 135.450 ;
        RECT 21.075 135.405 21.365 135.450 ;
        RECT 26.135 135.590 26.425 135.635 ;
        RECT 30.720 135.590 31.040 135.650 ;
        RECT 26.135 135.450 31.040 135.590 ;
        RECT 26.135 135.405 26.425 135.450 ;
        RECT 30.720 135.390 31.040 135.450 ;
        RECT 35.320 135.390 35.640 135.650 ;
        RECT 38.080 135.390 38.400 135.650 ;
        RECT 38.540 135.590 38.860 135.650 ;
        RECT 43.615 135.590 43.905 135.635 ;
        RECT 38.540 135.450 43.905 135.590 ;
        RECT 38.540 135.390 38.860 135.450 ;
        RECT 43.615 135.405 43.905 135.450 ;
        RECT 44.520 135.590 44.840 135.650 ;
        RECT 46.360 135.590 46.680 135.650 ;
        RECT 48.660 135.590 48.980 135.650 ;
        RECT 44.520 135.450 48.980 135.590 ;
        RECT 44.520 135.390 44.840 135.450 ;
        RECT 46.360 135.390 46.680 135.450 ;
        RECT 48.660 135.390 48.980 135.450 ;
        RECT 54.730 135.450 61.310 135.590 ;
        RECT 26.595 135.065 26.885 135.295 ;
        RECT 45.440 135.250 45.760 135.310 ;
        RECT 50.040 135.250 50.360 135.310 ;
        RECT 54.730 135.250 54.870 135.450 ;
        RECT 41.850 135.110 45.760 135.250 ;
        RECT 17.395 134.725 17.685 134.955 ;
        RECT 17.855 134.910 18.145 134.955 ;
        RECT 21.060 134.910 21.380 134.970 ;
        RECT 17.855 134.770 21.380 134.910 ;
        RECT 17.855 134.725 18.145 134.770 ;
        RECT 17.470 134.230 17.610 134.725 ;
        RECT 21.060 134.710 21.380 134.770 ;
        RECT 18.300 134.570 18.620 134.630 ;
        RECT 19.680 134.570 20.000 134.630 ;
        RECT 18.300 134.430 20.000 134.570 ;
        RECT 18.300 134.370 18.620 134.430 ;
        RECT 19.680 134.370 20.000 134.430 ;
        RECT 21.980 134.370 22.300 134.630 ;
        RECT 25.215 134.570 25.505 134.615 ;
        RECT 26.670 134.570 26.810 135.065 ;
        RECT 29.815 134.910 30.105 134.955 ;
        RECT 32.100 134.910 32.420 134.970 ;
        RECT 29.815 134.770 32.420 134.910 ;
        RECT 29.815 134.725 30.105 134.770 ;
        RECT 32.100 134.710 32.420 134.770 ;
        RECT 39.000 134.710 39.320 134.970 ;
        RECT 25.215 134.430 26.810 134.570 ;
        RECT 25.215 134.385 25.505 134.430 ;
        RECT 28.420 134.370 28.740 134.630 ;
        RECT 33.955 134.385 34.245 134.615 ;
        RECT 34.415 134.570 34.705 134.615 ;
        RECT 35.320 134.570 35.640 134.630 ;
        RECT 34.415 134.430 35.640 134.570 ;
        RECT 34.415 134.385 34.705 134.430 ;
        RECT 20.600 134.230 20.920 134.290 ;
        RECT 17.470 134.090 20.920 134.230 ;
        RECT 20.600 134.030 20.920 134.090 ;
        RECT 28.895 134.230 29.185 134.275 ;
        RECT 34.030 134.230 34.170 134.385 ;
        RECT 35.320 134.370 35.640 134.430 ;
        RECT 37.160 134.570 37.480 134.630 ;
        RECT 41.850 134.615 41.990 135.110 ;
        RECT 45.440 135.050 45.760 135.110 ;
        RECT 46.910 135.110 54.870 135.250 ;
        RECT 46.910 134.910 47.050 135.110 ;
        RECT 50.040 135.050 50.360 135.110 ;
        RECT 52.125 134.910 52.415 134.955 ;
        RECT 54.180 134.910 54.500 134.970 ;
        RECT 43.230 134.770 47.050 134.910 ;
        RECT 43.230 134.615 43.370 134.770 ;
        RECT 38.095 134.570 38.385 134.615 ;
        RECT 37.160 134.430 38.385 134.570 ;
        RECT 37.160 134.370 37.480 134.430 ;
        RECT 38.095 134.385 38.385 134.430 ;
        RECT 41.315 134.385 41.605 134.615 ;
        RECT 41.775 134.385 42.065 134.615 ;
        RECT 42.235 134.385 42.525 134.615 ;
        RECT 43.155 134.385 43.445 134.615 ;
        RECT 44.520 134.570 44.840 134.630 ;
        RECT 44.995 134.570 45.285 134.615 ;
        RECT 44.520 134.430 45.285 134.570 ;
        RECT 34.860 134.230 35.180 134.290 ;
        RECT 28.895 134.090 35.180 134.230 ;
        RECT 28.895 134.045 29.185 134.090 ;
        RECT 34.860 134.030 35.180 134.090 ;
        RECT 39.475 134.230 39.765 134.275 ;
        RECT 39.935 134.230 40.225 134.275 ;
        RECT 39.475 134.090 40.225 134.230 ;
        RECT 39.475 134.045 39.765 134.090 ;
        RECT 39.935 134.045 40.225 134.090 ;
        RECT 19.680 133.890 20.000 133.950 ;
        RECT 20.155 133.890 20.445 133.935 ;
        RECT 19.680 133.750 20.445 133.890 ;
        RECT 19.680 133.690 20.000 133.750 ;
        RECT 20.155 133.705 20.445 133.750 ;
        RECT 37.175 133.890 37.465 133.935 ;
        RECT 40.840 133.890 41.160 133.950 ;
        RECT 37.175 133.750 41.160 133.890 ;
        RECT 41.390 133.890 41.530 134.385 ;
        RECT 42.310 134.230 42.450 134.385 ;
        RECT 44.520 134.370 44.840 134.430 ;
        RECT 44.995 134.385 45.285 134.430 ;
        RECT 45.440 134.370 45.760 134.630 ;
        RECT 45.900 134.370 46.220 134.630 ;
        RECT 46.910 134.615 47.050 134.770 ;
        RECT 49.670 134.770 54.500 134.910 ;
        RECT 46.835 134.385 47.125 134.615 ;
        RECT 48.660 134.370 48.980 134.630 ;
        RECT 49.120 134.370 49.440 134.630 ;
        RECT 49.670 134.615 49.810 134.770 ;
        RECT 52.125 134.725 52.415 134.770 ;
        RECT 54.180 134.710 54.500 134.770 ;
        RECT 49.595 134.385 49.885 134.615 ;
        RECT 50.515 134.570 50.805 134.615 ;
        RECT 54.730 134.570 54.870 135.110 ;
        RECT 55.990 135.250 56.280 135.295 ;
        RECT 58.770 135.250 59.060 135.295 ;
        RECT 60.630 135.250 60.920 135.295 ;
        RECT 55.990 135.110 60.920 135.250 ;
        RECT 61.170 135.250 61.310 135.450 ;
        RECT 63.380 135.390 63.700 135.650 ;
        RECT 65.680 135.390 66.000 135.650 ;
        RECT 69.360 135.590 69.680 135.650 ;
        RECT 73.040 135.590 73.360 135.650 ;
        RECT 66.230 135.450 73.360 135.590 ;
        RECT 66.230 135.250 66.370 135.450 ;
        RECT 69.360 135.390 69.680 135.450 ;
        RECT 73.040 135.390 73.360 135.450 ;
        RECT 76.720 135.590 77.040 135.650 ;
        RECT 77.195 135.590 77.485 135.635 ;
        RECT 76.720 135.450 77.485 135.590 ;
        RECT 76.720 135.390 77.040 135.450 ;
        RECT 77.195 135.405 77.485 135.450 ;
        RECT 77.885 135.590 78.175 135.635 ;
        RECT 85.920 135.590 86.240 135.650 ;
        RECT 77.885 135.450 86.240 135.590 ;
        RECT 77.885 135.405 78.175 135.450 ;
        RECT 61.170 135.110 66.370 135.250 ;
        RECT 67.980 135.250 68.300 135.310 ;
        RECT 71.660 135.250 71.980 135.310 ;
        RECT 67.980 135.110 71.980 135.250 ;
        RECT 55.990 135.065 56.280 135.110 ;
        RECT 58.770 135.065 59.060 135.110 ;
        RECT 60.630 135.065 60.920 135.110 ;
        RECT 67.980 135.050 68.300 135.110 ;
        RECT 71.660 135.050 71.980 135.110 ;
        RECT 72.210 135.110 75.110 135.250 ;
        RECT 59.240 134.710 59.560 134.970 ;
        RECT 61.080 134.710 61.400 134.970 ;
        RECT 65.220 134.710 65.540 134.970 ;
        RECT 67.610 134.770 71.430 134.910 ;
        RECT 50.515 134.430 54.870 134.570 ;
        RECT 55.990 134.570 56.280 134.615 ;
        RECT 64.315 134.570 64.605 134.615 ;
        RECT 64.760 134.570 65.080 134.630 ;
        RECT 67.610 134.615 67.750 134.770 ;
        RECT 71.290 134.630 71.430 134.770 ;
        RECT 55.990 134.430 58.525 134.570 ;
        RECT 50.515 134.385 50.805 134.430 ;
        RECT 55.990 134.385 56.280 134.430 ;
        RECT 50.040 134.230 50.360 134.290 ;
        RECT 42.310 134.090 50.360 134.230 ;
        RECT 50.040 134.030 50.360 134.090 ;
        RECT 51.420 134.230 51.740 134.290 ;
        RECT 58.310 134.275 58.525 134.430 ;
        RECT 64.315 134.430 65.080 134.570 ;
        RECT 64.315 134.385 64.605 134.430 ;
        RECT 64.760 134.370 65.080 134.430 ;
        RECT 67.535 134.385 67.825 134.615 ;
        RECT 67.980 134.370 68.300 134.630 ;
        RECT 68.455 134.385 68.745 134.615 ;
        RECT 54.130 134.230 54.420 134.275 ;
        RECT 57.390 134.230 57.680 134.275 ;
        RECT 51.420 134.090 57.680 134.230 ;
        RECT 51.420 134.030 51.740 134.090 ;
        RECT 54.130 134.045 54.420 134.090 ;
        RECT 57.390 134.045 57.680 134.090 ;
        RECT 58.310 134.230 58.600 134.275 ;
        RECT 60.170 134.230 60.460 134.275 ;
        RECT 58.310 134.090 60.460 134.230 ;
        RECT 58.310 134.045 58.600 134.090 ;
        RECT 60.170 134.045 60.460 134.090 ;
        RECT 65.695 134.230 65.985 134.275 ;
        RECT 66.155 134.230 66.445 134.275 ;
        RECT 65.695 134.090 66.445 134.230 ;
        RECT 68.530 134.230 68.670 134.385 ;
        RECT 69.360 134.370 69.680 134.630 ;
        RECT 71.200 134.370 71.520 134.630 ;
        RECT 71.750 134.615 71.890 135.050 ;
        RECT 72.210 134.615 72.350 135.110 ;
        RECT 74.970 134.970 75.110 135.110 ;
        RECT 74.420 134.710 74.740 134.970 ;
        RECT 74.880 134.710 75.200 134.970 ;
        RECT 71.675 134.385 71.965 134.615 ;
        RECT 72.135 134.385 72.425 134.615 ;
        RECT 73.040 134.370 73.360 134.630 ;
        RECT 75.355 134.570 75.645 134.615 ;
        RECT 77.960 134.570 78.100 135.405 ;
        RECT 85.920 135.390 86.240 135.450 ;
        RECT 93.295 135.590 93.585 135.635 ;
        RECT 93.740 135.590 94.060 135.650 ;
        RECT 93.295 135.450 94.060 135.590 ;
        RECT 93.295 135.405 93.585 135.450 ;
        RECT 93.740 135.390 94.060 135.450 ;
        RECT 96.055 135.590 96.345 135.635 ;
        RECT 96.500 135.590 96.820 135.650 ;
        RECT 96.055 135.450 96.820 135.590 ;
        RECT 96.055 135.405 96.345 135.450 ;
        RECT 96.500 135.390 96.820 135.450 ;
        RECT 81.750 135.250 82.040 135.295 ;
        RECT 84.530 135.250 84.820 135.295 ;
        RECT 86.390 135.250 86.680 135.295 ;
        RECT 81.750 135.110 86.680 135.250 ;
        RECT 81.750 135.065 82.040 135.110 ;
        RECT 84.530 135.065 84.820 135.110 ;
        RECT 86.390 135.065 86.680 135.110 ;
        RECT 89.155 135.065 89.445 135.295 ;
        RECT 84.080 134.910 84.400 134.970 ;
        RECT 85.015 134.910 85.305 134.955 ;
        RECT 89.230 134.910 89.370 135.065 ;
        RECT 104.320 134.910 104.640 134.970 ;
        RECT 84.080 134.770 84.770 134.910 ;
        RECT 84.080 134.710 84.400 134.770 ;
        RECT 75.355 134.430 78.100 134.570 ;
        RECT 81.750 134.570 82.040 134.615 ;
        RECT 84.630 134.570 84.770 134.770 ;
        RECT 85.015 134.770 89.370 134.910 ;
        RECT 89.690 134.770 104.640 134.910 ;
        RECT 85.015 134.725 85.305 134.770 ;
        RECT 89.690 134.630 89.830 134.770 ;
        RECT 86.855 134.570 87.145 134.615 ;
        RECT 81.750 134.430 84.285 134.570 ;
        RECT 84.630 134.430 87.145 134.570 ;
        RECT 75.355 134.385 75.645 134.430 ;
        RECT 81.750 134.385 82.040 134.430 ;
        RECT 75.430 134.230 75.570 134.385 ;
        RECT 84.070 134.275 84.285 134.430 ;
        RECT 86.855 134.385 87.145 134.430 ;
        RECT 88.695 134.570 88.985 134.615 ;
        RECT 89.600 134.570 89.920 134.630 ;
        RECT 88.695 134.430 89.920 134.570 ;
        RECT 88.695 134.385 88.985 134.430 ;
        RECT 89.600 134.370 89.920 134.430 ;
        RECT 90.060 134.370 90.380 134.630 ;
        RECT 93.830 134.615 93.970 134.770 ;
        RECT 104.320 134.710 104.640 134.770 ;
        RECT 93.755 134.385 94.045 134.615 ;
        RECT 96.960 134.370 97.280 134.630 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 68.530 134.090 75.570 134.230 ;
        RECT 79.890 134.230 80.180 134.275 ;
        RECT 83.150 134.230 83.440 134.275 ;
        RECT 84.070 134.230 84.360 134.275 ;
        RECT 85.930 134.230 86.220 134.275 ;
        RECT 79.890 134.090 83.850 134.230 ;
        RECT 65.695 134.045 65.985 134.090 ;
        RECT 66.155 134.045 66.445 134.090 ;
        RECT 79.890 134.045 80.180 134.090 ;
        RECT 83.150 134.045 83.440 134.090 ;
        RECT 44.520 133.890 44.840 133.950 ;
        RECT 41.390 133.750 44.840 133.890 ;
        RECT 37.175 133.705 37.465 133.750 ;
        RECT 40.840 133.690 41.160 133.750 ;
        RECT 44.520 133.690 44.840 133.750 ;
        RECT 47.280 133.690 47.600 133.950 ;
        RECT 67.980 133.890 68.300 133.950 ;
        RECT 69.835 133.890 70.125 133.935 ;
        RECT 67.980 133.750 70.125 133.890 ;
        RECT 83.710 133.890 83.850 134.090 ;
        RECT 84.070 134.090 86.220 134.230 ;
        RECT 84.070 134.045 84.360 134.090 ;
        RECT 85.930 134.045 86.220 134.090 ;
        RECT 88.235 133.890 88.525 133.935 ;
        RECT 83.710 133.750 88.525 133.890 ;
        RECT 67.980 133.690 68.300 133.750 ;
        RECT 69.835 133.705 70.125 133.750 ;
        RECT 88.235 133.705 88.525 133.750 ;
        RECT 11.330 133.070 113.450 133.550 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 34.860 132.670 35.180 132.930 ;
        RECT 38.080 132.670 38.400 132.930 ;
        RECT 42.680 132.670 43.000 132.930 ;
        RECT 43.155 132.870 43.445 132.915 ;
        RECT 43.600 132.870 43.920 132.930 ;
        RECT 43.155 132.730 43.920 132.870 ;
        RECT 43.155 132.685 43.445 132.730 ;
        RECT 43.600 132.670 43.920 132.730 ;
        RECT 51.420 132.670 51.740 132.930 ;
        RECT 54.180 132.670 54.500 132.930 ;
        RECT 74.880 132.915 75.200 132.930 ;
        RECT 56.035 132.870 56.325 132.915 ;
        RECT 56.035 132.730 56.940 132.870 ;
        RECT 56.035 132.685 56.325 132.730 ;
        RECT 15.030 132.530 15.320 132.575 ;
        RECT 16.460 132.530 16.780 132.590 ;
        RECT 18.290 132.530 18.580 132.575 ;
        RECT 15.030 132.390 18.580 132.530 ;
        RECT 15.030 132.345 15.320 132.390 ;
        RECT 16.460 132.330 16.780 132.390 ;
        RECT 18.290 132.345 18.580 132.390 ;
        RECT 19.210 132.530 19.500 132.575 ;
        RECT 21.070 132.530 21.360 132.575 ;
        RECT 25.200 132.530 25.520 132.590 ;
        RECT 19.210 132.390 21.360 132.530 ;
        RECT 19.210 132.345 19.500 132.390 ;
        RECT 21.070 132.345 21.360 132.390 ;
        RECT 23.450 132.390 25.520 132.530 ;
        RECT 16.890 132.190 17.180 132.235 ;
        RECT 19.210 132.190 19.425 132.345 ;
        RECT 16.890 132.050 19.425 132.190 ;
        RECT 22.440 132.190 22.760 132.250 ;
        RECT 23.450 132.235 23.590 132.390 ;
        RECT 25.200 132.330 25.520 132.390 ;
        RECT 31.195 132.530 31.485 132.575 ;
        RECT 34.950 132.530 35.090 132.670 ;
        RECT 31.195 132.390 35.090 132.530 ;
        RECT 31.195 132.345 31.485 132.390 ;
        RECT 40.380 132.330 40.700 132.590 ;
        RECT 45.455 132.530 45.745 132.575 ;
        RECT 47.280 132.530 47.600 132.590 ;
        RECT 45.455 132.390 47.600 132.530 ;
        RECT 45.455 132.345 45.745 132.390 ;
        RECT 47.280 132.330 47.600 132.390 ;
        RECT 23.375 132.190 23.665 132.235 ;
        RECT 22.440 132.050 23.665 132.190 ;
        RECT 16.890 132.005 17.180 132.050 ;
        RECT 22.440 131.990 22.760 132.050 ;
        RECT 23.375 132.005 23.665 132.050 ;
        RECT 23.835 132.190 24.125 132.235 ;
        RECT 27.040 132.190 27.360 132.250 ;
        RECT 34.875 132.190 35.165 132.235 ;
        RECT 35.320 132.190 35.640 132.250 ;
        RECT 37.175 132.190 37.465 132.235 ;
        RECT 23.835 132.050 27.360 132.190 ;
        RECT 23.835 132.005 24.125 132.050 ;
        RECT 27.040 131.990 27.360 132.050 ;
        RECT 31.730 132.050 34.525 132.190 ;
        RECT 31.730 131.910 31.870 132.050 ;
        RECT 13.025 131.850 13.315 131.895 ;
        RECT 16.000 131.850 16.320 131.910 ;
        RECT 18.300 131.850 18.620 131.910 ;
        RECT 13.025 131.710 18.620 131.850 ;
        RECT 13.025 131.665 13.315 131.710 ;
        RECT 16.000 131.650 16.320 131.710 ;
        RECT 18.300 131.650 18.620 131.710 ;
        RECT 20.140 131.650 20.460 131.910 ;
        RECT 21.995 131.850 22.285 131.895 ;
        RECT 24.740 131.850 25.060 131.910 ;
        RECT 21.995 131.710 25.060 131.850 ;
        RECT 21.995 131.665 22.285 131.710 ;
        RECT 24.740 131.650 25.060 131.710 ;
        RECT 31.640 131.650 31.960 131.910 ;
        RECT 32.100 131.650 32.420 131.910 ;
        RECT 33.955 131.665 34.245 131.895 ;
        RECT 16.890 131.510 17.180 131.555 ;
        RECT 19.670 131.510 19.960 131.555 ;
        RECT 21.530 131.510 21.820 131.555 ;
        RECT 16.890 131.370 21.820 131.510 ;
        RECT 16.890 131.325 17.180 131.370 ;
        RECT 19.670 131.325 19.960 131.370 ;
        RECT 21.530 131.325 21.820 131.370 ;
        RECT 26.120 131.170 26.440 131.230 ;
        RECT 29.355 131.170 29.645 131.215 ;
        RECT 26.120 131.030 29.645 131.170 ;
        RECT 26.120 130.970 26.440 131.030 ;
        RECT 29.355 130.985 29.645 131.030 ;
        RECT 29.800 131.170 30.120 131.230 ;
        RECT 34.030 131.170 34.170 131.665 ;
        RECT 34.385 131.510 34.525 132.050 ;
        RECT 34.875 132.050 37.465 132.190 ;
        RECT 34.875 132.005 35.165 132.050 ;
        RECT 35.320 131.990 35.640 132.050 ;
        RECT 37.175 132.005 37.465 132.050 ;
        RECT 35.780 131.650 36.100 131.910 ;
        RECT 36.255 131.665 36.545 131.895 ;
        RECT 36.330 131.510 36.470 131.665 ;
        RECT 34.385 131.370 36.470 131.510 ;
        RECT 37.250 131.510 37.390 132.005 ;
        RECT 41.760 131.990 42.080 132.250 ;
        RECT 44.060 131.990 44.380 132.250 ;
        RECT 46.820 132.190 47.140 132.250 ;
        RECT 50.975 132.190 51.265 132.235 ;
        RECT 46.820 132.050 51.265 132.190 ;
        RECT 56.800 132.190 56.940 132.730 ;
        RECT 74.880 132.685 75.415 132.915 ;
        RECT 75.800 132.870 76.120 132.930 ;
        RECT 89.600 132.870 89.920 132.930 ;
        RECT 75.800 132.730 89.920 132.870 ;
        RECT 74.880 132.670 75.200 132.685 ;
        RECT 75.800 132.670 76.120 132.730 ;
        RECT 89.600 132.670 89.920 132.730 ;
        RECT 97.420 132.670 97.740 132.930 ;
        RECT 97.880 132.670 98.200 132.930 ;
        RECT 60.620 132.530 60.940 132.590 ;
        RECT 62.475 132.530 62.765 132.575 ;
        RECT 60.620 132.390 64.530 132.530 ;
        RECT 60.620 132.330 60.940 132.390 ;
        RECT 62.475 132.345 62.765 132.390 ;
        RECT 57.415 132.190 57.705 132.235 ;
        RECT 56.800 132.050 57.705 132.190 ;
        RECT 46.820 131.990 47.140 132.050 ;
        RECT 50.975 132.005 51.265 132.050 ;
        RECT 57.415 132.005 57.705 132.050 ;
        RECT 61.540 131.990 61.860 132.250 ;
        RECT 64.390 132.235 64.530 132.390 ;
        RECT 67.980 132.330 68.300 132.590 ;
        RECT 70.740 132.330 71.060 132.590 ;
        RECT 77.130 132.530 77.420 132.575 ;
        RECT 79.480 132.530 79.800 132.590 ;
        RECT 80.390 132.530 80.680 132.575 ;
        RECT 77.130 132.390 80.680 132.530 ;
        RECT 77.130 132.345 77.420 132.390 ;
        RECT 79.480 132.330 79.800 132.390 ;
        RECT 80.390 132.345 80.680 132.390 ;
        RECT 81.310 132.530 81.600 132.575 ;
        RECT 83.170 132.530 83.460 132.575 ;
        RECT 81.310 132.390 83.460 132.530 ;
        RECT 81.310 132.345 81.600 132.390 ;
        RECT 83.170 132.345 83.460 132.390 ;
        RECT 90.060 132.530 90.380 132.590 ;
        RECT 101.560 132.530 101.880 132.590 ;
        RECT 90.060 132.390 91.210 132.530 ;
        RECT 64.315 132.005 64.605 132.235 ;
        RECT 69.375 132.190 69.665 132.235 ;
        RECT 70.830 132.190 70.970 132.330 ;
        RECT 69.375 132.050 70.970 132.190 ;
        RECT 69.375 132.005 69.665 132.050 ;
        RECT 71.675 132.005 71.965 132.235 ;
        RECT 78.990 132.190 79.280 132.235 ;
        RECT 81.310 132.190 81.525 132.345 ;
        RECT 90.060 132.330 90.380 132.390 ;
        RECT 78.990 132.050 81.525 132.190 ;
        RECT 78.990 132.005 79.280 132.050 ;
        RECT 41.300 131.650 41.620 131.910 ;
        RECT 44.980 131.650 45.300 131.910 ;
        RECT 53.260 131.650 53.580 131.910 ;
        RECT 53.735 131.665 54.025 131.895 ;
        RECT 60.620 131.850 60.940 131.910 ;
        RECT 61.630 131.850 61.770 131.990 ;
        RECT 60.620 131.710 61.770 131.850 ;
        RECT 65.235 131.850 65.525 131.895 ;
        RECT 66.140 131.850 66.460 131.910 ;
        RECT 67.520 131.850 67.840 131.910 ;
        RECT 65.235 131.710 67.840 131.850 ;
        RECT 49.580 131.510 49.900 131.570 ;
        RECT 53.810 131.510 53.950 131.665 ;
        RECT 60.620 131.650 60.940 131.710 ;
        RECT 65.235 131.665 65.525 131.710 ;
        RECT 66.140 131.650 66.460 131.710 ;
        RECT 67.520 131.650 67.840 131.710 ;
        RECT 68.900 131.650 69.220 131.910 ;
        RECT 70.280 131.850 70.600 131.910 ;
        RECT 70.755 131.850 71.045 131.895 ;
        RECT 70.280 131.710 71.045 131.850 ;
        RECT 70.280 131.650 70.600 131.710 ;
        RECT 70.755 131.665 71.045 131.710 ;
        RECT 61.540 131.510 61.860 131.570 ;
        RECT 71.750 131.510 71.890 132.005 ;
        RECT 90.520 131.990 90.840 132.250 ;
        RECT 91.070 132.235 91.210 132.390 ;
        RECT 94.290 132.390 96.730 132.530 ;
        RECT 94.290 132.235 94.430 132.390 ;
        RECT 96.590 132.235 96.730 132.390 ;
        RECT 101.560 132.390 107.310 132.530 ;
        RECT 101.560 132.330 101.880 132.390 ;
        RECT 90.995 132.190 91.285 132.235 ;
        RECT 94.215 132.190 94.505 132.235 ;
        RECT 90.995 132.050 94.505 132.190 ;
        RECT 90.995 132.005 91.285 132.050 ;
        RECT 94.215 132.005 94.505 132.050 ;
        RECT 95.135 132.005 95.425 132.235 ;
        RECT 96.055 132.005 96.345 132.235 ;
        RECT 96.515 132.005 96.805 132.235 ;
        RECT 98.815 132.005 99.105 132.235 ;
        RECT 104.795 132.005 105.085 132.235 ;
        RECT 72.595 131.850 72.885 131.895 ;
        RECT 74.420 131.850 74.740 131.910 ;
        RECT 72.595 131.710 74.740 131.850 ;
        RECT 72.595 131.665 72.885 131.710 ;
        RECT 74.420 131.650 74.740 131.710 ;
        RECT 82.240 131.650 82.560 131.910 ;
        RECT 84.095 131.850 84.385 131.895 ;
        RECT 92.360 131.850 92.680 131.910 ;
        RECT 84.095 131.710 92.680 131.850 ;
        RECT 95.210 131.850 95.350 132.005 ;
        RECT 95.210 131.710 95.810 131.850 ;
        RECT 84.095 131.665 84.385 131.710 ;
        RECT 92.360 131.650 92.680 131.710 ;
        RECT 37.250 131.370 44.750 131.510 ;
        RECT 44.610 131.230 44.750 131.370 ;
        RECT 49.580 131.370 53.950 131.510 ;
        RECT 56.800 131.370 71.890 131.510 ;
        RECT 78.990 131.510 79.280 131.555 ;
        RECT 81.770 131.510 82.060 131.555 ;
        RECT 83.630 131.510 83.920 131.555 ;
        RECT 78.990 131.370 83.920 131.510 ;
        RECT 49.580 131.310 49.900 131.370 ;
        RECT 29.800 131.030 34.170 131.170 ;
        RECT 35.320 131.170 35.640 131.230 ;
        RECT 40.395 131.170 40.685 131.215 ;
        RECT 35.320 131.030 40.685 131.170 ;
        RECT 29.800 130.970 30.120 131.030 ;
        RECT 35.320 130.970 35.640 131.030 ;
        RECT 40.395 130.985 40.685 131.030 ;
        RECT 43.140 131.170 43.460 131.230 ;
        RECT 44.075 131.170 44.365 131.215 ;
        RECT 43.140 131.030 44.365 131.170 ;
        RECT 43.140 130.970 43.460 131.030 ;
        RECT 44.075 130.985 44.365 131.030 ;
        RECT 44.520 131.170 44.840 131.230 ;
        RECT 56.800 131.170 56.940 131.370 ;
        RECT 61.540 131.310 61.860 131.370 ;
        RECT 78.990 131.325 79.280 131.370 ;
        RECT 81.770 131.325 82.060 131.370 ;
        RECT 83.630 131.325 83.920 131.370 ;
        RECT 91.440 131.510 91.760 131.570 ;
        RECT 91.915 131.510 92.205 131.555 ;
        RECT 91.440 131.370 92.205 131.510 ;
        RECT 91.440 131.310 91.760 131.370 ;
        RECT 91.915 131.325 92.205 131.370 ;
        RECT 93.295 131.510 93.585 131.555 ;
        RECT 95.120 131.510 95.440 131.570 ;
        RECT 93.295 131.370 95.440 131.510 ;
        RECT 93.295 131.325 93.585 131.370 ;
        RECT 95.120 131.310 95.440 131.370 ;
        RECT 44.520 131.030 56.940 131.170 ;
        RECT 58.335 131.170 58.625 131.215 ;
        RECT 58.780 131.170 59.100 131.230 ;
        RECT 58.335 131.030 59.100 131.170 ;
        RECT 44.520 130.970 44.840 131.030 ;
        RECT 58.335 130.985 58.625 131.030 ;
        RECT 58.780 130.970 59.100 131.030 ;
        RECT 63.380 130.970 63.700 131.230 ;
        RECT 69.360 130.970 69.680 131.230 ;
        RECT 70.280 130.970 70.600 131.230 ;
        RECT 95.670 131.170 95.810 131.710 ;
        RECT 96.130 131.510 96.270 132.005 ;
        RECT 96.590 131.850 96.730 132.005 ;
        RECT 98.890 131.850 99.030 132.005 ;
        RECT 96.590 131.710 99.030 131.850 ;
        RECT 99.720 131.650 100.040 131.910 ;
        RECT 104.320 131.850 104.640 131.910 ;
        RECT 104.870 131.850 105.010 132.005 ;
        RECT 105.240 131.990 105.560 132.250 ;
        RECT 107.170 132.235 107.310 132.390 ;
        RECT 107.095 132.005 107.385 132.235 ;
        RECT 104.320 131.710 105.010 131.850 ;
        RECT 104.320 131.650 104.640 131.710 ;
        RECT 98.800 131.510 99.120 131.570 ;
        RECT 96.130 131.370 99.120 131.510 ;
        RECT 98.800 131.310 99.120 131.370 ;
        RECT 99.260 131.170 99.580 131.230 ;
        RECT 95.670 131.030 99.580 131.170 ;
        RECT 99.260 130.970 99.580 131.030 ;
        RECT 108.015 131.170 108.305 131.215 ;
        RECT 109.840 131.170 110.160 131.230 ;
        RECT 108.015 131.030 110.160 131.170 ;
        RECT 108.015 130.985 108.305 131.030 ;
        RECT 109.840 130.970 110.160 131.030 ;
        RECT 11.330 130.350 113.450 130.830 ;
        RECT 16.460 130.150 16.780 130.210 ;
        RECT 16.935 130.150 17.225 130.195 ;
        RECT 16.460 130.010 17.225 130.150 ;
        RECT 16.460 129.950 16.780 130.010 ;
        RECT 16.935 129.965 17.225 130.010 ;
        RECT 20.140 129.950 20.460 130.210 ;
        RECT 24.755 130.150 25.045 130.195 ;
        RECT 28.880 130.150 29.200 130.210 ;
        RECT 24.755 130.010 29.200 130.150 ;
        RECT 24.755 129.965 25.045 130.010 ;
        RECT 28.880 129.950 29.200 130.010 ;
        RECT 34.185 130.150 34.475 130.195 ;
        RECT 34.860 130.150 35.180 130.210 ;
        RECT 34.185 130.010 35.180 130.150 ;
        RECT 34.185 129.965 34.475 130.010 ;
        RECT 34.860 129.950 35.180 130.010 ;
        RECT 39.475 130.150 39.765 130.195 ;
        RECT 39.920 130.150 40.240 130.210 ;
        RECT 39.475 130.010 40.240 130.150 ;
        RECT 39.475 129.965 39.765 130.010 ;
        RECT 39.920 129.950 40.240 130.010 ;
        RECT 41.775 130.150 42.065 130.195 ;
        RECT 43.140 130.150 43.460 130.210 ;
        RECT 41.775 130.010 43.460 130.150 ;
        RECT 41.775 129.965 42.065 130.010 ;
        RECT 43.140 129.950 43.460 130.010 ;
        RECT 49.580 130.150 49.900 130.210 ;
        RECT 51.665 130.150 51.955 130.195 ;
        RECT 60.620 130.150 60.940 130.210 ;
        RECT 49.580 130.010 51.955 130.150 ;
        RECT 49.580 129.950 49.900 130.010 ;
        RECT 51.665 129.965 51.955 130.010 ;
        RECT 52.430 130.010 60.940 130.150 ;
        RECT 21.980 129.810 22.300 129.870 ;
        RECT 18.850 129.670 22.300 129.810 ;
        RECT 17.395 129.130 17.685 129.175 ;
        RECT 18.850 129.130 18.990 129.670 ;
        RECT 21.980 129.610 22.300 129.670 ;
        RECT 22.455 129.810 22.745 129.855 ;
        RECT 25.200 129.810 25.520 129.870 ;
        RECT 22.455 129.670 25.520 129.810 ;
        RECT 22.455 129.625 22.745 129.670 ;
        RECT 25.200 129.610 25.520 129.670 ;
        RECT 25.680 129.810 25.970 129.855 ;
        RECT 27.540 129.810 27.830 129.855 ;
        RECT 30.320 129.810 30.610 129.855 ;
        RECT 25.680 129.670 30.610 129.810 ;
        RECT 25.680 129.625 25.970 129.670 ;
        RECT 27.540 129.625 27.830 129.670 ;
        RECT 30.320 129.625 30.610 129.670 ;
        RECT 32.100 129.810 32.420 129.870 ;
        RECT 42.220 129.810 42.540 129.870 ;
        RECT 42.695 129.810 42.985 129.855 ;
        RECT 52.430 129.810 52.570 130.010 ;
        RECT 60.620 129.950 60.940 130.010 ;
        RECT 69.360 129.950 69.680 130.210 ;
        RECT 69.820 129.950 70.140 130.210 ;
        RECT 79.480 129.950 79.800 130.210 ;
        RECT 86.840 129.950 87.160 130.210 ;
        RECT 101.560 129.950 101.880 130.210 ;
        RECT 32.100 129.670 42.985 129.810 ;
        RECT 32.100 129.610 32.420 129.670 ;
        RECT 42.220 129.610 42.540 129.670 ;
        RECT 42.695 129.625 42.985 129.670 ;
        RECT 47.370 129.670 52.570 129.810 ;
        RECT 55.530 129.810 55.820 129.855 ;
        RECT 58.310 129.810 58.600 129.855 ;
        RECT 60.170 129.810 60.460 129.855 ;
        RECT 55.530 129.670 60.460 129.810 ;
        RECT 20.140 129.470 20.460 129.530 ;
        RECT 22.915 129.470 23.205 129.515 ;
        RECT 31.180 129.470 31.500 129.530 ;
        RECT 20.140 129.330 23.205 129.470 ;
        RECT 20.140 129.270 20.460 129.330 ;
        RECT 22.915 129.285 23.205 129.330 ;
        RECT 23.910 129.330 31.500 129.470 ;
        RECT 17.395 128.990 18.990 129.130 ;
        RECT 19.235 129.130 19.525 129.175 ;
        RECT 19.680 129.130 20.000 129.190 ;
        RECT 23.910 129.175 24.050 129.330 ;
        RECT 31.180 129.270 31.500 129.330 ;
        RECT 35.780 129.470 36.100 129.530 ;
        RECT 37.635 129.470 37.925 129.515 ;
        RECT 35.780 129.330 37.925 129.470 ;
        RECT 35.780 129.270 36.100 129.330 ;
        RECT 37.635 129.285 37.925 129.330 ;
        RECT 38.630 129.330 41.070 129.470 ;
        RECT 19.235 128.990 20.000 129.130 ;
        RECT 17.395 128.945 17.685 128.990 ;
        RECT 19.235 128.945 19.525 128.990 ;
        RECT 19.680 128.930 20.000 128.990 ;
        RECT 21.535 128.945 21.825 129.175 ;
        RECT 23.835 128.945 24.125 129.175 ;
        RECT 24.740 129.130 25.060 129.190 ;
        RECT 25.215 129.130 25.505 129.175 ;
        RECT 24.740 128.990 25.505 129.130 ;
        RECT 21.610 128.450 21.750 128.945 ;
        RECT 24.740 128.930 25.060 128.990 ;
        RECT 25.215 128.945 25.505 128.990 ;
        RECT 25.660 129.130 25.980 129.190 ;
        RECT 27.055 129.130 27.345 129.175 ;
        RECT 30.320 129.130 30.610 129.175 ;
        RECT 36.255 129.130 36.545 129.175 ;
        RECT 37.160 129.130 37.480 129.190 ;
        RECT 38.630 129.175 38.770 129.330 ;
        RECT 25.660 128.990 27.345 129.130 ;
        RECT 25.660 128.930 25.980 128.990 ;
        RECT 27.055 128.945 27.345 128.990 ;
        RECT 28.075 128.990 30.610 129.130 ;
        RECT 28.075 128.835 28.290 128.990 ;
        RECT 30.320 128.945 30.610 128.990 ;
        RECT 32.650 128.990 37.480 129.130 ;
        RECT 26.140 128.790 26.430 128.835 ;
        RECT 28.000 128.790 28.290 128.835 ;
        RECT 26.140 128.650 28.290 128.790 ;
        RECT 26.140 128.605 26.430 128.650 ;
        RECT 28.000 128.605 28.290 128.650 ;
        RECT 28.880 128.835 29.200 128.850 ;
        RECT 28.880 128.790 29.210 128.835 ;
        RECT 32.180 128.790 32.470 128.835 ;
        RECT 28.880 128.650 32.470 128.790 ;
        RECT 28.880 128.605 29.210 128.650 ;
        RECT 32.180 128.605 32.470 128.650 ;
        RECT 28.880 128.590 29.200 128.605 ;
        RECT 26.580 128.450 26.900 128.510 ;
        RECT 21.610 128.310 26.900 128.450 ;
        RECT 26.580 128.250 26.900 128.310 ;
        RECT 27.500 128.450 27.820 128.510 ;
        RECT 32.650 128.450 32.790 128.990 ;
        RECT 36.255 128.945 36.545 128.990 ;
        RECT 37.160 128.930 37.480 128.990 ;
        RECT 38.555 128.945 38.845 129.175 ;
        RECT 34.860 128.790 35.180 128.850 ;
        RECT 38.630 128.790 38.770 128.945 ;
        RECT 39.920 128.930 40.240 129.190 ;
        RECT 40.930 129.175 41.070 129.330 ;
        RECT 40.855 129.130 41.145 129.175 ;
        RECT 44.520 129.130 44.840 129.190 ;
        RECT 47.370 129.175 47.510 129.670 ;
        RECT 55.530 129.625 55.820 129.670 ;
        RECT 58.310 129.625 58.600 129.670 ;
        RECT 60.170 129.625 60.460 129.670 ;
        RECT 66.600 129.810 66.920 129.870 ;
        RECT 106.130 129.810 106.420 129.855 ;
        RECT 108.910 129.810 109.200 129.855 ;
        RECT 110.770 129.810 111.060 129.855 ;
        RECT 66.600 129.670 72.810 129.810 ;
        RECT 66.600 129.610 66.920 129.670 ;
        RECT 58.780 129.270 59.100 129.530 ;
        RECT 59.700 129.270 60.020 129.530 ;
        RECT 60.635 129.470 60.925 129.515 ;
        RECT 61.080 129.470 61.400 129.530 ;
        RECT 60.635 129.330 61.400 129.470 ;
        RECT 60.635 129.285 60.925 129.330 ;
        RECT 61.080 129.270 61.400 129.330 ;
        RECT 61.540 129.470 61.860 129.530 ;
        RECT 67.060 129.470 67.380 129.530 ;
        RECT 72.670 129.515 72.810 129.670 ;
        RECT 106.130 129.670 111.060 129.810 ;
        RECT 106.130 129.625 106.420 129.670 ;
        RECT 108.910 129.625 109.200 129.670 ;
        RECT 110.770 129.625 111.060 129.670 ;
        RECT 61.540 129.330 68.670 129.470 ;
        RECT 61.540 129.270 61.860 129.330 ;
        RECT 67.060 129.270 67.380 129.330 ;
        RECT 40.855 128.990 44.840 129.130 ;
        RECT 40.855 128.945 41.145 128.990 ;
        RECT 44.520 128.930 44.840 128.990 ;
        RECT 47.295 128.945 47.585 129.175 ;
        RECT 50.055 128.945 50.345 129.175 ;
        RECT 55.530 129.130 55.820 129.175 ;
        RECT 59.790 129.130 59.930 129.270 ;
        RECT 55.530 128.990 58.065 129.130 ;
        RECT 59.790 128.990 67.290 129.130 ;
        RECT 55.530 128.945 55.820 128.990 ;
        RECT 34.860 128.650 38.770 128.790 ;
        RECT 34.860 128.590 35.180 128.650 ;
        RECT 44.075 128.605 44.365 128.835 ;
        RECT 45.440 128.790 45.760 128.850 ;
        RECT 45.915 128.790 46.205 128.835 ;
        RECT 45.440 128.650 46.205 128.790 ;
        RECT 27.500 128.310 32.790 128.450 ;
        RECT 27.500 128.250 27.820 128.310 ;
        RECT 36.700 128.250 37.020 128.510 ;
        RECT 44.150 128.450 44.290 128.605 ;
        RECT 45.440 128.590 45.760 128.650 ;
        RECT 45.915 128.605 46.205 128.650 ;
        RECT 46.820 128.790 47.140 128.850 ;
        RECT 49.120 128.790 49.440 128.850 ;
        RECT 50.130 128.790 50.270 128.945 ;
        RECT 57.850 128.835 58.065 128.990 ;
        RECT 46.820 128.650 50.270 128.790 ;
        RECT 50.515 128.790 50.805 128.835 ;
        RECT 53.670 128.790 53.960 128.835 ;
        RECT 56.930 128.790 57.220 128.835 ;
        RECT 50.515 128.650 57.220 128.790 ;
        RECT 46.820 128.590 47.140 128.650 ;
        RECT 49.120 128.590 49.440 128.650 ;
        RECT 50.515 128.605 50.805 128.650 ;
        RECT 53.670 128.605 53.960 128.650 ;
        RECT 56.930 128.605 57.220 128.650 ;
        RECT 57.850 128.790 58.140 128.835 ;
        RECT 59.710 128.790 60.000 128.835 ;
        RECT 57.850 128.650 60.000 128.790 ;
        RECT 57.850 128.605 58.140 128.650 ;
        RECT 59.710 128.605 60.000 128.650 ;
        RECT 63.380 128.790 63.700 128.850 ;
        RECT 63.855 128.790 64.145 128.835 ;
        RECT 63.380 128.650 64.145 128.790 ;
        RECT 63.380 128.590 63.700 128.650 ;
        RECT 63.855 128.605 64.145 128.650 ;
        RECT 65.695 128.790 65.985 128.835 ;
        RECT 66.600 128.790 66.920 128.850 ;
        RECT 65.695 128.650 66.920 128.790 ;
        RECT 65.695 128.605 65.985 128.650 ;
        RECT 63.930 128.450 64.070 128.605 ;
        RECT 66.600 128.590 66.920 128.650 ;
        RECT 44.150 128.310 64.070 128.450 ;
        RECT 67.150 128.450 67.290 128.990 ;
        RECT 67.520 128.930 67.840 129.190 ;
        RECT 68.530 129.175 68.670 129.330 ;
        RECT 72.595 129.285 72.885 129.515 ;
        RECT 90.060 129.470 90.380 129.530 ;
        RECT 75.430 129.330 90.380 129.470 ;
        RECT 68.455 129.130 68.745 129.175 ;
        RECT 70.755 129.130 71.045 129.175 ;
        RECT 68.455 128.990 71.045 129.130 ;
        RECT 68.455 128.945 68.745 128.990 ;
        RECT 70.755 128.945 71.045 128.990 ;
        RECT 71.215 128.945 71.505 129.175 ;
        RECT 73.975 129.130 74.265 129.175 ;
        RECT 74.420 129.130 74.740 129.190 ;
        RECT 73.975 128.990 74.740 129.130 ;
        RECT 73.975 128.945 74.265 128.990 ;
        RECT 67.980 128.790 68.300 128.850 ;
        RECT 71.290 128.790 71.430 128.945 ;
        RECT 74.420 128.930 74.740 128.990 ;
        RECT 73.515 128.790 73.805 128.835 ;
        RECT 67.980 128.650 73.805 128.790 ;
        RECT 67.980 128.590 68.300 128.650 ;
        RECT 73.515 128.605 73.805 128.650 ;
        RECT 75.430 128.450 75.570 129.330 ;
        RECT 75.800 129.130 76.120 129.190 ;
        RECT 77.655 129.130 77.945 129.175 ;
        RECT 75.800 128.990 77.945 129.130 ;
        RECT 75.800 128.930 76.120 128.990 ;
        RECT 77.655 128.945 77.945 128.990 ;
        RECT 79.955 129.130 80.245 129.175 ;
        RECT 82.715 129.130 83.005 129.175 ;
        RECT 84.080 129.130 84.400 129.190 ;
        RECT 79.955 128.990 82.470 129.130 ;
        RECT 79.955 128.945 80.245 128.990 ;
        RECT 67.150 128.310 75.570 128.450 ;
        RECT 75.815 128.450 76.105 128.495 ;
        RECT 76.260 128.450 76.580 128.510 ;
        RECT 75.815 128.310 76.580 128.450 ;
        RECT 75.815 128.265 76.105 128.310 ;
        RECT 76.260 128.250 76.580 128.310 ;
        RECT 78.115 128.450 78.405 128.495 ;
        RECT 79.480 128.450 79.800 128.510 ;
        RECT 78.115 128.310 79.800 128.450 ;
        RECT 82.330 128.450 82.470 128.990 ;
        RECT 82.715 128.990 84.400 129.130 ;
        RECT 82.715 128.945 83.005 128.990 ;
        RECT 84.080 128.930 84.400 128.990 ;
        RECT 84.540 129.130 84.860 129.190 ;
        RECT 86.010 129.175 86.150 129.330 ;
        RECT 90.060 129.270 90.380 129.330 ;
        RECT 92.360 129.470 92.680 129.530 ;
        RECT 96.515 129.470 96.805 129.515 ;
        RECT 98.340 129.470 98.660 129.530 ;
        RECT 92.360 129.330 98.660 129.470 ;
        RECT 92.360 129.270 92.680 129.330 ;
        RECT 96.515 129.285 96.805 129.330 ;
        RECT 98.340 129.270 98.660 129.330 ;
        RECT 98.815 129.285 99.105 129.515 ;
        RECT 85.015 129.130 85.305 129.175 ;
        RECT 84.540 128.990 85.305 129.130 ;
        RECT 84.540 128.930 84.860 128.990 ;
        RECT 85.015 128.945 85.305 128.990 ;
        RECT 85.935 128.945 86.225 129.175 ;
        RECT 90.980 129.130 91.300 129.190 ;
        RECT 98.890 129.130 99.030 129.285 ;
        RECT 99.260 129.270 99.580 129.530 ;
        RECT 109.395 129.470 109.685 129.515 ;
        RECT 109.840 129.470 110.160 129.530 ;
        RECT 109.395 129.330 110.160 129.470 ;
        RECT 109.395 129.285 109.685 129.330 ;
        RECT 109.840 129.270 110.160 129.330 ;
        RECT 101.100 129.130 101.420 129.190 ;
        RECT 90.980 128.990 101.420 129.130 ;
        RECT 90.980 128.930 91.300 128.990 ;
        RECT 101.100 128.930 101.420 128.990 ;
        RECT 106.130 129.130 106.420 129.175 ;
        RECT 106.130 128.990 108.665 129.130 ;
        RECT 106.130 128.945 106.420 128.990 ;
        RECT 83.620 128.790 83.940 128.850 ;
        RECT 87.775 128.790 88.065 128.835 ;
        RECT 83.620 128.650 88.065 128.790 ;
        RECT 83.620 128.590 83.940 128.650 ;
        RECT 87.775 128.605 88.065 128.650 ;
        RECT 104.270 128.790 104.560 128.835 ;
        RECT 105.240 128.790 105.560 128.850 ;
        RECT 108.450 128.835 108.665 128.990 ;
        RECT 111.220 128.930 111.540 129.190 ;
        RECT 107.530 128.790 107.820 128.835 ;
        RECT 104.270 128.650 107.820 128.790 ;
        RECT 104.270 128.605 104.560 128.650 ;
        RECT 105.240 128.590 105.560 128.650 ;
        RECT 107.530 128.605 107.820 128.650 ;
        RECT 108.450 128.790 108.740 128.835 ;
        RECT 110.310 128.790 110.600 128.835 ;
        RECT 108.450 128.650 110.600 128.790 ;
        RECT 108.450 128.605 108.740 128.650 ;
        RECT 110.310 128.605 110.600 128.650 ;
        RECT 89.600 128.450 89.920 128.510 ;
        RECT 82.330 128.310 89.920 128.450 ;
        RECT 78.115 128.265 78.405 128.310 ;
        RECT 79.480 128.250 79.800 128.310 ;
        RECT 89.600 128.250 89.920 128.310 ;
        RECT 99.720 128.450 100.040 128.510 ;
        RECT 102.020 128.495 102.340 128.510 ;
        RECT 102.020 128.450 102.555 128.495 ;
        RECT 99.720 128.310 102.775 128.450 ;
        RECT 99.720 128.250 100.040 128.310 ;
        RECT 102.020 128.265 102.555 128.310 ;
        RECT 102.020 128.250 102.340 128.265 ;
        RECT 11.330 127.630 113.450 128.110 ;
        RECT 16.000 127.430 16.320 127.490 ;
        RECT 19.235 127.430 19.525 127.475 ;
        RECT 16.000 127.290 19.525 127.430 ;
        RECT 16.000 127.230 16.320 127.290 ;
        RECT 19.235 127.245 19.525 127.290 ;
        RECT 24.295 127.430 24.585 127.475 ;
        RECT 24.740 127.430 25.060 127.490 ;
        RECT 24.295 127.290 25.060 127.430 ;
        RECT 24.295 127.245 24.585 127.290 ;
        RECT 24.740 127.230 25.060 127.290 ;
        RECT 25.660 127.230 25.980 127.490 ;
        RECT 26.135 127.430 26.425 127.475 ;
        RECT 26.580 127.430 26.900 127.490 ;
        RECT 26.135 127.290 26.900 127.430 ;
        RECT 26.135 127.245 26.425 127.290 ;
        RECT 26.580 127.230 26.900 127.290 ;
        RECT 27.975 127.430 28.265 127.475 ;
        RECT 35.780 127.430 36.100 127.490 ;
        RECT 27.975 127.290 36.100 127.430 ;
        RECT 27.975 127.245 28.265 127.290 ;
        RECT 35.780 127.230 36.100 127.290 ;
        RECT 37.160 127.430 37.480 127.490 ;
        RECT 45.440 127.430 45.760 127.490 ;
        RECT 37.160 127.290 45.760 127.430 ;
        RECT 37.160 127.230 37.480 127.290 ;
        RECT 45.440 127.230 45.760 127.290 ;
        RECT 49.580 127.230 49.900 127.490 ;
        RECT 50.040 127.430 50.360 127.490 ;
        RECT 52.355 127.430 52.645 127.475 ;
        RECT 50.040 127.290 52.645 127.430 ;
        RECT 50.040 127.230 50.360 127.290 ;
        RECT 52.355 127.245 52.645 127.290 ;
        RECT 54.655 127.245 54.945 127.475 ;
        RECT 65.680 127.430 66.000 127.490 ;
        RECT 66.615 127.430 66.905 127.475 ;
        RECT 65.680 127.290 66.905 127.430 ;
        RECT 21.995 127.090 22.285 127.135 ;
        RECT 28.880 127.090 29.200 127.150 ;
        RECT 14.250 126.950 21.750 127.090 ;
        RECT 14.250 126.795 14.390 126.950 ;
        RECT 13.715 126.750 14.005 126.795 ;
        RECT 14.175 126.750 14.465 126.795 ;
        RECT 13.715 126.610 14.465 126.750 ;
        RECT 13.715 126.565 14.005 126.610 ;
        RECT 14.175 126.565 14.465 126.610 ;
        RECT 15.555 126.750 15.845 126.795 ;
        RECT 18.775 126.750 19.065 126.795 ;
        RECT 19.680 126.750 20.000 126.810 ;
        RECT 21.610 126.795 21.750 126.950 ;
        RECT 21.995 126.950 29.200 127.090 ;
        RECT 21.995 126.905 22.285 126.950 ;
        RECT 28.880 126.890 29.200 126.950 ;
        RECT 31.640 127.090 31.960 127.150 ;
        RECT 32.575 127.090 32.865 127.135 ;
        RECT 31.640 126.950 32.865 127.090 ;
        RECT 31.640 126.890 31.960 126.950 ;
        RECT 32.575 126.905 32.865 126.950 ;
        RECT 47.740 126.890 48.060 127.150 ;
        RECT 49.670 127.090 49.810 127.230 ;
        RECT 52.815 127.090 53.105 127.135 ;
        RECT 49.670 126.950 53.105 127.090 ;
        RECT 52.815 126.905 53.105 126.950 ;
        RECT 15.555 126.610 17.150 126.750 ;
        RECT 15.555 126.565 15.845 126.610 ;
        RECT 17.010 126.115 17.150 126.610 ;
        RECT 18.775 126.610 20.000 126.750 ;
        RECT 18.775 126.565 19.065 126.610 ;
        RECT 19.680 126.550 20.000 126.610 ;
        RECT 21.535 126.750 21.825 126.795 ;
        RECT 22.440 126.750 22.760 126.810 ;
        RECT 21.535 126.610 22.760 126.750 ;
        RECT 21.535 126.565 21.825 126.610 ;
        RECT 22.440 126.550 22.760 126.610 ;
        RECT 24.755 126.750 25.045 126.795 ;
        RECT 26.120 126.750 26.440 126.810 ;
        RECT 29.800 126.750 30.120 126.810 ;
        RECT 36.715 126.750 37.005 126.795 ;
        RECT 24.755 126.610 26.440 126.750 ;
        RECT 24.755 126.565 25.045 126.610 ;
        RECT 26.120 126.550 26.440 126.610 ;
        RECT 28.970 126.610 30.120 126.750 ;
        RECT 20.140 126.210 20.460 126.470 ;
        RECT 21.060 126.410 21.380 126.470 ;
        RECT 28.435 126.410 28.725 126.455 ;
        RECT 28.970 126.410 29.110 126.610 ;
        RECT 29.800 126.550 30.120 126.610 ;
        RECT 32.190 126.610 37.005 126.750 ;
        RECT 32.190 126.470 32.330 126.610 ;
        RECT 36.715 126.565 37.005 126.610 ;
        RECT 49.120 126.750 49.440 126.810 ;
        RECT 49.595 126.750 49.885 126.795 ;
        RECT 49.120 126.610 49.885 126.750 ;
        RECT 54.730 126.750 54.870 127.245 ;
        RECT 65.680 127.230 66.000 127.290 ;
        RECT 66.615 127.245 66.905 127.290 ;
        RECT 67.520 127.230 67.840 127.490 ;
        RECT 77.195 127.430 77.485 127.475 ;
        RECT 81.320 127.430 81.640 127.490 ;
        RECT 84.080 127.430 84.400 127.490 ;
        RECT 77.195 127.290 84.400 127.430 ;
        RECT 77.195 127.245 77.485 127.290 ;
        RECT 81.320 127.230 81.640 127.290 ;
        RECT 84.080 127.230 84.400 127.290 ;
        RECT 90.060 127.230 90.380 127.490 ;
        RECT 91.900 127.430 92.220 127.490 ;
        RECT 93.295 127.430 93.585 127.475 ;
        RECT 91.900 127.290 93.585 127.430 ;
        RECT 91.900 127.230 92.220 127.290 ;
        RECT 93.295 127.245 93.585 127.290 ;
        RECT 67.610 127.090 67.750 127.230 ;
        RECT 70.755 127.090 71.045 127.135 ;
        RECT 67.610 126.950 71.045 127.090 ;
        RECT 70.755 126.905 71.045 126.950 ;
        RECT 83.620 126.890 83.940 127.150 ;
        RECT 90.150 127.090 90.290 127.230 ;
        RECT 99.275 127.090 99.565 127.135 ;
        RECT 103.350 127.090 103.640 127.135 ;
        RECT 106.610 127.090 106.900 127.135 ;
        RECT 90.150 126.950 92.590 127.090 ;
        RECT 55.115 126.750 55.405 126.795 ;
        RECT 54.730 126.610 55.405 126.750 ;
        RECT 49.120 126.550 49.440 126.610 ;
        RECT 49.595 126.565 49.885 126.610 ;
        RECT 55.115 126.565 55.405 126.610 ;
        RECT 67.060 126.750 67.380 126.810 ;
        RECT 67.535 126.750 67.825 126.795 ;
        RECT 67.060 126.610 67.825 126.750 ;
        RECT 67.060 126.550 67.380 126.610 ;
        RECT 67.535 126.565 67.825 126.610 ;
        RECT 68.455 126.750 68.745 126.795 ;
        RECT 84.540 126.750 84.860 126.810 ;
        RECT 87.775 126.750 88.065 126.795 ;
        RECT 68.455 126.610 70.510 126.750 ;
        RECT 68.455 126.565 68.745 126.610 ;
        RECT 21.060 126.270 29.110 126.410 ;
        RECT 29.355 126.410 29.645 126.455 ;
        RECT 31.195 126.410 31.485 126.455 ;
        RECT 29.355 126.270 31.485 126.410 ;
        RECT 21.060 126.210 21.380 126.270 ;
        RECT 28.435 126.225 28.725 126.270 ;
        RECT 29.355 126.225 29.645 126.270 ;
        RECT 31.195 126.225 31.485 126.270 ;
        RECT 16.935 125.885 17.225 126.115 ;
        RECT 20.230 126.070 20.370 126.210 ;
        RECT 29.430 126.070 29.570 126.225 ;
        RECT 20.230 125.930 29.570 126.070 ;
        RECT 31.270 126.070 31.410 126.225 ;
        RECT 32.100 126.210 32.420 126.470 ;
        RECT 35.335 126.225 35.625 126.455 ;
        RECT 36.255 126.410 36.545 126.455 ;
        RECT 39.920 126.410 40.240 126.470 ;
        RECT 36.255 126.270 40.240 126.410 ;
        RECT 36.255 126.225 36.545 126.270 ;
        RECT 32.560 126.070 32.880 126.130 ;
        RECT 35.410 126.070 35.550 126.225 ;
        RECT 39.920 126.210 40.240 126.270 ;
        RECT 51.895 126.410 52.185 126.455 ;
        RECT 53.260 126.410 53.580 126.470 ;
        RECT 51.895 126.270 53.580 126.410 ;
        RECT 51.895 126.225 52.185 126.270 ;
        RECT 53.260 126.210 53.580 126.270 ;
        RECT 66.600 126.410 66.920 126.470 ;
        RECT 70.370 126.455 70.510 126.610 ;
        RECT 84.540 126.610 88.065 126.750 ;
        RECT 84.540 126.550 84.860 126.610 ;
        RECT 87.775 126.565 88.065 126.610 ;
        RECT 89.600 126.750 89.920 126.810 ;
        RECT 92.450 126.795 92.590 126.950 ;
        RECT 99.275 126.950 106.900 127.090 ;
        RECT 99.275 126.905 99.565 126.950 ;
        RECT 103.350 126.905 103.640 126.950 ;
        RECT 106.610 126.905 106.900 126.950 ;
        RECT 107.530 127.090 107.820 127.135 ;
        RECT 109.390 127.090 109.680 127.135 ;
        RECT 107.530 126.950 109.680 127.090 ;
        RECT 107.530 126.905 107.820 126.950 ;
        RECT 109.390 126.905 109.680 126.950 ;
        RECT 90.075 126.750 90.365 126.795 ;
        RECT 89.600 126.610 90.365 126.750 ;
        RECT 89.600 126.550 89.920 126.610 ;
        RECT 90.075 126.565 90.365 126.610 ;
        RECT 92.375 126.565 92.665 126.795 ;
        RECT 95.595 126.750 95.885 126.795 ;
        RECT 92.910 126.610 95.885 126.750 ;
        RECT 69.375 126.410 69.665 126.455 ;
        RECT 66.600 126.270 69.665 126.410 ;
        RECT 66.600 126.210 66.920 126.270 ;
        RECT 69.375 126.225 69.665 126.270 ;
        RECT 70.295 126.410 70.585 126.455 ;
        RECT 76.720 126.410 77.040 126.470 ;
        RECT 70.295 126.270 77.040 126.410 ;
        RECT 70.295 126.225 70.585 126.270 ;
        RECT 31.270 125.930 35.550 126.070 ;
        RECT 69.450 126.070 69.590 126.225 ;
        RECT 76.720 126.210 77.040 126.270 ;
        RECT 86.395 126.225 86.685 126.455 ;
        RECT 87.300 126.410 87.620 126.470 ;
        RECT 91.455 126.410 91.745 126.455 ;
        RECT 92.910 126.410 93.050 126.610 ;
        RECT 95.595 126.565 95.885 126.610 ;
        RECT 98.815 126.750 99.105 126.795 ;
        RECT 103.860 126.750 104.180 126.810 ;
        RECT 98.815 126.610 104.180 126.750 ;
        RECT 98.815 126.565 99.105 126.610 ;
        RECT 103.860 126.550 104.180 126.610 ;
        RECT 105.210 126.750 105.500 126.795 ;
        RECT 107.530 126.750 107.745 126.905 ;
        RECT 105.210 126.610 107.745 126.750 ;
        RECT 108.000 126.750 108.320 126.810 ;
        RECT 108.475 126.750 108.765 126.795 ;
        RECT 108.000 126.610 108.765 126.750 ;
        RECT 105.210 126.565 105.500 126.610 ;
        RECT 108.000 126.550 108.320 126.610 ;
        RECT 108.475 126.565 108.765 126.610 ;
        RECT 87.300 126.270 93.050 126.410 ;
        RECT 82.240 126.070 82.560 126.130 ;
        RECT 86.470 126.070 86.610 126.225 ;
        RECT 87.300 126.210 87.620 126.270 ;
        RECT 91.455 126.225 91.745 126.270 ;
        RECT 94.215 126.225 94.505 126.455 ;
        RECT 95.135 126.225 95.425 126.455 ;
        RECT 98.340 126.410 98.660 126.470 ;
        RECT 104.320 126.410 104.640 126.470 ;
        RECT 110.315 126.410 110.605 126.455 ;
        RECT 111.220 126.410 111.540 126.470 ;
        RECT 98.340 126.270 111.540 126.410 ;
        RECT 90.980 126.070 91.300 126.130 ;
        RECT 94.290 126.070 94.430 126.225 ;
        RECT 69.450 125.930 94.430 126.070 ;
        RECT 95.210 126.070 95.350 126.225 ;
        RECT 98.340 126.210 98.660 126.270 ;
        RECT 104.320 126.210 104.640 126.270 ;
        RECT 110.315 126.225 110.605 126.270 ;
        RECT 111.220 126.210 111.540 126.270 ;
        RECT 105.210 126.070 105.500 126.115 ;
        RECT 107.990 126.070 108.280 126.115 ;
        RECT 109.850 126.070 110.140 126.115 ;
        RECT 95.210 125.930 98.570 126.070 ;
        RECT 32.560 125.870 32.880 125.930 ;
        RECT 82.240 125.870 82.560 125.930 ;
        RECT 90.980 125.870 91.300 125.930 ;
        RECT 13.255 125.730 13.545 125.775 ;
        RECT 13.700 125.730 14.020 125.790 ;
        RECT 13.255 125.590 14.020 125.730 ;
        RECT 13.255 125.545 13.545 125.590 ;
        RECT 13.700 125.530 14.020 125.590 ;
        RECT 14.620 125.530 14.940 125.790 ;
        RECT 16.475 125.730 16.765 125.775 ;
        RECT 20.600 125.730 20.920 125.790 ;
        RECT 16.475 125.590 20.920 125.730 ;
        RECT 16.475 125.545 16.765 125.590 ;
        RECT 20.600 125.530 20.920 125.590 ;
        RECT 22.440 125.730 22.760 125.790 ;
        RECT 27.500 125.730 27.820 125.790 ;
        RECT 22.440 125.590 27.820 125.730 ;
        RECT 22.440 125.530 22.760 125.590 ;
        RECT 27.500 125.530 27.820 125.590 ;
        RECT 34.415 125.730 34.705 125.775 ;
        RECT 34.860 125.730 35.180 125.790 ;
        RECT 34.415 125.590 35.180 125.730 ;
        RECT 34.415 125.545 34.705 125.590 ;
        RECT 34.860 125.530 35.180 125.590 ;
        RECT 38.080 125.730 38.400 125.790 ;
        RECT 38.555 125.730 38.845 125.775 ;
        RECT 38.080 125.590 38.845 125.730 ;
        RECT 38.080 125.530 38.400 125.590 ;
        RECT 38.555 125.545 38.845 125.590 ;
        RECT 41.300 125.530 41.620 125.790 ;
        RECT 50.055 125.730 50.345 125.775 ;
        RECT 50.500 125.730 50.820 125.790 ;
        RECT 50.055 125.590 50.820 125.730 ;
        RECT 50.055 125.545 50.345 125.590 ;
        RECT 50.500 125.530 50.820 125.590 ;
        RECT 55.560 125.730 55.880 125.790 ;
        RECT 56.035 125.730 56.325 125.775 ;
        RECT 55.560 125.590 56.325 125.730 ;
        RECT 55.560 125.530 55.880 125.590 ;
        RECT 56.035 125.545 56.325 125.590 ;
        RECT 72.595 125.730 72.885 125.775 ;
        RECT 73.960 125.730 74.280 125.790 ;
        RECT 72.595 125.590 74.280 125.730 ;
        RECT 72.595 125.545 72.885 125.590 ;
        RECT 73.960 125.530 74.280 125.590 ;
        RECT 89.600 125.530 89.920 125.790 ;
        RECT 90.535 125.730 90.825 125.775 ;
        RECT 91.440 125.730 91.760 125.790 ;
        RECT 90.535 125.590 91.760 125.730 ;
        RECT 90.535 125.545 90.825 125.590 ;
        RECT 91.440 125.530 91.760 125.590 ;
        RECT 97.435 125.730 97.725 125.775 ;
        RECT 97.880 125.730 98.200 125.790 ;
        RECT 97.435 125.590 98.200 125.730 ;
        RECT 98.430 125.730 98.570 125.930 ;
        RECT 105.210 125.930 110.140 126.070 ;
        RECT 105.210 125.885 105.500 125.930 ;
        RECT 107.990 125.885 108.280 125.930 ;
        RECT 109.850 125.885 110.140 125.930 ;
        RECT 98.800 125.730 99.120 125.790 ;
        RECT 101.345 125.730 101.635 125.775 ;
        RECT 102.480 125.730 102.800 125.790 ;
        RECT 98.430 125.590 102.800 125.730 ;
        RECT 97.435 125.545 97.725 125.590 ;
        RECT 97.880 125.530 98.200 125.590 ;
        RECT 98.800 125.530 99.120 125.590 ;
        RECT 101.345 125.545 101.635 125.590 ;
        RECT 102.480 125.530 102.800 125.590 ;
        RECT 11.330 124.910 113.450 125.390 ;
        RECT 13.485 124.710 13.775 124.755 ;
        RECT 19.680 124.710 20.000 124.770 ;
        RECT 13.485 124.570 20.000 124.710 ;
        RECT 13.485 124.525 13.775 124.570 ;
        RECT 19.680 124.510 20.000 124.570 ;
        RECT 35.320 124.510 35.640 124.770 ;
        RECT 48.445 124.710 48.735 124.755 ;
        RECT 50.040 124.710 50.360 124.770 ;
        RECT 48.445 124.570 50.360 124.710 ;
        RECT 48.445 124.525 48.735 124.570 ;
        RECT 50.040 124.510 50.360 124.570 ;
        RECT 72.365 124.710 72.655 124.755 ;
        RECT 74.420 124.710 74.740 124.770 ;
        RECT 86.380 124.710 86.700 124.770 ;
        RECT 72.365 124.570 86.700 124.710 ;
        RECT 72.365 124.525 72.655 124.570 ;
        RECT 74.420 124.510 74.740 124.570 ;
        RECT 86.380 124.510 86.700 124.570 ;
        RECT 87.300 124.710 87.620 124.770 ;
        RECT 88.465 124.710 88.755 124.755 ;
        RECT 87.300 124.570 88.755 124.710 ;
        RECT 87.300 124.510 87.620 124.570 ;
        RECT 88.465 124.525 88.755 124.570 ;
        RECT 107.080 124.510 107.400 124.770 ;
        RECT 17.350 124.370 17.640 124.415 ;
        RECT 20.130 124.370 20.420 124.415 ;
        RECT 21.990 124.370 22.280 124.415 ;
        RECT 17.350 124.230 22.280 124.370 ;
        RECT 17.350 124.185 17.640 124.230 ;
        RECT 20.130 124.185 20.420 124.230 ;
        RECT 21.990 124.185 22.280 124.230 ;
        RECT 52.310 124.370 52.600 124.415 ;
        RECT 55.090 124.370 55.380 124.415 ;
        RECT 56.950 124.370 57.240 124.415 ;
        RECT 52.310 124.230 57.240 124.370 ;
        RECT 52.310 124.185 52.600 124.230 ;
        RECT 55.090 124.185 55.380 124.230 ;
        RECT 56.950 124.185 57.240 124.230 ;
        RECT 76.230 124.370 76.520 124.415 ;
        RECT 79.010 124.370 79.300 124.415 ;
        RECT 80.870 124.370 81.160 124.415 ;
        RECT 76.230 124.230 81.160 124.370 ;
        RECT 76.230 124.185 76.520 124.230 ;
        RECT 79.010 124.185 79.300 124.230 ;
        RECT 80.870 124.185 81.160 124.230 ;
        RECT 92.330 124.370 92.620 124.415 ;
        RECT 95.110 124.370 95.400 124.415 ;
        RECT 96.970 124.370 97.260 124.415 ;
        RECT 92.330 124.230 97.260 124.370 ;
        RECT 92.330 124.185 92.620 124.230 ;
        RECT 95.110 124.185 95.400 124.230 ;
        RECT 96.970 124.185 97.260 124.230 ;
        RECT 97.880 124.370 98.200 124.430 ;
        RECT 97.880 124.230 99.030 124.370 ;
        RECT 97.880 124.170 98.200 124.230 ;
        RECT 20.600 123.830 20.920 124.090 ;
        RECT 32.100 124.030 32.420 124.090 ;
        RECT 33.495 124.030 33.785 124.075 ;
        RECT 32.100 123.890 33.785 124.030 ;
        RECT 32.100 123.830 32.420 123.890 ;
        RECT 33.495 123.845 33.785 123.890 ;
        RECT 55.560 123.830 55.880 124.090 ;
        RECT 56.020 124.030 56.340 124.090 ;
        RECT 57.415 124.030 57.705 124.075 ;
        RECT 61.080 124.030 61.400 124.090 ;
        RECT 56.020 123.890 56.940 124.030 ;
        RECT 56.020 123.830 56.340 123.890 ;
        RECT 17.350 123.690 17.640 123.735 ;
        RECT 22.455 123.690 22.745 123.735 ;
        RECT 17.350 123.550 19.885 123.690 ;
        RECT 17.350 123.505 17.640 123.550 ;
        RECT 14.620 123.350 14.940 123.410 ;
        RECT 19.670 123.395 19.885 123.550 ;
        RECT 22.455 123.550 24.970 123.690 ;
        RECT 22.455 123.505 22.745 123.550 ;
        RECT 24.830 123.410 24.970 123.550 ;
        RECT 32.560 123.490 32.880 123.750 ;
        RECT 34.400 123.490 34.720 123.750 ;
        RECT 47.755 123.690 48.045 123.735 ;
        RECT 49.580 123.690 49.900 123.750 ;
        RECT 47.755 123.550 49.900 123.690 ;
        RECT 47.755 123.505 48.045 123.550 ;
        RECT 49.580 123.490 49.900 123.550 ;
        RECT 52.310 123.690 52.600 123.735 ;
        RECT 56.800 123.690 56.940 123.890 ;
        RECT 57.415 123.890 61.400 124.030 ;
        RECT 57.415 123.845 57.705 123.890 ;
        RECT 61.080 123.830 61.400 123.890 ;
        RECT 66.600 123.830 66.920 124.090 ;
        RECT 75.800 124.030 76.120 124.090 ;
        RECT 79.495 124.030 79.785 124.075 ;
        RECT 75.800 123.890 79.785 124.030 ;
        RECT 75.800 123.830 76.120 123.890 ;
        RECT 79.495 123.845 79.785 123.890 ;
        RECT 81.320 123.830 81.640 124.090 ;
        RECT 82.240 123.830 82.560 124.090 ;
        RECT 97.435 124.030 97.725 124.075 ;
        RECT 98.340 124.030 98.660 124.090 ;
        RECT 97.435 123.890 98.660 124.030 ;
        RECT 97.435 123.845 97.725 123.890 ;
        RECT 98.340 123.830 98.660 123.890 ;
        RECT 64.775 123.690 65.065 123.735 ;
        RECT 74.880 123.690 75.200 123.750 ;
        RECT 98.890 123.735 99.030 124.230 ;
        RECT 101.100 123.830 101.420 124.090 ;
        RECT 102.020 123.830 102.340 124.090 ;
        RECT 52.310 123.550 54.845 123.690 ;
        RECT 56.800 123.550 75.200 123.690 ;
        RECT 52.310 123.505 52.600 123.550 ;
        RECT 15.490 123.350 15.780 123.395 ;
        RECT 18.750 123.350 19.040 123.395 ;
        RECT 14.620 123.210 19.040 123.350 ;
        RECT 14.620 123.150 14.940 123.210 ;
        RECT 15.490 123.165 15.780 123.210 ;
        RECT 18.750 123.165 19.040 123.210 ;
        RECT 19.670 123.350 19.960 123.395 ;
        RECT 21.530 123.350 21.820 123.395 ;
        RECT 19.670 123.210 21.820 123.350 ;
        RECT 19.670 123.165 19.960 123.210 ;
        RECT 21.530 123.165 21.820 123.210 ;
        RECT 24.740 123.150 25.060 123.410 ;
        RECT 50.500 123.395 50.820 123.410 ;
        RECT 54.630 123.395 54.845 123.550 ;
        RECT 64.775 123.505 65.065 123.550 ;
        RECT 74.880 123.490 75.200 123.550 ;
        RECT 76.230 123.690 76.520 123.735 ;
        RECT 92.330 123.690 92.620 123.735 ;
        RECT 95.595 123.690 95.885 123.735 ;
        RECT 76.230 123.550 78.765 123.690 ;
        RECT 76.230 123.505 76.520 123.550 ;
        RECT 50.450 123.350 50.820 123.395 ;
        RECT 53.710 123.350 54.000 123.395 ;
        RECT 50.450 123.210 54.000 123.350 ;
        RECT 50.450 123.165 50.820 123.210 ;
        RECT 53.710 123.165 54.000 123.210 ;
        RECT 54.630 123.350 54.920 123.395 ;
        RECT 56.490 123.350 56.780 123.395 ;
        RECT 54.630 123.210 56.780 123.350 ;
        RECT 54.630 123.165 54.920 123.210 ;
        RECT 56.490 123.165 56.780 123.210 ;
        RECT 74.370 123.350 74.660 123.395 ;
        RECT 75.340 123.350 75.660 123.410 ;
        RECT 78.550 123.395 78.765 123.550 ;
        RECT 92.330 123.550 94.865 123.690 ;
        RECT 92.330 123.505 92.620 123.550 ;
        RECT 77.630 123.350 77.920 123.395 ;
        RECT 74.370 123.210 77.920 123.350 ;
        RECT 74.370 123.165 74.660 123.210 ;
        RECT 50.500 123.150 50.820 123.165 ;
        RECT 75.340 123.150 75.660 123.210 ;
        RECT 77.630 123.165 77.920 123.210 ;
        RECT 78.550 123.350 78.840 123.395 ;
        RECT 80.410 123.350 80.700 123.395 ;
        RECT 83.635 123.350 83.925 123.395 ;
        RECT 78.550 123.210 80.700 123.350 ;
        RECT 78.550 123.165 78.840 123.210 ;
        RECT 80.410 123.165 80.700 123.210 ;
        RECT 80.950 123.210 83.925 123.350 ;
        RECT 65.220 122.810 65.540 123.070 ;
        RECT 67.520 122.810 67.840 123.070 ;
        RECT 67.980 122.810 68.300 123.070 ;
        RECT 69.835 123.010 70.125 123.055 ;
        RECT 72.580 123.010 72.900 123.070 ;
        RECT 69.835 122.870 72.900 123.010 ;
        RECT 69.835 122.825 70.125 122.870 ;
        RECT 72.580 122.810 72.900 122.870 ;
        RECT 77.180 123.010 77.500 123.070 ;
        RECT 80.950 123.010 81.090 123.210 ;
        RECT 83.635 123.165 83.925 123.210 ;
        RECT 90.470 123.350 90.760 123.395 ;
        RECT 91.440 123.350 91.760 123.410 ;
        RECT 94.650 123.395 94.865 123.550 ;
        RECT 95.595 123.550 98.110 123.690 ;
        RECT 95.595 123.505 95.885 123.550 ;
        RECT 93.730 123.350 94.020 123.395 ;
        RECT 90.470 123.210 94.020 123.350 ;
        RECT 90.470 123.165 90.760 123.210 ;
        RECT 91.440 123.150 91.760 123.210 ;
        RECT 93.730 123.165 94.020 123.210 ;
        RECT 94.650 123.350 94.940 123.395 ;
        RECT 96.510 123.350 96.800 123.395 ;
        RECT 94.650 123.210 96.800 123.350 ;
        RECT 94.650 123.165 94.940 123.210 ;
        RECT 96.510 123.165 96.800 123.210 ;
        RECT 77.180 122.870 81.090 123.010 ;
        RECT 83.175 123.010 83.465 123.055 ;
        RECT 84.540 123.010 84.860 123.070 ;
        RECT 83.175 122.870 84.860 123.010 ;
        RECT 77.180 122.810 77.500 122.870 ;
        RECT 83.175 122.825 83.465 122.870 ;
        RECT 84.540 122.810 84.860 122.870 ;
        RECT 85.475 123.010 85.765 123.055 ;
        RECT 88.220 123.010 88.540 123.070 ;
        RECT 97.970 123.055 98.110 123.550 ;
        RECT 98.815 123.505 99.105 123.735 ;
        RECT 102.480 123.490 102.800 123.750 ;
        RECT 106.175 123.690 106.465 123.735 ;
        RECT 105.100 123.550 106.465 123.690 ;
        RECT 85.475 122.870 88.540 123.010 ;
        RECT 85.475 122.825 85.765 122.870 ;
        RECT 88.220 122.810 88.540 122.870 ;
        RECT 97.895 122.825 98.185 123.055 ;
        RECT 104.335 123.010 104.625 123.055 ;
        RECT 105.100 123.010 105.240 123.550 ;
        RECT 106.175 123.505 106.465 123.550 ;
        RECT 104.335 122.870 105.240 123.010 ;
        RECT 104.335 122.825 104.625 122.870 ;
        RECT 11.330 122.190 113.450 122.670 ;
        RECT 31.640 121.990 31.960 122.050 ;
        RECT 32.345 121.990 32.635 122.035 ;
        RECT 31.640 121.850 32.635 121.990 ;
        RECT 31.640 121.790 31.960 121.850 ;
        RECT 32.345 121.805 32.635 121.850 ;
        RECT 35.780 121.990 36.100 122.050 ;
        RECT 44.075 121.990 44.365 122.035 ;
        RECT 35.780 121.850 44.365 121.990 ;
        RECT 35.780 121.790 36.100 121.850 ;
        RECT 44.075 121.805 44.365 121.850 ;
        RECT 46.375 121.805 46.665 122.035 ;
        RECT 50.040 121.990 50.360 122.050 ;
        RECT 52.815 121.990 53.105 122.035 ;
        RECT 56.940 121.990 57.260 122.050 ;
        RECT 50.040 121.850 53.105 121.990 ;
        RECT 13.700 121.650 14.020 121.710 ;
        RECT 15.030 121.650 15.320 121.695 ;
        RECT 18.290 121.650 18.580 121.695 ;
        RECT 13.700 121.510 18.580 121.650 ;
        RECT 13.700 121.450 14.020 121.510 ;
        RECT 15.030 121.465 15.320 121.510 ;
        RECT 18.290 121.465 18.580 121.510 ;
        RECT 19.210 121.650 19.500 121.695 ;
        RECT 21.070 121.650 21.360 121.695 ;
        RECT 19.210 121.510 21.360 121.650 ;
        RECT 19.210 121.465 19.500 121.510 ;
        RECT 21.070 121.465 21.360 121.510 ;
        RECT 24.300 121.650 24.590 121.695 ;
        RECT 26.160 121.650 26.450 121.695 ;
        RECT 24.300 121.510 26.450 121.650 ;
        RECT 24.300 121.465 24.590 121.510 ;
        RECT 26.160 121.465 26.450 121.510 ;
        RECT 27.080 121.650 27.370 121.695 ;
        RECT 28.880 121.650 29.200 121.710 ;
        RECT 30.340 121.650 30.630 121.695 ;
        RECT 27.080 121.510 30.630 121.650 ;
        RECT 27.080 121.465 27.370 121.510 ;
        RECT 16.890 121.310 17.180 121.355 ;
        RECT 19.210 121.310 19.425 121.465 ;
        RECT 16.890 121.170 19.425 121.310 ;
        RECT 26.235 121.310 26.450 121.465 ;
        RECT 28.880 121.450 29.200 121.510 ;
        RECT 30.340 121.465 30.630 121.510 ;
        RECT 35.270 121.650 35.560 121.695 ;
        RECT 36.700 121.650 37.020 121.710 ;
        RECT 38.530 121.650 38.820 121.695 ;
        RECT 35.270 121.510 38.820 121.650 ;
        RECT 35.270 121.465 35.560 121.510 ;
        RECT 36.700 121.450 37.020 121.510 ;
        RECT 38.530 121.465 38.820 121.510 ;
        RECT 39.450 121.650 39.740 121.695 ;
        RECT 41.310 121.650 41.600 121.695 ;
        RECT 39.450 121.510 41.600 121.650 ;
        RECT 39.450 121.465 39.740 121.510 ;
        RECT 41.310 121.465 41.600 121.510 ;
        RECT 42.220 121.650 42.540 121.710 ;
        RECT 42.220 121.510 45.210 121.650 ;
        RECT 28.480 121.310 28.770 121.355 ;
        RECT 26.235 121.170 28.770 121.310 ;
        RECT 16.890 121.125 17.180 121.170 ;
        RECT 28.480 121.125 28.770 121.170 ;
        RECT 32.100 121.310 32.420 121.370 ;
        RECT 33.265 121.310 33.555 121.355 ;
        RECT 32.100 121.170 33.555 121.310 ;
        RECT 32.100 121.110 32.420 121.170 ;
        RECT 33.265 121.125 33.555 121.170 ;
        RECT 37.130 121.310 37.420 121.355 ;
        RECT 39.450 121.310 39.665 121.465 ;
        RECT 42.220 121.450 42.540 121.510 ;
        RECT 37.130 121.170 39.665 121.310 ;
        RECT 39.920 121.310 40.240 121.370 ;
        RECT 44.535 121.310 44.825 121.355 ;
        RECT 39.920 121.170 44.825 121.310 ;
        RECT 37.130 121.125 37.420 121.170 ;
        RECT 39.920 121.110 40.240 121.170 ;
        RECT 44.535 121.125 44.825 121.170 ;
        RECT 16.460 120.970 16.780 121.030 ;
        RECT 20.155 120.970 20.445 121.015 ;
        RECT 16.460 120.830 20.445 120.970 ;
        RECT 16.460 120.770 16.780 120.830 ;
        RECT 20.155 120.785 20.445 120.830 ;
        RECT 21.995 120.970 22.285 121.015 ;
        RECT 23.375 120.970 23.665 121.015 ;
        RECT 24.740 120.970 25.060 121.030 ;
        RECT 21.995 120.830 25.060 120.970 ;
        RECT 21.995 120.785 22.285 120.830 ;
        RECT 23.375 120.785 23.665 120.830 ;
        RECT 24.740 120.770 25.060 120.830 ;
        RECT 25.200 120.770 25.520 121.030 ;
        RECT 39.000 120.970 39.320 121.030 ;
        RECT 40.395 120.970 40.685 121.015 ;
        RECT 39.000 120.830 40.685 120.970 ;
        RECT 39.000 120.770 39.320 120.830 ;
        RECT 40.395 120.785 40.685 120.830 ;
        RECT 41.300 120.970 41.620 121.030 ;
        RECT 42.235 120.970 42.525 121.015 ;
        RECT 41.300 120.830 42.525 120.970 ;
        RECT 41.300 120.770 41.620 120.830 ;
        RECT 42.235 120.785 42.525 120.830 ;
        RECT 43.615 120.970 43.905 121.015 ;
        RECT 45.070 120.970 45.210 121.510 ;
        RECT 46.450 121.310 46.590 121.805 ;
        RECT 50.040 121.790 50.360 121.850 ;
        RECT 52.815 121.805 53.105 121.850 ;
        RECT 53.350 121.850 57.260 121.990 ;
        RECT 46.835 121.310 47.125 121.355 ;
        RECT 46.450 121.170 47.125 121.310 ;
        RECT 46.835 121.125 47.125 121.170 ;
        RECT 43.615 120.830 45.210 120.970 ;
        RECT 45.900 120.970 46.220 121.030 ;
        RECT 53.350 121.015 53.490 121.850 ;
        RECT 56.940 121.790 57.260 121.850 ;
        RECT 58.795 121.805 59.085 122.035 ;
        RECT 62.245 121.990 62.535 122.035 ;
        RECT 67.980 121.990 68.300 122.050 ;
        RECT 62.245 121.850 68.300 121.990 ;
        RECT 62.245 121.805 62.535 121.850 ;
        RECT 56.495 121.650 56.785 121.695 ;
        RECT 57.860 121.650 58.180 121.710 ;
        RECT 56.495 121.510 58.180 121.650 ;
        RECT 56.495 121.465 56.785 121.510 ;
        RECT 57.860 121.450 58.180 121.510 ;
        RECT 56.940 121.110 57.260 121.370 ;
        RECT 58.870 121.310 59.010 121.805 ;
        RECT 67.980 121.790 68.300 121.850 ;
        RECT 71.675 121.805 71.965 122.035 ;
        RECT 64.250 121.650 64.540 121.695 ;
        RECT 65.220 121.650 65.540 121.710 ;
        RECT 67.510 121.650 67.800 121.695 ;
        RECT 64.250 121.510 67.800 121.650 ;
        RECT 64.250 121.465 64.540 121.510 ;
        RECT 65.220 121.450 65.540 121.510 ;
        RECT 67.510 121.465 67.800 121.510 ;
        RECT 68.430 121.650 68.720 121.695 ;
        RECT 70.290 121.650 70.580 121.695 ;
        RECT 68.430 121.510 70.580 121.650 ;
        RECT 68.430 121.465 68.720 121.510 ;
        RECT 70.290 121.465 70.580 121.510 ;
        RECT 59.255 121.310 59.545 121.355 ;
        RECT 58.870 121.170 59.545 121.310 ;
        RECT 59.255 121.125 59.545 121.170 ;
        RECT 60.635 121.125 60.925 121.355 ;
        RECT 66.110 121.310 66.400 121.355 ;
        RECT 68.430 121.310 68.645 121.465 ;
        RECT 66.110 121.170 68.645 121.310 ;
        RECT 69.375 121.310 69.665 121.355 ;
        RECT 71.750 121.310 71.890 121.805 ;
        RECT 75.340 121.790 75.660 122.050 ;
        RECT 86.380 121.990 86.700 122.050 ;
        RECT 92.835 121.990 93.125 122.035 ;
        RECT 77.270 121.850 85.230 121.990 ;
        RECT 69.375 121.170 71.890 121.310 ;
        RECT 66.110 121.125 66.400 121.170 ;
        RECT 69.375 121.125 69.665 121.170 ;
        RECT 53.275 120.970 53.565 121.015 ;
        RECT 45.900 120.830 53.565 120.970 ;
        RECT 43.615 120.785 43.905 120.830 ;
        RECT 16.890 120.630 17.180 120.675 ;
        RECT 19.670 120.630 19.960 120.675 ;
        RECT 21.530 120.630 21.820 120.675 ;
        RECT 16.890 120.490 21.820 120.630 ;
        RECT 16.890 120.445 17.180 120.490 ;
        RECT 19.670 120.445 19.960 120.490 ;
        RECT 21.530 120.445 21.820 120.490 ;
        RECT 23.840 120.630 24.130 120.675 ;
        RECT 25.700 120.630 25.990 120.675 ;
        RECT 28.480 120.630 28.770 120.675 ;
        RECT 23.840 120.490 28.770 120.630 ;
        RECT 23.840 120.445 24.130 120.490 ;
        RECT 25.700 120.445 25.990 120.490 ;
        RECT 28.480 120.445 28.770 120.490 ;
        RECT 37.130 120.630 37.420 120.675 ;
        RECT 39.910 120.630 40.200 120.675 ;
        RECT 41.770 120.630 42.060 120.675 ;
        RECT 37.130 120.490 42.060 120.630 ;
        RECT 42.310 120.630 42.450 120.785 ;
        RECT 45.900 120.770 46.220 120.830 ;
        RECT 53.275 120.785 53.565 120.830 ;
        RECT 53.720 120.970 54.040 121.030 ;
        RECT 55.575 120.970 55.865 121.015 ;
        RECT 53.720 120.830 55.865 120.970 ;
        RECT 53.720 120.770 54.040 120.830 ;
        RECT 55.575 120.785 55.865 120.830 ;
        RECT 56.480 120.970 56.800 121.030 ;
        RECT 60.710 120.970 60.850 121.125 ;
        RECT 72.580 121.110 72.900 121.370 ;
        RECT 73.960 121.110 74.280 121.370 ;
        RECT 74.880 121.310 75.200 121.370 ;
        RECT 77.270 121.310 77.410 121.850 ;
        RECT 78.510 121.650 78.800 121.695 ;
        RECT 79.480 121.650 79.800 121.710 ;
        RECT 81.770 121.650 82.060 121.695 ;
        RECT 78.510 121.510 82.060 121.650 ;
        RECT 78.510 121.465 78.800 121.510 ;
        RECT 79.480 121.450 79.800 121.510 ;
        RECT 81.770 121.465 82.060 121.510 ;
        RECT 82.690 121.650 82.980 121.695 ;
        RECT 84.550 121.650 84.840 121.695 ;
        RECT 82.690 121.510 84.840 121.650 ;
        RECT 85.090 121.650 85.230 121.850 ;
        RECT 86.380 121.850 93.125 121.990 ;
        RECT 86.380 121.790 86.700 121.850 ;
        RECT 92.835 121.805 93.125 121.850 ;
        RECT 97.895 121.990 98.185 122.035 ;
        RECT 99.260 121.990 99.580 122.050 ;
        RECT 100.885 121.990 101.175 122.035 ;
        RECT 97.895 121.850 101.175 121.990 ;
        RECT 97.895 121.805 98.185 121.850 ;
        RECT 99.260 121.790 99.580 121.850 ;
        RECT 100.885 121.805 101.175 121.850 ;
        RECT 91.900 121.650 92.220 121.710 ;
        RECT 93.295 121.650 93.585 121.695 ;
        RECT 97.435 121.650 97.725 121.695 ;
        RECT 85.090 121.510 86.510 121.650 ;
        RECT 82.690 121.465 82.980 121.510 ;
        RECT 84.550 121.465 84.840 121.510 ;
        RECT 74.880 121.170 77.410 121.310 ;
        RECT 80.370 121.310 80.660 121.355 ;
        RECT 82.690 121.310 82.905 121.465 ;
        RECT 80.370 121.170 82.905 121.310 ;
        RECT 74.880 121.110 75.200 121.170 ;
        RECT 80.370 121.125 80.660 121.170 ;
        RECT 83.620 121.110 83.940 121.370 ;
        RECT 85.935 121.310 86.225 121.355 ;
        RECT 86.370 121.310 86.510 121.510 ;
        RECT 91.900 121.510 97.725 121.650 ;
        RECT 91.900 121.450 92.220 121.510 ;
        RECT 93.295 121.465 93.585 121.510 ;
        RECT 97.435 121.465 97.725 121.510 ;
        RECT 102.890 121.650 103.180 121.695 ;
        RECT 103.860 121.650 104.180 121.710 ;
        RECT 106.150 121.650 106.440 121.695 ;
        RECT 102.890 121.510 106.440 121.650 ;
        RECT 102.890 121.465 103.180 121.510 ;
        RECT 103.860 121.450 104.180 121.510 ;
        RECT 106.150 121.465 106.440 121.510 ;
        RECT 107.070 121.650 107.360 121.695 ;
        RECT 108.930 121.650 109.220 121.695 ;
        RECT 107.070 121.510 109.220 121.650 ;
        RECT 107.070 121.465 107.360 121.510 ;
        RECT 108.930 121.465 109.220 121.510 ;
        RECT 85.935 121.170 86.510 121.310 ;
        RECT 85.935 121.125 86.225 121.170 ;
        RECT 88.220 121.110 88.540 121.370 ;
        RECT 89.600 121.110 89.920 121.370 ;
        RECT 90.060 121.110 90.380 121.370 ;
        RECT 104.750 121.310 105.040 121.355 ;
        RECT 107.070 121.310 107.285 121.465 ;
        RECT 104.750 121.170 107.285 121.310 ;
        RECT 107.540 121.310 107.860 121.370 ;
        RECT 108.015 121.310 108.305 121.355 ;
        RECT 107.540 121.170 108.305 121.310 ;
        RECT 104.750 121.125 105.040 121.170 ;
        RECT 107.540 121.110 107.860 121.170 ;
        RECT 108.015 121.125 108.305 121.170 ;
        RECT 56.480 120.830 60.850 120.970 ;
        RECT 71.215 120.970 71.505 121.015 ;
        RECT 76.720 120.970 77.040 121.030 ;
        RECT 81.320 120.970 81.640 121.030 ;
        RECT 85.475 120.970 85.765 121.015 ;
        RECT 71.215 120.830 85.765 120.970 ;
        RECT 56.480 120.770 56.800 120.830 ;
        RECT 71.215 120.785 71.505 120.830 ;
        RECT 76.720 120.770 77.040 120.830 ;
        RECT 81.320 120.770 81.640 120.830 ;
        RECT 85.475 120.785 85.765 120.830 ;
        RECT 90.980 120.970 91.300 121.030 ;
        RECT 91.915 120.970 92.205 121.015 ;
        RECT 96.515 120.970 96.805 121.015 ;
        RECT 90.980 120.830 96.805 120.970 ;
        RECT 90.980 120.770 91.300 120.830 ;
        RECT 91.915 120.785 92.205 120.830 ;
        RECT 96.515 120.785 96.805 120.830 ;
        RECT 104.320 120.970 104.640 121.030 ;
        RECT 109.855 120.970 110.145 121.015 ;
        RECT 104.320 120.830 110.145 120.970 ;
        RECT 104.320 120.770 104.640 120.830 ;
        RECT 109.855 120.785 110.145 120.830 ;
        RECT 49.580 120.630 49.900 120.690 ;
        RECT 42.310 120.490 49.900 120.630 ;
        RECT 37.130 120.445 37.420 120.490 ;
        RECT 39.910 120.445 40.200 120.490 ;
        RECT 41.770 120.445 42.060 120.490 ;
        RECT 49.580 120.430 49.900 120.490 ;
        RECT 66.110 120.630 66.400 120.675 ;
        RECT 68.890 120.630 69.180 120.675 ;
        RECT 70.750 120.630 71.040 120.675 ;
        RECT 66.110 120.490 71.040 120.630 ;
        RECT 66.110 120.445 66.400 120.490 ;
        RECT 68.890 120.445 69.180 120.490 ;
        RECT 70.750 120.445 71.040 120.490 ;
        RECT 80.370 120.630 80.660 120.675 ;
        RECT 83.150 120.630 83.440 120.675 ;
        RECT 85.010 120.630 85.300 120.675 ;
        RECT 80.370 120.490 85.300 120.630 ;
        RECT 80.370 120.445 80.660 120.490 ;
        RECT 83.150 120.445 83.440 120.490 ;
        RECT 85.010 120.445 85.300 120.490 ;
        RECT 87.300 120.430 87.620 120.690 ;
        RECT 104.750 120.630 105.040 120.675 ;
        RECT 107.530 120.630 107.820 120.675 ;
        RECT 109.390 120.630 109.680 120.675 ;
        RECT 104.750 120.490 109.680 120.630 ;
        RECT 104.750 120.445 105.040 120.490 ;
        RECT 107.530 120.445 107.820 120.490 ;
        RECT 109.390 120.445 109.680 120.490 ;
        RECT 13.025 120.290 13.315 120.335 ;
        RECT 21.060 120.290 21.380 120.350 ;
        RECT 13.025 120.150 21.380 120.290 ;
        RECT 13.025 120.105 13.315 120.150 ;
        RECT 21.060 120.090 21.380 120.150 ;
        RECT 46.820 120.290 47.140 120.350 ;
        RECT 47.755 120.290 48.045 120.335 ;
        RECT 46.820 120.150 48.045 120.290 ;
        RECT 46.820 120.090 47.140 120.150 ;
        RECT 47.755 120.105 48.045 120.150 ;
        RECT 50.975 120.290 51.265 120.335 ;
        RECT 51.420 120.290 51.740 120.350 ;
        RECT 50.975 120.150 51.740 120.290 ;
        RECT 50.975 120.105 51.265 120.150 ;
        RECT 51.420 120.090 51.740 120.150 ;
        RECT 59.240 120.290 59.560 120.350 ;
        RECT 60.175 120.290 60.465 120.335 ;
        RECT 59.240 120.150 60.465 120.290 ;
        RECT 59.240 120.090 59.560 120.150 ;
        RECT 60.175 120.105 60.465 120.150 ;
        RECT 61.095 120.290 61.385 120.335 ;
        RECT 67.060 120.290 67.380 120.350 ;
        RECT 61.095 120.150 67.380 120.290 ;
        RECT 61.095 120.105 61.385 120.150 ;
        RECT 67.060 120.090 67.380 120.150 ;
        RECT 72.120 120.290 72.440 120.350 ;
        RECT 73.055 120.290 73.345 120.335 ;
        RECT 72.120 120.150 73.345 120.290 ;
        RECT 72.120 120.090 72.440 120.150 ;
        RECT 73.055 120.105 73.345 120.150 ;
        RECT 76.505 120.290 76.795 120.335 ;
        RECT 77.180 120.290 77.500 120.350 ;
        RECT 76.505 120.150 77.500 120.290 ;
        RECT 76.505 120.105 76.795 120.150 ;
        RECT 77.180 120.090 77.500 120.150 ;
        RECT 84.080 120.290 84.400 120.350 ;
        RECT 86.395 120.290 86.685 120.335 ;
        RECT 84.080 120.150 86.685 120.290 ;
        RECT 84.080 120.090 84.400 120.150 ;
        RECT 86.395 120.105 86.685 120.150 ;
        RECT 88.680 120.090 89.000 120.350 ;
        RECT 90.520 120.090 90.840 120.350 ;
        RECT 95.135 120.290 95.425 120.335 ;
        RECT 96.040 120.290 96.360 120.350 ;
        RECT 95.135 120.150 96.360 120.290 ;
        RECT 95.135 120.105 95.425 120.150 ;
        RECT 96.040 120.090 96.360 120.150 ;
        RECT 99.720 120.090 100.040 120.350 ;
        RECT 11.330 119.470 113.450 119.950 ;
        RECT 32.345 119.270 32.635 119.315 ;
        RECT 35.780 119.270 36.100 119.330 ;
        RECT 32.345 119.130 36.100 119.270 ;
        RECT 32.345 119.085 32.635 119.130 ;
        RECT 35.780 119.070 36.100 119.130 ;
        RECT 39.000 119.070 39.320 119.330 ;
        RECT 65.005 119.270 65.295 119.315 ;
        RECT 67.520 119.270 67.840 119.330 ;
        RECT 65.005 119.130 67.840 119.270 ;
        RECT 65.005 119.085 65.295 119.130 ;
        RECT 67.520 119.070 67.840 119.130 ;
        RECT 75.800 119.270 76.120 119.330 ;
        RECT 77.195 119.270 77.485 119.315 ;
        RECT 75.800 119.130 77.485 119.270 ;
        RECT 75.800 119.070 76.120 119.130 ;
        RECT 77.195 119.085 77.485 119.130 ;
        RECT 84.540 119.270 84.860 119.330 ;
        RECT 86.625 119.270 86.915 119.315 ;
        RECT 84.540 119.130 86.915 119.270 ;
        RECT 84.540 119.070 84.860 119.130 ;
        RECT 86.625 119.085 86.915 119.130 ;
        RECT 91.225 119.270 91.515 119.315 ;
        RECT 91.900 119.270 92.220 119.330 ;
        RECT 91.225 119.130 92.220 119.270 ;
        RECT 91.225 119.085 91.515 119.130 ;
        RECT 91.900 119.070 92.220 119.130 ;
        RECT 103.860 119.270 104.180 119.330 ;
        RECT 104.335 119.270 104.625 119.315 ;
        RECT 103.860 119.130 104.625 119.270 ;
        RECT 103.860 119.070 104.180 119.130 ;
        RECT 104.335 119.085 104.625 119.130 ;
        RECT 106.175 119.270 106.465 119.315 ;
        RECT 107.080 119.270 107.400 119.330 ;
        RECT 106.175 119.130 107.400 119.270 ;
        RECT 106.175 119.085 106.465 119.130 ;
        RECT 107.080 119.070 107.400 119.130 ;
        RECT 17.035 118.930 17.325 118.975 ;
        RECT 20.155 118.930 20.445 118.975 ;
        RECT 22.045 118.930 22.335 118.975 ;
        RECT 17.035 118.790 22.335 118.930 ;
        RECT 17.035 118.745 17.325 118.790 ;
        RECT 20.155 118.745 20.445 118.790 ;
        RECT 22.045 118.745 22.335 118.790 ;
        RECT 23.840 118.930 24.130 118.975 ;
        RECT 25.700 118.930 25.990 118.975 ;
        RECT 28.480 118.930 28.770 118.975 ;
        RECT 23.840 118.790 28.770 118.930 ;
        RECT 23.840 118.745 24.130 118.790 ;
        RECT 25.700 118.745 25.990 118.790 ;
        RECT 28.480 118.745 28.770 118.790 ;
        RECT 43.570 118.930 43.860 118.975 ;
        RECT 46.350 118.930 46.640 118.975 ;
        RECT 48.210 118.930 48.500 118.975 ;
        RECT 43.570 118.790 48.500 118.930 ;
        RECT 43.570 118.745 43.860 118.790 ;
        RECT 46.350 118.745 46.640 118.790 ;
        RECT 48.210 118.745 48.500 118.790 ;
        RECT 55.990 118.930 56.280 118.975 ;
        RECT 58.770 118.930 59.060 118.975 ;
        RECT 60.630 118.930 60.920 118.975 ;
        RECT 55.990 118.790 60.920 118.930 ;
        RECT 55.990 118.745 56.280 118.790 ;
        RECT 58.770 118.745 59.060 118.790 ;
        RECT 60.630 118.745 60.920 118.790 ;
        RECT 68.870 118.930 69.160 118.975 ;
        RECT 71.650 118.930 71.940 118.975 ;
        RECT 73.510 118.930 73.800 118.975 ;
        RECT 68.870 118.790 73.800 118.930 ;
        RECT 68.870 118.745 69.160 118.790 ;
        RECT 71.650 118.745 71.940 118.790 ;
        RECT 73.510 118.745 73.800 118.790 ;
        RECT 78.120 118.930 78.410 118.975 ;
        RECT 79.980 118.930 80.270 118.975 ;
        RECT 82.760 118.930 83.050 118.975 ;
        RECT 78.120 118.790 83.050 118.930 ;
        RECT 78.120 118.745 78.410 118.790 ;
        RECT 79.980 118.745 80.270 118.790 ;
        RECT 82.760 118.745 83.050 118.790 ;
        RECT 95.090 118.930 95.380 118.975 ;
        RECT 97.870 118.930 98.160 118.975 ;
        RECT 99.730 118.930 100.020 118.975 ;
        RECT 95.090 118.790 100.020 118.930 ;
        RECT 95.090 118.745 95.380 118.790 ;
        RECT 97.870 118.745 98.160 118.790 ;
        RECT 99.730 118.745 100.020 118.790 ;
        RECT 21.520 118.390 21.840 118.650 ;
        RECT 46.820 118.390 47.140 118.650 ;
        RECT 57.860 118.590 58.180 118.650 ;
        RECT 55.650 118.450 58.180 118.590 ;
        RECT 9.560 117.910 9.880 117.970 ;
        RECT 12.795 117.910 13.085 117.955 ;
        RECT 9.560 117.770 13.085 117.910 ;
        RECT 9.560 117.710 9.880 117.770 ;
        RECT 12.795 117.725 13.085 117.770 ;
        RECT 13.700 117.910 14.020 117.970 ;
        RECT 15.955 117.955 16.245 118.270 ;
        RECT 17.035 118.250 17.325 118.295 ;
        RECT 20.615 118.250 20.905 118.295 ;
        RECT 22.450 118.250 22.740 118.295 ;
        RECT 17.035 118.110 22.740 118.250 ;
        RECT 17.035 118.065 17.325 118.110 ;
        RECT 20.615 118.065 20.905 118.110 ;
        RECT 22.450 118.065 22.740 118.110 ;
        RECT 22.915 118.250 23.205 118.295 ;
        RECT 23.375 118.250 23.665 118.295 ;
        RECT 24.740 118.250 25.060 118.310 ;
        RECT 22.915 118.110 25.060 118.250 ;
        RECT 22.915 118.065 23.205 118.110 ;
        RECT 23.375 118.065 23.665 118.110 ;
        RECT 24.740 118.050 25.060 118.110 ;
        RECT 25.215 118.250 25.505 118.295 ;
        RECT 25.660 118.250 25.980 118.310 ;
        RECT 28.480 118.250 28.770 118.295 ;
        RECT 25.215 118.110 25.980 118.250 ;
        RECT 25.215 118.065 25.505 118.110 ;
        RECT 25.660 118.050 25.980 118.110 ;
        RECT 26.235 118.110 28.770 118.250 ;
        RECT 26.235 117.955 26.450 118.110 ;
        RECT 28.480 118.065 28.770 118.110 ;
        RECT 34.860 118.050 35.180 118.310 ;
        RECT 38.080 118.050 38.400 118.310 ;
        RECT 39.920 118.295 40.240 118.310 ;
        RECT 39.705 118.065 40.240 118.295 ;
        RECT 43.570 118.250 43.860 118.295 ;
        RECT 48.675 118.250 48.965 118.295 ;
        RECT 49.580 118.250 49.900 118.310 ;
        RECT 43.570 118.110 46.105 118.250 ;
        RECT 43.570 118.065 43.860 118.110 ;
        RECT 39.920 118.050 40.240 118.065 ;
        RECT 15.655 117.910 16.245 117.955 ;
        RECT 18.895 117.910 19.545 117.955 ;
        RECT 13.700 117.770 19.545 117.910 ;
        RECT 13.700 117.710 14.020 117.770 ;
        RECT 15.655 117.725 15.945 117.770 ;
        RECT 18.895 117.725 19.545 117.770 ;
        RECT 24.300 117.910 24.590 117.955 ;
        RECT 26.160 117.910 26.450 117.955 ;
        RECT 24.300 117.770 26.450 117.910 ;
        RECT 24.300 117.725 24.590 117.770 ;
        RECT 26.160 117.725 26.450 117.770 ;
        RECT 27.040 117.955 27.360 117.970 ;
        RECT 27.040 117.910 27.370 117.955 ;
        RECT 30.340 117.910 30.630 117.955 ;
        RECT 27.040 117.770 30.630 117.910 ;
        RECT 27.040 117.725 27.370 117.770 ;
        RECT 30.340 117.725 30.630 117.770 ;
        RECT 41.710 117.910 42.000 117.955 ;
        RECT 44.060 117.910 44.380 117.970 ;
        RECT 45.890 117.955 46.105 118.110 ;
        RECT 48.675 118.110 49.900 118.250 ;
        RECT 48.675 118.065 48.965 118.110 ;
        RECT 49.580 118.050 49.900 118.110 ;
        RECT 51.420 118.050 51.740 118.310 ;
        RECT 52.125 118.250 52.415 118.295 ;
        RECT 55.650 118.250 55.790 118.450 ;
        RECT 57.860 118.390 58.180 118.450 ;
        RECT 59.240 118.390 59.560 118.650 ;
        RECT 61.080 118.390 61.400 118.650 ;
        RECT 72.120 118.390 72.440 118.650 ;
        RECT 73.040 118.590 73.360 118.650 ;
        RECT 73.975 118.590 74.265 118.635 ;
        RECT 76.720 118.590 77.040 118.650 ;
        RECT 77.655 118.590 77.945 118.635 ;
        RECT 73.040 118.450 77.945 118.590 ;
        RECT 73.040 118.390 73.360 118.450 ;
        RECT 73.975 118.405 74.265 118.450 ;
        RECT 76.720 118.390 77.040 118.450 ;
        RECT 77.655 118.405 77.945 118.450 ;
        RECT 79.495 118.590 79.785 118.635 ;
        RECT 88.680 118.590 89.000 118.650 ;
        RECT 101.560 118.590 101.880 118.650 ;
        RECT 104.320 118.590 104.640 118.650 ;
        RECT 79.495 118.450 89.000 118.590 ;
        RECT 79.495 118.405 79.785 118.450 ;
        RECT 88.680 118.390 89.000 118.450 ;
        RECT 100.270 118.450 104.640 118.590 ;
        RECT 52.125 118.110 55.790 118.250 ;
        RECT 55.990 118.250 56.280 118.295 ;
        RECT 60.620 118.250 60.940 118.310 ;
        RECT 62.935 118.250 63.225 118.295 ;
        RECT 68.870 118.250 69.160 118.295 ;
        RECT 55.990 118.110 58.525 118.250 ;
        RECT 52.125 118.065 52.415 118.110 ;
        RECT 55.990 118.065 56.280 118.110 ;
        RECT 58.310 117.955 58.525 118.110 ;
        RECT 60.620 118.110 63.610 118.250 ;
        RECT 60.620 118.050 60.940 118.110 ;
        RECT 62.935 118.065 63.225 118.110 ;
        RECT 44.970 117.910 45.260 117.955 ;
        RECT 41.710 117.770 45.260 117.910 ;
        RECT 41.710 117.725 42.000 117.770 ;
        RECT 27.040 117.710 27.360 117.725 ;
        RECT 44.060 117.710 44.380 117.770 ;
        RECT 44.970 117.725 45.260 117.770 ;
        RECT 45.890 117.910 46.180 117.955 ;
        RECT 47.750 117.910 48.040 117.955 ;
        RECT 45.890 117.770 48.040 117.910 ;
        RECT 45.890 117.725 46.180 117.770 ;
        RECT 47.750 117.725 48.040 117.770 ;
        RECT 54.130 117.910 54.420 117.955 ;
        RECT 57.390 117.910 57.680 117.955 ;
        RECT 58.310 117.910 58.600 117.955 ;
        RECT 60.170 117.910 60.460 117.955 ;
        RECT 54.130 117.770 58.090 117.910 ;
        RECT 54.130 117.725 54.420 117.770 ;
        RECT 57.390 117.725 57.680 117.770 ;
        RECT 25.200 117.570 25.520 117.630 ;
        RECT 33.955 117.570 34.245 117.615 ;
        RECT 25.200 117.430 34.245 117.570 ;
        RECT 25.200 117.370 25.520 117.430 ;
        RECT 33.955 117.385 34.245 117.430 ;
        RECT 50.500 117.370 50.820 117.630 ;
        RECT 57.950 117.570 58.090 117.770 ;
        RECT 58.310 117.770 60.460 117.910 ;
        RECT 58.310 117.725 58.600 117.770 ;
        RECT 60.170 117.725 60.460 117.770 ;
        RECT 62.475 117.570 62.765 117.615 ;
        RECT 57.950 117.430 62.765 117.570 ;
        RECT 63.470 117.570 63.610 118.110 ;
        RECT 68.870 118.110 71.405 118.250 ;
        RECT 68.870 118.065 69.160 118.110 ;
        RECT 67.060 117.955 67.380 117.970 ;
        RECT 71.190 117.955 71.405 118.110 ;
        RECT 76.260 118.050 76.580 118.310 ;
        RECT 82.760 118.250 83.050 118.295 ;
        RECT 80.515 118.110 83.050 118.250 ;
        RECT 80.515 117.955 80.730 118.110 ;
        RECT 82.760 118.065 83.050 118.110 ;
        RECT 95.090 118.250 95.380 118.295 ;
        RECT 95.090 118.110 97.625 118.250 ;
        RECT 95.090 118.065 95.380 118.110 ;
        RECT 67.010 117.910 67.380 117.955 ;
        RECT 70.270 117.910 70.560 117.955 ;
        RECT 67.010 117.770 70.560 117.910 ;
        RECT 67.010 117.725 67.380 117.770 ;
        RECT 70.270 117.725 70.560 117.770 ;
        RECT 71.190 117.910 71.480 117.955 ;
        RECT 73.050 117.910 73.340 117.955 ;
        RECT 71.190 117.770 73.340 117.910 ;
        RECT 71.190 117.725 71.480 117.770 ;
        RECT 73.050 117.725 73.340 117.770 ;
        RECT 78.580 117.910 78.870 117.955 ;
        RECT 80.440 117.910 80.730 117.955 ;
        RECT 78.580 117.770 80.730 117.910 ;
        RECT 78.580 117.725 78.870 117.770 ;
        RECT 80.440 117.725 80.730 117.770 ;
        RECT 81.360 117.910 81.650 117.955 ;
        RECT 84.080 117.910 84.400 117.970 ;
        RECT 84.620 117.910 84.910 117.955 ;
        RECT 81.360 117.770 84.910 117.910 ;
        RECT 81.360 117.725 81.650 117.770 ;
        RECT 67.060 117.710 67.380 117.725 ;
        RECT 84.080 117.710 84.400 117.770 ;
        RECT 84.620 117.725 84.910 117.770 ;
        RECT 90.520 117.910 90.840 117.970 ;
        RECT 97.410 117.955 97.625 118.110 ;
        RECT 98.340 118.050 98.660 118.310 ;
        RECT 100.270 118.295 100.410 118.450 ;
        RECT 101.560 118.390 101.880 118.450 ;
        RECT 104.320 118.390 104.640 118.450 ;
        RECT 100.195 118.065 100.485 118.295 ;
        RECT 103.400 118.250 103.720 118.310 ;
        RECT 103.875 118.250 104.165 118.295 ;
        RECT 105.215 118.260 105.505 118.295 ;
        RECT 103.400 118.110 104.165 118.250 ;
        RECT 103.400 118.050 103.720 118.110 ;
        RECT 103.875 118.065 104.165 118.110 ;
        RECT 104.870 118.120 105.505 118.260 ;
        RECT 93.230 117.910 93.520 117.955 ;
        RECT 96.490 117.910 96.780 117.955 ;
        RECT 90.520 117.770 96.780 117.910 ;
        RECT 90.520 117.710 90.840 117.770 ;
        RECT 93.230 117.725 93.520 117.770 ;
        RECT 96.490 117.725 96.780 117.770 ;
        RECT 97.410 117.910 97.700 117.955 ;
        RECT 99.270 117.910 99.560 117.955 ;
        RECT 97.410 117.770 99.560 117.910 ;
        RECT 97.410 117.725 97.700 117.770 ;
        RECT 99.270 117.725 99.560 117.770 ;
        RECT 99.720 117.910 100.040 117.970 ;
        RECT 104.870 117.910 105.010 118.120 ;
        RECT 105.215 118.065 105.505 118.120 ;
        RECT 99.720 117.770 105.010 117.910 ;
        RECT 99.720 117.710 100.040 117.770 ;
        RECT 70.740 117.570 71.060 117.630 ;
        RECT 63.470 117.430 71.060 117.570 ;
        RECT 62.475 117.385 62.765 117.430 ;
        RECT 70.740 117.370 71.060 117.430 ;
        RECT 11.330 116.750 113.450 117.230 ;
        RECT 16.460 116.350 16.780 116.610 ;
        RECT 19.235 116.550 19.525 116.595 ;
        RECT 19.680 116.550 20.000 116.610 ;
        RECT 19.235 116.410 20.000 116.550 ;
        RECT 19.235 116.365 19.525 116.410 ;
        RECT 19.680 116.350 20.000 116.410 ;
        RECT 28.880 116.550 29.200 116.610 ;
        RECT 30.735 116.550 31.025 116.595 ;
        RECT 28.880 116.410 31.025 116.550 ;
        RECT 28.880 116.350 29.200 116.410 ;
        RECT 30.735 116.365 31.025 116.410 ;
        RECT 43.615 116.550 43.905 116.595 ;
        RECT 44.060 116.550 44.380 116.610 ;
        RECT 43.615 116.410 44.380 116.550 ;
        RECT 43.615 116.365 43.905 116.410 ;
        RECT 44.060 116.350 44.380 116.410 ;
        RECT 56.940 116.550 57.260 116.610 ;
        RECT 58.105 116.550 58.395 116.595 ;
        RECT 56.940 116.410 58.395 116.550 ;
        RECT 56.940 116.350 57.260 116.410 ;
        RECT 58.105 116.365 58.395 116.410 ;
        RECT 96.975 116.550 97.265 116.595 ;
        RECT 98.340 116.550 98.660 116.610 ;
        RECT 96.975 116.410 98.660 116.550 ;
        RECT 96.975 116.365 97.265 116.410 ;
        RECT 98.340 116.350 98.660 116.410 ;
        RECT 18.775 116.210 19.065 116.255 ;
        RECT 21.060 116.210 21.380 116.270 ;
        RECT 52.800 116.255 53.120 116.270 ;
        RECT 18.775 116.070 21.380 116.210 ;
        RECT 18.775 116.025 19.065 116.070 ;
        RECT 21.060 116.010 21.380 116.070 ;
        RECT 50.060 116.210 50.350 116.255 ;
        RECT 51.920 116.210 52.210 116.255 ;
        RECT 50.060 116.070 52.210 116.210 ;
        RECT 50.060 116.025 50.350 116.070 ;
        RECT 51.920 116.025 52.210 116.070 ;
        RECT 15.555 115.870 15.845 115.915 ;
        RECT 31.195 115.870 31.485 115.915 ;
        RECT 44.075 115.870 44.365 115.915 ;
        RECT 45.440 115.870 45.760 115.930 ;
        RECT 15.555 115.730 17.150 115.870 ;
        RECT 15.555 115.685 15.845 115.730 ;
        RECT 17.010 115.235 17.150 115.730 ;
        RECT 31.195 115.730 45.760 115.870 ;
        RECT 31.195 115.685 31.485 115.730 ;
        RECT 44.075 115.685 44.365 115.730 ;
        RECT 45.440 115.670 45.760 115.730 ;
        RECT 49.135 115.870 49.425 115.915 ;
        RECT 49.580 115.870 49.900 115.930 ;
        RECT 49.135 115.730 49.900 115.870 ;
        RECT 49.135 115.685 49.425 115.730 ;
        RECT 49.580 115.670 49.900 115.730 ;
        RECT 50.500 115.870 50.820 115.930 ;
        RECT 50.975 115.870 51.265 115.915 ;
        RECT 50.500 115.730 51.265 115.870 ;
        RECT 51.995 115.870 52.210 116.025 ;
        RECT 52.800 116.210 53.130 116.255 ;
        RECT 56.100 116.210 56.390 116.255 ;
        RECT 52.800 116.070 56.390 116.210 ;
        RECT 52.800 116.025 53.130 116.070 ;
        RECT 56.100 116.025 56.390 116.070 ;
        RECT 89.140 116.210 89.460 116.270 ;
        RECT 89.140 116.070 105.470 116.210 ;
        RECT 52.800 116.010 53.120 116.025 ;
        RECT 89.140 116.010 89.460 116.070 ;
        RECT 54.240 115.870 54.530 115.915 ;
        RECT 51.995 115.730 54.530 115.870 ;
        RECT 50.500 115.670 50.820 115.730 ;
        RECT 50.975 115.685 51.265 115.730 ;
        RECT 54.240 115.685 54.530 115.730 ;
        RECT 96.040 115.670 96.360 115.930 ;
        RECT 105.330 115.915 105.470 116.070 ;
        RECT 105.255 115.685 105.545 115.915 ;
        RECT 105.700 115.670 106.020 115.930 ;
        RECT 106.160 115.870 106.480 115.930 ;
        RECT 108.935 115.870 109.225 115.915 ;
        RECT 106.160 115.730 109.225 115.870 ;
        RECT 106.160 115.670 106.480 115.730 ;
        RECT 108.935 115.685 109.225 115.730 ;
        RECT 20.140 115.330 20.460 115.590 ;
        RECT 16.935 115.005 17.225 115.235 ;
        RECT 49.600 115.190 49.890 115.235 ;
        RECT 51.460 115.190 51.750 115.235 ;
        RECT 54.240 115.190 54.530 115.235 ;
        RECT 49.600 115.050 54.530 115.190 ;
        RECT 49.600 115.005 49.890 115.050 ;
        RECT 51.460 115.005 51.750 115.050 ;
        RECT 54.240 115.005 54.530 115.050 ;
        RECT 102.940 114.850 103.260 114.910 ;
        RECT 104.335 114.850 104.625 114.895 ;
        RECT 102.940 114.710 104.625 114.850 ;
        RECT 102.940 114.650 103.260 114.710 ;
        RECT 104.335 114.665 104.625 114.710 ;
        RECT 106.160 114.650 106.480 114.910 ;
        RECT 106.620 114.850 106.940 114.910 ;
        RECT 108.015 114.850 108.305 114.895 ;
        RECT 106.620 114.710 108.305 114.850 ;
        RECT 106.620 114.650 106.940 114.710 ;
        RECT 108.015 114.665 108.305 114.710 ;
        RECT 11.330 114.030 113.450 114.510 ;
        RECT 50.515 113.830 50.805 113.875 ;
        RECT 52.800 113.830 53.120 113.890 ;
        RECT 50.515 113.690 53.120 113.830 ;
        RECT 50.515 113.645 50.805 113.690 ;
        RECT 52.800 113.630 53.120 113.690 ;
        RECT 66.140 113.830 66.460 113.890 ;
        RECT 69.835 113.830 70.125 113.875 ;
        RECT 66.140 113.690 70.125 113.830 ;
        RECT 66.140 113.630 66.460 113.690 ;
        RECT 69.835 113.645 70.125 113.690 ;
        RECT 96.960 113.630 97.280 113.890 ;
        RECT 18.415 113.490 18.705 113.535 ;
        RECT 21.535 113.490 21.825 113.535 ;
        RECT 23.425 113.490 23.715 113.535 ;
        RECT 18.415 113.350 23.715 113.490 ;
        RECT 18.415 113.305 18.705 113.350 ;
        RECT 21.535 113.305 21.825 113.350 ;
        RECT 23.425 113.305 23.715 113.350 ;
        RECT 31.640 113.490 31.960 113.550 ;
        RECT 39.935 113.490 40.225 113.535 ;
        RECT 31.640 113.350 40.225 113.490 ;
        RECT 31.640 113.290 31.960 113.350 ;
        RECT 39.935 113.305 40.225 113.350 ;
        RECT 65.220 113.490 65.540 113.550 ;
        RECT 67.995 113.490 68.285 113.535 ;
        RECT 65.220 113.350 68.285 113.490 ;
        RECT 65.220 113.290 65.540 113.350 ;
        RECT 67.995 113.305 68.285 113.350 ;
        RECT 96.500 113.490 96.820 113.550 ;
        RECT 97.435 113.490 97.725 113.535 ;
        RECT 96.500 113.350 97.725 113.490 ;
        RECT 96.500 113.290 96.820 113.350 ;
        RECT 97.435 113.305 97.725 113.350 ;
        RECT 102.445 113.490 102.735 113.535 ;
        RECT 104.335 113.490 104.625 113.535 ;
        RECT 107.455 113.490 107.745 113.535 ;
        RECT 102.445 113.350 107.745 113.490 ;
        RECT 102.445 113.305 102.735 113.350 ;
        RECT 104.335 113.305 104.625 113.350 ;
        RECT 107.455 113.305 107.745 113.350 ;
        RECT 60.620 113.150 60.940 113.210 ;
        RECT 71.660 113.150 71.980 113.210 ;
        RECT 52.890 113.010 60.940 113.150 ;
        RECT 14.160 112.270 14.480 112.530 ;
        RECT 17.335 112.515 17.625 112.830 ;
        RECT 18.415 112.810 18.705 112.855 ;
        RECT 21.995 112.810 22.285 112.855 ;
        RECT 23.830 112.810 24.120 112.855 ;
        RECT 18.415 112.670 24.120 112.810 ;
        RECT 18.415 112.625 18.705 112.670 ;
        RECT 21.995 112.625 22.285 112.670 ;
        RECT 23.830 112.625 24.120 112.670 ;
        RECT 24.295 112.810 24.585 112.855 ;
        RECT 25.200 112.810 25.520 112.870 ;
        RECT 24.295 112.670 25.520 112.810 ;
        RECT 24.295 112.625 24.585 112.670 ;
        RECT 25.200 112.610 25.520 112.670 ;
        RECT 27.040 112.810 27.360 112.870 ;
        RECT 28.435 112.810 28.725 112.855 ;
        RECT 27.040 112.670 28.725 112.810 ;
        RECT 27.040 112.610 27.360 112.670 ;
        RECT 28.435 112.625 28.725 112.670 ;
        RECT 36.240 112.810 36.560 112.870 ;
        RECT 37.175 112.810 37.465 112.855 ;
        RECT 36.240 112.670 37.465 112.810 ;
        RECT 36.240 112.610 36.560 112.670 ;
        RECT 37.175 112.625 37.465 112.670 ;
        RECT 40.840 112.610 41.160 112.870 ;
        RECT 42.680 112.810 43.000 112.870 ;
        RECT 44.075 112.810 44.365 112.855 ;
        RECT 42.680 112.670 44.365 112.810 ;
        RECT 42.680 112.610 43.000 112.670 ;
        RECT 44.075 112.625 44.365 112.670 ;
        RECT 50.055 112.810 50.345 112.855 ;
        RECT 51.435 112.810 51.725 112.855 ;
        RECT 52.890 112.810 53.030 113.010 ;
        RECT 60.620 112.950 60.940 113.010 ;
        RECT 67.610 113.010 71.980 113.150 ;
        RECT 50.055 112.670 53.030 112.810 ;
        RECT 56.955 112.810 57.245 112.855 ;
        RECT 57.400 112.810 57.720 112.870 ;
        RECT 56.955 112.670 57.720 112.810 ;
        RECT 50.055 112.625 50.345 112.670 ;
        RECT 51.435 112.625 51.725 112.670 ;
        RECT 56.955 112.625 57.245 112.670 ;
        RECT 57.400 112.610 57.720 112.670 ;
        RECT 60.160 112.610 60.480 112.870 ;
        RECT 67.610 112.855 67.750 113.010 ;
        RECT 71.660 112.950 71.980 113.010 ;
        RECT 95.580 113.150 95.900 113.210 ;
        RECT 95.580 113.010 98.570 113.150 ;
        RECT 95.580 112.950 95.900 113.010 ;
        RECT 67.535 112.625 67.825 112.855 ;
        RECT 68.440 112.810 68.760 112.870 ;
        RECT 68.915 112.810 69.205 112.855 ;
        RECT 68.440 112.670 69.205 112.810 ;
        RECT 68.440 112.610 68.760 112.670 ;
        RECT 68.915 112.625 69.205 112.670 ;
        RECT 70.280 112.610 70.600 112.870 ;
        RECT 70.740 112.610 71.060 112.870 ;
        RECT 83.175 112.625 83.465 112.855 ;
        RECT 85.460 112.810 85.780 112.870 ;
        RECT 88.235 112.810 88.525 112.855 ;
        RECT 85.460 112.670 88.525 112.810 ;
        RECT 17.035 112.470 17.625 112.515 ;
        RECT 19.220 112.470 19.540 112.530 ;
        RECT 20.275 112.470 20.925 112.515 ;
        RECT 17.035 112.330 20.925 112.470 ;
        RECT 17.035 112.285 17.325 112.330 ;
        RECT 19.220 112.270 19.540 112.330 ;
        RECT 20.275 112.285 20.925 112.330 ;
        RECT 22.915 112.470 23.205 112.515 ;
        RECT 23.360 112.470 23.680 112.530 ;
        RECT 22.915 112.330 23.680 112.470 ;
        RECT 22.915 112.285 23.205 112.330 ;
        RECT 23.360 112.270 23.680 112.330 ;
        RECT 50.500 112.470 50.820 112.530 ;
        RECT 52.815 112.470 53.105 112.515 ;
        RECT 50.500 112.330 53.105 112.470 ;
        RECT 50.500 112.270 50.820 112.330 ;
        RECT 52.815 112.285 53.105 112.330 ;
        RECT 62.000 112.470 62.320 112.530 ;
        RECT 83.250 112.470 83.390 112.625 ;
        RECT 85.460 112.610 85.780 112.670 ;
        RECT 88.235 112.625 88.525 112.670 ;
        RECT 93.755 112.810 94.045 112.855 ;
        RECT 94.660 112.810 94.980 112.870 ;
        RECT 98.430 112.855 98.570 113.010 ;
        RECT 101.560 112.950 101.880 113.210 ;
        RECT 102.955 113.150 103.245 113.195 ;
        RECT 106.620 113.150 106.940 113.210 ;
        RECT 102.955 113.010 106.940 113.150 ;
        RECT 102.955 112.965 103.245 113.010 ;
        RECT 106.620 112.950 106.940 113.010 ;
        RECT 93.755 112.670 94.980 112.810 ;
        RECT 93.755 112.625 94.045 112.670 ;
        RECT 94.660 112.610 94.980 112.670 ;
        RECT 96.055 112.625 96.345 112.855 ;
        RECT 98.355 112.625 98.645 112.855 ;
        RECT 102.040 112.810 102.330 112.855 ;
        RECT 103.875 112.810 104.165 112.855 ;
        RECT 107.455 112.810 107.745 112.855 ;
        RECT 102.040 112.670 107.745 112.810 ;
        RECT 102.040 112.625 102.330 112.670 ;
        RECT 103.875 112.625 104.165 112.670 ;
        RECT 107.455 112.625 107.745 112.670 ;
        RECT 62.000 112.330 83.390 112.470 ;
        RECT 96.130 112.470 96.270 112.625 ;
        RECT 100.180 112.470 100.500 112.530 ;
        RECT 96.130 112.330 100.500 112.470 ;
        RECT 62.000 112.270 62.320 112.330 ;
        RECT 100.180 112.270 100.500 112.330 ;
        RECT 105.235 112.470 105.885 112.515 ;
        RECT 106.160 112.470 106.480 112.530 ;
        RECT 108.535 112.515 108.825 112.830 ;
        RECT 108.535 112.470 109.125 112.515 ;
        RECT 105.235 112.330 109.125 112.470 ;
        RECT 105.235 112.285 105.885 112.330 ;
        RECT 106.160 112.270 106.480 112.330 ;
        RECT 108.835 112.285 109.125 112.330 ;
        RECT 111.695 112.470 111.985 112.515 ;
        RECT 114.440 112.470 114.760 112.530 ;
        RECT 111.695 112.330 114.760 112.470 ;
        RECT 111.695 112.285 111.985 112.330 ;
        RECT 114.440 112.270 114.760 112.330 ;
        RECT 27.975 112.130 28.265 112.175 ;
        RECT 28.420 112.130 28.740 112.190 ;
        RECT 27.975 111.990 28.740 112.130 ;
        RECT 27.975 111.945 28.265 111.990 ;
        RECT 28.420 111.930 28.740 111.990 ;
        RECT 36.240 111.930 36.560 112.190 ;
        RECT 44.995 112.130 45.285 112.175 ;
        RECT 46.820 112.130 47.140 112.190 ;
        RECT 44.995 111.990 47.140 112.130 ;
        RECT 44.995 111.945 45.285 111.990 ;
        RECT 46.820 111.930 47.140 111.990 ;
        RECT 57.875 112.130 58.165 112.175 ;
        RECT 60.160 112.130 60.480 112.190 ;
        RECT 57.875 111.990 60.480 112.130 ;
        RECT 57.875 111.945 58.165 111.990 ;
        RECT 60.160 111.930 60.480 111.990 ;
        RECT 61.095 112.130 61.385 112.175 ;
        RECT 61.540 112.130 61.860 112.190 ;
        RECT 61.095 111.990 61.860 112.130 ;
        RECT 61.095 111.945 61.385 111.990 ;
        RECT 61.540 111.930 61.860 111.990 ;
        RECT 66.600 112.130 66.920 112.190 ;
        RECT 67.075 112.130 67.365 112.175 ;
        RECT 66.600 111.990 67.365 112.130 ;
        RECT 66.600 111.930 66.920 111.990 ;
        RECT 67.075 111.945 67.365 111.990 ;
        RECT 83.620 112.130 83.940 112.190 ;
        RECT 84.095 112.130 84.385 112.175 ;
        RECT 83.620 111.990 84.385 112.130 ;
        RECT 83.620 111.930 83.940 111.990 ;
        RECT 84.095 111.945 84.385 111.990 ;
        RECT 89.140 111.930 89.460 112.190 ;
        RECT 94.675 112.130 94.965 112.175 ;
        RECT 97.420 112.130 97.740 112.190 ;
        RECT 94.675 111.990 97.740 112.130 ;
        RECT 94.675 111.945 94.965 111.990 ;
        RECT 97.420 111.930 97.740 111.990 ;
        RECT 11.330 111.310 113.450 111.790 ;
        RECT 18.775 111.110 19.065 111.155 ;
        RECT 19.220 111.110 19.540 111.170 ;
        RECT 18.775 110.970 19.540 111.110 ;
        RECT 18.775 110.925 19.065 110.970 ;
        RECT 19.220 110.910 19.540 110.970 ;
        RECT 21.520 110.910 21.840 111.170 ;
        RECT 23.360 110.910 23.680 111.170 ;
        RECT 43.600 111.110 43.920 111.170 ;
        RECT 43.600 110.970 49.350 111.110 ;
        RECT 43.600 110.910 43.920 110.970 ;
        RECT 23.820 110.770 24.140 110.830 ;
        RECT 33.940 110.815 34.260 110.830 ;
        RECT 30.375 110.770 30.665 110.815 ;
        RECT 33.615 110.770 34.265 110.815 ;
        RECT 23.820 110.630 25.890 110.770 ;
        RECT 23.820 110.570 24.140 110.630 ;
        RECT 16.920 110.430 17.240 110.490 ;
        RECT 19.235 110.430 19.525 110.475 ;
        RECT 16.920 110.290 19.525 110.430 ;
        RECT 16.920 110.230 17.240 110.290 ;
        RECT 19.235 110.245 19.525 110.290 ;
        RECT 22.455 110.430 22.745 110.475 ;
        RECT 22.900 110.430 23.220 110.490 ;
        RECT 22.455 110.290 23.220 110.430 ;
        RECT 22.455 110.245 22.745 110.290 ;
        RECT 19.310 110.090 19.450 110.245 ;
        RECT 22.900 110.230 23.220 110.290 ;
        RECT 24.280 110.230 24.600 110.490 ;
        RECT 25.750 110.475 25.890 110.630 ;
        RECT 30.375 110.630 34.265 110.770 ;
        RECT 30.375 110.585 30.965 110.630 ;
        RECT 33.615 110.585 34.265 110.630 ;
        RECT 25.675 110.245 25.965 110.475 ;
        RECT 26.135 110.430 26.425 110.475 ;
        RECT 27.960 110.430 28.280 110.490 ;
        RECT 26.135 110.290 28.280 110.430 ;
        RECT 26.135 110.245 26.425 110.290 ;
        RECT 27.960 110.230 28.280 110.290 ;
        RECT 30.675 110.270 30.965 110.585 ;
        RECT 33.940 110.570 34.260 110.585 ;
        RECT 36.240 110.570 36.560 110.830 ;
        RECT 44.060 110.815 44.380 110.830 ;
        RECT 40.955 110.770 41.245 110.815 ;
        RECT 44.060 110.770 44.845 110.815 ;
        RECT 40.955 110.630 44.845 110.770 ;
        RECT 40.955 110.585 41.545 110.630 ;
        RECT 31.755 110.430 32.045 110.475 ;
        RECT 35.335 110.430 35.625 110.475 ;
        RECT 37.170 110.430 37.460 110.475 ;
        RECT 31.755 110.290 37.460 110.430 ;
        RECT 31.755 110.245 32.045 110.290 ;
        RECT 35.335 110.245 35.625 110.290 ;
        RECT 37.170 110.245 37.460 110.290 ;
        RECT 41.255 110.270 41.545 110.585 ;
        RECT 44.060 110.585 44.845 110.630 ;
        RECT 44.060 110.570 44.380 110.585 ;
        RECT 46.820 110.570 47.140 110.830 ;
        RECT 49.210 110.475 49.350 110.970 ;
        RECT 61.080 110.910 61.400 111.170 ;
        RECT 69.820 110.910 70.140 111.170 ;
        RECT 83.620 111.110 83.940 111.170 ;
        RECT 83.620 110.970 87.070 111.110 ;
        RECT 83.620 110.910 83.940 110.970 ;
        RECT 54.295 110.770 54.585 110.815 ;
        RECT 56.480 110.770 56.800 110.830 ;
        RECT 57.535 110.770 58.185 110.815 ;
        RECT 54.295 110.630 58.185 110.770 ;
        RECT 54.295 110.585 54.885 110.630 ;
        RECT 42.335 110.430 42.625 110.475 ;
        RECT 45.915 110.430 46.205 110.475 ;
        RECT 47.750 110.430 48.040 110.475 ;
        RECT 42.335 110.290 48.040 110.430 ;
        RECT 42.335 110.245 42.625 110.290 ;
        RECT 45.915 110.245 46.205 110.290 ;
        RECT 47.750 110.245 48.040 110.290 ;
        RECT 49.135 110.245 49.425 110.475 ;
        RECT 51.435 110.430 51.725 110.475 ;
        RECT 53.720 110.430 54.040 110.490 ;
        RECT 51.435 110.290 54.040 110.430 ;
        RECT 51.435 110.245 51.725 110.290 ;
        RECT 53.720 110.230 54.040 110.290 ;
        RECT 54.595 110.270 54.885 110.585 ;
        RECT 56.480 110.570 56.800 110.630 ;
        RECT 57.535 110.585 58.185 110.630 ;
        RECT 60.160 110.570 60.480 110.830 ;
        RECT 61.170 110.770 61.310 110.910 ;
        RECT 65.795 110.770 66.085 110.815 ;
        RECT 66.600 110.770 66.920 110.830 ;
        RECT 69.035 110.770 69.685 110.815 ;
        RECT 61.170 110.630 61.770 110.770 ;
        RECT 61.630 110.475 61.770 110.630 ;
        RECT 65.795 110.630 69.685 110.770 ;
        RECT 69.910 110.770 70.050 110.910 ;
        RECT 84.540 110.815 84.860 110.830 ;
        RECT 86.930 110.815 87.070 110.970 ;
        RECT 80.975 110.770 81.265 110.815 ;
        RECT 84.215 110.770 84.865 110.815 ;
        RECT 69.910 110.630 76.950 110.770 ;
        RECT 65.795 110.585 66.385 110.630 ;
        RECT 55.675 110.430 55.965 110.475 ;
        RECT 59.255 110.430 59.545 110.475 ;
        RECT 61.090 110.430 61.380 110.475 ;
        RECT 55.675 110.290 61.380 110.430 ;
        RECT 55.675 110.245 55.965 110.290 ;
        RECT 59.255 110.245 59.545 110.290 ;
        RECT 61.090 110.245 61.380 110.290 ;
        RECT 61.555 110.245 61.845 110.475 ;
        RECT 66.095 110.270 66.385 110.585 ;
        RECT 66.600 110.570 66.920 110.630 ;
        RECT 69.035 110.585 69.685 110.630 ;
        RECT 67.175 110.430 67.465 110.475 ;
        RECT 70.755 110.430 71.045 110.475 ;
        RECT 72.590 110.430 72.880 110.475 ;
        RECT 67.175 110.290 72.880 110.430 ;
        RECT 67.175 110.245 67.465 110.290 ;
        RECT 70.755 110.245 71.045 110.290 ;
        RECT 72.590 110.245 72.880 110.290 ;
        RECT 27.040 110.090 27.360 110.150 ;
        RECT 19.310 109.950 27.360 110.090 ;
        RECT 27.040 109.890 27.360 109.950 ;
        RECT 27.515 110.090 27.805 110.135 ;
        RECT 30.260 110.090 30.580 110.150 ;
        RECT 27.515 109.950 30.580 110.090 ;
        RECT 27.515 109.905 27.805 109.950 ;
        RECT 30.260 109.890 30.580 109.950 ;
        RECT 37.620 109.890 37.940 110.150 ;
        RECT 38.095 110.090 38.385 110.135 ;
        RECT 41.760 110.090 42.080 110.150 ;
        RECT 38.095 109.950 42.080 110.090 ;
        RECT 38.095 109.905 38.385 109.950 ;
        RECT 41.760 109.890 42.080 109.950 ;
        RECT 48.215 110.090 48.505 110.135 ;
        RECT 49.580 110.090 49.900 110.150 ;
        RECT 56.940 110.090 57.260 110.150 ;
        RECT 61.630 110.090 61.770 110.245 ;
        RECT 73.040 110.230 73.360 110.490 ;
        RECT 73.500 110.430 73.820 110.490 ;
        RECT 76.810 110.475 76.950 110.630 ;
        RECT 80.975 110.630 84.865 110.770 ;
        RECT 80.975 110.585 81.565 110.630 ;
        RECT 84.215 110.585 84.865 110.630 ;
        RECT 86.855 110.585 87.145 110.815 ;
        RECT 91.555 110.770 91.845 110.815 ;
        RECT 94.795 110.770 95.445 110.815 ;
        RECT 91.555 110.630 95.445 110.770 ;
        RECT 91.555 110.585 92.145 110.630 ;
        RECT 94.795 110.585 95.445 110.630 ;
        RECT 75.815 110.430 76.105 110.475 ;
        RECT 73.500 110.290 76.105 110.430 ;
        RECT 73.500 110.230 73.820 110.290 ;
        RECT 75.815 110.245 76.105 110.290 ;
        RECT 76.735 110.245 77.025 110.475 ;
        RECT 78.115 110.430 78.405 110.475 ;
        RECT 80.400 110.430 80.720 110.490 ;
        RECT 78.115 110.290 80.720 110.430 ;
        RECT 78.115 110.245 78.405 110.290 ;
        RECT 80.400 110.230 80.720 110.290 ;
        RECT 81.275 110.270 81.565 110.585 ;
        RECT 84.540 110.570 84.860 110.585 ;
        RECT 91.855 110.490 92.145 110.585 ;
        RECT 97.420 110.570 97.740 110.830 ;
        RECT 102.940 110.570 103.260 110.830 ;
        RECT 105.235 110.770 105.885 110.815 ;
        RECT 106.160 110.770 106.480 110.830 ;
        RECT 108.835 110.770 109.125 110.815 ;
        RECT 105.235 110.630 109.125 110.770 ;
        RECT 105.235 110.585 105.885 110.630 ;
        RECT 106.160 110.570 106.480 110.630 ;
        RECT 108.535 110.585 109.125 110.630 ;
        RECT 82.355 110.430 82.645 110.475 ;
        RECT 85.935 110.430 86.225 110.475 ;
        RECT 87.770 110.430 88.060 110.475 ;
        RECT 82.355 110.290 88.060 110.430 ;
        RECT 82.355 110.245 82.645 110.290 ;
        RECT 85.935 110.245 86.225 110.290 ;
        RECT 87.770 110.245 88.060 110.290 ;
        RECT 91.855 110.270 92.220 110.490 ;
        RECT 91.900 110.230 92.220 110.270 ;
        RECT 92.935 110.430 93.225 110.475 ;
        RECT 96.515 110.430 96.805 110.475 ;
        RECT 98.350 110.430 98.640 110.475 ;
        RECT 92.935 110.290 98.640 110.430 ;
        RECT 92.935 110.245 93.225 110.290 ;
        RECT 96.515 110.245 96.805 110.290 ;
        RECT 98.350 110.245 98.640 110.290 ;
        RECT 98.815 110.430 99.105 110.475 ;
        RECT 99.260 110.430 99.580 110.490 ;
        RECT 101.560 110.430 101.880 110.490 ;
        RECT 98.815 110.290 101.880 110.430 ;
        RECT 98.815 110.245 99.105 110.290 ;
        RECT 99.260 110.230 99.580 110.290 ;
        RECT 101.560 110.230 101.880 110.290 ;
        RECT 102.040 110.430 102.330 110.475 ;
        RECT 103.875 110.430 104.165 110.475 ;
        RECT 107.455 110.430 107.745 110.475 ;
        RECT 102.040 110.290 107.745 110.430 ;
        RECT 102.040 110.245 102.330 110.290 ;
        RECT 103.875 110.245 104.165 110.290 ;
        RECT 107.455 110.245 107.745 110.290 ;
        RECT 108.535 110.270 108.825 110.585 ;
        RECT 48.215 109.950 61.770 110.090 ;
        RECT 62.935 110.090 63.225 110.135 ;
        RECT 64.760 110.090 65.080 110.150 ;
        RECT 62.935 109.950 65.080 110.090 ;
        RECT 48.215 109.905 48.505 109.950 ;
        RECT 49.580 109.890 49.900 109.950 ;
        RECT 56.940 109.890 57.260 109.950 ;
        RECT 62.935 109.905 63.225 109.950 ;
        RECT 64.760 109.890 65.080 109.950 ;
        RECT 71.675 110.090 71.965 110.135 ;
        RECT 73.130 110.090 73.270 110.230 ;
        RECT 83.620 110.090 83.940 110.150 ;
        RECT 88.235 110.090 88.525 110.135 ;
        RECT 71.675 109.950 72.810 110.090 ;
        RECT 73.130 109.950 88.525 110.090 ;
        RECT 71.675 109.905 71.965 109.950 ;
        RECT 31.755 109.750 32.045 109.795 ;
        RECT 34.875 109.750 35.165 109.795 ;
        RECT 36.765 109.750 37.055 109.795 ;
        RECT 31.755 109.610 37.055 109.750 ;
        RECT 31.755 109.565 32.045 109.610 ;
        RECT 34.875 109.565 35.165 109.610 ;
        RECT 36.765 109.565 37.055 109.610 ;
        RECT 42.335 109.750 42.625 109.795 ;
        RECT 45.455 109.750 45.745 109.795 ;
        RECT 47.345 109.750 47.635 109.795 ;
        RECT 42.335 109.610 47.635 109.750 ;
        RECT 42.335 109.565 42.625 109.610 ;
        RECT 45.455 109.565 45.745 109.610 ;
        RECT 47.345 109.565 47.635 109.610 ;
        RECT 55.675 109.750 55.965 109.795 ;
        RECT 58.795 109.750 59.085 109.795 ;
        RECT 60.685 109.750 60.975 109.795 ;
        RECT 55.675 109.610 60.975 109.750 ;
        RECT 55.675 109.565 55.965 109.610 ;
        RECT 58.795 109.565 59.085 109.610 ;
        RECT 60.685 109.565 60.975 109.610 ;
        RECT 67.175 109.750 67.465 109.795 ;
        RECT 70.295 109.750 70.585 109.795 ;
        RECT 72.185 109.750 72.475 109.795 ;
        RECT 67.175 109.610 72.475 109.750 ;
        RECT 72.670 109.750 72.810 109.950 ;
        RECT 83.620 109.890 83.940 109.950 ;
        RECT 88.235 109.905 88.525 109.950 ;
        RECT 88.695 110.090 88.985 110.135 ;
        RECT 91.440 110.090 91.760 110.150 ;
        RECT 88.695 109.950 91.760 110.090 ;
        RECT 88.695 109.905 88.985 109.950 ;
        RECT 91.440 109.890 91.760 109.950 ;
        RECT 109.840 110.090 110.160 110.150 ;
        RECT 111.695 110.090 111.985 110.135 ;
        RECT 109.840 109.950 111.985 110.090 ;
        RECT 109.840 109.890 110.160 109.950 ;
        RECT 111.695 109.905 111.985 109.950 ;
        RECT 74.895 109.750 75.185 109.795 ;
        RECT 72.670 109.610 75.185 109.750 ;
        RECT 67.175 109.565 67.465 109.610 ;
        RECT 70.295 109.565 70.585 109.610 ;
        RECT 72.185 109.565 72.475 109.610 ;
        RECT 74.895 109.565 75.185 109.610 ;
        RECT 82.355 109.750 82.645 109.795 ;
        RECT 85.475 109.750 85.765 109.795 ;
        RECT 87.365 109.750 87.655 109.795 ;
        RECT 82.355 109.610 87.655 109.750 ;
        RECT 82.355 109.565 82.645 109.610 ;
        RECT 85.475 109.565 85.765 109.610 ;
        RECT 87.365 109.565 87.655 109.610 ;
        RECT 92.935 109.750 93.225 109.795 ;
        RECT 96.055 109.750 96.345 109.795 ;
        RECT 97.945 109.750 98.235 109.795 ;
        RECT 92.935 109.610 98.235 109.750 ;
        RECT 92.935 109.565 93.225 109.610 ;
        RECT 96.055 109.565 96.345 109.610 ;
        RECT 97.945 109.565 98.235 109.610 ;
        RECT 102.445 109.750 102.735 109.795 ;
        RECT 104.335 109.750 104.625 109.795 ;
        RECT 107.455 109.750 107.745 109.795 ;
        RECT 102.445 109.610 107.745 109.750 ;
        RECT 102.445 109.565 102.735 109.610 ;
        RECT 104.335 109.565 104.625 109.610 ;
        RECT 107.455 109.565 107.745 109.610 ;
        RECT 23.360 109.410 23.680 109.470 ;
        RECT 24.755 109.410 25.045 109.455 ;
        RECT 23.360 109.270 25.045 109.410 ;
        RECT 23.360 109.210 23.680 109.270 ;
        RECT 24.755 109.225 25.045 109.270 ;
        RECT 27.040 109.210 27.360 109.470 ;
        RECT 50.040 109.210 50.360 109.470 ;
        RECT 77.655 109.410 77.945 109.455 ;
        RECT 79.480 109.410 79.800 109.470 ;
        RECT 77.655 109.270 79.800 109.410 ;
        RECT 77.655 109.225 77.945 109.270 ;
        RECT 79.480 109.210 79.800 109.270 ;
        RECT 11.330 108.590 113.450 109.070 ;
        RECT 13.700 108.190 14.020 108.450 ;
        RECT 33.940 108.390 34.260 108.450 ;
        RECT 36.715 108.390 37.005 108.435 ;
        RECT 33.940 108.250 37.005 108.390 ;
        RECT 33.940 108.190 34.260 108.250 ;
        RECT 36.715 108.205 37.005 108.250 ;
        RECT 44.060 108.190 44.380 108.450 ;
        RECT 56.035 108.390 56.325 108.435 ;
        RECT 56.480 108.390 56.800 108.450 ;
        RECT 56.035 108.250 56.800 108.390 ;
        RECT 56.035 108.205 56.325 108.250 ;
        RECT 56.480 108.190 56.800 108.250 ;
        RECT 70.280 108.390 70.600 108.450 ;
        RECT 70.280 108.250 84.310 108.390 ;
        RECT 70.280 108.190 70.600 108.250 ;
        RECT 18.875 108.050 19.165 108.095 ;
        RECT 21.995 108.050 22.285 108.095 ;
        RECT 23.885 108.050 24.175 108.095 ;
        RECT 18.875 107.910 24.175 108.050 ;
        RECT 18.875 107.865 19.165 107.910 ;
        RECT 21.995 107.865 22.285 107.910 ;
        RECT 23.885 107.865 24.175 107.910 ;
        RECT 26.085 108.050 26.375 108.095 ;
        RECT 27.975 108.050 28.265 108.095 ;
        RECT 31.095 108.050 31.385 108.095 ;
        RECT 26.085 107.910 31.385 108.050 ;
        RECT 26.085 107.865 26.375 107.910 ;
        RECT 27.975 107.865 28.265 107.910 ;
        RECT 31.095 107.865 31.385 107.910 ;
        RECT 49.235 108.050 49.525 108.095 ;
        RECT 52.355 108.050 52.645 108.095 ;
        RECT 54.245 108.050 54.535 108.095 ;
        RECT 49.235 107.910 54.535 108.050 ;
        RECT 49.235 107.865 49.525 107.910 ;
        RECT 52.355 107.865 52.645 107.910 ;
        RECT 54.245 107.865 54.535 107.910 ;
        RECT 66.255 108.050 66.545 108.095 ;
        RECT 69.375 108.050 69.665 108.095 ;
        RECT 71.265 108.050 71.555 108.095 ;
        RECT 66.255 107.910 71.555 108.050 ;
        RECT 66.255 107.865 66.545 107.910 ;
        RECT 69.375 107.865 69.665 107.910 ;
        RECT 71.265 107.865 71.555 107.910 ;
        RECT 77.755 108.050 78.045 108.095 ;
        RECT 80.875 108.050 81.165 108.095 ;
        RECT 82.765 108.050 83.055 108.095 ;
        RECT 77.755 107.910 83.055 108.050 ;
        RECT 84.170 108.050 84.310 108.250 ;
        RECT 84.540 108.190 84.860 108.450 ;
        RECT 110.775 108.390 111.065 108.435 ;
        RECT 87.850 108.250 111.065 108.390 ;
        RECT 87.850 108.050 87.990 108.250 ;
        RECT 110.775 108.205 111.065 108.250 ;
        RECT 84.170 107.910 87.990 108.050 ;
        RECT 92.015 108.050 92.305 108.095 ;
        RECT 95.135 108.050 95.425 108.095 ;
        RECT 97.025 108.050 97.315 108.095 ;
        RECT 92.015 107.910 97.315 108.050 ;
        RECT 77.755 107.865 78.045 107.910 ;
        RECT 80.875 107.865 81.165 107.910 ;
        RECT 82.765 107.865 83.055 107.910 ;
        RECT 92.015 107.865 92.305 107.910 ;
        RECT 95.135 107.865 95.425 107.910 ;
        RECT 97.025 107.865 97.315 107.910 ;
        RECT 100.145 108.050 100.435 108.095 ;
        RECT 102.035 108.050 102.325 108.095 ;
        RECT 105.155 108.050 105.445 108.095 ;
        RECT 100.145 107.910 105.445 108.050 ;
        RECT 100.145 107.865 100.435 107.910 ;
        RECT 102.035 107.865 102.325 107.910 ;
        RECT 105.155 107.865 105.445 107.910 ;
        RECT 14.635 107.710 14.925 107.755 ;
        RECT 20.600 107.710 20.920 107.770 ;
        RECT 14.635 107.570 20.920 107.710 ;
        RECT 14.635 107.525 14.925 107.570 ;
        RECT 20.600 107.510 20.920 107.570 ;
        RECT 23.360 107.510 23.680 107.770 ;
        RECT 26.595 107.710 26.885 107.755 ;
        RECT 31.640 107.710 31.960 107.770 ;
        RECT 38.555 107.710 38.845 107.755 ;
        RECT 26.595 107.570 31.960 107.710 ;
        RECT 26.595 107.525 26.885 107.570 ;
        RECT 31.640 107.510 31.960 107.570 ;
        RECT 32.190 107.570 38.845 107.710 ;
        RECT 14.175 107.370 14.465 107.415 ;
        RECT 16.920 107.370 17.240 107.430 ;
        RECT 14.175 107.230 17.240 107.370 ;
        RECT 14.175 107.185 14.465 107.230 ;
        RECT 16.920 107.170 17.240 107.230 ;
        RECT 17.795 107.075 18.085 107.390 ;
        RECT 18.875 107.370 19.165 107.415 ;
        RECT 22.455 107.370 22.745 107.415 ;
        RECT 24.290 107.370 24.580 107.415 ;
        RECT 18.875 107.230 24.580 107.370 ;
        RECT 18.875 107.185 19.165 107.230 ;
        RECT 22.455 107.185 22.745 107.230 ;
        RECT 24.290 107.185 24.580 107.230 ;
        RECT 24.755 107.370 25.045 107.415 ;
        RECT 25.200 107.370 25.520 107.430 ;
        RECT 24.755 107.230 25.520 107.370 ;
        RECT 24.755 107.185 25.045 107.230 ;
        RECT 25.200 107.170 25.520 107.230 ;
        RECT 25.680 107.370 25.970 107.415 ;
        RECT 27.515 107.370 27.805 107.415 ;
        RECT 31.095 107.370 31.385 107.415 ;
        RECT 32.190 107.390 32.330 107.570 ;
        RECT 38.555 107.525 38.845 107.570 ;
        RECT 50.040 107.710 50.360 107.770 ;
        RECT 53.735 107.710 54.025 107.755 ;
        RECT 50.040 107.570 54.025 107.710 ;
        RECT 50.040 107.510 50.360 107.570 ;
        RECT 53.735 107.525 54.025 107.570 ;
        RECT 55.115 107.710 55.405 107.755 ;
        RECT 56.940 107.710 57.260 107.770 ;
        RECT 55.115 107.570 57.260 107.710 ;
        RECT 55.115 107.525 55.405 107.570 ;
        RECT 56.940 107.510 57.260 107.570 ;
        RECT 61.540 107.710 61.860 107.770 ;
        RECT 70.755 107.710 71.045 107.755 ;
        RECT 61.540 107.570 71.045 107.710 ;
        RECT 61.540 107.510 61.860 107.570 ;
        RECT 70.755 107.525 71.045 107.570 ;
        RECT 72.135 107.710 72.425 107.755 ;
        RECT 73.040 107.710 73.360 107.770 ;
        RECT 72.135 107.570 73.360 107.710 ;
        RECT 72.135 107.525 72.425 107.570 ;
        RECT 73.040 107.510 73.360 107.570 ;
        RECT 79.480 107.710 79.800 107.770 ;
        RECT 82.255 107.710 82.545 107.755 ;
        RECT 79.480 107.570 82.545 107.710 ;
        RECT 79.480 107.510 79.800 107.570 ;
        RECT 82.255 107.525 82.545 107.570 ;
        RECT 83.620 107.510 83.940 107.770 ;
        RECT 89.140 107.710 89.460 107.770 ;
        RECT 96.515 107.710 96.805 107.755 ;
        RECT 89.140 107.570 96.805 107.710 ;
        RECT 89.140 107.510 89.460 107.570 ;
        RECT 96.515 107.525 96.805 107.570 ;
        RECT 97.895 107.710 98.185 107.755 ;
        RECT 99.260 107.710 99.580 107.770 ;
        RECT 97.895 107.570 99.580 107.710 ;
        RECT 97.895 107.525 98.185 107.570 ;
        RECT 99.260 107.510 99.580 107.570 ;
        RECT 103.400 107.710 103.720 107.770 ;
        RECT 109.395 107.710 109.685 107.755 ;
        RECT 103.400 107.570 109.685 107.710 ;
        RECT 103.400 107.510 103.720 107.570 ;
        RECT 109.395 107.525 109.685 107.570 ;
        RECT 25.680 107.230 31.385 107.370 ;
        RECT 25.680 107.185 25.970 107.230 ;
        RECT 27.515 107.185 27.805 107.230 ;
        RECT 31.095 107.185 31.385 107.230 ;
        RECT 17.495 107.030 18.085 107.075 ;
        RECT 20.735 107.030 21.385 107.075 ;
        RECT 21.980 107.030 22.300 107.090 ;
        RECT 32.175 107.075 32.465 107.390 ;
        RECT 37.175 107.370 37.465 107.415 ;
        RECT 39.015 107.370 39.305 107.415 ;
        RECT 44.535 107.370 44.825 107.415 ;
        RECT 34.965 107.230 44.825 107.370 ;
        RECT 17.495 106.890 22.300 107.030 ;
        RECT 17.495 106.845 17.785 106.890 ;
        RECT 20.735 106.845 21.385 106.890 ;
        RECT 21.980 106.830 22.300 106.890 ;
        RECT 28.875 107.030 29.525 107.075 ;
        RECT 32.175 107.030 32.765 107.075 ;
        RECT 28.875 106.890 32.765 107.030 ;
        RECT 28.875 106.845 29.525 106.890 ;
        RECT 32.475 106.845 32.765 106.890 ;
        RECT 27.500 106.690 27.820 106.750 ;
        RECT 34.965 106.690 35.105 107.230 ;
        RECT 37.175 107.185 37.465 107.230 ;
        RECT 39.015 107.185 39.305 107.230 ;
        RECT 44.535 107.185 44.825 107.230 ;
        RECT 35.335 106.845 35.625 107.075 ;
        RECT 27.500 106.550 35.105 106.690 ;
        RECT 35.410 106.690 35.550 106.845 ;
        RECT 37.160 106.690 37.480 106.750 ;
        RECT 35.410 106.550 37.480 106.690 ;
        RECT 44.610 106.690 44.750 107.185 ;
        RECT 44.995 107.030 45.285 107.075 ;
        RECT 46.820 107.030 47.140 107.090 ;
        RECT 48.155 107.075 48.445 107.390 ;
        RECT 49.235 107.370 49.525 107.415 ;
        RECT 52.815 107.370 53.105 107.415 ;
        RECT 54.650 107.370 54.940 107.415 ;
        RECT 49.235 107.230 54.940 107.370 ;
        RECT 49.235 107.185 49.525 107.230 ;
        RECT 52.815 107.185 53.105 107.230 ;
        RECT 54.650 107.185 54.940 107.230 ;
        RECT 56.495 107.370 56.785 107.415 ;
        RECT 57.415 107.370 57.705 107.415 ;
        RECT 56.495 107.230 57.705 107.370 ;
        RECT 56.495 107.185 56.785 107.230 ;
        RECT 57.415 107.185 57.705 107.230 ;
        RECT 57.875 107.370 58.165 107.415 ;
        RECT 65.175 107.370 65.465 107.390 ;
        RECT 57.875 107.230 65.465 107.370 ;
        RECT 57.875 107.185 58.165 107.230 ;
        RECT 44.995 106.890 47.140 107.030 ;
        RECT 44.995 106.845 45.285 106.890 ;
        RECT 46.820 106.830 47.140 106.890 ;
        RECT 47.855 107.030 48.445 107.075 ;
        RECT 48.660 107.030 48.980 107.090 ;
        RECT 51.095 107.030 51.745 107.075 ;
        RECT 47.855 106.890 51.745 107.030 ;
        RECT 47.855 106.845 48.145 106.890 ;
        RECT 48.660 106.830 48.980 106.890 ;
        RECT 51.095 106.845 51.745 106.890 ;
        RECT 50.040 106.690 50.360 106.750 ;
        RECT 56.570 106.690 56.710 107.185 ;
        RECT 59.240 107.030 59.560 107.090 ;
        RECT 65.175 107.075 65.465 107.230 ;
        RECT 66.255 107.370 66.545 107.415 ;
        RECT 69.835 107.370 70.125 107.415 ;
        RECT 71.670 107.370 71.960 107.415 ;
        RECT 66.255 107.230 71.960 107.370 ;
        RECT 66.255 107.185 66.545 107.230 ;
        RECT 69.835 107.185 70.125 107.230 ;
        RECT 71.670 107.185 71.960 107.230 ;
        RECT 62.015 107.030 62.305 107.075 ;
        RECT 59.240 106.890 62.305 107.030 ;
        RECT 59.240 106.830 59.560 106.890 ;
        RECT 62.015 106.845 62.305 106.890 ;
        RECT 64.875 107.030 65.465 107.075 ;
        RECT 68.115 107.030 68.765 107.075 ;
        RECT 64.875 106.890 68.765 107.030 ;
        RECT 64.875 106.845 65.165 106.890 ;
        RECT 68.115 106.845 68.765 106.890 ;
        RECT 73.515 107.030 73.805 107.075 ;
        RECT 75.800 107.030 76.120 107.090 ;
        RECT 76.675 107.075 76.965 107.390 ;
        RECT 77.755 107.370 78.045 107.415 ;
        RECT 81.335 107.370 81.625 107.415 ;
        RECT 83.170 107.370 83.460 107.415 ;
        RECT 77.755 107.230 83.460 107.370 ;
        RECT 77.755 107.185 78.045 107.230 ;
        RECT 81.335 107.185 81.625 107.230 ;
        RECT 83.170 107.185 83.460 107.230 ;
        RECT 85.015 107.370 85.305 107.415 ;
        RECT 85.920 107.370 86.240 107.430 ;
        RECT 85.015 107.230 86.240 107.370 ;
        RECT 85.015 107.185 85.305 107.230 ;
        RECT 85.920 107.170 86.240 107.230 ;
        RECT 86.395 107.370 86.685 107.415 ;
        RECT 90.935 107.370 91.225 107.390 ;
        RECT 86.395 107.230 91.225 107.370 ;
        RECT 86.395 107.185 86.685 107.230 ;
        RECT 73.515 106.890 76.120 107.030 ;
        RECT 73.515 106.845 73.805 106.890 ;
        RECT 75.800 106.830 76.120 106.890 ;
        RECT 76.375 107.030 76.965 107.075 ;
        RECT 78.560 107.030 78.880 107.090 ;
        RECT 79.615 107.030 80.265 107.075 ;
        RECT 76.375 106.890 80.265 107.030 ;
        RECT 76.375 106.845 76.665 106.890 ;
        RECT 78.560 106.830 78.880 106.890 ;
        RECT 79.615 106.845 80.265 106.890 ;
        RECT 86.840 107.030 87.160 107.090 ;
        RECT 90.935 107.075 91.225 107.230 ;
        RECT 92.015 107.370 92.305 107.415 ;
        RECT 95.595 107.370 95.885 107.415 ;
        RECT 97.430 107.370 97.720 107.415 ;
        RECT 92.015 107.230 97.720 107.370 ;
        RECT 92.015 107.185 92.305 107.230 ;
        RECT 95.595 107.185 95.885 107.230 ;
        RECT 97.430 107.185 97.720 107.230 ;
        RECT 99.740 107.370 100.030 107.415 ;
        RECT 101.575 107.370 101.865 107.415 ;
        RECT 105.155 107.370 105.445 107.415 ;
        RECT 99.740 107.230 105.445 107.370 ;
        RECT 99.740 107.185 100.030 107.230 ;
        RECT 101.575 107.185 101.865 107.230 ;
        RECT 105.155 107.185 105.445 107.230 ;
        RECT 87.775 107.030 88.065 107.075 ;
        RECT 86.840 106.890 88.065 107.030 ;
        RECT 86.840 106.830 87.160 106.890 ;
        RECT 87.775 106.845 88.065 106.890 ;
        RECT 90.635 107.030 91.225 107.075 ;
        RECT 93.875 107.030 94.525 107.075 ;
        RECT 90.635 106.890 94.525 107.030 ;
        RECT 90.635 106.845 90.925 106.890 ;
        RECT 93.875 106.845 94.525 106.890 ;
        RECT 96.960 107.030 97.280 107.090 ;
        RECT 100.655 107.030 100.945 107.075 ;
        RECT 96.960 106.890 100.945 107.030 ;
        RECT 96.960 106.830 97.280 106.890 ;
        RECT 100.655 106.845 100.945 106.890 ;
        RECT 102.935 107.030 103.585 107.075 ;
        RECT 103.860 107.030 104.180 107.090 ;
        RECT 106.235 107.075 106.525 107.390 ;
        RECT 111.695 107.370 111.985 107.415 ;
        RECT 114.900 107.370 115.220 107.430 ;
        RECT 111.695 107.230 115.220 107.370 ;
        RECT 111.695 107.185 111.985 107.230 ;
        RECT 114.900 107.170 115.220 107.230 ;
        RECT 106.235 107.030 106.825 107.075 ;
        RECT 102.935 106.890 106.825 107.030 ;
        RECT 102.935 106.845 103.585 106.890 ;
        RECT 103.860 106.830 104.180 106.890 ;
        RECT 106.535 106.845 106.825 106.890 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 44.610 106.550 56.710 106.690 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 27.500 106.490 27.820 106.550 ;
        RECT 37.160 106.490 37.480 106.550 ;
        RECT 50.040 106.490 50.360 106.550 ;
        RECT 11.330 105.870 113.450 106.350 ;
        RECT 21.980 105.470 22.300 105.730 ;
        RECT 25.200 105.670 25.520 105.730 ;
        RECT 48.660 105.670 48.980 105.730 ;
        RECT 49.595 105.670 49.885 105.715 ;
        RECT 25.200 105.530 33.710 105.670 ;
        RECT 25.200 105.470 25.520 105.530 ;
        RECT 26.235 105.330 26.525 105.375 ;
        RECT 28.420 105.330 28.740 105.390 ;
        RECT 29.475 105.330 30.125 105.375 ;
        RECT 26.235 105.190 30.125 105.330 ;
        RECT 26.235 105.145 26.825 105.190 ;
        RECT 16.920 104.990 17.240 105.050 ;
        RECT 22.455 104.990 22.745 105.035 ;
        RECT 16.920 104.850 22.745 104.990 ;
        RECT 16.920 104.790 17.240 104.850 ;
        RECT 22.455 104.805 22.745 104.850 ;
        RECT 26.535 104.830 26.825 105.145 ;
        RECT 28.420 105.130 28.740 105.190 ;
        RECT 29.475 105.145 30.125 105.190 ;
        RECT 33.570 105.035 33.710 105.530 ;
        RECT 48.660 105.530 49.885 105.670 ;
        RECT 48.660 105.470 48.980 105.530 ;
        RECT 49.595 105.485 49.885 105.530 ;
        RECT 78.115 105.670 78.405 105.715 ;
        RECT 78.560 105.670 78.880 105.730 ;
        RECT 78.115 105.530 78.880 105.670 ;
        RECT 78.115 105.485 78.405 105.530 ;
        RECT 78.560 105.470 78.880 105.530 ;
        RECT 88.695 105.670 88.985 105.715 ;
        RECT 91.900 105.670 92.220 105.730 ;
        RECT 88.695 105.530 92.220 105.670 ;
        RECT 88.695 105.485 88.985 105.530 ;
        RECT 91.900 105.470 92.220 105.530 ;
        RECT 92.910 105.530 101.790 105.670 ;
        RECT 65.220 105.130 65.540 105.390 ;
        RECT 67.515 105.330 68.165 105.375 ;
        RECT 71.115 105.330 71.405 105.375 ;
        RECT 67.515 105.190 71.405 105.330 ;
        RECT 67.515 105.145 68.165 105.190 ;
        RECT 70.815 105.145 71.405 105.190 ;
        RECT 71.660 105.330 71.980 105.390 ;
        RECT 92.910 105.330 93.050 105.530 ;
        RECT 71.660 105.190 76.030 105.330 ;
        RECT 27.615 104.990 27.905 105.035 ;
        RECT 31.195 104.990 31.485 105.035 ;
        RECT 33.030 104.990 33.320 105.035 ;
        RECT 27.615 104.850 33.320 104.990 ;
        RECT 27.615 104.805 27.905 104.850 ;
        RECT 31.195 104.805 31.485 104.850 ;
        RECT 33.030 104.805 33.320 104.850 ;
        RECT 33.495 104.990 33.785 105.035 ;
        RECT 37.620 104.990 37.940 105.050 ;
        RECT 33.495 104.850 37.940 104.990 ;
        RECT 33.495 104.805 33.785 104.850 ;
        RECT 37.620 104.790 37.940 104.850 ;
        RECT 50.040 104.790 50.360 105.050 ;
        RECT 56.940 104.990 57.260 105.050 ;
        RECT 63.855 104.990 64.145 105.035 ;
        RECT 56.940 104.850 64.145 104.990 ;
        RECT 56.940 104.790 57.260 104.850 ;
        RECT 63.855 104.805 64.145 104.850 ;
        RECT 64.320 104.990 64.610 105.035 ;
        RECT 66.155 104.990 66.445 105.035 ;
        RECT 69.735 104.990 70.025 105.035 ;
        RECT 64.320 104.850 70.025 104.990 ;
        RECT 64.320 104.805 64.610 104.850 ;
        RECT 66.155 104.805 66.445 104.850 ;
        RECT 69.735 104.805 70.025 104.850 ;
        RECT 70.815 104.990 71.105 105.145 ;
        RECT 71.660 105.130 71.980 105.190 ;
        RECT 75.890 105.035 76.030 105.190 ;
        RECT 88.310 105.190 93.050 105.330 ;
        RECT 93.275 105.330 93.925 105.375 ;
        RECT 96.875 105.330 97.165 105.375 ;
        RECT 101.115 105.330 101.405 105.375 ;
        RECT 93.275 105.190 101.405 105.330 ;
        RECT 75.355 104.990 75.645 105.035 ;
        RECT 70.815 104.850 75.645 104.990 ;
        RECT 70.815 104.830 71.105 104.850 ;
        RECT 75.355 104.805 75.645 104.850 ;
        RECT 75.815 104.990 76.105 105.035 ;
        RECT 78.575 104.990 78.865 105.035 ;
        RECT 85.920 104.990 86.240 105.050 ;
        RECT 88.310 105.035 88.450 105.190 ;
        RECT 93.275 105.145 93.925 105.190 ;
        RECT 96.575 105.145 97.165 105.190 ;
        RECT 101.115 105.145 101.405 105.190 ;
        RECT 88.235 104.990 88.525 105.035 ;
        RECT 75.815 104.850 88.525 104.990 ;
        RECT 75.815 104.805 76.105 104.850 ;
        RECT 78.575 104.805 78.865 104.850 ;
        RECT 85.920 104.790 86.240 104.850 ;
        RECT 88.235 104.805 88.525 104.850 ;
        RECT 90.080 104.990 90.370 105.035 ;
        RECT 91.915 104.990 92.205 105.035 ;
        RECT 95.495 104.990 95.785 105.035 ;
        RECT 90.080 104.850 95.785 104.990 ;
        RECT 90.080 104.805 90.370 104.850 ;
        RECT 91.915 104.805 92.205 104.850 ;
        RECT 95.495 104.805 95.785 104.850 ;
        RECT 96.575 104.830 96.865 105.145 ;
        RECT 97.880 104.990 98.200 105.050 ;
        RECT 101.650 105.035 101.790 105.530 ;
        RECT 103.860 105.470 104.180 105.730 ;
        RECT 106.160 105.470 106.480 105.730 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 99.735 104.990 100.025 105.035 ;
        RECT 97.880 104.850 100.025 104.990 ;
        RECT 97.880 104.790 98.200 104.850 ;
        RECT 99.735 104.805 100.025 104.850 ;
        RECT 101.575 104.990 101.865 105.035 ;
        RECT 104.335 104.990 104.625 105.035 ;
        RECT 105.700 104.990 106.020 105.050 ;
        RECT 101.575 104.850 106.020 104.990 ;
        RECT 101.575 104.805 101.865 104.850 ;
        RECT 104.335 104.805 104.625 104.850 ;
        RECT 105.700 104.790 106.020 104.850 ;
        RECT 23.375 104.650 23.665 104.695 ;
        RECT 26.120 104.650 26.440 104.710 ;
        RECT 23.375 104.510 26.440 104.650 ;
        RECT 23.375 104.465 23.665 104.510 ;
        RECT 26.120 104.450 26.440 104.510 ;
        RECT 70.280 104.650 70.600 104.710 ;
        RECT 73.975 104.650 74.265 104.695 ;
        RECT 70.280 104.510 74.265 104.650 ;
        RECT 70.280 104.450 70.600 104.510 ;
        RECT 73.975 104.465 74.265 104.510 ;
        RECT 89.615 104.650 89.905 104.695 ;
        RECT 99.260 104.650 99.580 104.710 ;
        RECT 89.615 104.510 99.580 104.650 ;
        RECT 89.615 104.465 89.905 104.510 ;
        RECT 99.260 104.450 99.580 104.510 ;
        RECT 27.615 104.310 27.905 104.355 ;
        RECT 30.735 104.310 31.025 104.355 ;
        RECT 32.625 104.310 32.915 104.355 ;
        RECT 27.615 104.170 32.915 104.310 ;
        RECT 27.615 104.125 27.905 104.170 ;
        RECT 30.735 104.125 31.025 104.170 ;
        RECT 32.625 104.125 32.915 104.170 ;
        RECT 64.725 104.310 65.015 104.355 ;
        RECT 66.615 104.310 66.905 104.355 ;
        RECT 69.735 104.310 70.025 104.355 ;
        RECT 64.725 104.170 70.025 104.310 ;
        RECT 64.725 104.125 65.015 104.170 ;
        RECT 66.615 104.125 66.905 104.170 ;
        RECT 69.735 104.125 70.025 104.170 ;
        RECT 90.485 104.310 90.775 104.355 ;
        RECT 92.375 104.310 92.665 104.355 ;
        RECT 95.495 104.310 95.785 104.355 ;
        RECT 90.485 104.170 95.785 104.310 ;
        RECT 90.485 104.125 90.775 104.170 ;
        RECT 92.375 104.125 92.665 104.170 ;
        RECT 95.495 104.125 95.785 104.170 ;
        RECT 27.040 103.970 27.360 104.030 ;
        RECT 32.180 103.970 32.470 104.015 ;
        RECT 27.040 103.830 32.470 103.970 ;
        RECT 27.040 103.770 27.360 103.830 ;
        RECT 32.180 103.785 32.470 103.830 ;
        RECT 90.935 103.970 91.225 104.015 ;
        RECT 96.500 103.970 96.820 104.030 ;
        RECT 90.935 103.830 96.820 103.970 ;
        RECT 90.935 103.785 91.225 103.830 ;
        RECT 96.500 103.770 96.820 103.830 ;
        RECT 11.330 103.150 113.450 103.630 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 32.510 203.845 34.390 204.215 ;
        RECT 62.510 203.845 64.390 204.215 ;
        RECT 92.510 203.845 94.390 204.215 ;
        RECT 17.510 201.125 19.390 201.495 ;
        RECT 47.510 201.125 49.390 201.495 ;
        RECT 77.510 201.125 79.390 201.495 ;
        RECT 107.510 201.125 109.390 201.495 ;
        RECT 58.350 199.620 58.610 199.940 ;
        RECT 70.770 199.620 71.030 199.940 ;
        RECT 71.690 199.620 71.950 199.940 ;
        RECT 56.510 198.940 56.770 199.260 ;
        RECT 32.510 198.405 34.390 198.775 ;
        RECT 56.570 197.900 56.710 198.940 ;
        RECT 56.510 197.580 56.770 197.900 ;
        RECT 58.410 197.810 58.550 199.620 ;
        RECT 69.390 199.280 69.650 199.600 ;
        RECT 60.190 198.940 60.450 199.260 ;
        RECT 64.790 198.940 65.050 199.260 ;
        RECT 59.270 197.810 59.530 197.900 ;
        RECT 58.410 197.670 59.530 197.810 ;
        RECT 50.070 196.900 50.330 197.220 ;
        RECT 52.830 196.900 53.090 197.220 ;
        RECT 17.510 195.685 19.390 196.055 ;
        RECT 47.510 195.685 49.390 196.055 ;
        RECT 32.510 192.965 34.390 193.335 ;
        RECT 34.890 192.140 35.150 192.460 ;
        RECT 40.410 192.140 40.670 192.460 ;
        RECT 30.290 190.780 30.550 191.100 ;
        RECT 17.510 190.245 19.390 190.615 ;
        RECT 20.630 188.740 20.890 189.060 ;
        RECT 17.510 184.805 19.390 185.175 ;
        RECT 17.510 179.365 19.390 179.735 ;
        RECT 20.690 178.520 20.830 188.740 ;
        RECT 23.850 188.400 24.110 188.720 ;
        RECT 24.310 188.400 24.570 188.720 ;
        RECT 23.910 184.640 24.050 188.400 ;
        RECT 24.370 187.360 24.510 188.400 ;
        RECT 28.450 188.060 28.710 188.380 ;
        RECT 28.510 187.360 28.650 188.060 ;
        RECT 24.310 187.040 24.570 187.360 ;
        RECT 28.450 187.040 28.710 187.360 ;
        RECT 24.770 186.360 25.030 186.680 ;
        RECT 23.850 184.320 24.110 184.640 ;
        RECT 24.830 183.620 24.970 186.360 ;
        RECT 30.350 183.960 30.490 190.780 ;
        RECT 30.750 189.420 31.010 189.740 ;
        RECT 30.810 186.000 30.950 189.420 ;
        RECT 31.210 189.080 31.470 189.400 ;
        RECT 32.130 189.080 32.390 189.400 ;
        RECT 31.270 186.340 31.410 189.080 ;
        RECT 31.210 186.020 31.470 186.340 ;
        RECT 30.750 185.680 31.010 186.000 ;
        RECT 30.290 183.640 30.550 183.960 ;
        RECT 22.930 183.300 23.190 183.620 ;
        RECT 24.770 183.300 25.030 183.620 ;
        RECT 22.990 181.920 23.130 183.300 ;
        RECT 27.070 182.960 27.330 183.280 ;
        RECT 24.770 182.620 25.030 182.940 ;
        RECT 26.610 182.620 26.870 182.940 ;
        RECT 22.930 181.600 23.190 181.920 ;
        RECT 20.630 178.430 20.890 178.520 ;
        RECT 19.770 178.290 20.890 178.430 ;
        RECT 17.510 173.925 19.390 174.295 ;
        RECT 17.510 168.485 19.390 168.855 ;
        RECT 19.770 167.300 19.910 178.290 ;
        RECT 20.630 178.200 20.890 178.290 ;
        RECT 24.830 177.840 24.970 182.620 ;
        RECT 26.670 181.580 26.810 182.620 ;
        RECT 26.610 181.260 26.870 181.580 ;
        RECT 25.230 180.580 25.490 180.900 ;
        RECT 22.010 177.520 22.270 177.840 ;
        RECT 24.770 177.520 25.030 177.840 ;
        RECT 22.070 176.480 22.210 177.520 ;
        RECT 25.290 177.500 25.430 180.580 ;
        RECT 25.230 177.180 25.490 177.500 ;
        RECT 22.010 176.160 22.270 176.480 ;
        RECT 26.610 175.710 26.870 175.800 ;
        RECT 27.130 175.710 27.270 182.960 ;
        RECT 28.910 182.620 29.170 182.940 ;
        RECT 28.970 180.220 29.110 182.620 ;
        RECT 29.370 180.920 29.630 181.240 ;
        RECT 28.910 179.900 29.170 180.220 ;
        RECT 28.970 176.480 29.110 179.900 ;
        RECT 29.430 178.860 29.570 180.920 ;
        RECT 29.830 180.240 30.090 180.560 ;
        RECT 29.370 178.540 29.630 178.860 ;
        RECT 29.370 177.180 29.630 177.500 ;
        RECT 28.910 176.160 29.170 176.480 ;
        RECT 29.430 175.880 29.570 177.180 ;
        RECT 26.610 175.570 27.270 175.710 ;
        RECT 26.610 175.480 26.870 175.570 ;
        RECT 28.450 175.480 28.710 175.800 ;
        RECT 28.970 175.740 29.570 175.880 ;
        RECT 25.690 174.460 25.950 174.780 ;
        RECT 25.750 172.400 25.890 174.460 ;
        RECT 25.690 172.080 25.950 172.400 ;
        RECT 26.670 170.360 26.810 175.480 ;
        RECT 28.510 173.420 28.650 175.480 ;
        RECT 28.450 173.100 28.710 173.420 ;
        RECT 28.970 170.360 29.110 175.740 ;
        RECT 29.890 170.360 30.030 180.240 ;
        RECT 30.350 178.520 30.490 183.640 ;
        RECT 30.810 181.580 30.950 185.680 ;
        RECT 31.270 183.620 31.410 186.020 ;
        RECT 32.190 184.300 32.330 189.080 ;
        RECT 32.510 187.525 34.390 187.895 ;
        RECT 34.430 186.700 34.690 187.020 ;
        RECT 34.490 184.300 34.630 186.700 ;
        RECT 34.950 184.640 35.090 192.140 ;
        RECT 37.650 191.460 37.910 191.780 ;
        RECT 36.270 189.080 36.530 189.400 ;
        RECT 35.350 185.400 35.610 185.660 ;
        RECT 35.350 185.340 36.010 185.400 ;
        RECT 35.410 185.260 36.010 185.340 ;
        RECT 34.890 184.320 35.150 184.640 ;
        RECT 32.130 183.980 32.390 184.300 ;
        RECT 34.430 183.980 34.690 184.300 ;
        RECT 35.870 183.960 36.010 185.260 ;
        RECT 35.810 183.640 36.070 183.960 ;
        RECT 31.210 183.300 31.470 183.620 ;
        RECT 30.750 181.260 31.010 181.580 ;
        RECT 31.270 179.200 31.410 183.300 ;
        RECT 32.130 182.620 32.390 182.940 ;
        RECT 32.190 181.920 32.330 182.620 ;
        RECT 32.510 182.085 34.390 182.455 ;
        RECT 32.130 181.600 32.390 181.920 ;
        RECT 31.210 178.880 31.470 179.200 ;
        RECT 30.750 178.540 31.010 178.860 ;
        RECT 30.290 178.200 30.550 178.520 ;
        RECT 30.290 177.180 30.550 177.500 ;
        RECT 30.350 170.700 30.490 177.180 ;
        RECT 30.810 171.040 30.950 178.540 ;
        RECT 32.190 176.480 32.330 181.600 ;
        RECT 35.870 180.900 36.010 183.640 ;
        RECT 33.970 180.580 34.230 180.900 ;
        RECT 35.810 180.580 36.070 180.900 ;
        RECT 34.030 178.860 34.170 180.580 ;
        RECT 33.970 178.540 34.230 178.860 ;
        RECT 34.030 178.180 34.170 178.540 ;
        RECT 33.970 177.860 34.230 178.180 ;
        RECT 34.030 177.500 34.170 177.860 ;
        RECT 33.970 177.180 34.230 177.500 ;
        RECT 35.350 177.355 35.610 177.500 ;
        RECT 32.510 176.645 34.390 177.015 ;
        RECT 35.340 176.985 35.620 177.355 ;
        RECT 32.130 176.160 32.390 176.480 ;
        RECT 35.870 175.460 36.010 180.580 ;
        RECT 36.330 175.800 36.470 189.080 ;
        RECT 37.710 184.640 37.850 191.460 ;
        RECT 39.490 190.780 39.750 191.100 ;
        RECT 39.550 189.400 39.690 190.780 ;
        RECT 40.470 190.080 40.610 192.140 ;
        RECT 50.130 191.780 50.270 196.900 ;
        RECT 52.890 195.520 53.030 196.900 ;
        RECT 52.830 195.200 53.090 195.520 ;
        RECT 57.890 194.180 58.150 194.500 ;
        RECT 57.950 192.800 58.090 194.180 ;
        RECT 57.890 192.480 58.150 192.800 ;
        RECT 58.410 192.120 58.550 197.670 ;
        RECT 59.270 197.580 59.530 197.670 ;
        RECT 60.250 194.840 60.390 198.940 ;
        RECT 62.510 198.405 64.390 198.775 ;
        RECT 64.850 198.240 64.990 198.940 ;
        RECT 69.450 198.240 69.590 199.280 ;
        RECT 70.310 198.940 70.570 199.260 ;
        RECT 64.790 197.920 65.050 198.240 ;
        RECT 69.390 197.920 69.650 198.240 ;
        RECT 66.170 197.240 66.430 197.560 ;
        RECT 63.410 196.900 63.670 197.220 ;
        RECT 65.250 196.900 65.510 197.220 ;
        RECT 61.110 196.220 61.370 196.540 ;
        RECT 59.730 194.520 59.990 194.840 ;
        RECT 60.190 194.520 60.450 194.840 ;
        RECT 58.350 191.800 58.610 192.120 ;
        RECT 50.070 191.460 50.330 191.780 ;
        RECT 44.090 190.780 44.350 191.100 ;
        RECT 44.150 190.080 44.290 190.780 ;
        RECT 47.510 190.245 49.390 190.615 ;
        RECT 40.410 189.760 40.670 190.080 ;
        RECT 44.090 189.760 44.350 190.080 ;
        RECT 42.250 189.420 42.510 189.740 ;
        RECT 39.490 189.080 39.750 189.400 ;
        RECT 39.030 188.060 39.290 188.380 ;
        RECT 39.090 186.680 39.230 188.060 ;
        RECT 42.310 187.360 42.450 189.420 ;
        RECT 43.170 188.740 43.430 189.060 ;
        RECT 42.710 188.060 42.970 188.380 ;
        RECT 42.250 187.040 42.510 187.360 ;
        RECT 42.770 187.020 42.910 188.060 ;
        RECT 43.230 187.360 43.370 188.740 ;
        RECT 44.090 188.400 44.350 188.720 ;
        RECT 45.010 188.400 45.270 188.720 ;
        RECT 43.170 187.040 43.430 187.360 ;
        RECT 42.710 186.700 42.970 187.020 ;
        RECT 38.570 186.360 38.830 186.680 ;
        RECT 39.030 186.360 39.290 186.680 ;
        RECT 38.630 186.000 38.770 186.360 ;
        RECT 43.170 186.020 43.430 186.340 ;
        RECT 38.570 185.680 38.830 186.000 ;
        RECT 37.650 184.320 37.910 184.640 ;
        RECT 39.030 183.300 39.290 183.620 ;
        RECT 39.090 181.920 39.230 183.300 ;
        RECT 39.030 181.600 39.290 181.920 ;
        RECT 38.110 180.580 38.370 180.900 ;
        RECT 41.790 180.580 42.050 180.900 ;
        RECT 37.190 177.860 37.450 178.180 ;
        RECT 37.250 175.800 37.390 177.860 ;
        RECT 36.270 175.480 36.530 175.800 ;
        RECT 37.190 175.480 37.450 175.800 ;
        RECT 35.810 175.140 36.070 175.460 ;
        RECT 35.350 174.460 35.610 174.780 ;
        RECT 35.410 172.740 35.550 174.460 ;
        RECT 37.250 173.420 37.390 175.480 ;
        RECT 37.190 173.100 37.450 173.420 ;
        RECT 34.890 172.420 35.150 172.740 ;
        RECT 35.350 172.420 35.610 172.740 ;
        RECT 32.130 171.740 32.390 172.060 ;
        RECT 32.190 171.040 32.330 171.740 ;
        RECT 32.510 171.205 34.390 171.575 ;
        RECT 30.750 170.720 31.010 171.040 ;
        RECT 31.670 170.720 31.930 171.040 ;
        RECT 32.130 170.720 32.390 171.040 ;
        RECT 30.290 170.380 30.550 170.700 ;
        RECT 26.610 170.040 26.870 170.360 ;
        RECT 28.910 170.040 29.170 170.360 ;
        RECT 29.830 170.040 30.090 170.360 ;
        RECT 26.150 169.020 26.410 169.340 ;
        RECT 25.230 167.320 25.490 167.640 ;
        RECT 13.730 166.980 13.990 167.300 ;
        RECT 14.190 166.980 14.450 167.300 ;
        RECT 19.710 166.980 19.970 167.300 ;
        RECT 20.170 166.980 20.430 167.300 ;
        RECT 12.810 164.260 13.070 164.580 ;
        RECT 12.870 159.480 13.010 164.260 ;
        RECT 13.790 162.880 13.930 166.980 ;
        RECT 13.730 162.560 13.990 162.880 ;
        RECT 14.250 161.860 14.390 166.980 ;
        RECT 15.110 166.640 15.370 166.960 ;
        RECT 14.650 166.300 14.910 166.620 ;
        RECT 14.710 164.920 14.850 166.300 ;
        RECT 15.170 165.600 15.310 166.640 ;
        RECT 15.110 165.280 15.370 165.600 ;
        RECT 14.650 164.600 14.910 164.920 ;
        RECT 19.770 164.580 19.910 166.980 ;
        RECT 19.710 164.260 19.970 164.580 ;
        RECT 17.510 163.045 19.390 163.415 ;
        RECT 19.770 162.280 19.910 164.260 ;
        RECT 20.230 164.240 20.370 166.980 ;
        RECT 24.310 165.280 24.570 165.600 ;
        RECT 20.170 163.920 20.430 164.240 ;
        RECT 23.390 163.580 23.650 163.900 ;
        RECT 19.310 162.140 19.910 162.280 ;
        RECT 19.310 161.860 19.450 162.140 ;
        RECT 20.170 161.880 20.430 162.200 ;
        RECT 14.190 161.540 14.450 161.860 ;
        RECT 19.250 161.540 19.510 161.860 ;
        RECT 12.810 159.160 13.070 159.480 ;
        RECT 12.870 152.880 13.010 159.160 ;
        RECT 14.250 154.040 14.390 161.540 ;
        RECT 16.950 160.860 17.210 161.180 ;
        RECT 19.710 160.860 19.970 161.180 ;
        RECT 17.010 159.820 17.150 160.860 ;
        RECT 16.950 159.500 17.210 159.820 ;
        RECT 15.110 158.820 15.370 159.140 ;
        RECT 15.170 157.440 15.310 158.820 ;
        RECT 19.770 158.460 19.910 160.860 ;
        RECT 19.710 158.140 19.970 158.460 ;
        RECT 17.510 157.605 19.390 157.975 ;
        RECT 15.110 157.120 15.370 157.440 ;
        RECT 19.770 157.100 19.910 158.140 ;
        RECT 19.710 156.780 19.970 157.100 ;
        RECT 20.230 156.760 20.370 161.880 ;
        RECT 22.470 161.200 22.730 161.520 ;
        RECT 22.530 157.440 22.670 161.200 ;
        RECT 23.450 159.480 23.590 163.580 ;
        RECT 24.370 161.860 24.510 165.280 ;
        RECT 25.290 164.920 25.430 167.320 ;
        RECT 24.770 164.600 25.030 164.920 ;
        RECT 25.230 164.600 25.490 164.920 ;
        RECT 24.830 162.880 24.970 164.600 ;
        RECT 24.770 162.560 25.030 162.880 ;
        RECT 25.290 161.860 25.430 164.600 ;
        RECT 25.690 163.920 25.950 164.240 ;
        RECT 25.750 162.200 25.890 163.920 ;
        RECT 25.690 161.880 25.950 162.200 ;
        RECT 24.310 161.540 24.570 161.860 ;
        RECT 25.230 161.540 25.490 161.860 ;
        RECT 24.310 160.860 24.570 161.180 ;
        RECT 24.370 160.160 24.510 160.860 ;
        RECT 24.310 159.840 24.570 160.160 ;
        RECT 25.290 159.820 25.430 161.540 ;
        RECT 25.230 159.500 25.490 159.820 ;
        RECT 23.390 159.160 23.650 159.480 ;
        RECT 22.470 157.120 22.730 157.440 ;
        RECT 22.930 156.780 23.190 157.100 ;
        RECT 18.330 156.440 18.590 156.760 ;
        RECT 20.170 156.440 20.430 156.760 ;
        RECT 17.870 155.420 18.130 155.740 ;
        RECT 17.930 154.720 18.070 155.420 ;
        RECT 17.870 154.400 18.130 154.720 ;
        RECT 18.390 154.380 18.530 156.440 ;
        RECT 18.330 154.060 18.590 154.380 ;
        RECT 14.190 153.720 14.450 154.040 ;
        RECT 12.870 152.740 13.470 152.880 ;
        RECT 13.330 150.980 13.470 152.740 ;
        RECT 13.270 150.660 13.530 150.980 ;
        RECT 13.330 148.600 13.470 150.660 ;
        RECT 13.270 148.280 13.530 148.600 ;
        RECT 14.250 145.540 14.390 153.720 ;
        RECT 20.230 153.700 20.370 156.440 ;
        RECT 21.550 154.400 21.810 154.720 ;
        RECT 21.090 153.720 21.350 154.040 ;
        RECT 20.170 153.380 20.430 153.700 ;
        RECT 14.650 152.700 14.910 153.020 ;
        RECT 15.570 152.700 15.830 153.020 ;
        RECT 14.710 150.300 14.850 152.700 ;
        RECT 15.630 151.320 15.770 152.700 ;
        RECT 17.510 152.165 19.390 152.535 ;
        RECT 15.570 151.000 15.830 151.320 ;
        RECT 14.650 149.980 14.910 150.300 ;
        RECT 14.650 148.960 14.910 149.280 ;
        RECT 14.710 146.560 14.850 148.960 ;
        RECT 15.110 147.940 15.370 148.260 ;
        RECT 15.170 146.560 15.310 147.940 ;
        RECT 20.230 147.920 20.370 153.380 ;
        RECT 21.150 151.320 21.290 153.720 ;
        RECT 21.610 152.000 21.750 154.400 ;
        RECT 21.550 151.680 21.810 152.000 ;
        RECT 21.090 151.000 21.350 151.320 ;
        RECT 21.150 149.280 21.290 151.000 ;
        RECT 22.470 149.980 22.730 150.300 ;
        RECT 21.090 148.960 21.350 149.280 ;
        RECT 20.170 147.600 20.430 147.920 ;
        RECT 17.510 146.725 19.390 147.095 ;
        RECT 14.650 146.240 14.910 146.560 ;
        RECT 15.110 146.240 15.370 146.560 ;
        RECT 20.230 146.220 20.370 147.600 ;
        RECT 20.170 145.900 20.430 146.220 ;
        RECT 21.150 145.880 21.290 148.960 ;
        RECT 22.530 146.560 22.670 149.980 ;
        RECT 22.470 146.240 22.730 146.560 ;
        RECT 21.090 145.560 21.350 145.880 ;
        RECT 14.190 145.220 14.450 145.540 ;
        RECT 17.510 141.285 19.390 141.655 ;
        RECT 21.550 140.120 21.810 140.440 ;
        RECT 21.090 139.780 21.350 140.100 ;
        RECT 17.870 139.100 18.130 139.420 ;
        RECT 17.930 138.060 18.070 139.100 ;
        RECT 21.150 138.400 21.290 139.780 ;
        RECT 21.090 138.080 21.350 138.400 ;
        RECT 17.870 137.740 18.130 138.060 ;
        RECT 20.630 137.060 20.890 137.380 ;
        RECT 19.710 136.380 19.970 136.700 ;
        RECT 17.510 135.845 19.390 136.215 ;
        RECT 19.770 134.660 19.910 136.380 ;
        RECT 20.690 135.680 20.830 137.060 ;
        RECT 20.630 135.360 20.890 135.680 ;
        RECT 21.150 135.000 21.290 138.080 ;
        RECT 21.090 134.680 21.350 135.000 ;
        RECT 18.330 134.340 18.590 134.660 ;
        RECT 19.710 134.340 19.970 134.660 ;
        RECT 21.610 134.400 21.750 140.120 ;
        RECT 22.470 139.440 22.730 139.760 ;
        RECT 22.010 139.100 22.270 139.420 ;
        RECT 22.070 134.660 22.210 139.100 ;
        RECT 22.530 138.400 22.670 139.440 ;
        RECT 22.470 138.080 22.730 138.400 ;
        RECT 16.490 132.300 16.750 132.620 ;
        RECT 16.030 131.620 16.290 131.940 ;
        RECT 16.090 127.520 16.230 131.620 ;
        RECT 16.550 130.240 16.690 132.300 ;
        RECT 18.390 131.940 18.530 134.340 ;
        RECT 20.690 134.320 21.750 134.400 ;
        RECT 22.010 134.340 22.270 134.660 ;
        RECT 20.630 134.260 21.750 134.320 ;
        RECT 20.630 134.000 20.890 134.260 ;
        RECT 19.710 133.660 19.970 133.980 ;
        RECT 18.330 131.620 18.590 131.940 ;
        RECT 17.510 130.405 19.390 130.775 ;
        RECT 16.490 129.920 16.750 130.240 ;
        RECT 19.770 129.220 19.910 133.660 ;
        RECT 20.170 131.620 20.430 131.940 ;
        RECT 20.230 130.240 20.370 131.620 ;
        RECT 20.170 129.920 20.430 130.240 ;
        RECT 20.170 129.240 20.430 129.560 ;
        RECT 19.710 128.900 19.970 129.220 ;
        RECT 20.230 128.280 20.370 129.240 ;
        RECT 19.770 128.140 20.370 128.280 ;
        RECT 16.030 127.200 16.290 127.520 ;
        RECT 19.770 126.840 19.910 128.140 ;
        RECT 20.690 127.600 20.830 134.000 ;
        RECT 22.470 131.960 22.730 132.280 ;
        RECT 22.010 129.640 22.270 129.900 ;
        RECT 22.530 129.640 22.670 131.960 ;
        RECT 22.010 129.580 22.670 129.640 ;
        RECT 22.070 129.500 22.670 129.580 ;
        RECT 20.230 127.460 20.830 127.600 ;
        RECT 19.710 126.520 19.970 126.840 ;
        RECT 13.730 125.500 13.990 125.820 ;
        RECT 14.650 125.500 14.910 125.820 ;
        RECT 13.790 121.740 13.930 125.500 ;
        RECT 14.710 123.440 14.850 125.500 ;
        RECT 17.510 124.965 19.390 125.335 ;
        RECT 19.770 124.800 19.910 126.520 ;
        RECT 20.230 126.500 20.370 127.460 ;
        RECT 22.530 126.840 22.670 129.500 ;
        RECT 22.470 126.520 22.730 126.840 ;
        RECT 20.170 126.180 20.430 126.500 ;
        RECT 21.090 126.180 21.350 126.500 ;
        RECT 19.710 124.480 19.970 124.800 ;
        RECT 14.650 123.120 14.910 123.440 ;
        RECT 13.730 121.420 13.990 121.740 ;
        RECT 16.490 120.740 16.750 121.060 ;
        RECT 9.590 117.680 9.850 118.000 ;
        RECT 13.730 117.680 13.990 118.000 ;
        RECT 9.650 92.720 9.790 117.680 ;
        RECT 13.790 108.480 13.930 117.680 ;
        RECT 16.550 116.640 16.690 120.740 ;
        RECT 17.510 119.525 19.390 119.895 ;
        RECT 19.770 116.640 19.910 124.480 ;
        RECT 16.490 116.320 16.750 116.640 ;
        RECT 19.710 116.320 19.970 116.640 ;
        RECT 20.230 115.620 20.370 126.180 ;
        RECT 20.630 125.500 20.890 125.820 ;
        RECT 20.690 124.120 20.830 125.500 ;
        RECT 20.630 123.800 20.890 124.120 ;
        RECT 21.150 120.380 21.290 126.180 ;
        RECT 22.530 125.820 22.670 126.520 ;
        RECT 22.470 125.500 22.730 125.820 ;
        RECT 21.090 120.060 21.350 120.380 ;
        RECT 21.150 116.300 21.290 120.060 ;
        RECT 21.550 118.360 21.810 118.680 ;
        RECT 21.090 115.980 21.350 116.300 ;
        RECT 20.170 115.300 20.430 115.620 ;
        RECT 17.510 114.085 19.390 114.455 ;
        RECT 14.190 112.240 14.450 112.560 ;
        RECT 19.250 112.240 19.510 112.560 ;
        RECT 13.730 108.160 13.990 108.480 ;
        RECT 9.580 90.720 9.860 92.720 ;
        RECT 14.250 92.240 14.390 112.240 ;
        RECT 19.310 111.200 19.450 112.240 ;
        RECT 21.610 111.200 21.750 118.360 ;
        RECT 19.250 110.880 19.510 111.200 ;
        RECT 21.550 110.880 21.810 111.200 ;
        RECT 22.990 110.520 23.130 156.780 ;
        RECT 24.770 155.760 25.030 156.080 ;
        RECT 24.310 155.420 24.570 155.740 ;
        RECT 23.850 152.700 24.110 153.020 ;
        RECT 23.910 150.640 24.050 152.700 ;
        RECT 23.850 150.320 24.110 150.640 ;
        RECT 23.850 147.260 24.110 147.580 ;
        RECT 23.390 112.240 23.650 112.560 ;
        RECT 23.450 111.200 23.590 112.240 ;
        RECT 23.390 110.880 23.650 111.200 ;
        RECT 23.910 110.860 24.050 147.260 ;
        RECT 23.850 110.540 24.110 110.860 ;
        RECT 24.370 110.520 24.510 155.420 ;
        RECT 24.830 154.040 24.970 155.760 ;
        RECT 24.770 153.720 25.030 154.040 ;
        RECT 25.230 152.700 25.490 153.020 ;
        RECT 25.290 148.600 25.430 152.700 ;
        RECT 25.230 148.280 25.490 148.600 ;
        RECT 26.210 148.260 26.350 169.020 ;
        RECT 26.670 156.080 26.810 170.040 ;
        RECT 30.810 170.020 30.950 170.720 ;
        RECT 31.730 170.440 31.870 170.720 ;
        RECT 31.730 170.360 32.330 170.440 ;
        RECT 31.730 170.300 32.390 170.360 ;
        RECT 32.130 170.040 32.390 170.300 ;
        RECT 30.750 169.700 31.010 170.020 ;
        RECT 29.830 169.020 30.090 169.340 ;
        RECT 30.750 169.020 31.010 169.340 ;
        RECT 31.670 169.020 31.930 169.340 ;
        RECT 27.070 166.640 27.330 166.960 ;
        RECT 27.130 165.600 27.270 166.640 ;
        RECT 27.070 165.280 27.330 165.600 ;
        RECT 29.370 164.600 29.630 164.920 ;
        RECT 27.530 164.260 27.790 164.580 ;
        RECT 27.590 162.280 27.730 164.260 ;
        RECT 27.590 162.200 28.190 162.280 ;
        RECT 27.590 162.140 28.250 162.200 ;
        RECT 27.590 160.160 27.730 162.140 ;
        RECT 27.990 161.880 28.250 162.140 ;
        RECT 27.530 159.840 27.790 160.160 ;
        RECT 29.430 159.730 29.570 164.600 ;
        RECT 29.890 161.430 30.030 169.020 ;
        RECT 30.290 161.430 30.550 161.520 ;
        RECT 29.890 161.290 30.550 161.430 ;
        RECT 30.290 161.200 30.550 161.290 ;
        RECT 28.970 159.590 29.570 159.730 ;
        RECT 28.450 159.160 28.710 159.480 ;
        RECT 27.070 157.120 27.330 157.440 ;
        RECT 26.610 155.760 26.870 156.080 ;
        RECT 27.130 152.000 27.270 157.120 ;
        RECT 28.510 156.955 28.650 159.160 ;
        RECT 28.440 156.585 28.720 156.955 ;
        RECT 28.510 154.040 28.650 156.585 ;
        RECT 28.970 156.420 29.110 159.590 ;
        RECT 29.830 159.160 30.090 159.480 ;
        RECT 30.290 159.160 30.550 159.480 ;
        RECT 29.370 156.440 29.630 156.760 ;
        RECT 28.910 156.275 29.170 156.420 ;
        RECT 28.900 155.905 29.180 156.275 ;
        RECT 29.430 155.480 29.570 156.440 ;
        RECT 28.970 155.340 29.570 155.480 ;
        RECT 28.450 153.720 28.710 154.040 ;
        RECT 28.450 153.040 28.710 153.360 ;
        RECT 27.070 151.680 27.330 152.000 ;
        RECT 27.130 148.600 27.270 151.680 ;
        RECT 28.510 150.300 28.650 153.040 ;
        RECT 28.450 149.980 28.710 150.300 ;
        RECT 28.510 149.280 28.650 149.980 ;
        RECT 28.450 148.960 28.710 149.280 ;
        RECT 27.070 148.280 27.330 148.600 ;
        RECT 26.150 147.940 26.410 148.260 ;
        RECT 26.150 147.260 26.410 147.580 ;
        RECT 27.530 147.260 27.790 147.580 ;
        RECT 26.210 141.120 26.350 147.260 ;
        RECT 27.590 145.880 27.730 147.260 ;
        RECT 27.530 145.560 27.790 145.880 ;
        RECT 27.990 141.820 28.250 142.140 ;
        RECT 26.150 140.800 26.410 141.120 ;
        RECT 25.230 140.460 25.490 140.780 ;
        RECT 25.290 140.100 25.430 140.460 ;
        RECT 25.230 139.780 25.490 140.100 ;
        RECT 24.770 139.100 25.030 139.420 ;
        RECT 24.830 138.060 24.970 139.100 ;
        RECT 24.770 137.740 25.030 138.060 ;
        RECT 24.770 137.060 25.030 137.380 ;
        RECT 24.830 131.940 24.970 137.060 ;
        RECT 25.290 132.620 25.430 139.780 ;
        RECT 25.230 132.300 25.490 132.620 ;
        RECT 27.070 131.960 27.330 132.280 ;
        RECT 24.770 131.620 25.030 131.940 ;
        RECT 24.830 129.220 24.970 131.620 ;
        RECT 26.150 130.940 26.410 131.260 ;
        RECT 25.230 129.580 25.490 129.900 ;
        RECT 24.770 128.900 25.030 129.220 ;
        RECT 24.830 127.520 24.970 128.900 ;
        RECT 24.770 127.200 25.030 127.520 ;
        RECT 24.830 123.440 24.970 127.200 ;
        RECT 25.290 126.920 25.430 129.580 ;
        RECT 25.690 128.900 25.950 129.220 ;
        RECT 25.750 127.520 25.890 128.900 ;
        RECT 25.690 127.200 25.950 127.520 ;
        RECT 25.290 126.780 25.890 126.920 ;
        RECT 26.210 126.840 26.350 130.940 ;
        RECT 26.610 128.220 26.870 128.540 ;
        RECT 26.670 127.520 26.810 128.220 ;
        RECT 26.610 127.200 26.870 127.520 ;
        RECT 24.770 123.120 25.030 123.440 ;
        RECT 24.830 121.060 24.970 123.120 ;
        RECT 24.770 120.740 25.030 121.060 ;
        RECT 25.230 120.740 25.490 121.060 ;
        RECT 24.830 118.340 24.970 120.740 ;
        RECT 24.770 118.020 25.030 118.340 ;
        RECT 24.830 112.810 24.970 118.020 ;
        RECT 25.290 117.660 25.430 120.740 ;
        RECT 25.750 118.340 25.890 126.780 ;
        RECT 26.150 126.520 26.410 126.840 ;
        RECT 25.690 118.020 25.950 118.340 ;
        RECT 27.130 118.000 27.270 131.960 ;
        RECT 27.530 128.220 27.790 128.540 ;
        RECT 27.590 125.820 27.730 128.220 ;
        RECT 27.530 125.500 27.790 125.820 ;
        RECT 27.070 117.680 27.330 118.000 ;
        RECT 25.230 117.340 25.490 117.660 ;
        RECT 25.230 112.810 25.490 112.900 ;
        RECT 24.830 112.670 25.490 112.810 ;
        RECT 25.230 112.580 25.490 112.670 ;
        RECT 27.070 112.580 27.330 112.900 ;
        RECT 16.950 110.200 17.210 110.520 ;
        RECT 22.930 110.200 23.190 110.520 ;
        RECT 24.310 110.200 24.570 110.520 ;
        RECT 17.010 107.460 17.150 110.200 ;
        RECT 23.390 109.180 23.650 109.500 ;
        RECT 17.510 108.645 19.390 109.015 ;
        RECT 23.450 107.800 23.590 109.180 ;
        RECT 20.630 107.480 20.890 107.800 ;
        RECT 23.390 107.480 23.650 107.800 ;
        RECT 16.950 107.140 17.210 107.460 ;
        RECT 17.010 105.080 17.150 107.140 ;
        RECT 16.950 104.760 17.210 105.080 ;
        RECT 17.510 103.205 19.390 103.575 ;
        RECT 20.690 92.720 20.830 107.480 ;
        RECT 25.290 107.460 25.430 112.580 ;
        RECT 27.130 110.180 27.270 112.580 ;
        RECT 28.050 110.520 28.190 141.820 ;
        RECT 28.450 139.780 28.710 140.100 ;
        RECT 28.510 138.400 28.650 139.780 ;
        RECT 28.450 138.080 28.710 138.400 ;
        RECT 28.510 134.660 28.650 138.080 ;
        RECT 28.450 134.340 28.710 134.660 ;
        RECT 28.970 130.240 29.110 155.340 ;
        RECT 29.890 154.235 30.030 159.160 ;
        RECT 29.820 153.865 30.100 154.235 ;
        RECT 30.350 154.040 30.490 159.160 ;
        RECT 29.830 153.720 30.090 153.865 ;
        RECT 30.290 153.720 30.550 154.040 ;
        RECT 30.350 153.440 30.490 153.720 ;
        RECT 29.890 153.300 30.490 153.440 ;
        RECT 29.890 153.020 30.030 153.300 ;
        RECT 29.830 152.700 30.090 153.020 ;
        RECT 30.290 152.700 30.550 153.020 ;
        RECT 29.370 149.980 29.630 150.300 ;
        RECT 29.430 146.560 29.570 149.980 ;
        RECT 29.370 146.240 29.630 146.560 ;
        RECT 30.350 143.160 30.490 152.700 ;
        RECT 30.810 143.160 30.950 169.020 ;
        RECT 31.210 166.640 31.470 166.960 ;
        RECT 31.270 156.420 31.410 166.640 ;
        RECT 31.730 156.420 31.870 169.020 ;
        RECT 32.590 166.870 32.850 166.960 ;
        RECT 32.190 166.730 32.850 166.870 ;
        RECT 32.190 158.800 32.330 166.730 ;
        RECT 32.590 166.640 32.850 166.730 ;
        RECT 34.950 166.620 35.090 172.420 ;
        RECT 38.170 170.440 38.310 180.580 ;
        RECT 40.410 178.880 40.670 179.200 ;
        RECT 38.570 177.520 38.830 177.840 ;
        RECT 39.030 177.520 39.290 177.840 ;
        RECT 38.630 176.140 38.770 177.520 ;
        RECT 38.570 175.820 38.830 176.140 ;
        RECT 38.630 172.740 38.770 175.820 ;
        RECT 39.090 175.460 39.230 177.520 ;
        RECT 39.490 177.355 39.750 177.500 ;
        RECT 39.480 176.985 39.760 177.355 ;
        RECT 39.030 175.140 39.290 175.460 ;
        RECT 39.090 173.080 39.230 175.140 ;
        RECT 39.950 174.460 40.210 174.780 ;
        RECT 39.030 172.990 39.290 173.080 ;
        RECT 39.030 172.850 39.690 172.990 ;
        RECT 39.030 172.760 39.290 172.850 ;
        RECT 38.570 172.420 38.830 172.740 ;
        RECT 38.630 171.040 38.770 172.420 ;
        RECT 38.570 170.720 38.830 171.040 ;
        RECT 38.170 170.300 38.770 170.440 ;
        RECT 39.550 170.360 39.690 172.850 ;
        RECT 38.110 169.700 38.370 170.020 ;
        RECT 38.170 169.340 38.310 169.700 ;
        RECT 38.110 169.020 38.370 169.340 ;
        RECT 36.270 167.320 36.530 167.640 ;
        RECT 34.890 166.300 35.150 166.620 ;
        RECT 32.510 165.765 34.390 166.135 ;
        RECT 34.950 165.600 35.090 166.300 ;
        RECT 34.890 165.280 35.150 165.600 ;
        RECT 35.350 164.940 35.610 165.260 ;
        RECT 34.890 161.200 35.150 161.520 ;
        RECT 32.510 160.325 34.390 160.695 ;
        RECT 34.950 159.820 35.090 161.200 ;
        RECT 34.890 159.500 35.150 159.820 ;
        RECT 33.050 159.160 33.310 159.480 ;
        RECT 32.130 158.480 32.390 158.800 ;
        RECT 32.130 157.120 32.390 157.440 ;
        RECT 32.580 157.265 32.860 157.635 ;
        RECT 31.210 156.100 31.470 156.420 ;
        RECT 31.670 156.100 31.930 156.420 ;
        RECT 31.670 155.420 31.930 155.740 ;
        RECT 31.730 154.040 31.870 155.420 ;
        RECT 31.210 153.720 31.470 154.040 ;
        RECT 31.670 153.720 31.930 154.040 ;
        RECT 31.270 150.835 31.410 153.720 ;
        RECT 31.730 153.555 31.870 153.720 ;
        RECT 31.660 153.185 31.940 153.555 ;
        RECT 31.670 151.680 31.930 152.000 ;
        RECT 31.730 151.320 31.870 151.680 ;
        RECT 31.670 151.000 31.930 151.320 ;
        RECT 31.200 150.465 31.480 150.835 ;
        RECT 31.210 148.960 31.470 149.280 ;
        RECT 31.270 145.880 31.410 148.960 ;
        RECT 31.210 145.560 31.470 145.880 ;
        RECT 30.290 142.840 30.550 143.160 ;
        RECT 30.750 142.840 31.010 143.160 ;
        RECT 30.290 141.820 30.550 142.140 ;
        RECT 30.350 141.120 30.490 141.820 ;
        RECT 30.290 140.800 30.550 141.120 ;
        RECT 31.210 139.780 31.470 140.100 ;
        RECT 31.270 137.720 31.410 139.780 ;
        RECT 32.190 138.400 32.330 157.120 ;
        RECT 32.650 156.760 32.790 157.265 ;
        RECT 32.590 156.440 32.850 156.760 ;
        RECT 33.110 155.740 33.250 159.160 ;
        RECT 34.890 158.480 35.150 158.800 ;
        RECT 33.050 155.420 33.310 155.740 ;
        RECT 32.510 154.885 34.390 155.255 ;
        RECT 33.500 153.865 33.780 154.235 ;
        RECT 34.950 154.040 35.090 158.480 ;
        RECT 35.410 154.720 35.550 164.940 ;
        RECT 36.330 162.880 36.470 167.320 ;
        RECT 38.170 167.300 38.310 169.020 ;
        RECT 38.110 166.980 38.370 167.300 ;
        RECT 36.270 162.560 36.530 162.880 ;
        RECT 35.810 162.220 36.070 162.540 ;
        RECT 35.870 159.140 36.010 162.220 ;
        RECT 35.810 158.820 36.070 159.140 ;
        RECT 35.810 155.420 36.070 155.740 ;
        RECT 35.350 154.400 35.610 154.720 ;
        RECT 32.590 153.040 32.850 153.360 ;
        RECT 33.040 153.185 33.320 153.555 ;
        RECT 32.650 150.980 32.790 153.040 ;
        RECT 33.110 151.660 33.250 153.185 ;
        RECT 33.050 151.340 33.310 151.660 ;
        RECT 33.570 150.980 33.710 153.865 ;
        RECT 33.970 153.720 34.230 154.040 ;
        RECT 34.890 153.720 35.150 154.040 ;
        RECT 34.030 153.360 34.170 153.720 ;
        RECT 33.970 153.040 34.230 153.360 ;
        RECT 34.890 151.680 35.150 152.000 ;
        RECT 32.590 150.660 32.850 150.980 ;
        RECT 33.510 150.660 33.770 150.980 ;
        RECT 33.970 150.835 34.230 150.980 ;
        RECT 33.960 150.465 34.240 150.835 ;
        RECT 32.510 149.445 34.390 149.815 ;
        RECT 33.970 148.960 34.230 149.280 ;
        RECT 34.030 148.680 34.170 148.960 ;
        RECT 34.950 148.680 35.090 151.680 ;
        RECT 35.870 150.640 36.010 155.420 ;
        RECT 36.330 154.040 36.470 162.560 ;
        RECT 37.650 160.860 37.910 161.180 ;
        RECT 37.710 159.820 37.850 160.860 ;
        RECT 37.650 159.500 37.910 159.820 ;
        RECT 38.110 159.160 38.370 159.480 ;
        RECT 37.640 158.625 37.920 158.995 ;
        RECT 37.190 158.140 37.450 158.460 ;
        RECT 37.250 156.420 37.390 158.140 ;
        RECT 37.190 156.100 37.450 156.420 ;
        RECT 37.710 156.080 37.850 158.625 ;
        RECT 37.650 155.760 37.910 156.080 ;
        RECT 38.170 154.040 38.310 159.160 ;
        RECT 38.630 156.760 38.770 170.300 ;
        RECT 39.490 170.040 39.750 170.360 ;
        RECT 39.030 166.640 39.290 166.960 ;
        RECT 39.090 164.580 39.230 166.640 ;
        RECT 39.030 164.260 39.290 164.580 ;
        RECT 39.090 162.200 39.230 164.260 ;
        RECT 39.490 162.220 39.750 162.540 ;
        RECT 39.030 161.880 39.290 162.200 ;
        RECT 39.090 159.140 39.230 161.880 ;
        RECT 39.030 158.820 39.290 159.140 ;
        RECT 39.550 157.440 39.690 162.220 ;
        RECT 39.490 157.120 39.750 157.440 ;
        RECT 38.570 156.440 38.830 156.760 ;
        RECT 39.030 156.440 39.290 156.760 ;
        RECT 38.570 154.400 38.830 154.720 ;
        RECT 38.630 154.040 38.770 154.400 ;
        RECT 36.270 153.720 36.530 154.040 ;
        RECT 38.110 153.720 38.370 154.040 ;
        RECT 38.570 153.720 38.830 154.040 ;
        RECT 37.190 152.700 37.450 153.020 ;
        RECT 35.810 150.320 36.070 150.640 ;
        RECT 35.350 149.980 35.610 150.300 ;
        RECT 36.270 149.980 36.530 150.300 ;
        RECT 34.030 148.540 35.090 148.680 ;
        RECT 32.590 147.940 32.850 148.260 ;
        RECT 32.650 144.860 32.790 147.940 ;
        RECT 32.590 144.540 32.850 144.860 ;
        RECT 32.510 144.005 34.390 144.375 ;
        RECT 32.510 138.565 34.390 138.935 ;
        RECT 32.130 138.080 32.390 138.400 ;
        RECT 35.410 137.720 35.550 149.980 ;
        RECT 36.330 148.940 36.470 149.980 ;
        RECT 36.270 148.620 36.530 148.940 ;
        RECT 35.810 140.800 36.070 141.120 ;
        RECT 30.750 137.400 31.010 137.720 ;
        RECT 31.210 137.400 31.470 137.720 ;
        RECT 35.350 137.400 35.610 137.720 ;
        RECT 30.810 135.680 30.950 137.400 ;
        RECT 30.750 135.360 31.010 135.680 ;
        RECT 29.830 130.940 30.090 131.260 ;
        RECT 28.910 129.920 29.170 130.240 ;
        RECT 28.910 128.560 29.170 128.880 ;
        RECT 28.970 127.180 29.110 128.560 ;
        RECT 28.910 126.860 29.170 127.180 ;
        RECT 29.890 126.840 30.030 130.940 ;
        RECT 31.270 129.560 31.410 137.400 ;
        RECT 35.350 136.380 35.610 136.700 ;
        RECT 35.410 135.680 35.550 136.380 ;
        RECT 35.350 135.360 35.610 135.680 ;
        RECT 32.130 134.680 32.390 135.000 ;
        RECT 32.190 131.940 32.330 134.680 ;
        RECT 35.350 134.340 35.610 134.660 ;
        RECT 34.890 134.000 35.150 134.320 ;
        RECT 32.510 133.125 34.390 133.495 ;
        RECT 34.950 132.960 35.090 134.000 ;
        RECT 34.890 132.640 35.150 132.960 ;
        RECT 31.670 131.620 31.930 131.940 ;
        RECT 32.130 131.620 32.390 131.940 ;
        RECT 31.210 129.240 31.470 129.560 ;
        RECT 31.730 127.180 31.870 131.620 ;
        RECT 32.190 129.900 32.330 131.620 ;
        RECT 34.950 130.240 35.090 132.640 ;
        RECT 35.410 132.280 35.550 134.340 ;
        RECT 35.350 131.960 35.610 132.280 ;
        RECT 35.870 131.940 36.010 140.800 ;
        RECT 36.270 136.720 36.530 137.040 ;
        RECT 35.810 131.620 36.070 131.940 ;
        RECT 35.350 130.940 35.610 131.260 ;
        RECT 34.890 129.920 35.150 130.240 ;
        RECT 32.130 129.580 32.390 129.900 ;
        RECT 31.670 126.860 31.930 127.180 ;
        RECT 32.190 126.920 32.330 129.580 ;
        RECT 34.890 128.560 35.150 128.880 ;
        RECT 32.510 127.685 34.390 128.055 ;
        RECT 34.950 126.920 35.090 128.560 ;
        RECT 29.830 126.520 30.090 126.840 ;
        RECT 31.730 122.080 31.870 126.860 ;
        RECT 32.190 126.780 32.790 126.920 ;
        RECT 32.130 126.180 32.390 126.500 ;
        RECT 32.190 124.120 32.330 126.180 ;
        RECT 32.650 126.160 32.790 126.780 ;
        RECT 34.490 126.780 35.090 126.920 ;
        RECT 32.590 125.840 32.850 126.160 ;
        RECT 32.580 124.625 32.860 124.995 ;
        RECT 32.130 123.800 32.390 124.120 ;
        RECT 31.670 121.760 31.930 122.080 ;
        RECT 28.910 121.420 29.170 121.740 ;
        RECT 28.970 116.640 29.110 121.420 ;
        RECT 32.190 121.400 32.330 123.800 ;
        RECT 32.650 123.780 32.790 124.625 ;
        RECT 34.490 123.780 34.630 126.780 ;
        RECT 34.890 125.500 35.150 125.820 ;
        RECT 32.590 123.460 32.850 123.780 ;
        RECT 34.430 123.460 34.690 123.780 ;
        RECT 32.510 122.245 34.390 122.615 ;
        RECT 32.130 121.080 32.390 121.400 ;
        RECT 34.950 118.340 35.090 125.500 ;
        RECT 35.410 124.800 35.550 130.940 ;
        RECT 35.810 129.240 36.070 129.560 ;
        RECT 35.870 127.520 36.010 129.240 ;
        RECT 35.810 127.200 36.070 127.520 ;
        RECT 35.350 124.480 35.610 124.800 ;
        RECT 35.870 122.080 36.010 127.200 ;
        RECT 35.810 121.760 36.070 122.080 ;
        RECT 35.870 119.360 36.010 121.760 ;
        RECT 35.810 119.040 36.070 119.360 ;
        RECT 34.890 118.020 35.150 118.340 ;
        RECT 32.510 116.805 34.390 117.175 ;
        RECT 28.910 116.320 29.170 116.640 ;
        RECT 31.670 113.260 31.930 113.580 ;
        RECT 28.450 111.900 28.710 112.220 ;
        RECT 27.990 110.200 28.250 110.520 ;
        RECT 27.070 109.920 27.330 110.180 ;
        RECT 27.070 109.860 27.730 109.920 ;
        RECT 27.130 109.780 27.730 109.860 ;
        RECT 27.070 109.180 27.330 109.500 ;
        RECT 25.230 107.140 25.490 107.460 ;
        RECT 22.010 106.800 22.270 107.120 ;
        RECT 22.070 105.760 22.210 106.800 ;
        RECT 25.290 105.760 25.430 107.140 ;
        RECT 22.010 105.440 22.270 105.760 ;
        RECT 25.230 105.440 25.490 105.760 ;
        RECT 26.150 104.420 26.410 104.740 ;
        RECT 26.210 92.720 26.350 104.420 ;
        RECT 27.130 104.060 27.270 109.180 ;
        RECT 27.590 106.780 27.730 109.780 ;
        RECT 27.530 106.460 27.790 106.780 ;
        RECT 28.510 105.420 28.650 111.900 ;
        RECT 30.290 109.860 30.550 110.180 ;
        RECT 28.450 105.100 28.710 105.420 ;
        RECT 27.070 103.740 27.330 104.060 ;
        RECT 15.100 92.240 15.380 92.720 ;
        RECT 14.250 92.100 15.380 92.240 ;
        RECT 15.100 90.720 15.380 92.100 ;
        RECT 20.620 90.720 20.900 92.720 ;
        RECT 26.140 90.720 26.420 92.720 ;
        RECT 30.350 92.240 30.490 109.860 ;
        RECT 31.730 107.800 31.870 113.260 ;
        RECT 36.330 112.900 36.470 136.720 ;
        RECT 37.250 134.660 37.390 152.700 ;
        RECT 38.630 150.980 38.770 153.720 ;
        RECT 38.570 150.660 38.830 150.980 ;
        RECT 38.110 149.980 38.370 150.300 ;
        RECT 38.170 145.540 38.310 149.980 ;
        RECT 39.090 148.000 39.230 156.440 ;
        RECT 39.490 156.100 39.750 156.420 ;
        RECT 39.550 154.380 39.690 156.100 ;
        RECT 39.490 154.060 39.750 154.380 ;
        RECT 39.550 148.260 39.690 154.060 ;
        RECT 38.630 147.860 39.230 148.000 ;
        RECT 39.490 147.940 39.750 148.260 ;
        RECT 38.110 145.220 38.370 145.540 ;
        RECT 38.630 145.280 38.770 147.860 ;
        RECT 39.030 147.260 39.290 147.580 ;
        RECT 40.010 147.490 40.150 174.460 ;
        RECT 40.470 170.360 40.610 178.880 ;
        RECT 41.850 178.180 41.990 180.580 ;
        RECT 41.790 177.860 42.050 178.180 ;
        RECT 42.710 177.860 42.970 178.180 ;
        RECT 41.850 176.480 41.990 177.860 ;
        RECT 41.790 176.160 42.050 176.480 ;
        RECT 41.330 173.100 41.590 173.420 ;
        RECT 41.390 170.700 41.530 173.100 ;
        RECT 41.790 171.740 42.050 172.060 ;
        RECT 41.330 170.380 41.590 170.700 ;
        RECT 40.410 170.040 40.670 170.360 ;
        RECT 41.330 169.195 41.590 169.340 ;
        RECT 41.320 168.825 41.600 169.195 ;
        RECT 41.850 166.680 41.990 171.740 ;
        RECT 42.770 171.040 42.910 177.860 ;
        RECT 43.230 177.840 43.370 186.020 ;
        RECT 44.150 183.620 44.290 188.400 ;
        RECT 45.070 184.640 45.210 188.400 ;
        RECT 45.470 188.120 45.730 188.380 ;
        RECT 45.470 188.060 46.130 188.120 ;
        RECT 45.530 187.980 46.130 188.060 ;
        RECT 45.990 186.340 46.130 187.980 ;
        RECT 49.610 186.360 49.870 186.680 ;
        RECT 45.930 186.020 46.190 186.340 ;
        RECT 45.010 184.320 45.270 184.640 ;
        RECT 44.090 183.300 44.350 183.620 ;
        RECT 43.630 182.620 43.890 182.940 ;
        RECT 43.690 181.580 43.830 182.620 ;
        RECT 43.630 181.260 43.890 181.580 ;
        RECT 45.010 177.860 45.270 178.180 ;
        RECT 43.170 177.520 43.430 177.840 ;
        RECT 43.230 175.460 43.370 177.520 ;
        RECT 45.070 176.480 45.210 177.860 ;
        RECT 45.010 176.160 45.270 176.480 ;
        RECT 44.090 175.480 44.350 175.800 ;
        RECT 43.170 175.140 43.430 175.460 ;
        RECT 43.230 173.080 43.370 175.140 ;
        RECT 43.630 174.460 43.890 174.780 ;
        RECT 43.690 173.080 43.830 174.460 ;
        RECT 43.170 172.760 43.430 173.080 ;
        RECT 43.630 172.760 43.890 173.080 ;
        RECT 42.710 170.720 42.970 171.040 ;
        RECT 42.310 170.360 43.370 170.440 ;
        RECT 44.150 170.360 44.290 175.480 ;
        RECT 45.990 172.740 46.130 186.020 ;
        RECT 46.390 185.340 46.650 185.660 ;
        RECT 46.450 183.960 46.590 185.340 ;
        RECT 47.510 184.805 49.390 185.175 ;
        RECT 49.670 184.640 49.810 186.360 ;
        RECT 50.130 186.000 50.270 191.460 ;
        RECT 56.970 190.780 57.230 191.100 ;
        RECT 53.290 188.740 53.550 189.060 ;
        RECT 51.910 188.400 52.170 188.720 ;
        RECT 51.970 187.360 52.110 188.400 ;
        RECT 53.350 187.440 53.490 188.740 ;
        RECT 54.210 188.060 54.470 188.380 ;
        RECT 51.910 187.040 52.170 187.360 ;
        RECT 52.890 187.300 53.490 187.440 ;
        RECT 52.890 186.340 53.030 187.300 ;
        RECT 54.270 187.020 54.410 188.060 ;
        RECT 57.030 187.020 57.170 190.780 ;
        RECT 54.210 186.700 54.470 187.020 ;
        RECT 56.970 186.700 57.230 187.020 ;
        RECT 52.830 186.020 53.090 186.340 ;
        RECT 50.070 185.680 50.330 186.000 ;
        RECT 49.610 184.320 49.870 184.640 ;
        RECT 46.390 183.640 46.650 183.960 ;
        RECT 46.390 182.960 46.650 183.280 ;
        RECT 46.450 175.710 46.590 182.960 ;
        RECT 50.130 180.900 50.270 185.680 ;
        RECT 57.890 183.300 58.150 183.620 ;
        RECT 57.950 180.900 58.090 183.300 ;
        RECT 50.070 180.580 50.330 180.900 ;
        RECT 57.890 180.580 58.150 180.900 ;
        RECT 46.850 179.900 47.110 180.220 ;
        RECT 46.910 179.200 47.050 179.900 ;
        RECT 47.510 179.365 49.390 179.735 ;
        RECT 46.850 178.880 47.110 179.200 ;
        RECT 49.610 177.860 49.870 178.180 ;
        RECT 46.850 175.710 47.110 175.800 ;
        RECT 46.450 175.570 47.110 175.710 ;
        RECT 46.850 175.480 47.110 175.570 ;
        RECT 46.390 173.100 46.650 173.420 ;
        RECT 46.910 173.160 47.050 175.480 ;
        RECT 47.510 173.925 49.390 174.295 ;
        RECT 49.670 173.760 49.810 177.860 ;
        RECT 50.130 175.460 50.270 180.580 ;
        RECT 51.450 178.540 51.710 178.860 ;
        RECT 51.510 176.480 51.650 178.540 ;
        RECT 58.410 178.520 58.550 191.800 ;
        RECT 59.790 189.400 59.930 194.520 ;
        RECT 59.730 189.080 59.990 189.400 ;
        RECT 59.270 183.980 59.530 184.300 ;
        RECT 58.810 182.620 59.070 182.940 ;
        RECT 58.870 181.240 59.010 182.620 ;
        RECT 59.330 181.240 59.470 183.980 ;
        RECT 60.190 183.640 60.450 183.960 ;
        RECT 60.250 181.920 60.390 183.640 ;
        RECT 60.190 181.600 60.450 181.920 ;
        RECT 60.650 181.600 60.910 181.920 ;
        RECT 60.250 181.240 60.390 181.600 ;
        RECT 58.810 180.920 59.070 181.240 ;
        RECT 59.270 180.920 59.530 181.240 ;
        RECT 60.190 180.920 60.450 181.240 ;
        RECT 58.810 179.900 59.070 180.220 ;
        RECT 58.350 178.200 58.610 178.520 ;
        RECT 56.970 177.860 57.230 178.180 ;
        RECT 56.510 177.180 56.770 177.500 ;
        RECT 51.450 176.160 51.710 176.480 ;
        RECT 56.570 176.140 56.710 177.180 ;
        RECT 56.510 175.820 56.770 176.140 ;
        RECT 50.070 175.140 50.330 175.460 ;
        RECT 49.610 173.440 49.870 173.760 ;
        RECT 57.030 173.160 57.170 177.860 ;
        RECT 58.870 175.800 59.010 179.900 ;
        RECT 58.810 175.480 59.070 175.800 ;
        RECT 57.890 175.140 58.150 175.460 ;
        RECT 45.930 172.420 46.190 172.740 ;
        RECT 45.930 171.740 46.190 172.060 ;
        RECT 42.250 170.300 43.370 170.360 ;
        RECT 42.250 170.040 42.510 170.300 ;
        RECT 43.230 167.980 43.370 170.300 ;
        RECT 44.090 170.040 44.350 170.360 ;
        RECT 45.010 169.020 45.270 169.340 ;
        RECT 43.170 167.660 43.430 167.980 ;
        RECT 44.090 167.660 44.350 167.980 ;
        RECT 41.850 166.540 42.450 166.680 ;
        RECT 41.790 165.280 42.050 165.600 ;
        RECT 40.410 160.860 40.670 161.180 ;
        RECT 40.470 159.480 40.610 160.860 ;
        RECT 41.850 159.480 41.990 165.280 ;
        RECT 40.410 159.160 40.670 159.480 ;
        RECT 41.790 159.160 42.050 159.480 ;
        RECT 41.320 157.520 41.600 157.635 ;
        RECT 41.850 157.520 41.990 159.160 ;
        RECT 41.320 157.380 41.990 157.520 ;
        RECT 41.320 157.265 41.600 157.380 ;
        RECT 40.870 156.330 41.130 156.420 ;
        RECT 40.470 156.190 41.130 156.330 ;
        RECT 40.470 154.040 40.610 156.190 ;
        RECT 40.870 156.100 41.130 156.190 ;
        RECT 40.870 155.420 41.130 155.740 ;
        RECT 40.930 154.720 41.070 155.420 ;
        RECT 40.870 154.400 41.130 154.720 ;
        RECT 40.410 153.720 40.670 154.040 ;
        RECT 40.470 150.980 40.610 153.720 ;
        RECT 40.870 153.380 41.130 153.700 ;
        RECT 40.410 150.660 40.670 150.980 ;
        RECT 40.470 148.260 40.610 150.660 ;
        RECT 40.930 148.510 41.070 153.380 ;
        RECT 41.390 152.080 41.530 157.265 ;
        RECT 41.790 155.760 42.050 156.080 ;
        RECT 41.850 153.360 41.990 155.760 ;
        RECT 42.310 155.740 42.450 166.540 ;
        RECT 43.630 159.050 43.890 159.140 ;
        RECT 43.230 158.910 43.890 159.050 ;
        RECT 42.250 155.420 42.510 155.740 ;
        RECT 41.790 153.040 42.050 153.360 ;
        RECT 42.710 152.700 42.970 153.020 ;
        RECT 41.390 151.940 41.990 152.080 ;
        RECT 41.850 148.600 41.990 151.940 ;
        RECT 42.250 151.680 42.510 152.000 ;
        RECT 41.330 148.510 41.590 148.600 ;
        RECT 40.930 148.370 41.590 148.510 ;
        RECT 41.330 148.280 41.590 148.370 ;
        RECT 41.790 148.280 42.050 148.600 ;
        RECT 40.410 147.940 40.670 148.260 ;
        RECT 39.550 147.350 40.150 147.490 ;
        RECT 39.090 145.880 39.230 147.260 ;
        RECT 39.030 145.560 39.290 145.880 ;
        RECT 38.630 145.140 39.230 145.280 ;
        RECT 38.570 141.820 38.830 142.140 ;
        RECT 38.630 140.100 38.770 141.820 ;
        RECT 39.090 140.100 39.230 145.140 ;
        RECT 39.550 140.440 39.690 147.350 ;
        RECT 39.950 145.450 40.210 145.540 ;
        RECT 40.470 145.450 40.610 147.940 ;
        RECT 40.870 147.600 41.130 147.920 ;
        RECT 40.930 145.540 41.070 147.600 ;
        RECT 39.950 145.310 40.610 145.450 ;
        RECT 39.950 145.220 40.210 145.310 ;
        RECT 40.870 145.220 41.130 145.540 ;
        RECT 41.390 145.200 41.530 148.280 ;
        RECT 41.330 144.880 41.590 145.200 ;
        RECT 41.790 144.540 42.050 144.860 ;
        RECT 39.950 140.800 40.210 141.120 ;
        RECT 39.490 140.120 39.750 140.440 ;
        RECT 38.570 139.780 38.830 140.100 ;
        RECT 39.030 139.780 39.290 140.100 ;
        RECT 39.020 138.225 39.300 138.595 ;
        RECT 37.640 137.545 37.920 137.915 ;
        RECT 37.650 137.400 37.910 137.545 ;
        RECT 38.570 137.400 38.830 137.720 ;
        RECT 38.630 135.680 38.770 137.400 ;
        RECT 38.110 135.360 38.370 135.680 ;
        RECT 38.570 135.360 38.830 135.680 ;
        RECT 37.190 134.340 37.450 134.660 ;
        RECT 38.170 132.960 38.310 135.360 ;
        RECT 39.090 135.000 39.230 138.225 ;
        RECT 39.030 134.680 39.290 135.000 ;
        RECT 38.110 132.640 38.370 132.960 ;
        RECT 40.010 130.240 40.150 140.800 ;
        RECT 40.410 136.380 40.670 136.700 ;
        RECT 40.470 132.620 40.610 136.380 ;
        RECT 40.870 133.660 41.130 133.980 ;
        RECT 40.410 132.300 40.670 132.620 ;
        RECT 39.950 129.920 40.210 130.240 ;
        RECT 37.190 128.900 37.450 129.220 ;
        RECT 39.950 128.900 40.210 129.220 ;
        RECT 36.730 128.220 36.990 128.540 ;
        RECT 36.790 121.740 36.930 128.220 ;
        RECT 37.250 127.520 37.390 128.900 ;
        RECT 37.190 127.200 37.450 127.520 ;
        RECT 40.010 126.500 40.150 128.900 ;
        RECT 39.950 126.180 40.210 126.500 ;
        RECT 38.110 125.500 38.370 125.820 ;
        RECT 36.730 121.420 36.990 121.740 ;
        RECT 38.170 118.340 38.310 125.500 ;
        RECT 40.010 121.400 40.150 126.180 ;
        RECT 39.950 121.080 40.210 121.400 ;
        RECT 39.030 120.740 39.290 121.060 ;
        RECT 39.090 119.360 39.230 120.740 ;
        RECT 39.030 119.040 39.290 119.360 ;
        RECT 40.010 118.340 40.150 121.080 ;
        RECT 38.110 118.020 38.370 118.340 ;
        RECT 39.950 118.020 40.210 118.340 ;
        RECT 40.930 112.900 41.070 133.660 ;
        RECT 41.850 132.280 41.990 144.540 ;
        RECT 42.310 140.440 42.450 151.680 ;
        RECT 42.250 140.120 42.510 140.440 ;
        RECT 42.770 140.100 42.910 152.700 ;
        RECT 43.230 151.320 43.370 158.910 ;
        RECT 43.630 158.820 43.890 158.910 ;
        RECT 43.630 158.140 43.890 158.460 ;
        RECT 43.690 156.420 43.830 158.140 ;
        RECT 43.630 156.100 43.890 156.420 ;
        RECT 43.630 155.420 43.890 155.740 ;
        RECT 43.690 152.000 43.830 155.420 ;
        RECT 44.150 154.040 44.290 167.660 ;
        RECT 44.550 158.995 44.810 159.140 ;
        RECT 44.540 158.625 44.820 158.995 ;
        RECT 44.090 153.720 44.350 154.040 ;
        RECT 44.150 152.000 44.290 153.720 ;
        RECT 43.630 151.680 43.890 152.000 ;
        RECT 44.090 151.680 44.350 152.000 ;
        RECT 43.170 151.000 43.430 151.320 ;
        RECT 44.090 147.260 44.350 147.580 ;
        RECT 42.710 139.780 42.970 140.100 ;
        RECT 42.710 132.640 42.970 132.960 ;
        RECT 43.630 132.640 43.890 132.960 ;
        RECT 41.790 131.960 42.050 132.280 ;
        RECT 41.330 131.795 41.590 131.940 ;
        RECT 41.320 131.425 41.600 131.795 ;
        RECT 42.250 129.580 42.510 129.900 ;
        RECT 41.330 125.500 41.590 125.820 ;
        RECT 41.390 121.060 41.530 125.500 ;
        RECT 42.310 121.740 42.450 129.580 ;
        RECT 42.250 121.420 42.510 121.740 ;
        RECT 41.330 120.740 41.590 121.060 ;
        RECT 42.770 112.900 42.910 132.640 ;
        RECT 43.170 130.940 43.430 131.260 ;
        RECT 43.230 130.240 43.370 130.940 ;
        RECT 43.170 129.920 43.430 130.240 ;
        RECT 36.270 112.580 36.530 112.900 ;
        RECT 40.870 112.580 41.130 112.900 ;
        RECT 42.710 112.580 42.970 112.900 ;
        RECT 36.270 111.900 36.530 112.220 ;
        RECT 32.510 111.365 34.390 111.735 ;
        RECT 36.330 110.860 36.470 111.900 ;
        RECT 43.690 111.200 43.830 132.640 ;
        RECT 44.150 132.280 44.290 147.260 ;
        RECT 44.550 145.560 44.810 145.880 ;
        RECT 44.610 143.160 44.750 145.560 ;
        RECT 44.550 142.840 44.810 143.160 ;
        RECT 44.610 140.100 44.750 142.840 ;
        RECT 44.550 139.780 44.810 140.100 ;
        RECT 44.550 135.360 44.810 135.680 ;
        RECT 44.610 134.660 44.750 135.360 ;
        RECT 44.550 134.340 44.810 134.660 ;
        RECT 44.610 133.980 44.750 134.340 ;
        RECT 44.550 133.660 44.810 133.980 ;
        RECT 44.090 131.960 44.350 132.280 ;
        RECT 45.070 131.940 45.210 169.020 ;
        RECT 45.990 168.320 46.130 171.740 ;
        RECT 46.450 170.360 46.590 173.100 ;
        RECT 46.910 173.080 47.510 173.160 ;
        RECT 46.910 173.020 47.570 173.080 ;
        RECT 47.310 172.760 47.570 173.020 ;
        RECT 54.670 172.760 54.930 173.080 ;
        RECT 56.050 172.760 56.310 173.080 ;
        RECT 56.570 173.020 57.170 173.160 ;
        RECT 48.690 172.080 48.950 172.400 ;
        RECT 54.210 172.080 54.470 172.400 ;
        RECT 48.750 171.040 48.890 172.080 ;
        RECT 50.070 171.740 50.330 172.060 ;
        RECT 50.530 171.740 50.790 172.060 ;
        RECT 48.690 170.720 48.950 171.040 ;
        RECT 48.750 170.360 48.890 170.720 ;
        RECT 50.130 170.360 50.270 171.740 ;
        RECT 50.590 170.700 50.730 171.740 ;
        RECT 54.270 171.040 54.410 172.080 ;
        RECT 54.210 170.720 54.470 171.040 ;
        RECT 50.530 170.380 50.790 170.700 ;
        RECT 46.390 170.040 46.650 170.360 ;
        RECT 48.690 170.040 48.950 170.360 ;
        RECT 50.070 170.040 50.330 170.360 ;
        RECT 47.510 168.485 49.390 168.855 ;
        RECT 45.930 168.000 46.190 168.320 ;
        RECT 50.590 167.640 50.730 170.380 ;
        RECT 54.730 170.360 54.870 172.760 ;
        RECT 56.110 171.040 56.250 172.760 ;
        RECT 56.050 170.720 56.310 171.040 ;
        RECT 54.670 170.040 54.930 170.360 ;
        RECT 46.390 167.320 46.650 167.640 ;
        RECT 50.530 167.320 50.790 167.640 ;
        RECT 50.990 167.320 51.250 167.640 ;
        RECT 45.930 164.260 46.190 164.580 ;
        RECT 45.470 159.160 45.730 159.480 ;
        RECT 45.530 157.440 45.670 159.160 ;
        RECT 45.470 157.120 45.730 157.440 ;
        RECT 45.990 157.100 46.130 164.260 ;
        RECT 45.930 156.780 46.190 157.100 ;
        RECT 45.930 153.380 46.190 153.700 ;
        RECT 45.990 150.300 46.130 153.380 ;
        RECT 46.450 152.880 46.590 167.320 ;
        RECT 47.310 166.300 47.570 166.620 ;
        RECT 47.370 164.920 47.510 166.300 ;
        RECT 47.310 164.600 47.570 164.920 ;
        RECT 49.610 164.600 49.870 164.920 ;
        RECT 47.510 163.045 49.390 163.415 ;
        RECT 49.670 162.200 49.810 164.600 ;
        RECT 49.610 161.880 49.870 162.200 ;
        RECT 51.050 160.160 51.190 167.320 ;
        RECT 54.730 164.580 54.870 170.040 ;
        RECT 56.570 169.340 56.710 173.020 ;
        RECT 57.950 172.400 58.090 175.140 ;
        RECT 57.890 172.080 58.150 172.400 ;
        RECT 55.590 169.020 55.850 169.340 ;
        RECT 56.510 169.020 56.770 169.340 ;
        RECT 55.130 166.980 55.390 167.300 ;
        RECT 55.190 165.260 55.330 166.980 ;
        RECT 55.130 164.940 55.390 165.260 ;
        RECT 54.670 164.260 54.930 164.580 ;
        RECT 55.650 164.320 55.790 169.020 ;
        RECT 55.190 164.180 55.790 164.320 ;
        RECT 56.510 164.260 56.770 164.580 ;
        RECT 55.190 163.900 55.330 164.180 ;
        RECT 55.130 163.580 55.390 163.900 ;
        RECT 55.190 161.860 55.330 163.580 ;
        RECT 55.130 161.540 55.390 161.860 ;
        RECT 50.990 159.840 51.250 160.160 ;
        RECT 53.750 159.840 54.010 160.160 ;
        RECT 52.370 159.500 52.630 159.820 ;
        RECT 46.850 159.160 47.110 159.480 ;
        RECT 46.910 158.995 47.050 159.160 ;
        RECT 46.840 158.625 47.120 158.995 ;
        RECT 49.610 158.140 49.870 158.460 ;
        RECT 50.530 158.140 50.790 158.460 ;
        RECT 47.510 157.605 49.390 157.975 ;
        RECT 49.670 157.100 49.810 158.140 ;
        RECT 49.610 156.780 49.870 157.100 ;
        RECT 47.770 156.100 48.030 156.420 ;
        RECT 47.830 154.380 47.970 156.100 ;
        RECT 50.590 156.080 50.730 158.140 ;
        RECT 50.530 155.760 50.790 156.080 ;
        RECT 47.770 154.060 48.030 154.380 ;
        RECT 52.430 153.700 52.570 159.500 ;
        RECT 52.830 159.160 53.090 159.480 ;
        RECT 53.290 159.160 53.550 159.480 ;
        RECT 52.890 154.720 53.030 159.160 ;
        RECT 52.830 154.400 53.090 154.720 ;
        RECT 53.350 154.040 53.490 159.160 ;
        RECT 53.810 157.440 53.950 159.840 ;
        RECT 54.210 159.160 54.470 159.480 ;
        RECT 53.750 157.120 54.010 157.440 ;
        RECT 53.810 156.955 53.950 157.120 ;
        RECT 53.740 156.585 54.020 156.955 ;
        RECT 53.290 153.950 53.550 154.040 ;
        RECT 53.290 153.810 53.950 153.950 ;
        RECT 53.290 153.720 53.550 153.810 ;
        RECT 51.910 153.380 52.170 153.700 ;
        RECT 52.370 153.380 52.630 153.700 ;
        RECT 46.450 152.740 47.050 152.880 ;
        RECT 45.930 149.980 46.190 150.300 ;
        RECT 45.990 143.160 46.130 149.980 ;
        RECT 46.910 148.600 47.050 152.740 ;
        RECT 49.610 152.700 49.870 153.020 ;
        RECT 47.510 152.165 49.390 152.535 ;
        RECT 47.310 150.320 47.570 150.640 ;
        RECT 47.370 149.280 47.510 150.320 ;
        RECT 47.310 148.960 47.570 149.280 ;
        RECT 49.670 148.600 49.810 152.700 ;
        RECT 51.450 149.980 51.710 150.300 ;
        RECT 51.510 149.280 51.650 149.980 ;
        RECT 51.450 148.960 51.710 149.280 ;
        RECT 46.850 148.280 47.110 148.600 ;
        RECT 49.610 148.280 49.870 148.600 ;
        RECT 45.470 142.840 45.730 143.160 ;
        RECT 45.930 142.840 46.190 143.160 ;
        RECT 45.530 139.670 45.670 142.840 ;
        RECT 46.390 139.780 46.650 140.100 ;
        RECT 45.930 139.670 46.190 139.760 ;
        RECT 45.530 139.530 46.190 139.670 ;
        RECT 45.930 139.440 46.190 139.530 ;
        RECT 45.470 137.290 45.730 137.380 ;
        RECT 45.990 137.290 46.130 139.440 ;
        RECT 46.450 137.720 46.590 139.780 ;
        RECT 46.910 138.400 47.050 148.280 ;
        RECT 47.510 146.725 49.390 147.095 ;
        RECT 50.990 144.540 51.250 144.860 ;
        RECT 51.050 143.500 51.190 144.540 ;
        RECT 50.990 143.180 51.250 143.500 ;
        RECT 51.970 143.160 52.110 153.380 ;
        RECT 53.290 151.680 53.550 152.000 ;
        RECT 53.350 149.280 53.490 151.680 ;
        RECT 53.810 150.640 53.950 153.810 ;
        RECT 54.270 150.980 54.410 159.160 ;
        RECT 55.190 158.880 55.330 161.540 ;
        RECT 54.730 158.800 55.330 158.880 ;
        RECT 54.670 158.740 55.330 158.800 ;
        RECT 54.670 158.480 54.930 158.740 ;
        RECT 54.670 154.400 54.930 154.720 ;
        RECT 54.730 152.000 54.870 154.400 ;
        RECT 55.190 152.880 55.330 158.740 ;
        RECT 55.580 154.545 55.860 154.915 ;
        RECT 55.590 154.400 55.850 154.545 ;
        RECT 56.570 154.120 56.710 164.260 ;
        RECT 57.950 161.520 58.090 172.080 ;
        RECT 60.190 170.040 60.450 170.360 ;
        RECT 60.250 167.300 60.390 170.040 ;
        RECT 60.190 166.980 60.450 167.300 ;
        RECT 57.890 161.200 58.150 161.520 ;
        RECT 57.430 160.860 57.690 161.180 ;
        RECT 57.490 159.820 57.630 160.860 ;
        RECT 57.430 159.500 57.690 159.820 ;
        RECT 57.950 156.420 58.090 161.200 ;
        RECT 58.350 160.860 58.610 161.180 ;
        RECT 59.730 160.860 59.990 161.180 ;
        RECT 57.890 156.100 58.150 156.420 ;
        RECT 56.110 153.980 56.710 154.120 ;
        RECT 55.190 152.740 55.790 152.880 ;
        RECT 54.670 151.680 54.930 152.000 ;
        RECT 54.210 150.660 54.470 150.980 ;
        RECT 53.750 150.320 54.010 150.640 ;
        RECT 53.290 148.960 53.550 149.280 ;
        RECT 53.810 148.600 53.950 150.320 ;
        RECT 54.210 148.960 54.470 149.280 ;
        RECT 52.370 148.280 52.630 148.600 ;
        RECT 53.750 148.510 54.010 148.600 ;
        RECT 52.890 148.370 54.010 148.510 ;
        RECT 52.430 145.540 52.570 148.280 ;
        RECT 52.890 145.540 53.030 148.370 ;
        RECT 53.750 148.280 54.010 148.370 ;
        RECT 54.270 145.540 54.410 148.960 ;
        RECT 54.730 148.940 54.870 151.680 ;
        RECT 54.670 148.620 54.930 148.940 ;
        RECT 55.650 145.880 55.790 152.740 ;
        RECT 55.590 145.560 55.850 145.880 ;
        RECT 52.370 145.220 52.630 145.540 ;
        RECT 52.830 145.220 53.090 145.540 ;
        RECT 54.210 145.450 54.470 145.540 ;
        RECT 54.210 145.310 54.870 145.450 ;
        RECT 54.210 145.220 54.470 145.310 ;
        RECT 54.730 143.840 54.870 145.310 ;
        RECT 52.370 143.520 52.630 143.840 ;
        RECT 54.670 143.520 54.930 143.840 ;
        RECT 50.070 142.840 50.330 143.160 ;
        RECT 51.910 142.840 52.170 143.160 ;
        RECT 47.510 141.285 49.390 141.655 ;
        RECT 50.130 140.100 50.270 142.840 ;
        RECT 50.070 139.780 50.330 140.100 ;
        RECT 46.850 138.080 47.110 138.400 ;
        RECT 46.390 137.400 46.650 137.720 ;
        RECT 45.470 137.150 46.130 137.290 ;
        RECT 45.470 137.060 45.730 137.150 ;
        RECT 45.530 135.340 45.670 137.060 ;
        RECT 46.450 135.680 46.590 137.400 ;
        RECT 46.390 135.360 46.650 135.680 ;
        RECT 45.470 135.020 45.730 135.340 ;
        RECT 45.530 134.660 45.670 135.020 ;
        RECT 45.470 134.515 45.730 134.660 ;
        RECT 45.460 134.145 45.740 134.515 ;
        RECT 45.930 134.340 46.190 134.660 ;
        RECT 45.010 131.620 45.270 131.940 ;
        RECT 44.550 130.940 44.810 131.260 ;
        RECT 44.610 129.220 44.750 130.940 ;
        RECT 44.550 128.900 44.810 129.220 ;
        RECT 45.470 128.560 45.730 128.880 ;
        RECT 45.530 127.520 45.670 128.560 ;
        RECT 45.470 127.200 45.730 127.520 ;
        RECT 44.090 117.680 44.350 118.000 ;
        RECT 44.150 116.640 44.290 117.680 ;
        RECT 44.090 116.320 44.350 116.640 ;
        RECT 45.530 115.960 45.670 127.200 ;
        RECT 45.990 121.060 46.130 134.340 ;
        RECT 46.910 132.280 47.050 138.080 ;
        RECT 50.130 137.720 50.270 139.780 ;
        RECT 51.910 139.440 52.170 139.760 ;
        RECT 51.970 138.400 52.110 139.440 ;
        RECT 52.430 139.420 52.570 143.520 ;
        RECT 53.750 142.500 54.010 142.820 ;
        RECT 52.370 139.100 52.630 139.420 ;
        RECT 52.430 138.400 52.570 139.100 ;
        RECT 51.910 138.080 52.170 138.400 ;
        RECT 52.370 138.080 52.630 138.400 ;
        RECT 50.070 137.400 50.330 137.720 ;
        RECT 49.610 137.060 49.870 137.380 ;
        RECT 47.510 135.845 49.390 136.215 ;
        RECT 48.690 135.360 48.950 135.680 ;
        RECT 48.750 134.660 48.890 135.360 ;
        RECT 48.690 134.340 48.950 134.660 ;
        RECT 49.150 134.515 49.410 134.660 ;
        RECT 49.140 134.145 49.420 134.515 ;
        RECT 47.310 133.660 47.570 133.980 ;
        RECT 47.370 132.620 47.510 133.660 ;
        RECT 47.310 132.300 47.570 132.620 ;
        RECT 46.850 131.960 47.110 132.280 ;
        RECT 46.910 128.880 47.050 131.960 ;
        RECT 49.670 131.600 49.810 137.060 ;
        RECT 50.130 135.340 50.270 137.400 ;
        RECT 53.810 137.380 53.950 142.500 ;
        RECT 53.750 137.060 54.010 137.380 ;
        RECT 54.210 137.060 54.470 137.380 ;
        RECT 53.810 136.440 53.950 137.060 ;
        RECT 53.350 136.300 53.950 136.440 ;
        RECT 50.070 135.020 50.330 135.340 ;
        RECT 50.070 134.000 50.330 134.320 ;
        RECT 51.450 134.000 51.710 134.320 ;
        RECT 49.610 131.280 49.870 131.600 ;
        RECT 47.510 130.405 49.390 130.775 ;
        RECT 49.670 130.240 49.810 131.280 ;
        RECT 49.610 129.920 49.870 130.240 ;
        RECT 46.850 128.560 47.110 128.880 ;
        RECT 49.150 128.560 49.410 128.880 ;
        RECT 47.760 127.345 48.040 127.715 ;
        RECT 47.830 127.180 47.970 127.345 ;
        RECT 47.770 126.860 48.030 127.180 ;
        RECT 49.210 126.840 49.350 128.560 ;
        RECT 49.670 127.520 49.810 129.920 ;
        RECT 50.130 127.520 50.270 134.000 ;
        RECT 51.510 132.960 51.650 134.000 ;
        RECT 51.450 132.640 51.710 132.960 ;
        RECT 53.350 131.940 53.490 136.300 ;
        RECT 54.270 135.000 54.410 137.060 ;
        RECT 54.210 134.680 54.470 135.000 ;
        RECT 54.270 132.960 54.410 134.680 ;
        RECT 54.210 132.640 54.470 132.960 ;
        RECT 53.290 131.620 53.550 131.940 ;
        RECT 49.610 127.200 49.870 127.520 ;
        RECT 50.070 127.200 50.330 127.520 ;
        RECT 49.150 126.520 49.410 126.840 ;
        RECT 47.510 124.965 49.390 125.335 ;
        RECT 50.130 124.800 50.270 127.200 ;
        RECT 53.350 126.500 53.490 131.620 ;
        RECT 53.290 126.180 53.550 126.500 ;
        RECT 50.530 125.500 50.790 125.820 ;
        RECT 50.070 124.480 50.330 124.800 ;
        RECT 49.610 123.460 49.870 123.780 ;
        RECT 45.930 120.740 46.190 121.060 ;
        RECT 49.670 120.720 49.810 123.460 ;
        RECT 50.130 122.080 50.270 124.480 ;
        RECT 50.590 123.440 50.730 125.500 ;
        RECT 50.530 123.120 50.790 123.440 ;
        RECT 50.070 121.760 50.330 122.080 ;
        RECT 53.350 121.480 53.490 126.180 ;
        RECT 55.590 125.500 55.850 125.820 ;
        RECT 55.650 124.120 55.790 125.500 ;
        RECT 56.110 124.120 56.250 153.980 ;
        RECT 56.510 153.380 56.770 153.700 ;
        RECT 56.570 151.320 56.710 153.380 ;
        RECT 57.950 151.660 58.090 156.100 ;
        RECT 57.890 151.340 58.150 151.660 ;
        RECT 56.510 151.000 56.770 151.320 ;
        RECT 56.570 145.880 56.710 151.000 ;
        RECT 58.410 150.835 58.550 160.860 ;
        RECT 59.790 154.235 59.930 160.860 ;
        RECT 60.190 156.100 60.450 156.420 ;
        RECT 59.720 153.865 60.000 154.235 ;
        RECT 60.250 152.000 60.390 156.100 ;
        RECT 60.190 151.680 60.450 152.000 ;
        RECT 58.340 150.465 58.620 150.835 ;
        RECT 57.430 149.980 57.690 150.300 ;
        RECT 57.490 148.260 57.630 149.980 ;
        RECT 60.190 148.620 60.450 148.940 ;
        RECT 57.430 147.940 57.690 148.260 ;
        RECT 57.490 145.880 57.630 147.940 ;
        RECT 60.250 145.880 60.390 148.620 ;
        RECT 56.510 145.560 56.770 145.880 ;
        RECT 57.430 145.560 57.690 145.880 ;
        RECT 60.190 145.560 60.450 145.880 ;
        RECT 56.570 142.820 56.710 145.560 ;
        RECT 57.890 144.880 58.150 145.200 ;
        RECT 56.510 142.500 56.770 142.820 ;
        RECT 56.510 141.820 56.770 142.140 ;
        RECT 56.570 140.440 56.710 141.820 ;
        RECT 57.430 140.800 57.690 141.120 ;
        RECT 56.510 140.120 56.770 140.440 ;
        RECT 55.590 123.800 55.850 124.120 ;
        RECT 56.050 123.800 56.310 124.120 ;
        RECT 56.110 121.480 56.250 123.800 ;
        RECT 56.970 121.760 57.230 122.080 ;
        RECT 53.350 121.340 53.950 121.480 ;
        RECT 56.110 121.340 56.710 121.480 ;
        RECT 57.030 121.400 57.170 121.760 ;
        RECT 53.810 121.060 53.950 121.340 ;
        RECT 56.570 121.060 56.710 121.340 ;
        RECT 56.970 121.080 57.230 121.400 ;
        RECT 53.750 120.740 54.010 121.060 ;
        RECT 56.510 120.740 56.770 121.060 ;
        RECT 49.610 120.400 49.870 120.720 ;
        RECT 46.850 120.060 47.110 120.380 ;
        RECT 46.910 118.680 47.050 120.060 ;
        RECT 47.510 119.525 49.390 119.895 ;
        RECT 46.850 118.360 47.110 118.680 ;
        RECT 49.670 118.340 49.810 120.400 ;
        RECT 51.450 120.060 51.710 120.380 ;
        RECT 51.510 118.340 51.650 120.060 ;
        RECT 49.610 118.020 49.870 118.340 ;
        RECT 51.450 118.020 51.710 118.340 ;
        RECT 49.670 115.960 49.810 118.020 ;
        RECT 50.530 117.340 50.790 117.660 ;
        RECT 50.590 115.960 50.730 117.340 ;
        RECT 57.030 116.640 57.170 121.080 ;
        RECT 56.970 116.320 57.230 116.640 ;
        RECT 52.830 115.980 53.090 116.300 ;
        RECT 45.470 115.640 45.730 115.960 ;
        RECT 49.610 115.640 49.870 115.960 ;
        RECT 50.530 115.640 50.790 115.960 ;
        RECT 47.510 114.085 49.390 114.455 ;
        RECT 46.850 111.900 47.110 112.220 ;
        RECT 43.630 110.880 43.890 111.200 ;
        RECT 46.910 110.860 47.050 111.900 ;
        RECT 33.970 110.540 34.230 110.860 ;
        RECT 36.270 110.540 36.530 110.860 ;
        RECT 44.090 110.540 44.350 110.860 ;
        RECT 46.850 110.540 47.110 110.860 ;
        RECT 34.030 108.480 34.170 110.540 ;
        RECT 37.650 109.860 37.910 110.180 ;
        RECT 41.790 109.860 42.050 110.180 ;
        RECT 33.970 108.160 34.230 108.480 ;
        RECT 31.670 107.480 31.930 107.800 ;
        RECT 37.190 106.460 37.450 106.780 ;
        RECT 32.510 105.925 34.390 106.295 ;
        RECT 37.250 92.720 37.390 106.460 ;
        RECT 37.710 105.080 37.850 109.860 ;
        RECT 37.650 104.760 37.910 105.080 ;
        RECT 31.660 92.240 31.940 92.720 ;
        RECT 30.350 92.100 31.940 92.240 ;
        RECT 31.660 90.720 31.940 92.100 ;
        RECT 37.180 90.720 37.460 92.720 ;
        RECT 41.850 92.240 41.990 109.860 ;
        RECT 44.150 108.480 44.290 110.540 ;
        RECT 49.670 110.180 49.810 115.640 ;
        RECT 52.890 113.920 53.030 115.980 ;
        RECT 52.830 113.600 53.090 113.920 ;
        RECT 57.490 112.900 57.630 140.800 ;
        RECT 57.950 121.740 58.090 144.880 ;
        RECT 59.730 144.540 59.990 144.860 ;
        RECT 59.790 143.160 59.930 144.540 ;
        RECT 59.730 142.840 59.990 143.160 ;
        RECT 60.190 139.440 60.450 139.760 ;
        RECT 59.730 137.740 59.990 138.060 ;
        RECT 59.270 136.380 59.530 136.700 ;
        RECT 59.330 135.000 59.470 136.380 ;
        RECT 59.270 134.680 59.530 135.000 ;
        RECT 58.810 130.940 59.070 131.260 ;
        RECT 58.870 129.560 59.010 130.940 ;
        RECT 59.790 129.560 59.930 137.740 ;
        RECT 58.810 129.240 59.070 129.560 ;
        RECT 59.730 129.240 59.990 129.560 ;
        RECT 57.890 121.420 58.150 121.740 ;
        RECT 57.950 118.680 58.090 121.420 ;
        RECT 59.270 120.060 59.530 120.380 ;
        RECT 59.330 118.680 59.470 120.060 ;
        RECT 57.890 118.360 58.150 118.680 ;
        RECT 59.270 118.360 59.530 118.680 ;
        RECT 60.250 112.900 60.390 139.440 ;
        RECT 60.710 138.060 60.850 181.600 ;
        RECT 61.170 170.700 61.310 196.220 ;
        RECT 62.030 195.200 62.290 195.520 ;
        RECT 62.090 194.500 62.230 195.200 ;
        RECT 63.470 194.840 63.610 196.900 ;
        RECT 64.790 194.860 65.050 195.180 ;
        RECT 63.410 194.520 63.670 194.840 ;
        RECT 62.030 194.180 62.290 194.500 ;
        RECT 62.030 193.500 62.290 193.820 ;
        RECT 62.090 192.800 62.230 193.500 ;
        RECT 62.510 192.965 64.390 193.335 ;
        RECT 62.030 192.480 62.290 192.800 ;
        RECT 64.850 192.200 64.990 194.860 ;
        RECT 65.310 194.160 65.450 196.900 ;
        RECT 66.230 195.180 66.370 197.240 ;
        RECT 67.550 196.900 67.810 197.220 ;
        RECT 69.390 196.900 69.650 197.220 ;
        RECT 66.170 194.860 66.430 195.180 ;
        RECT 65.250 193.840 65.510 194.160 ;
        RECT 64.390 192.060 64.990 192.200 ;
        RECT 65.310 192.120 65.450 193.840 ;
        RECT 67.610 193.820 67.750 196.900 ;
        RECT 68.470 195.200 68.730 195.520 ;
        RECT 68.000 194.665 68.280 195.035 ;
        RECT 68.010 194.520 68.270 194.665 ;
        RECT 68.530 194.500 68.670 195.200 ;
        RECT 68.470 194.180 68.730 194.500 ;
        RECT 67.550 193.500 67.810 193.820 ;
        RECT 64.390 191.100 64.530 192.060 ;
        RECT 65.250 191.800 65.510 192.120 ;
        RECT 64.790 191.460 65.050 191.780 ;
        RECT 62.030 190.780 62.290 191.100 ;
        RECT 64.330 190.780 64.590 191.100 ;
        RECT 61.570 189.760 61.830 190.080 ;
        RECT 61.630 189.060 61.770 189.760 ;
        RECT 62.090 189.740 62.230 190.780 ;
        RECT 62.030 189.420 62.290 189.740 ;
        RECT 61.570 188.800 61.830 189.060 ;
        RECT 61.570 188.740 62.230 188.800 ;
        RECT 61.630 188.660 62.230 188.740 ;
        RECT 64.390 188.720 64.530 190.780 ;
        RECT 64.850 190.080 64.990 191.460 ;
        RECT 64.790 189.760 65.050 190.080 ;
        RECT 65.310 189.060 65.450 191.800 ;
        RECT 66.170 190.780 66.430 191.100 ;
        RECT 66.230 189.060 66.370 190.780 ;
        RECT 65.250 188.740 65.510 189.060 ;
        RECT 66.170 188.740 66.430 189.060 ;
        RECT 62.090 185.660 62.230 188.660 ;
        RECT 64.330 188.630 64.590 188.720 ;
        RECT 64.330 188.490 64.990 188.630 ;
        RECT 64.330 188.400 64.590 188.490 ;
        RECT 62.510 187.525 64.390 187.895 ;
        RECT 62.030 185.340 62.290 185.660 ;
        RECT 61.570 182.960 61.830 183.280 ;
        RECT 61.110 170.380 61.370 170.700 ;
        RECT 61.170 161.860 61.310 170.380 ;
        RECT 61.630 167.300 61.770 182.960 ;
        RECT 62.090 181.320 62.230 185.340 ;
        RECT 64.330 183.870 64.590 183.960 ;
        RECT 64.850 183.870 64.990 188.490 ;
        RECT 64.330 183.730 64.990 183.870 ;
        RECT 64.330 183.640 64.590 183.730 ;
        RECT 62.510 182.085 64.390 182.455 ;
        RECT 64.850 181.920 64.990 183.730 ;
        RECT 65.310 183.530 65.450 188.740 ;
        RECT 67.610 188.720 67.750 193.500 ;
        RECT 68.530 192.460 68.670 194.180 ;
        RECT 68.470 192.140 68.730 192.460 ;
        RECT 68.010 190.780 68.270 191.100 ;
        RECT 68.070 190.080 68.210 190.780 ;
        RECT 68.010 189.760 68.270 190.080 ;
        RECT 68.530 189.400 68.670 192.140 ;
        RECT 69.450 190.080 69.590 196.900 ;
        RECT 70.370 194.500 70.510 198.940 ;
        RECT 70.830 195.520 70.970 199.620 ;
        RECT 71.750 197.560 71.890 199.620 ;
        RECT 73.530 198.940 73.790 199.260 ;
        RECT 82.270 198.940 82.530 199.260 ;
        RECT 73.590 197.900 73.730 198.940 ;
        RECT 82.330 197.900 82.470 198.940 ;
        RECT 92.510 198.405 94.390 198.775 ;
        RECT 73.530 197.580 73.790 197.900 ;
        RECT 82.270 197.580 82.530 197.900 ;
        RECT 71.690 197.240 71.950 197.560 ;
        RECT 98.830 197.240 99.090 197.560 ;
        RECT 70.770 195.200 71.030 195.520 ;
        RECT 70.310 194.180 70.570 194.500 ;
        RECT 70.370 192.800 70.510 194.180 ;
        RECT 70.770 193.840 71.030 194.160 ;
        RECT 70.310 192.480 70.570 192.800 ;
        RECT 69.390 189.760 69.650 190.080 ;
        RECT 68.470 189.080 68.730 189.400 ;
        RECT 67.550 188.400 67.810 188.720 ;
        RECT 66.170 188.060 66.430 188.380 ;
        RECT 66.230 184.300 66.370 188.060 ;
        RECT 66.170 183.980 66.430 184.300 ;
        RECT 65.710 183.530 65.970 183.620 ;
        RECT 65.310 183.390 65.970 183.530 ;
        RECT 65.710 183.300 65.970 183.390 ;
        RECT 64.790 181.600 65.050 181.920 ;
        RECT 62.090 181.180 62.690 181.320 ;
        RECT 62.550 180.560 62.690 181.180 ;
        RECT 62.490 180.240 62.750 180.560 ;
        RECT 62.030 178.540 62.290 178.860 ;
        RECT 62.090 175.800 62.230 178.540 ;
        RECT 62.550 178.180 62.690 180.240 ;
        RECT 64.330 178.430 64.590 178.520 ;
        RECT 64.850 178.430 64.990 181.600 ;
        RECT 65.770 181.580 65.910 183.300 ;
        RECT 65.710 181.260 65.970 181.580 ;
        RECT 65.770 178.520 65.910 181.260 ;
        RECT 66.230 180.560 66.370 183.980 ;
        RECT 68.530 183.960 68.670 189.080 ;
        RECT 70.370 188.380 70.510 192.480 ;
        RECT 70.830 192.460 70.970 193.840 ;
        RECT 70.770 192.140 71.030 192.460 ;
        RECT 71.750 191.780 71.890 197.240 ;
        RECT 84.570 196.900 84.830 197.220 ;
        RECT 72.150 196.220 72.410 196.540 ;
        RECT 73.990 196.220 74.250 196.540 ;
        RECT 74.910 196.220 75.170 196.540 ;
        RECT 72.210 194.160 72.350 196.220 ;
        RECT 74.050 194.840 74.190 196.220 ;
        RECT 73.990 194.520 74.250 194.840 ;
        RECT 72.150 193.840 72.410 194.160 ;
        RECT 74.970 192.460 75.110 196.220 ;
        RECT 77.510 195.685 79.390 196.055 ;
        RECT 84.630 195.520 84.770 196.900 ;
        RECT 84.570 195.200 84.830 195.520 ;
        RECT 96.530 195.200 96.790 195.520 ;
        RECT 74.910 192.140 75.170 192.460 ;
        RECT 79.510 191.800 79.770 192.120 ;
        RECT 71.690 191.460 71.950 191.780 ;
        RECT 77.510 190.245 79.390 190.615 ;
        RECT 70.310 188.060 70.570 188.380 ;
        RECT 79.570 187.360 79.710 191.800 ;
        RECT 81.350 190.780 81.610 191.100 ;
        RECT 81.410 189.400 81.550 190.780 ;
        RECT 84.630 189.400 84.770 195.200 ;
        RECT 90.090 194.180 90.350 194.500 ;
        RECT 88.710 191.460 88.970 191.780 ;
        RECT 85.030 190.780 85.290 191.100 ;
        RECT 81.350 189.080 81.610 189.400 ;
        RECT 84.570 189.080 84.830 189.400 ;
        RECT 84.110 188.740 84.370 189.060 ;
        RECT 80.890 188.400 81.150 188.720 ;
        RECT 79.970 188.060 80.230 188.380 ;
        RECT 79.510 187.040 79.770 187.360 ;
        RECT 71.690 186.700 71.950 187.020 ;
        RECT 69.390 186.360 69.650 186.680 ;
        RECT 66.630 183.640 66.890 183.960 ;
        RECT 68.470 183.640 68.730 183.960 ;
        RECT 66.690 182.940 66.830 183.640 ;
        RECT 66.630 182.620 66.890 182.940 ;
        RECT 66.690 181.920 66.830 182.620 ;
        RECT 66.630 181.600 66.890 181.920 ;
        RECT 66.170 180.240 66.430 180.560 ;
        RECT 66.230 179.200 66.370 180.240 ;
        RECT 66.170 178.880 66.430 179.200 ;
        RECT 66.690 178.860 66.830 181.600 ;
        RECT 69.450 181.240 69.590 186.360 ;
        RECT 71.750 182.940 71.890 186.700 ;
        RECT 80.030 186.340 80.170 188.060 ;
        RECT 80.950 187.360 81.090 188.400 ;
        RECT 80.890 187.040 81.150 187.360 ;
        RECT 84.170 186.760 84.310 188.740 ;
        RECT 83.710 186.620 84.310 186.760 ;
        RECT 76.750 186.020 77.010 186.340 ;
        RECT 79.970 186.020 80.230 186.340 ;
        RECT 73.530 185.340 73.790 185.660 ;
        RECT 73.590 183.280 73.730 185.340 ;
        RECT 76.810 184.040 76.950 186.020 ;
        RECT 77.510 184.805 79.390 185.175 ;
        RECT 76.810 183.900 77.870 184.040 ;
        RECT 73.530 182.960 73.790 183.280 ;
        RECT 71.690 182.620 71.950 182.940 ;
        RECT 76.750 182.620 77.010 182.940 ;
        RECT 69.390 180.920 69.650 181.240 ;
        RECT 71.750 180.900 71.890 182.620 ;
        RECT 76.810 181.920 76.950 182.620 ;
        RECT 76.750 181.600 77.010 181.920 ;
        RECT 76.290 181.260 76.550 181.580 ;
        RECT 73.070 180.920 73.330 181.240 ;
        RECT 67.090 180.580 67.350 180.900 ;
        RECT 70.770 180.580 71.030 180.900 ;
        RECT 71.230 180.580 71.490 180.900 ;
        RECT 71.690 180.580 71.950 180.900 ;
        RECT 66.630 178.540 66.890 178.860 ;
        RECT 64.330 178.290 64.990 178.430 ;
        RECT 64.330 178.200 64.590 178.290 ;
        RECT 65.710 178.200 65.970 178.520 ;
        RECT 62.490 177.860 62.750 178.180 ;
        RECT 66.630 177.860 66.890 178.180 ;
        RECT 64.790 177.180 65.050 177.500 ;
        RECT 62.510 176.645 64.390 177.015 ;
        RECT 64.850 176.140 64.990 177.180 ;
        RECT 64.790 175.820 65.050 176.140 ;
        RECT 62.030 175.480 62.290 175.800 ;
        RECT 62.030 174.460 62.290 174.780 ;
        RECT 63.410 174.460 63.670 174.780 ;
        RECT 62.090 173.080 62.230 174.460 ;
        RECT 63.470 173.760 63.610 174.460 ;
        RECT 63.410 173.440 63.670 173.760 ;
        RECT 62.030 172.760 62.290 173.080 ;
        RECT 62.090 170.020 62.230 172.760 ;
        RECT 64.850 172.740 64.990 175.820 ;
        RECT 65.250 175.480 65.510 175.800 ;
        RECT 64.790 172.420 65.050 172.740 ;
        RECT 62.510 171.205 64.390 171.575 ;
        RECT 62.950 170.720 63.210 171.040 ;
        RECT 62.030 169.700 62.290 170.020 ;
        RECT 63.010 169.340 63.150 170.720 ;
        RECT 63.410 170.380 63.670 170.700 ;
        RECT 62.950 169.020 63.210 169.340 ;
        RECT 63.470 167.640 63.610 170.380 ;
        RECT 64.850 170.360 64.990 172.420 ;
        RECT 65.310 170.950 65.450 175.480 ;
        RECT 66.690 172.740 66.830 177.860 ;
        RECT 66.630 172.420 66.890 172.740 ;
        RECT 65.310 170.810 66.370 170.950 ;
        RECT 64.790 170.040 65.050 170.360 ;
        RECT 65.310 169.760 65.450 170.810 ;
        RECT 65.710 170.040 65.970 170.360 ;
        RECT 64.390 169.620 65.450 169.760 ;
        RECT 64.390 167.640 64.530 169.620 ;
        RECT 65.250 169.020 65.510 169.340 ;
        RECT 63.410 167.320 63.670 167.640 ;
        RECT 64.330 167.320 64.590 167.640 ;
        RECT 61.570 166.980 61.830 167.300 ;
        RECT 61.630 162.200 61.770 166.980 ;
        RECT 62.030 166.640 62.290 166.960 ;
        RECT 62.090 165.260 62.230 166.640 ;
        RECT 62.510 165.765 64.390 166.135 ;
        RECT 62.030 164.940 62.290 165.260 ;
        RECT 61.570 161.880 61.830 162.200 ;
        RECT 61.110 161.540 61.370 161.860 ;
        RECT 64.790 160.860 65.050 161.180 ;
        RECT 62.510 160.325 64.390 160.695 ;
        RECT 62.490 158.820 62.750 159.140 ;
        RECT 62.550 157.440 62.690 158.820 ;
        RECT 64.330 158.140 64.590 158.460 ;
        RECT 62.490 157.120 62.750 157.440 ;
        RECT 64.390 156.420 64.530 158.140 ;
        RECT 64.850 156.760 64.990 160.860 ;
        RECT 64.790 156.440 65.050 156.760 ;
        RECT 64.330 156.100 64.590 156.420 ;
        RECT 62.510 154.885 64.390 155.255 ;
        RECT 64.850 154.720 64.990 156.440 ;
        RECT 64.790 154.400 65.050 154.720 ;
        RECT 62.030 153.720 62.290 154.040 ;
        RECT 62.090 153.555 62.230 153.720 ;
        RECT 62.020 153.185 62.300 153.555 ;
        RECT 64.790 152.700 65.050 153.020 ;
        RECT 62.510 149.445 64.390 149.815 ;
        RECT 62.030 147.940 62.290 148.260 ;
        RECT 61.570 145.220 61.830 145.540 ;
        RECT 61.110 139.780 61.370 140.100 ;
        RECT 60.650 137.740 60.910 138.060 ;
        RECT 60.710 132.620 60.850 137.740 ;
        RECT 61.170 135.000 61.310 139.780 ;
        RECT 61.110 134.680 61.370 135.000 ;
        RECT 60.650 132.300 60.910 132.620 ;
        RECT 60.650 131.620 60.910 131.940 ;
        RECT 60.710 130.240 60.850 131.620 ;
        RECT 60.650 129.920 60.910 130.240 ;
        RECT 60.710 118.340 60.850 129.920 ;
        RECT 61.170 129.560 61.310 134.680 ;
        RECT 61.630 132.280 61.770 145.220 ;
        RECT 62.090 143.840 62.230 147.940 ;
        RECT 62.510 144.005 64.390 144.375 ;
        RECT 62.030 143.520 62.290 143.840 ;
        RECT 62.510 138.565 64.390 138.935 ;
        RECT 63.410 135.360 63.670 135.680 ;
        RECT 63.470 134.400 63.610 135.360 ;
        RECT 64.850 134.660 64.990 152.700 ;
        RECT 65.310 135.000 65.450 169.020 ;
        RECT 65.770 167.300 65.910 170.040 ;
        RECT 65.710 166.980 65.970 167.300 ;
        RECT 65.770 158.460 65.910 166.980 ;
        RECT 66.230 158.995 66.370 170.810 ;
        RECT 66.160 158.625 66.440 158.995 ;
        RECT 65.710 158.140 65.970 158.460 ;
        RECT 66.230 151.230 66.370 158.625 ;
        RECT 66.630 158.140 66.890 158.460 ;
        RECT 66.690 152.875 66.830 158.140 ;
        RECT 66.620 152.505 66.900 152.875 ;
        RECT 67.150 151.320 67.290 180.580 ;
        RECT 68.010 178.200 68.270 178.520 ;
        RECT 67.550 177.520 67.810 177.840 ;
        RECT 67.610 176.140 67.750 177.520 ;
        RECT 67.550 175.820 67.810 176.140 ;
        RECT 68.070 175.120 68.210 178.200 ;
        RECT 70.830 177.840 70.970 180.580 ;
        RECT 71.290 179.200 71.430 180.580 ;
        RECT 71.230 178.880 71.490 179.200 ;
        RECT 70.770 177.520 71.030 177.840 ;
        RECT 70.770 175.480 71.030 175.800 ;
        RECT 68.010 174.800 68.270 175.120 ;
        RECT 67.550 174.460 67.810 174.780 ;
        RECT 70.310 174.460 70.570 174.780 ;
        RECT 67.610 172.740 67.750 174.460 ;
        RECT 67.550 172.420 67.810 172.740 ;
        RECT 68.930 171.915 69.190 172.060 ;
        RECT 68.920 171.545 69.200 171.915 ;
        RECT 69.390 171.740 69.650 172.060 ;
        RECT 67.550 163.580 67.810 163.900 ;
        RECT 67.610 161.180 67.750 163.580 ;
        RECT 68.010 162.560 68.270 162.880 ;
        RECT 67.550 160.860 67.810 161.180 ;
        RECT 67.610 160.160 67.750 160.860 ;
        RECT 67.550 159.840 67.810 160.160 ;
        RECT 67.610 157.100 67.750 159.840 ;
        RECT 67.550 156.780 67.810 157.100 ;
        RECT 67.550 156.330 67.810 156.420 ;
        RECT 68.070 156.330 68.210 162.560 ;
        RECT 68.470 159.500 68.730 159.820 ;
        RECT 68.530 156.760 68.670 159.500 ;
        RECT 69.450 158.315 69.590 171.740 ;
        RECT 69.850 166.980 70.110 167.300 ;
        RECT 69.910 162.540 70.050 166.980 ;
        RECT 69.850 162.220 70.110 162.540 ;
        RECT 69.850 161.540 70.110 161.860 ;
        RECT 69.910 160.160 70.050 161.540 ;
        RECT 69.850 159.840 70.110 160.160 ;
        RECT 69.380 157.945 69.660 158.315 ;
        RECT 68.930 156.780 69.190 157.100 ;
        RECT 70.370 156.955 70.510 174.460 ;
        RECT 70.830 172.740 70.970 175.480 ;
        RECT 71.750 172.740 71.890 180.580 ;
        RECT 73.130 179.200 73.270 180.920 ;
        RECT 73.070 178.880 73.330 179.200 ;
        RECT 76.350 175.800 76.490 181.260 ;
        RECT 77.730 180.900 77.870 183.900 ;
        RECT 79.510 180.920 79.770 181.240 ;
        RECT 77.670 180.580 77.930 180.900 ;
        RECT 77.510 179.365 79.390 179.735 ;
        RECT 79.570 177.500 79.710 180.920 ;
        RECT 79.510 177.180 79.770 177.500 ;
        RECT 72.150 175.480 72.410 175.800 ;
        RECT 73.070 175.480 73.330 175.800 ;
        RECT 76.290 175.480 76.550 175.800 ;
        RECT 72.210 173.080 72.350 175.480 ;
        RECT 72.150 172.760 72.410 173.080 ;
        RECT 70.770 172.420 71.030 172.740 ;
        RECT 71.690 172.420 71.950 172.740 ;
        RECT 70.830 170.360 70.970 172.420 ;
        RECT 72.210 170.360 72.350 172.760 ;
        RECT 73.130 172.400 73.270 175.480 ;
        RECT 77.510 173.925 79.390 174.295 ;
        RECT 74.910 172.420 75.170 172.740 ;
        RECT 77.670 172.420 77.930 172.740 ;
        RECT 73.070 172.080 73.330 172.400 ;
        RECT 73.130 170.360 73.270 172.080 ;
        RECT 74.970 171.040 75.110 172.420 ;
        RECT 74.910 170.720 75.170 171.040 ;
        RECT 77.730 170.360 77.870 172.420 ;
        RECT 79.570 170.700 79.710 177.180 ;
        RECT 80.030 175.460 80.170 186.020 ;
        RECT 82.270 183.640 82.530 183.960 ;
        RECT 82.330 180.900 82.470 183.640 ;
        RECT 82.270 180.580 82.530 180.900 ;
        RECT 82.330 178.520 82.470 180.580 ;
        RECT 83.710 180.560 83.850 186.620 ;
        RECT 84.110 186.020 84.370 186.340 ;
        RECT 84.170 183.620 84.310 186.020 ;
        RECT 84.630 183.960 84.770 189.080 ;
        RECT 85.090 186.340 85.230 190.780 ;
        RECT 88.770 189.060 88.910 191.460 ;
        RECT 90.150 190.080 90.290 194.180 ;
        RECT 94.690 193.840 94.950 194.160 ;
        RECT 91.010 193.500 91.270 193.820 ;
        RECT 91.070 192.460 91.210 193.500 ;
        RECT 92.510 192.965 94.390 193.335 ;
        RECT 91.010 192.140 91.270 192.460 ;
        RECT 94.750 190.080 94.890 193.840 ;
        RECT 96.590 191.780 96.730 195.200 ;
        RECT 96.990 193.500 97.250 193.820 ;
        RECT 97.050 192.120 97.190 193.500 ;
        RECT 96.990 191.800 97.250 192.120 ;
        RECT 96.530 191.460 96.790 191.780 ;
        RECT 90.090 189.760 90.350 190.080 ;
        RECT 94.690 189.760 94.950 190.080 ;
        RECT 88.710 188.740 88.970 189.060 ;
        RECT 90.550 188.060 90.810 188.380 ;
        RECT 90.610 187.360 90.750 188.060 ;
        RECT 92.510 187.525 94.390 187.895 ;
        RECT 90.550 187.040 90.810 187.360 ;
        RECT 91.930 186.360 92.190 186.680 ;
        RECT 85.030 186.020 85.290 186.340 ;
        RECT 88.250 186.020 88.510 186.340 ;
        RECT 84.570 183.640 84.830 183.960 ;
        RECT 84.110 183.300 84.370 183.620 ;
        RECT 83.650 180.240 83.910 180.560 ;
        RECT 83.710 178.520 83.850 180.240 ;
        RECT 82.270 178.200 82.530 178.520 ;
        RECT 83.650 178.200 83.910 178.520 ;
        RECT 80.890 177.520 81.150 177.840 ;
        RECT 80.950 176.480 81.090 177.520 ;
        RECT 80.890 176.160 81.150 176.480 ;
        RECT 79.970 175.140 80.230 175.460 ;
        RECT 82.330 172.060 82.470 178.200 ;
        RECT 83.190 177.180 83.450 177.500 ;
        RECT 83.250 175.800 83.390 177.180 ;
        RECT 83.190 175.480 83.450 175.800 ;
        RECT 82.270 171.740 82.530 172.060 ;
        RECT 82.330 171.040 82.470 171.740 ;
        RECT 82.270 170.720 82.530 171.040 ;
        RECT 79.510 170.380 79.770 170.700 ;
        RECT 70.770 170.040 71.030 170.360 ;
        RECT 72.150 170.040 72.410 170.360 ;
        RECT 73.070 170.040 73.330 170.360 ;
        RECT 75.830 170.040 76.090 170.360 ;
        RECT 77.670 170.040 77.930 170.360 ;
        RECT 75.890 169.875 76.030 170.040 ;
        RECT 75.820 169.505 76.100 169.875 ;
        RECT 77.510 168.485 79.390 168.855 ;
        RECT 82.330 167.640 82.470 170.720 ;
        RECT 84.170 170.360 84.310 183.300 ;
        RECT 85.030 182.620 85.290 182.940 ;
        RECT 87.790 182.620 88.050 182.940 ;
        RECT 85.090 181.580 85.230 182.620 ;
        RECT 85.030 181.260 85.290 181.580 ;
        RECT 87.850 178.520 87.990 182.620 ;
        RECT 87.790 178.200 88.050 178.520 ;
        RECT 87.330 177.860 87.590 178.180 ;
        RECT 87.390 176.480 87.530 177.860 ;
        RECT 87.330 176.160 87.590 176.480 ;
        RECT 88.310 176.140 88.450 186.020 ;
        RECT 91.990 181.920 92.130 186.360 ;
        RECT 95.150 186.020 95.410 186.340 ;
        RECT 92.850 185.340 93.110 185.660 ;
        RECT 94.690 185.340 94.950 185.660 ;
        RECT 92.910 183.960 93.050 185.340 ;
        RECT 92.850 183.640 93.110 183.960 ;
        RECT 92.510 182.085 94.390 182.455 ;
        RECT 91.930 181.600 92.190 181.920 ;
        RECT 94.750 181.580 94.890 185.340 ;
        RECT 94.690 181.260 94.950 181.580 ;
        RECT 91.010 180.580 91.270 180.900 ;
        RECT 93.770 180.580 94.030 180.900 ;
        RECT 90.550 178.200 90.810 178.520 ;
        RECT 86.410 175.820 86.670 176.140 ;
        RECT 88.250 175.820 88.510 176.140 ;
        RECT 85.950 175.140 86.210 175.460 ;
        RECT 85.490 172.990 85.750 173.080 ;
        RECT 86.010 172.990 86.150 175.140 ;
        RECT 86.470 173.760 86.610 175.820 ;
        RECT 90.610 175.800 90.750 178.200 ;
        RECT 91.070 177.840 91.210 180.580 ;
        RECT 91.470 179.900 91.730 180.220 ;
        RECT 91.530 179.200 91.670 179.900 ;
        RECT 91.470 178.880 91.730 179.200 ;
        RECT 93.830 178.860 93.970 180.580 ;
        RECT 95.210 180.560 95.350 186.020 ;
        RECT 96.590 183.960 96.730 191.460 ;
        RECT 96.530 183.640 96.790 183.960 ;
        RECT 96.530 182.960 96.790 183.280 ;
        RECT 95.150 180.240 95.410 180.560 ;
        RECT 93.770 178.540 94.030 178.860 ;
        RECT 95.210 178.180 95.350 180.240 ;
        RECT 94.230 177.920 94.490 178.180 ;
        RECT 94.230 177.860 94.890 177.920 ;
        RECT 95.150 177.860 95.410 178.180 ;
        RECT 96.070 177.860 96.330 178.180 ;
        RECT 91.010 177.520 91.270 177.840 ;
        RECT 94.290 177.780 94.890 177.860 ;
        RECT 92.510 176.645 94.390 177.015 ;
        RECT 91.470 176.160 91.730 176.480 ;
        RECT 91.530 175.800 91.670 176.160 ;
        RECT 94.750 176.050 94.890 177.780 ;
        RECT 95.150 177.180 95.410 177.500 ;
        RECT 94.290 175.910 94.890 176.050 ;
        RECT 89.630 175.480 89.890 175.800 ;
        RECT 90.550 175.480 90.810 175.800 ;
        RECT 91.470 175.480 91.730 175.800 ;
        RECT 93.310 175.480 93.570 175.800 ;
        RECT 89.170 174.800 89.430 175.120 ;
        RECT 86.870 174.460 87.130 174.780 ;
        RECT 86.410 173.440 86.670 173.760 ;
        RECT 85.490 172.850 86.150 172.990 ;
        RECT 85.490 172.760 85.750 172.850 ;
        RECT 85.490 172.080 85.750 172.400 ;
        RECT 84.110 170.040 84.370 170.360 ;
        RECT 85.550 168.320 85.690 172.080 ;
        RECT 85.490 168.000 85.750 168.320 ;
        RECT 78.590 167.320 78.850 167.640 ;
        RECT 82.270 167.320 82.530 167.640 ;
        RECT 76.750 166.640 77.010 166.960 ;
        RECT 75.830 165.280 76.090 165.600 ;
        RECT 70.770 164.260 71.030 164.580 ;
        RECT 70.830 162.880 70.970 164.260 ;
        RECT 74.450 163.580 74.710 163.900 ;
        RECT 70.770 162.560 71.030 162.880 ;
        RECT 74.510 162.200 74.650 163.580 ;
        RECT 75.890 162.880 76.030 165.280 ;
        RECT 76.810 162.880 76.950 166.640 ;
        RECT 77.670 164.600 77.930 164.920 ;
        RECT 77.730 163.900 77.870 164.600 ;
        RECT 78.650 164.580 78.790 167.320 ;
        RECT 79.970 166.300 80.230 166.620 ;
        RECT 78.590 164.260 78.850 164.580 ;
        RECT 77.670 163.580 77.930 163.900 ;
        RECT 77.510 163.045 79.390 163.415 ;
        RECT 75.830 162.560 76.090 162.880 ;
        RECT 76.750 162.560 77.010 162.880 ;
        RECT 74.450 161.880 74.710 162.200 ;
        RECT 73.530 160.860 73.790 161.180 ;
        RECT 72.150 159.500 72.410 159.820 ;
        RECT 72.210 158.800 72.350 159.500 ;
        RECT 72.150 158.480 72.410 158.800 ;
        RECT 68.470 156.440 68.730 156.760 ;
        RECT 67.550 156.190 68.210 156.330 ;
        RECT 67.550 156.100 67.810 156.190 ;
        RECT 67.550 155.420 67.810 155.740 ;
        RECT 67.610 154.720 67.750 155.420 ;
        RECT 67.550 154.400 67.810 154.720 ;
        RECT 67.610 154.040 67.750 154.400 ;
        RECT 67.550 153.720 67.810 154.040 ;
        RECT 68.070 153.020 68.210 156.190 ;
        RECT 68.530 154.040 68.670 156.440 ;
        RECT 68.470 153.720 68.730 154.040 ;
        RECT 67.540 152.505 67.820 152.875 ;
        RECT 68.010 152.760 68.270 153.020 ;
        RECT 68.010 152.700 68.670 152.760 ;
        RECT 68.070 152.620 68.670 152.700 ;
        RECT 67.090 151.230 67.350 151.320 ;
        RECT 65.770 151.090 66.370 151.230 ;
        RECT 66.690 151.090 67.350 151.230 ;
        RECT 65.770 148.940 65.910 151.090 ;
        RECT 65.710 148.620 65.970 148.940 ;
        RECT 66.160 148.425 66.440 148.795 ;
        RECT 66.690 148.600 66.830 151.090 ;
        RECT 67.090 151.000 67.350 151.090 ;
        RECT 67.090 150.320 67.350 150.640 ;
        RECT 67.150 149.280 67.290 150.320 ;
        RECT 67.610 149.360 67.750 152.505 ;
        RECT 68.010 151.680 68.270 152.000 ;
        RECT 68.070 150.300 68.210 151.680 ;
        RECT 68.530 150.980 68.670 152.620 ;
        RECT 68.470 150.660 68.730 150.980 ;
        RECT 68.010 149.980 68.270 150.300 ;
        RECT 68.470 149.980 68.730 150.300 ;
        RECT 67.090 148.960 67.350 149.280 ;
        RECT 67.610 149.220 68.210 149.360 ;
        RECT 68.070 148.600 68.210 149.220 ;
        RECT 66.170 148.280 66.430 148.425 ;
        RECT 66.630 148.280 66.890 148.600 ;
        RECT 68.010 148.280 68.270 148.600 ;
        RECT 66.230 146.220 66.370 148.280 ;
        RECT 66.170 145.900 66.430 146.220 ;
        RECT 66.170 145.450 66.430 145.540 ;
        RECT 66.690 145.450 66.830 148.280 ;
        RECT 67.080 147.745 67.360 148.115 ;
        RECT 67.550 147.940 67.810 148.260 ;
        RECT 66.170 145.310 66.830 145.450 ;
        RECT 66.170 145.220 66.430 145.310 ;
        RECT 67.150 142.820 67.290 147.745 ;
        RECT 67.090 142.500 67.350 142.820 ;
        RECT 65.710 135.360 65.970 135.680 ;
        RECT 65.250 134.680 65.510 135.000 ;
        RECT 62.090 134.260 63.610 134.400 ;
        RECT 64.790 134.340 65.050 134.660 ;
        RECT 61.570 131.960 61.830 132.280 ;
        RECT 61.570 131.280 61.830 131.600 ;
        RECT 61.630 129.560 61.770 131.280 ;
        RECT 61.110 129.240 61.370 129.560 ;
        RECT 61.570 129.240 61.830 129.560 ;
        RECT 61.170 124.120 61.310 129.240 ;
        RECT 61.110 123.800 61.370 124.120 ;
        RECT 61.170 118.680 61.310 123.800 ;
        RECT 61.110 118.360 61.370 118.680 ;
        RECT 60.650 118.020 60.910 118.340 ;
        RECT 60.710 113.240 60.850 118.020 ;
        RECT 60.650 112.920 60.910 113.240 ;
        RECT 57.430 112.580 57.690 112.900 ;
        RECT 60.190 112.580 60.450 112.900 ;
        RECT 50.530 112.240 50.790 112.560 ;
        RECT 49.610 109.860 49.870 110.180 ;
        RECT 50.070 109.180 50.330 109.500 ;
        RECT 47.510 108.645 49.390 109.015 ;
        RECT 44.090 108.160 44.350 108.480 ;
        RECT 50.130 107.800 50.270 109.180 ;
        RECT 50.070 107.480 50.330 107.800 ;
        RECT 50.590 107.200 50.730 112.240 ;
        RECT 60.190 111.900 60.450 112.220 ;
        RECT 60.250 110.860 60.390 111.900 ;
        RECT 61.170 111.200 61.310 118.360 ;
        RECT 62.090 112.560 62.230 134.260 ;
        RECT 62.510 133.125 64.390 133.495 ;
        RECT 63.410 130.940 63.670 131.260 ;
        RECT 63.470 128.880 63.610 130.940 ;
        RECT 63.410 128.560 63.670 128.880 ;
        RECT 62.510 127.685 64.390 128.055 ;
        RECT 65.770 127.520 65.910 135.360 ;
        RECT 67.610 131.940 67.750 147.940 ;
        RECT 68.070 145.200 68.210 148.280 ;
        RECT 68.010 144.880 68.270 145.200 ;
        RECT 68.530 143.160 68.670 149.980 ;
        RECT 68.470 142.840 68.730 143.160 ;
        RECT 68.990 137.720 69.130 156.780 ;
        RECT 70.300 156.585 70.580 156.955 ;
        RECT 71.690 154.400 71.950 154.720 ;
        RECT 69.850 153.720 70.110 154.040 ;
        RECT 69.390 152.700 69.650 153.020 ;
        RECT 69.450 151.320 69.590 152.700 ;
        RECT 69.390 151.000 69.650 151.320 ;
        RECT 69.910 150.980 70.050 153.720 ;
        RECT 70.310 152.700 70.570 153.020 ;
        RECT 70.770 152.700 71.030 153.020 ;
        RECT 69.850 150.660 70.110 150.980 ;
        RECT 70.370 150.835 70.510 152.700 ;
        RECT 70.300 150.465 70.580 150.835 ;
        RECT 69.850 149.980 70.110 150.300 ;
        RECT 69.910 148.795 70.050 149.980 ;
        RECT 69.840 148.425 70.120 148.795 ;
        RECT 69.850 141.820 70.110 142.140 ;
        RECT 69.380 138.225 69.660 138.595 ;
        RECT 69.450 137.720 69.590 138.225 ;
        RECT 68.930 137.400 69.190 137.720 ;
        RECT 69.390 137.400 69.650 137.720 ;
        RECT 69.910 137.120 70.050 141.820 ;
        RECT 70.310 139.100 70.570 139.420 ;
        RECT 70.370 138.060 70.510 139.100 ;
        RECT 70.310 137.740 70.570 138.060 ;
        RECT 69.910 136.980 70.510 137.120 ;
        RECT 68.470 136.380 68.730 136.700 ;
        RECT 69.850 136.380 70.110 136.700 ;
        RECT 68.010 135.020 68.270 135.340 ;
        RECT 68.070 134.660 68.210 135.020 ;
        RECT 68.010 134.515 68.270 134.660 ;
        RECT 68.000 134.145 68.280 134.515 ;
        RECT 68.010 133.660 68.270 133.980 ;
        RECT 68.070 132.620 68.210 133.660 ;
        RECT 68.010 132.300 68.270 132.620 ;
        RECT 66.170 131.620 66.430 131.940 ;
        RECT 67.550 131.620 67.810 131.940 ;
        RECT 65.710 127.200 65.970 127.520 ;
        RECT 65.250 122.780 65.510 123.100 ;
        RECT 62.510 122.245 64.390 122.615 ;
        RECT 65.310 121.740 65.450 122.780 ;
        RECT 65.250 121.420 65.510 121.740 ;
        RECT 62.510 116.805 64.390 117.175 ;
        RECT 66.230 113.920 66.370 131.620 ;
        RECT 66.630 129.580 66.890 129.900 ;
        RECT 66.690 128.880 66.830 129.580 ;
        RECT 67.090 129.240 67.350 129.560 ;
        RECT 66.630 128.560 66.890 128.880 ;
        RECT 66.690 126.500 66.830 128.560 ;
        RECT 67.150 126.840 67.290 129.240 ;
        RECT 67.550 128.900 67.810 129.220 ;
        RECT 67.610 127.520 67.750 128.900 ;
        RECT 68.010 128.560 68.270 128.880 ;
        RECT 67.550 127.200 67.810 127.520 ;
        RECT 67.090 126.520 67.350 126.840 ;
        RECT 66.630 126.180 66.890 126.500 ;
        RECT 66.690 124.120 66.830 126.180 ;
        RECT 66.630 123.800 66.890 124.120 ;
        RECT 67.610 123.100 67.750 127.200 ;
        RECT 68.070 123.100 68.210 128.560 ;
        RECT 67.550 122.780 67.810 123.100 ;
        RECT 68.010 122.780 68.270 123.100 ;
        RECT 67.090 120.060 67.350 120.380 ;
        RECT 67.150 118.000 67.290 120.060 ;
        RECT 67.610 119.360 67.750 122.780 ;
        RECT 68.070 122.080 68.210 122.780 ;
        RECT 68.010 121.760 68.270 122.080 ;
        RECT 67.550 119.040 67.810 119.360 ;
        RECT 67.090 117.680 67.350 118.000 ;
        RECT 66.170 113.600 66.430 113.920 ;
        RECT 65.250 113.260 65.510 113.580 ;
        RECT 62.030 112.240 62.290 112.560 ;
        RECT 61.570 111.900 61.830 112.220 ;
        RECT 61.110 110.880 61.370 111.200 ;
        RECT 56.510 110.540 56.770 110.860 ;
        RECT 60.190 110.540 60.450 110.860 ;
        RECT 53.750 110.200 54.010 110.520 ;
        RECT 46.850 106.800 47.110 107.120 ;
        RECT 48.690 106.800 48.950 107.120 ;
        RECT 50.130 107.060 50.730 107.200 ;
        RECT 42.700 92.240 42.980 92.720 ;
        RECT 41.850 92.100 42.980 92.240 ;
        RECT 46.910 92.240 47.050 106.800 ;
        RECT 48.750 105.760 48.890 106.800 ;
        RECT 50.130 106.780 50.270 107.060 ;
        RECT 50.070 106.460 50.330 106.780 ;
        RECT 48.690 105.440 48.950 105.760 ;
        RECT 50.130 105.080 50.270 106.460 ;
        RECT 50.070 104.760 50.330 105.080 ;
        RECT 47.510 103.205 49.390 103.575 ;
        RECT 53.810 92.720 53.950 110.200 ;
        RECT 56.570 108.480 56.710 110.540 ;
        RECT 56.970 109.860 57.230 110.180 ;
        RECT 56.510 108.160 56.770 108.480 ;
        RECT 57.030 107.800 57.170 109.860 ;
        RECT 61.630 107.800 61.770 111.900 ;
        RECT 62.510 111.365 64.390 111.735 ;
        RECT 64.790 109.860 65.050 110.180 ;
        RECT 56.970 107.480 57.230 107.800 ;
        RECT 61.570 107.480 61.830 107.800 ;
        RECT 57.030 105.080 57.170 107.480 ;
        RECT 59.270 106.800 59.530 107.120 ;
        RECT 56.970 104.760 57.230 105.080 ;
        RECT 59.330 92.720 59.470 106.800 ;
        RECT 62.510 105.925 64.390 106.295 ;
        RECT 64.850 92.720 64.990 109.860 ;
        RECT 65.310 105.420 65.450 113.260 ;
        RECT 68.530 112.900 68.670 136.380 ;
        RECT 69.390 135.360 69.650 135.680 ;
        RECT 69.450 134.660 69.590 135.360 ;
        RECT 69.390 134.340 69.650 134.660 ;
        RECT 68.930 131.795 69.190 131.940 ;
        RECT 68.920 131.425 69.200 131.795 ;
        RECT 69.390 130.940 69.650 131.260 ;
        RECT 69.450 130.240 69.590 130.940 ;
        RECT 69.910 130.240 70.050 136.380 ;
        RECT 70.370 131.940 70.510 136.980 ;
        RECT 70.830 132.620 70.970 152.700 ;
        RECT 71.750 150.980 71.890 154.400 ;
        RECT 72.210 154.380 72.350 158.480 ;
        RECT 72.150 154.060 72.410 154.380 ;
        RECT 72.610 151.515 72.870 151.660 ;
        RECT 72.600 151.145 72.880 151.515 ;
        RECT 73.590 151.320 73.730 160.860 ;
        RECT 74.510 159.140 74.650 161.880 ;
        RECT 79.050 161.540 79.310 161.860 ;
        RECT 79.110 160.920 79.250 161.540 ;
        RECT 80.030 161.180 80.170 166.300 ;
        RECT 81.810 161.880 82.070 162.200 ;
        RECT 79.110 160.780 79.710 160.920 ;
        RECT 79.970 160.860 80.230 161.180 ;
        RECT 74.450 158.820 74.710 159.140 ;
        RECT 76.750 158.140 77.010 158.460 ;
        RECT 74.450 157.120 74.710 157.440 ;
        RECT 73.990 155.760 74.250 156.080 ;
        RECT 74.050 154.720 74.190 155.760 ;
        RECT 73.990 154.400 74.250 154.720 ;
        RECT 74.510 154.380 74.650 157.120 ;
        RECT 76.810 156.760 76.950 158.140 ;
        RECT 77.510 157.605 79.390 157.975 ;
        RECT 76.750 156.440 77.010 156.760 ;
        RECT 79.570 156.420 79.710 160.780 ;
        RECT 79.970 159.500 80.230 159.820 ;
        RECT 80.030 157.440 80.170 159.500 ;
        RECT 80.430 158.480 80.690 158.800 ;
        RECT 79.970 157.120 80.230 157.440 ;
        RECT 80.490 156.420 80.630 158.480 ;
        RECT 81.870 156.760 82.010 161.880 ;
        RECT 82.330 159.140 82.470 167.320 ;
        RECT 84.110 166.640 84.370 166.960 ;
        RECT 82.730 164.940 82.990 165.260 ;
        RECT 82.270 158.820 82.530 159.140 ;
        RECT 82.330 157.100 82.470 158.820 ;
        RECT 82.790 158.460 82.930 164.940 ;
        RECT 84.170 162.880 84.310 166.640 ;
        RECT 84.570 163.920 84.830 164.240 ;
        RECT 84.110 162.560 84.370 162.880 ;
        RECT 84.630 161.180 84.770 163.920 ;
        RECT 84.570 160.860 84.830 161.180 ;
        RECT 82.730 158.140 82.990 158.460 ;
        RECT 82.270 156.780 82.530 157.100 ;
        RECT 81.810 156.440 82.070 156.760 ;
        RECT 79.510 156.100 79.770 156.420 ;
        RECT 80.430 156.100 80.690 156.420 ;
        RECT 74.450 154.060 74.710 154.380 ;
        RECT 79.570 154.040 79.710 156.100 ;
        RECT 84.110 155.760 84.370 156.080 ;
        RECT 79.510 153.720 79.770 154.040 ;
        RECT 77.510 152.165 79.390 152.535 ;
        RECT 73.530 151.000 73.790 151.320 ;
        RECT 84.170 150.980 84.310 155.760 ;
        RECT 84.630 155.740 84.770 160.860 ;
        RECT 86.010 159.820 86.150 172.850 ;
        RECT 86.470 161.860 86.610 173.440 ;
        RECT 86.410 161.540 86.670 161.860 ;
        RECT 85.950 159.500 86.210 159.820 ;
        RECT 85.030 159.160 85.290 159.480 ;
        RECT 85.090 157.440 85.230 159.160 ;
        RECT 85.030 157.120 85.290 157.440 ;
        RECT 84.570 155.420 84.830 155.740 ;
        RECT 85.950 152.700 86.210 153.020 ;
        RECT 71.690 150.660 71.950 150.980 ;
        RECT 72.150 150.660 72.410 150.980 ;
        RECT 84.110 150.660 84.370 150.980 ;
        RECT 72.210 148.600 72.350 150.660 ;
        RECT 79.970 150.320 80.230 150.640 ;
        RECT 80.030 149.280 80.170 150.320 ;
        RECT 84.110 149.980 84.370 150.300 ;
        RECT 79.970 148.960 80.230 149.280 ;
        RECT 84.170 148.940 84.310 149.980 ;
        RECT 84.110 148.620 84.370 148.940 ;
        RECT 72.150 148.280 72.410 148.600 ;
        RECT 76.750 148.280 77.010 148.600 ;
        RECT 75.830 147.940 76.090 148.260 ;
        RECT 72.150 145.560 72.410 145.880 ;
        RECT 71.690 144.540 71.950 144.860 ;
        RECT 71.750 143.160 71.890 144.540 ;
        RECT 72.210 143.160 72.350 145.560 ;
        RECT 72.610 145.450 72.870 145.540 ;
        RECT 73.530 145.450 73.790 145.540 ;
        RECT 72.610 145.310 73.270 145.450 ;
        RECT 72.610 145.220 72.870 145.310 ;
        RECT 73.130 143.160 73.270 145.310 ;
        RECT 73.530 145.310 74.190 145.450 ;
        RECT 73.530 145.220 73.790 145.310 ;
        RECT 71.690 142.840 71.950 143.160 ;
        RECT 72.150 142.840 72.410 143.160 ;
        RECT 73.070 142.840 73.330 143.160 ;
        RECT 71.750 140.780 71.890 142.840 ;
        RECT 71.690 140.520 71.950 140.780 ;
        RECT 71.290 140.460 71.950 140.520 ;
        RECT 71.290 140.380 71.890 140.460 ;
        RECT 71.290 134.660 71.430 140.380 ;
        RECT 72.210 139.840 72.350 142.840 ;
        RECT 73.130 140.100 73.270 142.840 ;
        RECT 73.530 142.160 73.790 142.480 ;
        RECT 71.750 139.700 72.350 139.840 ;
        RECT 73.070 139.780 73.330 140.100 ;
        RECT 71.750 139.420 71.890 139.700 ;
        RECT 71.690 139.100 71.950 139.420 ;
        RECT 71.750 135.340 71.890 139.100 ;
        RECT 73.130 135.680 73.270 139.780 ;
        RECT 73.070 135.360 73.330 135.680 ;
        RECT 71.690 135.020 71.950 135.340 ;
        RECT 73.130 134.660 73.270 135.360 ;
        RECT 71.230 134.340 71.490 134.660 ;
        RECT 73.070 134.340 73.330 134.660 ;
        RECT 70.770 132.300 71.030 132.620 ;
        RECT 70.310 131.620 70.570 131.940 ;
        RECT 70.310 130.940 70.570 131.260 ;
        RECT 69.390 129.920 69.650 130.240 ;
        RECT 69.850 129.920 70.110 130.240 ;
        RECT 70.370 121.480 70.510 130.940 ;
        RECT 72.610 122.780 72.870 123.100 ;
        RECT 69.910 121.340 70.510 121.480 ;
        RECT 72.670 121.400 72.810 122.780 ;
        RECT 68.470 112.580 68.730 112.900 ;
        RECT 66.630 111.900 66.890 112.220 ;
        RECT 66.690 110.860 66.830 111.900 ;
        RECT 69.910 111.200 70.050 121.340 ;
        RECT 72.610 121.080 72.870 121.400 ;
        RECT 72.150 120.060 72.410 120.380 ;
        RECT 72.210 118.680 72.350 120.060 ;
        RECT 72.150 118.360 72.410 118.680 ;
        RECT 73.070 118.360 73.330 118.680 ;
        RECT 70.770 117.340 71.030 117.660 ;
        RECT 70.830 112.900 70.970 117.340 ;
        RECT 71.690 112.920 71.950 113.240 ;
        RECT 70.310 112.580 70.570 112.900 ;
        RECT 70.770 112.580 71.030 112.900 ;
        RECT 69.850 110.880 70.110 111.200 ;
        RECT 66.630 110.540 66.890 110.860 ;
        RECT 70.370 108.480 70.510 112.580 ;
        RECT 70.310 108.160 70.570 108.480 ;
        RECT 71.750 105.420 71.890 112.920 ;
        RECT 73.130 110.520 73.270 118.360 ;
        RECT 73.590 110.520 73.730 142.160 ;
        RECT 74.050 137.720 74.190 145.310 ;
        RECT 75.890 142.820 76.030 147.940 ;
        RECT 76.810 145.540 76.950 148.280 ;
        RECT 82.270 147.600 82.530 147.920 ;
        RECT 77.510 146.725 79.390 147.095 ;
        RECT 82.330 145.880 82.470 147.600 ;
        RECT 82.270 145.560 82.530 145.880 ;
        RECT 84.110 145.560 84.370 145.880 ;
        RECT 76.750 145.220 77.010 145.540 ;
        RECT 81.350 145.220 81.610 145.540 ;
        RECT 76.810 143.840 76.950 145.220 ;
        RECT 81.410 143.840 81.550 145.220 ;
        RECT 76.750 143.520 77.010 143.840 ;
        RECT 81.350 143.520 81.610 143.840 ;
        RECT 76.750 143.070 77.010 143.160 ;
        RECT 76.350 142.930 77.010 143.070 ;
        RECT 75.830 142.500 76.090 142.820 ;
        RECT 75.890 140.440 76.030 142.500 ;
        RECT 76.350 140.440 76.490 142.930 ;
        RECT 76.750 142.840 77.010 142.930 ;
        RECT 77.510 141.285 79.390 141.655 ;
        RECT 74.450 140.120 74.710 140.440 ;
        RECT 75.830 140.120 76.090 140.440 ;
        RECT 76.290 140.120 76.550 140.440 ;
        RECT 77.210 140.350 77.470 140.440 ;
        RECT 76.810 140.210 77.470 140.350 ;
        RECT 73.990 137.400 74.250 137.720 ;
        RECT 74.510 136.700 74.650 140.120 ;
        RECT 76.350 139.760 76.490 140.120 ;
        RECT 76.290 139.440 76.550 139.760 ;
        RECT 74.910 139.100 75.170 139.420 ;
        RECT 74.450 136.380 74.710 136.700 ;
        RECT 74.510 135.000 74.650 136.380 ;
        RECT 74.970 135.000 75.110 139.100 ;
        RECT 76.350 138.400 76.490 139.440 ;
        RECT 76.290 138.080 76.550 138.400 ;
        RECT 75.830 137.400 76.090 137.720 ;
        RECT 74.450 134.680 74.710 135.000 ;
        RECT 74.910 134.680 75.170 135.000 ;
        RECT 74.970 132.960 75.110 134.680 ;
        RECT 75.890 132.960 76.030 137.400 ;
        RECT 76.810 135.680 76.950 140.210 ;
        RECT 77.210 140.120 77.470 140.210 ;
        RECT 80.430 139.100 80.690 139.420 ;
        RECT 82.270 139.100 82.530 139.420 ;
        RECT 80.490 137.380 80.630 139.100 ;
        RECT 80.430 137.060 80.690 137.380 ;
        RECT 77.510 135.845 79.390 136.215 ;
        RECT 76.750 135.360 77.010 135.680 ;
        RECT 74.910 132.640 75.170 132.960 ;
        RECT 75.830 132.640 76.090 132.960 ;
        RECT 79.510 132.300 79.770 132.620 ;
        RECT 74.450 131.620 74.710 131.940 ;
        RECT 74.510 129.220 74.650 131.620 ;
        RECT 77.510 130.405 79.390 130.775 ;
        RECT 79.570 130.240 79.710 132.300 ;
        RECT 82.330 131.940 82.470 139.100 ;
        RECT 84.170 137.720 84.310 145.560 ;
        RECT 86.010 143.160 86.150 152.700 ;
        RECT 86.410 149.980 86.670 150.300 ;
        RECT 86.470 148.940 86.610 149.980 ;
        RECT 86.410 148.620 86.670 148.940 ;
        RECT 85.950 142.840 86.210 143.160 ;
        RECT 86.930 142.820 87.070 174.460 ;
        RECT 89.230 172.740 89.370 174.800 ;
        RECT 89.690 173.760 89.830 175.480 ;
        RECT 89.630 173.440 89.890 173.760 ;
        RECT 89.690 172.740 89.830 173.440 ;
        RECT 91.530 172.740 91.670 175.480 ;
        RECT 92.850 175.140 93.110 175.460 ;
        RECT 91.930 174.460 92.190 174.780 ;
        RECT 87.330 172.420 87.590 172.740 ;
        RECT 89.170 172.420 89.430 172.740 ;
        RECT 89.630 172.420 89.890 172.740 ;
        RECT 91.470 172.420 91.730 172.740 ;
        RECT 87.390 169.680 87.530 172.420 ;
        RECT 91.010 171.740 91.270 172.060 ;
        RECT 87.330 169.360 87.590 169.680 ;
        RECT 87.780 169.505 88.060 169.875 ;
        RECT 87.850 167.300 87.990 169.505 ;
        RECT 88.250 169.020 88.510 169.340 ;
        RECT 87.790 166.980 88.050 167.300 ;
        RECT 88.310 162.200 88.450 169.020 ;
        RECT 88.250 161.880 88.510 162.200 ;
        RECT 90.550 161.880 90.810 162.200 ;
        RECT 88.710 159.160 88.970 159.480 ;
        RECT 90.090 159.160 90.350 159.480 ;
        RECT 88.770 157.440 88.910 159.160 ;
        RECT 88.710 157.120 88.970 157.440 ;
        RECT 90.150 156.160 90.290 159.160 ;
        RECT 90.610 156.760 90.750 161.880 ;
        RECT 90.550 156.440 90.810 156.760 ;
        RECT 90.150 156.080 90.750 156.160 ;
        RECT 90.150 156.020 90.810 156.080 ;
        RECT 90.550 155.760 90.810 156.020 ;
        RECT 87.330 155.420 87.590 155.740 ;
        RECT 87.790 155.420 88.050 155.740 ;
        RECT 87.390 154.040 87.530 155.420 ;
        RECT 87.850 154.235 87.990 155.420 ;
        RECT 87.330 153.720 87.590 154.040 ;
        RECT 87.780 153.865 88.060 154.235 ;
        RECT 87.850 153.700 87.990 153.865 ;
        RECT 90.610 153.700 90.750 155.760 ;
        RECT 87.790 153.380 88.050 153.700 ;
        RECT 90.550 153.380 90.810 153.700 ;
        RECT 89.170 152.700 89.430 153.020 ;
        RECT 86.870 142.500 87.130 142.820 ;
        RECT 85.490 141.820 85.750 142.140 ;
        RECT 86.870 141.820 87.130 142.140 ;
        RECT 84.110 137.400 84.370 137.720 ;
        RECT 84.170 135.000 84.310 137.400 ;
        RECT 84.110 134.680 84.370 135.000 ;
        RECT 82.270 131.620 82.530 131.940 ;
        RECT 79.510 129.920 79.770 130.240 ;
        RECT 84.170 129.220 84.310 134.680 ;
        RECT 74.450 128.900 74.710 129.220 ;
        RECT 75.830 129.130 76.090 129.220 ;
        RECT 74.970 128.990 76.090 129.130 ;
        RECT 73.990 125.500 74.250 125.820 ;
        RECT 74.050 121.400 74.190 125.500 ;
        RECT 74.510 124.800 74.650 128.900 ;
        RECT 74.450 124.480 74.710 124.800 ;
        RECT 74.970 123.780 75.110 128.990 ;
        RECT 75.830 128.900 76.090 128.990 ;
        RECT 84.110 128.900 84.370 129.220 ;
        RECT 84.570 128.900 84.830 129.220 ;
        RECT 83.650 128.560 83.910 128.880 ;
        RECT 76.290 128.220 76.550 128.540 ;
        RECT 79.510 128.220 79.770 128.540 ;
        RECT 75.830 123.800 76.090 124.120 ;
        RECT 74.910 123.460 75.170 123.780 ;
        RECT 74.970 121.400 75.110 123.460 ;
        RECT 75.370 123.120 75.630 123.440 ;
        RECT 75.430 122.080 75.570 123.120 ;
        RECT 75.370 121.760 75.630 122.080 ;
        RECT 73.990 121.080 74.250 121.400 ;
        RECT 74.910 121.080 75.170 121.400 ;
        RECT 75.890 119.360 76.030 123.800 ;
        RECT 75.830 119.040 76.090 119.360 ;
        RECT 76.350 118.340 76.490 128.220 ;
        RECT 76.750 126.180 77.010 126.500 ;
        RECT 76.810 124.710 76.950 126.180 ;
        RECT 77.510 124.965 79.390 125.335 ;
        RECT 76.810 124.570 77.410 124.710 ;
        RECT 77.270 123.100 77.410 124.570 ;
        RECT 77.210 122.780 77.470 123.100 ;
        RECT 76.750 120.740 77.010 121.060 ;
        RECT 76.810 118.680 76.950 120.740 ;
        RECT 77.270 120.380 77.410 122.780 ;
        RECT 79.570 121.740 79.710 128.220 ;
        RECT 81.350 127.200 81.610 127.520 ;
        RECT 81.410 124.120 81.550 127.200 ;
        RECT 83.710 127.180 83.850 128.560 ;
        RECT 84.170 127.520 84.310 128.900 ;
        RECT 84.110 127.200 84.370 127.520 ;
        RECT 83.650 127.035 83.910 127.180 ;
        RECT 83.640 126.665 83.920 127.035 ;
        RECT 84.630 126.840 84.770 128.900 ;
        RECT 84.570 126.520 84.830 126.840 ;
        RECT 82.270 125.840 82.530 126.160 ;
        RECT 82.330 124.120 82.470 125.840 ;
        RECT 81.350 123.800 81.610 124.120 ;
        RECT 82.270 123.800 82.530 124.120 ;
        RECT 79.510 121.420 79.770 121.740 ;
        RECT 81.410 121.060 81.550 123.800 ;
        RECT 84.630 123.100 84.770 126.520 ;
        RECT 84.570 122.780 84.830 123.100 ;
        RECT 83.650 121.080 83.910 121.400 ;
        RECT 81.350 120.740 81.610 121.060 ;
        RECT 83.710 120.915 83.850 121.080 ;
        RECT 83.640 120.545 83.920 120.915 ;
        RECT 77.210 120.060 77.470 120.380 ;
        RECT 84.110 120.060 84.370 120.380 ;
        RECT 77.510 119.525 79.390 119.895 ;
        RECT 76.750 118.360 77.010 118.680 ;
        RECT 76.290 118.020 76.550 118.340 ;
        RECT 84.170 118.000 84.310 120.060 ;
        RECT 84.630 119.360 84.770 122.780 ;
        RECT 84.570 119.040 84.830 119.360 ;
        RECT 84.110 117.680 84.370 118.000 ;
        RECT 77.510 114.085 79.390 114.455 ;
        RECT 85.550 112.900 85.690 141.820 ;
        RECT 85.950 137.060 86.210 137.380 ;
        RECT 86.010 135.680 86.150 137.060 ;
        RECT 85.950 135.360 86.210 135.680 ;
        RECT 86.930 130.240 87.070 141.820 ;
        RECT 86.870 129.920 87.130 130.240 ;
        RECT 87.330 126.180 87.590 126.500 ;
        RECT 87.390 124.800 87.530 126.180 ;
        RECT 86.410 124.480 86.670 124.800 ;
        RECT 87.330 124.480 87.590 124.800 ;
        RECT 86.470 122.080 86.610 124.480 ;
        RECT 88.250 122.780 88.510 123.100 ;
        RECT 86.410 121.760 86.670 122.080 ;
        RECT 88.310 121.400 88.450 122.780 ;
        RECT 88.250 121.080 88.510 121.400 ;
        RECT 87.320 120.545 87.600 120.915 ;
        RECT 87.330 120.400 87.590 120.545 ;
        RECT 88.710 120.060 88.970 120.380 ;
        RECT 88.770 118.680 88.910 120.060 ;
        RECT 88.710 118.360 88.970 118.680 ;
        RECT 89.230 116.300 89.370 152.700 ;
        RECT 90.540 151.145 90.820 151.515 ;
        RECT 89.630 149.980 89.890 150.300 ;
        RECT 89.690 142.480 89.830 149.980 ;
        RECT 90.610 148.600 90.750 151.145 ;
        RECT 91.070 148.795 91.210 171.740 ;
        RECT 91.470 163.580 91.730 163.900 ;
        RECT 91.530 162.880 91.670 163.580 ;
        RECT 91.470 162.560 91.730 162.880 ;
        RECT 91.470 158.140 91.730 158.460 ;
        RECT 91.530 154.040 91.670 158.140 ;
        RECT 91.470 153.720 91.730 154.040 ;
        RECT 91.470 151.680 91.730 152.000 ;
        RECT 90.550 148.280 90.810 148.600 ;
        RECT 91.000 148.425 91.280 148.795 ;
        RECT 90.610 143.840 90.750 148.280 ;
        RECT 90.550 143.520 90.810 143.840 ;
        RECT 90.090 142.840 90.350 143.160 ;
        RECT 89.630 142.160 89.890 142.480 ;
        RECT 90.150 140.100 90.290 142.840 ;
        RECT 90.610 142.390 90.750 143.520 ;
        RECT 91.010 142.390 91.270 142.480 ;
        RECT 90.610 142.250 91.270 142.390 ;
        RECT 91.010 142.160 91.270 142.250 ;
        RECT 90.090 139.780 90.350 140.100 ;
        RECT 90.150 138.400 90.290 139.780 ;
        RECT 90.090 138.080 90.350 138.400 ;
        RECT 90.090 136.380 90.350 136.700 ;
        RECT 90.150 134.660 90.290 136.380 ;
        RECT 89.630 134.340 89.890 134.660 ;
        RECT 90.090 134.340 90.350 134.660 ;
        RECT 89.690 132.960 89.830 134.340 ;
        RECT 89.630 132.640 89.890 132.960 ;
        RECT 89.690 128.540 89.830 132.640 ;
        RECT 90.090 132.300 90.350 132.620 ;
        RECT 90.150 129.560 90.290 132.300 ;
        RECT 90.550 131.960 90.810 132.280 ;
        RECT 90.610 131.000 90.750 131.960 ;
        RECT 91.530 131.600 91.670 151.680 ;
        RECT 91.990 151.320 92.130 174.460 ;
        RECT 92.910 172.740 93.050 175.140 ;
        RECT 93.370 175.120 93.510 175.480 ;
        RECT 94.290 175.120 94.430 175.910 ;
        RECT 93.310 174.800 93.570 175.120 ;
        RECT 94.230 174.800 94.490 175.120 ;
        RECT 93.370 173.760 93.510 174.800 ;
        RECT 94.690 174.460 94.950 174.780 ;
        RECT 93.310 173.440 93.570 173.760 ;
        RECT 93.370 172.740 93.510 173.440 ;
        RECT 92.850 172.420 93.110 172.740 ;
        RECT 93.310 172.420 93.570 172.740 ;
        RECT 92.510 171.205 94.390 171.575 ;
        RECT 92.510 165.765 94.390 166.135 ;
        RECT 92.510 160.325 94.390 160.695 ;
        RECT 92.380 159.305 92.660 159.675 ;
        RECT 92.390 159.160 92.650 159.305 ;
        RECT 92.850 159.160 93.110 159.480 ;
        RECT 92.450 156.420 92.590 159.160 ;
        RECT 92.910 156.420 93.050 159.160 ;
        RECT 94.750 159.140 94.890 174.460 ;
        RECT 94.690 158.820 94.950 159.140 ;
        RECT 94.690 158.140 94.950 158.460 ;
        RECT 92.390 156.100 92.650 156.420 ;
        RECT 92.850 156.100 93.110 156.420 ;
        RECT 92.510 154.885 94.390 155.255 ;
        RECT 93.770 153.720 94.030 154.040 ;
        RECT 94.220 153.865 94.500 154.235 ;
        RECT 94.230 153.720 94.490 153.865 ;
        RECT 93.830 153.020 93.970 153.720 ;
        RECT 92.390 152.700 92.650 153.020 ;
        RECT 93.770 152.700 94.030 153.020 ;
        RECT 94.750 152.880 94.890 158.140 ;
        RECT 94.290 152.740 94.890 152.880 ;
        RECT 91.930 151.000 92.190 151.320 ;
        RECT 92.450 150.835 92.590 152.700 ;
        RECT 94.290 150.980 94.430 152.740 ;
        RECT 91.930 150.320 92.190 150.640 ;
        RECT 92.380 150.465 92.660 150.835 ;
        RECT 94.230 150.660 94.490 150.980 ;
        RECT 91.990 148.940 92.130 150.320 ;
        RECT 94.690 149.980 94.950 150.300 ;
        RECT 92.510 149.445 94.390 149.815 ;
        RECT 94.750 149.280 94.890 149.980 ;
        RECT 94.690 148.960 94.950 149.280 ;
        RECT 91.930 148.620 92.190 148.940 ;
        RECT 91.930 146.240 92.190 146.560 ;
        RECT 91.470 131.280 91.730 131.600 ;
        RECT 90.610 130.860 91.670 131.000 ;
        RECT 90.090 129.240 90.350 129.560 ;
        RECT 89.630 128.220 89.890 128.540 ;
        RECT 89.690 126.840 89.830 128.220 ;
        RECT 90.150 127.520 90.290 129.240 ;
        RECT 91.010 128.900 91.270 129.220 ;
        RECT 90.090 127.200 90.350 127.520 ;
        RECT 89.630 126.750 89.890 126.840 ;
        RECT 89.630 126.610 90.290 126.750 ;
        RECT 89.630 126.520 89.890 126.610 ;
        RECT 89.630 125.500 89.890 125.820 ;
        RECT 89.690 121.400 89.830 125.500 ;
        RECT 90.150 121.400 90.290 126.610 ;
        RECT 91.070 126.160 91.210 128.900 ;
        RECT 91.530 126.240 91.670 130.860 ;
        RECT 91.990 127.520 92.130 146.240 ;
        RECT 95.210 145.880 95.350 177.180 ;
        RECT 96.130 175.800 96.270 177.860 ;
        RECT 96.070 175.480 96.330 175.800 ;
        RECT 96.590 173.080 96.730 182.960 ;
        RECT 97.050 175.800 97.190 191.800 ;
        RECT 98.370 191.460 98.630 191.780 ;
        RECT 97.450 190.780 97.710 191.100 ;
        RECT 97.510 189.060 97.650 190.780 ;
        RECT 97.450 188.740 97.710 189.060 ;
        RECT 98.430 188.720 98.570 191.460 ;
        RECT 98.890 190.080 99.030 197.240 ;
        RECT 99.750 196.220 100.010 196.540 ;
        RECT 99.810 194.840 99.950 196.220 ;
        RECT 107.510 195.685 109.390 196.055 ;
        RECT 99.750 194.520 100.010 194.840 ;
        RECT 109.410 193.840 109.670 194.160 ;
        RECT 109.470 192.120 109.610 193.840 ;
        RECT 109.410 191.800 109.670 192.120 ;
        RECT 110.790 191.800 111.050 192.120 ;
        RECT 104.810 191.460 105.070 191.780 ;
        RECT 99.290 190.780 99.550 191.100 ;
        RECT 98.830 189.760 99.090 190.080 ;
        RECT 98.370 188.400 98.630 188.720 ;
        RECT 98.430 186.590 98.570 188.400 ;
        RECT 99.350 188.380 99.490 190.780 ;
        RECT 104.870 190.080 105.010 191.460 ;
        RECT 107.510 190.245 109.390 190.615 ;
        RECT 104.810 189.760 105.070 190.080 ;
        RECT 104.350 188.740 104.610 189.060 ;
        RECT 99.290 188.060 99.550 188.380 ;
        RECT 102.970 188.060 103.230 188.380 ;
        RECT 98.830 186.590 99.090 186.680 ;
        RECT 98.430 186.450 99.090 186.590 ;
        RECT 98.830 186.360 99.090 186.450 ;
        RECT 98.890 183.620 99.030 186.360 ;
        RECT 99.350 186.340 99.490 188.060 ;
        RECT 103.030 186.680 103.170 188.060 ;
        RECT 104.410 187.360 104.550 188.740 ;
        RECT 104.350 187.040 104.610 187.360 ;
        RECT 102.970 186.360 103.230 186.680 ;
        RECT 99.290 186.020 99.550 186.340 ;
        RECT 98.830 183.300 99.090 183.620 ;
        RECT 97.450 177.520 97.710 177.840 ;
        RECT 97.510 175.800 97.650 177.520 ;
        RECT 96.990 175.480 97.250 175.800 ;
        RECT 97.450 175.480 97.710 175.800 ;
        RECT 96.530 172.760 96.790 173.080 ;
        RECT 97.450 172.990 97.710 173.080 ;
        RECT 97.450 172.850 98.570 172.990 ;
        RECT 97.450 172.760 97.710 172.850 ;
        RECT 96.070 171.740 96.330 172.060 ;
        RECT 97.450 171.740 97.710 172.060 ;
        RECT 95.610 166.300 95.870 166.620 ;
        RECT 95.670 164.580 95.810 166.300 ;
        RECT 95.610 164.260 95.870 164.580 ;
        RECT 96.130 164.320 96.270 171.740 ;
        RECT 96.990 169.700 97.250 170.020 ;
        RECT 97.050 167.640 97.190 169.700 ;
        RECT 96.990 167.320 97.250 167.640 ;
        RECT 97.050 165.260 97.190 167.320 ;
        RECT 96.990 164.940 97.250 165.260 ;
        RECT 95.670 159.820 95.810 164.260 ;
        RECT 96.130 164.180 97.190 164.320 ;
        RECT 95.610 159.500 95.870 159.820 ;
        RECT 96.070 159.160 96.330 159.480 ;
        RECT 96.520 159.305 96.800 159.675 ;
        RECT 96.530 159.160 96.790 159.305 ;
        RECT 96.130 156.420 96.270 159.160 ;
        RECT 96.590 157.100 96.730 159.160 ;
        RECT 96.530 156.780 96.790 157.100 ;
        RECT 96.070 156.100 96.330 156.420 ;
        RECT 95.610 155.420 95.870 155.740 ;
        RECT 95.670 153.440 95.810 155.420 ;
        RECT 96.130 154.040 96.270 156.100 ;
        RECT 96.530 155.420 96.790 155.740 ;
        RECT 96.590 154.380 96.730 155.420 ;
        RECT 96.530 154.060 96.790 154.380 ;
        RECT 96.070 153.720 96.330 154.040 ;
        RECT 95.670 153.300 96.730 153.440 ;
        RECT 96.070 152.700 96.330 153.020 ;
        RECT 95.600 149.785 95.880 150.155 ;
        RECT 95.150 145.560 95.410 145.880 ;
        RECT 95.670 145.280 95.810 149.785 ;
        RECT 96.130 149.280 96.270 152.700 ;
        RECT 96.070 148.960 96.330 149.280 ;
        RECT 96.590 145.540 96.730 153.300 ;
        RECT 94.690 144.880 94.950 145.200 ;
        RECT 95.210 145.140 95.810 145.280 ;
        RECT 96.530 145.220 96.790 145.540 ;
        RECT 92.510 144.005 94.390 144.375 ;
        RECT 94.750 143.840 94.890 144.880 ;
        RECT 94.690 143.520 94.950 143.840 ;
        RECT 94.690 142.160 94.950 142.480 ;
        RECT 92.510 138.565 94.390 138.935 ;
        RECT 93.770 137.740 94.030 138.060 ;
        RECT 93.830 135.680 93.970 137.740 ;
        RECT 93.770 135.360 94.030 135.680 ;
        RECT 92.510 133.125 94.390 133.495 ;
        RECT 92.390 131.620 92.650 131.940 ;
        RECT 92.450 129.560 92.590 131.620 ;
        RECT 92.390 129.240 92.650 129.560 ;
        RECT 92.510 127.685 94.390 128.055 ;
        RECT 91.930 127.200 92.190 127.520 ;
        RECT 91.010 125.840 91.270 126.160 ;
        RECT 91.530 126.100 92.130 126.240 ;
        RECT 89.630 121.080 89.890 121.400 ;
        RECT 90.090 121.080 90.350 121.400 ;
        RECT 91.070 121.060 91.210 125.840 ;
        RECT 91.470 125.500 91.730 125.820 ;
        RECT 91.530 123.440 91.670 125.500 ;
        RECT 91.470 123.120 91.730 123.440 ;
        RECT 91.990 121.740 92.130 126.100 ;
        RECT 92.510 122.245 94.390 122.615 ;
        RECT 91.930 121.420 92.190 121.740 ;
        RECT 91.010 120.740 91.270 121.060 ;
        RECT 90.550 120.060 90.810 120.380 ;
        RECT 90.610 118.000 90.750 120.060 ;
        RECT 91.990 119.360 92.130 121.420 ;
        RECT 91.930 119.040 92.190 119.360 ;
        RECT 90.550 117.680 90.810 118.000 ;
        RECT 92.510 116.805 94.390 117.175 ;
        RECT 89.170 115.980 89.430 116.300 ;
        RECT 94.750 112.900 94.890 142.160 ;
        RECT 95.210 131.600 95.350 145.140 ;
        RECT 96.070 144.540 96.330 144.860 ;
        RECT 96.530 144.540 96.790 144.860 ;
        RECT 95.610 143.520 95.870 143.840 ;
        RECT 95.150 131.280 95.410 131.600 ;
        RECT 95.670 113.240 95.810 143.520 ;
        RECT 96.130 142.480 96.270 144.540 ;
        RECT 96.590 143.160 96.730 144.540 ;
        RECT 96.530 142.840 96.790 143.160 ;
        RECT 96.070 142.160 96.330 142.480 ;
        RECT 96.590 142.140 96.730 142.840 ;
        RECT 97.050 142.480 97.190 164.180 ;
        RECT 97.510 162.880 97.650 171.740 ;
        RECT 97.910 170.040 98.170 170.360 ;
        RECT 97.450 162.560 97.710 162.880 ;
        RECT 97.970 162.540 98.110 170.040 ;
        RECT 98.430 164.580 98.570 172.850 ;
        RECT 99.350 172.400 99.490 186.020 ;
        RECT 101.130 185.340 101.390 185.660 ;
        RECT 101.590 185.340 101.850 185.660 ;
        RECT 100.210 182.620 100.470 182.940 ;
        RECT 100.270 181.580 100.410 182.620 ;
        RECT 101.190 181.580 101.330 185.340 ;
        RECT 100.210 181.260 100.470 181.580 ;
        RECT 101.130 181.260 101.390 181.580 ;
        RECT 100.270 178.180 100.410 181.260 ;
        RECT 101.650 178.180 101.790 185.340 ;
        RECT 107.510 184.805 109.390 185.175 ;
        RECT 110.850 183.960 110.990 191.800 ;
        RECT 110.790 183.640 111.050 183.960 ;
        RECT 109.870 182.960 110.130 183.280 ;
        RECT 104.350 179.900 104.610 180.220 ;
        RECT 105.270 179.900 105.530 180.220 ;
        RECT 104.410 178.180 104.550 179.900 ;
        RECT 105.330 179.200 105.470 179.900 ;
        RECT 107.510 179.365 109.390 179.735 ;
        RECT 109.930 179.200 110.070 182.960 ;
        RECT 110.850 181.240 110.990 183.640 ;
        RECT 110.790 180.920 111.050 181.240 ;
        RECT 110.850 180.480 110.990 180.920 ;
        RECT 110.850 180.340 111.910 180.480 ;
        RECT 105.270 178.880 105.530 179.200 ;
        RECT 109.870 178.880 110.130 179.200 ;
        RECT 100.210 177.860 100.470 178.180 ;
        RECT 101.590 177.860 101.850 178.180 ;
        RECT 104.350 177.860 104.610 178.180 ;
        RECT 99.750 175.480 100.010 175.800 ;
        RECT 99.810 173.760 99.950 175.480 ;
        RECT 109.870 174.460 110.130 174.780 ;
        RECT 107.510 173.925 109.390 174.295 ;
        RECT 99.750 173.440 100.010 173.760 ;
        RECT 109.930 173.080 110.070 174.460 ;
        RECT 109.870 172.760 110.130 173.080 ;
        RECT 111.770 172.740 111.910 180.340 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 101.130 172.420 101.390 172.740 ;
        RECT 111.710 172.420 111.970 172.740 ;
        RECT 99.290 172.080 99.550 172.400 ;
        RECT 100.670 171.740 100.930 172.060 ;
        RECT 98.370 164.260 98.630 164.580 ;
        RECT 97.910 162.220 98.170 162.540 ;
        RECT 98.430 162.200 98.570 164.260 ;
        RECT 99.750 163.580 100.010 163.900 ;
        RECT 98.370 161.880 98.630 162.200 ;
        RECT 99.810 161.860 99.950 163.580 ;
        RECT 100.730 162.200 100.870 171.740 ;
        RECT 101.190 171.040 101.330 172.420 ;
        RECT 101.130 170.720 101.390 171.040 ;
        RECT 106.650 170.720 106.910 171.040 ;
        RECT 101.130 169.020 101.390 169.340 ;
        RECT 102.050 169.020 102.310 169.340 ;
        RECT 101.190 166.960 101.330 169.020 ;
        RECT 101.130 166.640 101.390 166.960 ;
        RECT 102.110 165.260 102.250 169.020 ;
        RECT 106.710 167.300 106.850 170.720 ;
        RECT 107.110 170.380 107.370 170.700 ;
        RECT 109.870 170.380 110.130 170.700 ;
        RECT 107.170 168.320 107.310 170.380 ;
        RECT 107.510 168.485 109.390 168.855 ;
        RECT 109.930 168.320 110.070 170.380 ;
        RECT 111.770 170.020 111.910 172.420 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 111.710 169.700 111.970 170.020 ;
        RECT 107.110 168.000 107.370 168.320 ;
        RECT 109.870 168.000 110.130 168.320 ;
        RECT 107.570 167.660 107.830 167.980 ;
        RECT 106.650 166.980 106.910 167.300 ;
        RECT 104.810 166.640 105.070 166.960 ;
        RECT 104.870 165.600 105.010 166.640 ;
        RECT 104.810 165.280 105.070 165.600 ;
        RECT 102.050 164.940 102.310 165.260 ;
        RECT 101.590 164.260 101.850 164.580 ;
        RECT 101.650 162.200 101.790 164.260 ;
        RECT 100.670 161.880 100.930 162.200 ;
        RECT 101.590 161.880 101.850 162.200 ;
        RECT 99.750 161.540 100.010 161.860 ;
        RECT 102.110 161.180 102.250 164.940 ;
        RECT 107.630 164.320 107.770 167.660 ;
        RECT 111.770 167.640 111.910 169.700 ;
        RECT 113.540 168.145 113.820 168.515 ;
        RECT 111.710 167.320 111.970 167.640 ;
        RECT 110.790 166.980 111.050 167.300 ;
        RECT 107.170 164.180 107.770 164.320 ;
        RECT 102.510 162.220 102.770 162.540 ;
        RECT 102.050 160.860 102.310 161.180 ;
        RECT 99.290 158.480 99.550 158.800 ;
        RECT 97.910 156.330 98.170 156.420 ;
        RECT 97.910 156.190 98.570 156.330 ;
        RECT 97.910 156.100 98.170 156.190 ;
        RECT 97.450 155.760 97.710 156.080 ;
        RECT 97.510 152.000 97.650 155.760 ;
        RECT 98.430 152.930 98.570 156.190 ;
        RECT 98.830 156.100 99.090 156.420 ;
        RECT 98.890 153.700 99.030 156.100 ;
        RECT 98.830 153.380 99.090 153.700 ;
        RECT 98.430 152.790 99.030 152.930 ;
        RECT 97.450 151.680 97.710 152.000 ;
        RECT 98.370 151.680 98.630 152.000 ;
        RECT 97.450 150.660 97.710 150.980 ;
        RECT 97.510 147.580 97.650 150.660 ;
        RECT 98.430 148.940 98.570 151.680 ;
        RECT 98.890 151.515 99.030 152.790 ;
        RECT 98.820 151.145 99.100 151.515 ;
        RECT 98.830 151.000 99.090 151.145 ;
        RECT 98.830 149.980 99.090 150.300 ;
        RECT 97.900 148.425 98.180 148.795 ;
        RECT 98.370 148.620 98.630 148.940 ;
        RECT 97.970 148.260 98.110 148.425 ;
        RECT 97.910 147.940 98.170 148.260 ;
        RECT 98.370 147.600 98.630 147.920 ;
        RECT 97.450 147.260 97.710 147.580 ;
        RECT 97.910 147.260 98.170 147.580 ;
        RECT 96.990 142.160 97.250 142.480 ;
        RECT 96.530 141.820 96.790 142.140 ;
        RECT 97.450 141.820 97.710 142.140 ;
        RECT 96.070 140.120 96.330 140.440 ;
        RECT 96.130 138.400 96.270 140.120 ;
        RECT 96.990 139.100 97.250 139.420 ;
        RECT 96.070 138.080 96.330 138.400 ;
        RECT 96.530 137.060 96.790 137.380 ;
        RECT 96.590 135.680 96.730 137.060 ;
        RECT 96.530 135.360 96.790 135.680 ;
        RECT 97.050 134.660 97.190 139.100 ;
        RECT 96.990 134.340 97.250 134.660 ;
        RECT 97.510 132.960 97.650 141.820 ;
        RECT 97.970 132.960 98.110 147.260 ;
        RECT 98.430 140.440 98.570 147.600 ;
        RECT 98.890 146.220 99.030 149.980 ;
        RECT 98.830 145.900 99.090 146.220 ;
        RECT 98.890 143.500 99.030 145.900 ;
        RECT 99.350 143.500 99.490 158.480 ;
        RECT 100.670 156.100 100.930 156.420 ;
        RECT 100.210 155.420 100.470 155.740 ;
        RECT 100.270 154.720 100.410 155.420 ;
        RECT 100.210 154.400 100.470 154.720 ;
        RECT 99.750 152.700 100.010 153.020 ;
        RECT 99.810 151.230 99.950 152.700 ;
        RECT 99.810 151.090 100.410 151.230 ;
        RECT 100.270 150.300 100.410 151.090 ;
        RECT 100.210 149.980 100.470 150.300 ;
        RECT 100.270 148.940 100.410 149.980 ;
        RECT 100.210 148.620 100.470 148.940 ;
        RECT 100.210 148.170 100.470 148.260 ;
        RECT 100.730 148.170 100.870 156.100 ;
        RECT 102.110 153.360 102.250 160.860 ;
        RECT 102.570 156.420 102.710 162.220 ;
        RECT 107.170 161.860 107.310 164.180 ;
        RECT 107.510 163.045 109.390 163.415 ;
        RECT 110.850 162.880 110.990 166.980 ;
        RECT 110.790 162.560 111.050 162.880 ;
        RECT 107.110 161.540 107.370 161.860 ;
        RECT 105.730 161.200 105.990 161.520 ;
        RECT 102.970 158.820 103.230 159.140 ;
        RECT 104.350 158.820 104.610 159.140 ;
        RECT 103.030 156.420 103.170 158.820 ;
        RECT 102.510 156.100 102.770 156.420 ;
        RECT 102.970 156.100 103.230 156.420 ;
        RECT 103.890 155.760 104.150 156.080 ;
        RECT 102.050 153.040 102.310 153.360 ;
        RECT 103.950 151.660 104.090 155.760 ;
        RECT 101.120 151.145 101.400 151.515 ;
        RECT 103.890 151.340 104.150 151.660 ;
        RECT 100.210 148.030 100.870 148.170 ;
        RECT 100.210 147.940 100.470 148.030 ;
        RECT 99.750 147.260 100.010 147.580 ;
        RECT 98.830 143.180 99.090 143.500 ;
        RECT 99.290 143.180 99.550 143.500 ;
        RECT 98.830 142.500 99.090 142.820 ;
        RECT 98.890 140.780 99.030 142.500 ;
        RECT 98.830 140.460 99.090 140.780 ;
        RECT 98.370 140.120 98.630 140.440 ;
        RECT 98.430 137.720 98.570 140.120 ;
        RECT 98.370 137.400 98.630 137.720 ;
        RECT 97.450 132.640 97.710 132.960 ;
        RECT 97.910 132.640 98.170 132.960 ;
        RECT 98.430 129.560 98.570 137.400 ;
        RECT 99.810 132.360 99.950 147.260 ;
        RECT 100.270 146.560 100.410 147.940 ;
        RECT 100.210 146.240 100.470 146.560 ;
        RECT 101.190 145.540 101.330 151.145 ;
        RECT 102.050 150.660 102.310 150.980 ;
        RECT 102.110 148.260 102.250 150.660 ;
        RECT 103.890 150.320 104.150 150.640 ;
        RECT 103.950 149.280 104.090 150.320 ;
        RECT 103.890 148.960 104.150 149.280 ;
        RECT 102.050 147.940 102.310 148.260 ;
        RECT 102.110 146.220 102.250 147.940 ;
        RECT 102.050 145.900 102.310 146.220 ;
        RECT 101.130 145.220 101.390 145.540 ;
        RECT 100.210 144.540 100.470 144.860 ;
        RECT 100.270 143.500 100.410 144.540 ;
        RECT 100.210 143.180 100.470 143.500 ;
        RECT 101.590 141.820 101.850 142.140 ;
        RECT 101.650 139.760 101.790 141.820 ;
        RECT 101.590 139.440 101.850 139.760 ;
        RECT 102.110 138.400 102.250 145.900 ;
        RECT 103.950 145.540 104.090 148.960 ;
        RECT 103.890 145.220 104.150 145.540 ;
        RECT 102.970 144.540 103.230 144.860 ;
        RECT 103.030 143.500 103.170 144.540 ;
        RECT 102.970 143.180 103.230 143.500 ;
        RECT 102.510 140.460 102.770 140.780 ;
        RECT 102.570 138.400 102.710 140.460 ;
        RECT 103.030 138.400 103.170 143.180 ;
        RECT 102.050 138.080 102.310 138.400 ;
        RECT 102.510 138.080 102.770 138.400 ;
        RECT 102.970 138.080 103.230 138.400 ;
        RECT 104.410 135.000 104.550 158.820 ;
        RECT 105.790 156.420 105.930 161.200 ;
        RECT 107.170 160.160 107.310 161.540 ;
        RECT 107.110 159.840 107.370 160.160 ;
        RECT 107.510 157.605 109.390 157.975 ;
        RECT 105.730 156.100 105.990 156.420 ;
        RECT 107.110 156.100 107.370 156.420 ;
        RECT 104.810 155.420 105.070 155.740 ;
        RECT 106.190 155.420 106.450 155.740 ;
        RECT 104.870 154.380 105.010 155.420 ;
        RECT 104.810 154.060 105.070 154.380 ;
        RECT 105.730 151.680 105.990 152.000 ;
        RECT 105.790 150.040 105.930 151.680 ;
        RECT 106.250 150.640 106.390 155.420 ;
        RECT 106.190 150.320 106.450 150.640 ;
        RECT 105.790 149.900 106.390 150.040 ;
        RECT 105.730 145.220 105.990 145.540 ;
        RECT 105.790 143.160 105.930 145.220 ;
        RECT 105.730 142.840 105.990 143.160 ;
        RECT 104.350 134.680 104.610 135.000 ;
        RECT 99.810 132.220 100.410 132.360 ;
        RECT 101.590 132.300 101.850 132.620 ;
        RECT 99.750 131.620 100.010 131.940 ;
        RECT 98.830 131.280 99.090 131.600 ;
        RECT 98.370 129.240 98.630 129.560 ;
        RECT 98.430 126.500 98.570 129.240 ;
        RECT 98.370 126.180 98.630 126.500 ;
        RECT 97.910 125.500 98.170 125.820 ;
        RECT 97.970 124.460 98.110 125.500 ;
        RECT 97.910 124.140 98.170 124.460 ;
        RECT 98.430 124.120 98.570 126.180 ;
        RECT 98.890 125.820 99.030 131.280 ;
        RECT 99.290 130.940 99.550 131.260 ;
        RECT 99.350 129.560 99.490 130.940 ;
        RECT 99.290 129.240 99.550 129.560 ;
        RECT 98.830 125.500 99.090 125.820 ;
        RECT 98.370 123.800 98.630 124.120 ;
        RECT 99.350 122.080 99.490 129.240 ;
        RECT 99.810 128.540 99.950 131.620 ;
        RECT 99.750 128.220 100.010 128.540 ;
        RECT 99.290 121.760 99.550 122.080 ;
        RECT 96.070 120.060 96.330 120.380 ;
        RECT 99.750 120.060 100.010 120.380 ;
        RECT 96.130 115.960 96.270 120.060 ;
        RECT 98.370 118.020 98.630 118.340 ;
        RECT 98.430 116.640 98.570 118.020 ;
        RECT 99.810 118.000 99.950 120.060 ;
        RECT 99.750 117.680 100.010 118.000 ;
        RECT 98.370 116.320 98.630 116.640 ;
        RECT 96.070 115.640 96.330 115.960 ;
        RECT 96.990 113.600 97.250 113.920 ;
        RECT 96.530 113.260 96.790 113.580 ;
        RECT 95.610 112.920 95.870 113.240 ;
        RECT 85.490 112.580 85.750 112.900 ;
        RECT 94.690 112.580 94.950 112.900 ;
        RECT 83.650 111.900 83.910 112.220 ;
        RECT 89.170 111.900 89.430 112.220 ;
        RECT 83.710 111.200 83.850 111.900 ;
        RECT 83.650 110.880 83.910 111.200 ;
        RECT 84.570 110.540 84.830 110.860 ;
        RECT 73.070 110.200 73.330 110.520 ;
        RECT 73.530 110.200 73.790 110.520 ;
        RECT 80.430 110.200 80.690 110.520 ;
        RECT 73.130 107.800 73.270 110.200 ;
        RECT 79.510 109.180 79.770 109.500 ;
        RECT 77.510 108.645 79.390 109.015 ;
        RECT 79.570 107.800 79.710 109.180 ;
        RECT 73.070 107.480 73.330 107.800 ;
        RECT 79.510 107.480 79.770 107.800 ;
        RECT 75.830 106.800 76.090 107.120 ;
        RECT 78.590 106.800 78.850 107.120 ;
        RECT 65.250 105.100 65.510 105.420 ;
        RECT 71.690 105.100 71.950 105.420 ;
        RECT 70.310 104.420 70.570 104.740 ;
        RECT 70.370 92.720 70.510 104.420 ;
        RECT 75.890 92.720 76.030 106.800 ;
        RECT 78.650 105.760 78.790 106.800 ;
        RECT 78.590 105.440 78.850 105.760 ;
        RECT 80.490 104.580 80.630 110.200 ;
        RECT 83.650 109.860 83.910 110.180 ;
        RECT 83.710 107.800 83.850 109.860 ;
        RECT 84.630 108.480 84.770 110.540 ;
        RECT 84.570 108.160 84.830 108.480 ;
        RECT 89.230 107.800 89.370 111.900 ;
        RECT 92.510 111.365 94.390 111.735 ;
        RECT 91.930 110.200 92.190 110.520 ;
        RECT 91.470 109.860 91.730 110.180 ;
        RECT 83.650 107.480 83.910 107.800 ;
        RECT 89.170 107.480 89.430 107.800 ;
        RECT 85.950 107.140 86.210 107.460 ;
        RECT 86.010 105.080 86.150 107.140 ;
        RECT 86.870 106.800 87.130 107.120 ;
        RECT 85.950 104.760 86.210 105.080 ;
        RECT 80.490 104.440 81.550 104.580 ;
        RECT 77.510 103.205 79.390 103.575 ;
        RECT 81.410 92.720 81.550 104.440 ;
        RECT 86.930 92.720 87.070 106.800 ;
        RECT 91.530 101.760 91.670 109.860 ;
        RECT 91.990 105.760 92.130 110.200 ;
        RECT 92.510 105.925 94.390 106.295 ;
        RECT 91.930 105.440 92.190 105.760 ;
        RECT 96.590 104.060 96.730 113.260 ;
        RECT 97.050 107.120 97.190 113.600 ;
        RECT 100.270 112.560 100.410 132.220 ;
        RECT 101.650 130.240 101.790 132.300 ;
        RECT 104.410 131.940 104.550 134.680 ;
        RECT 105.270 131.960 105.530 132.280 ;
        RECT 104.350 131.620 104.610 131.940 ;
        RECT 101.590 129.920 101.850 130.240 ;
        RECT 101.130 128.900 101.390 129.220 ;
        RECT 101.190 124.120 101.330 128.900 ;
        RECT 102.050 128.220 102.310 128.540 ;
        RECT 102.110 124.120 102.250 128.220 ;
        RECT 104.410 126.920 104.550 131.620 ;
        RECT 105.330 128.880 105.470 131.960 ;
        RECT 105.270 128.560 105.530 128.880 ;
        RECT 103.950 126.840 104.550 126.920 ;
        RECT 103.890 126.780 104.550 126.840 ;
        RECT 103.890 126.750 104.150 126.780 ;
        RECT 103.490 126.610 104.150 126.750 ;
        RECT 102.510 125.500 102.770 125.820 ;
        RECT 101.130 123.800 101.390 124.120 ;
        RECT 102.050 123.800 102.310 124.120 ;
        RECT 102.570 123.780 102.710 125.500 ;
        RECT 102.510 123.460 102.770 123.780 ;
        RECT 101.590 118.360 101.850 118.680 ;
        RECT 101.650 113.240 101.790 118.360 ;
        RECT 103.490 118.340 103.630 126.610 ;
        RECT 103.890 126.520 104.150 126.610 ;
        RECT 104.350 126.180 104.610 126.500 ;
        RECT 103.890 121.420 104.150 121.740 ;
        RECT 103.950 119.360 104.090 121.420 ;
        RECT 104.410 121.060 104.550 126.180 ;
        RECT 104.350 120.740 104.610 121.060 ;
        RECT 103.890 119.040 104.150 119.360 ;
        RECT 104.410 118.680 104.550 120.740 ;
        RECT 104.350 118.360 104.610 118.680 ;
        RECT 103.430 118.020 103.690 118.340 ;
        RECT 106.250 115.960 106.390 149.900 ;
        RECT 107.170 145.540 107.310 156.100 ;
        RECT 108.490 155.420 108.750 155.740 ;
        RECT 108.550 154.380 108.690 155.420 ;
        RECT 108.490 154.060 108.750 154.380 ;
        RECT 111.770 153.700 111.910 167.320 ;
        RECT 113.610 166.960 113.750 168.145 ;
        RECT 113.550 166.640 113.810 166.960 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 111.710 153.380 111.970 153.700 ;
        RECT 107.510 152.165 109.390 152.535 ;
        RECT 111.770 151.320 111.910 153.380 ;
        RECT 111.710 151.000 111.970 151.320 ;
        RECT 109.870 150.660 110.130 150.980 ;
        RECT 109.930 149.280 110.070 150.660 ;
        RECT 109.870 148.960 110.130 149.280 ;
        RECT 107.510 146.725 109.390 147.095 ;
        RECT 107.110 145.220 107.370 145.540 ;
        RECT 107.110 144.540 107.370 144.860 ;
        RECT 109.870 144.540 110.130 144.860 ;
        RECT 107.170 143.500 107.310 144.540 ;
        RECT 107.110 143.180 107.370 143.500 ;
        RECT 109.930 143.160 110.070 144.540 ;
        RECT 109.870 142.840 110.130 143.160 ;
        RECT 111.710 142.500 111.970 142.820 ;
        RECT 107.510 141.285 109.390 141.655 ;
        RECT 108.030 140.120 108.290 140.440 ;
        RECT 108.090 138.400 108.230 140.120 ;
        RECT 111.770 140.100 111.910 142.500 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 111.710 139.780 111.970 140.100 ;
        RECT 108.030 138.080 108.290 138.400 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 107.510 135.845 109.390 136.215 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 109.870 130.940 110.130 131.260 ;
        RECT 107.510 130.405 109.390 130.775 ;
        RECT 109.930 129.560 110.070 130.940 ;
        RECT 109.870 129.240 110.130 129.560 ;
        RECT 111.250 128.900 111.510 129.220 ;
        RECT 108.030 126.750 108.290 126.840 ;
        RECT 107.170 126.610 108.290 126.750 ;
        RECT 107.170 124.800 107.310 126.610 ;
        RECT 108.030 126.520 108.290 126.610 ;
        RECT 111.310 126.500 111.450 128.900 ;
        RECT 111.250 126.180 111.510 126.500 ;
        RECT 107.510 124.965 109.390 125.335 ;
        RECT 107.110 124.480 107.370 124.800 ;
        RECT 107.570 121.080 107.830 121.400 ;
        RECT 107.630 120.800 107.770 121.080 ;
        RECT 107.170 120.660 107.770 120.800 ;
        RECT 107.170 119.360 107.310 120.660 ;
        RECT 107.510 119.525 109.390 119.895 ;
        RECT 107.110 119.040 107.370 119.360 ;
        RECT 105.730 115.640 105.990 115.960 ;
        RECT 106.190 115.640 106.450 115.960 ;
        RECT 102.970 114.620 103.230 114.940 ;
        RECT 101.590 112.920 101.850 113.240 ;
        RECT 100.210 112.240 100.470 112.560 ;
        RECT 97.450 111.900 97.710 112.220 ;
        RECT 97.510 110.860 97.650 111.900 ;
        RECT 97.450 110.540 97.710 110.860 ;
        RECT 101.650 110.520 101.790 112.920 ;
        RECT 103.030 110.860 103.170 114.620 ;
        RECT 102.970 110.540 103.230 110.860 ;
        RECT 99.290 110.200 99.550 110.520 ;
        RECT 101.590 110.200 101.850 110.520 ;
        RECT 99.350 107.800 99.490 110.200 ;
        RECT 99.290 107.480 99.550 107.800 ;
        RECT 103.430 107.480 103.690 107.800 ;
        RECT 96.990 106.800 97.250 107.120 ;
        RECT 97.910 104.760 98.170 105.080 ;
        RECT 96.530 103.740 96.790 104.060 ;
        RECT 91.530 101.620 92.590 101.760 ;
        RECT 92.450 92.720 92.590 101.620 ;
        RECT 97.970 92.720 98.110 104.760 ;
        RECT 99.350 104.740 99.490 107.480 ;
        RECT 99.290 104.420 99.550 104.740 ;
        RECT 103.490 92.720 103.630 107.480 ;
        RECT 103.890 106.800 104.150 107.120 ;
        RECT 103.950 105.760 104.090 106.800 ;
        RECT 103.890 105.440 104.150 105.760 ;
        RECT 105.790 105.080 105.930 115.640 ;
        RECT 106.190 114.620 106.450 114.940 ;
        RECT 106.650 114.620 106.910 114.940 ;
        RECT 106.250 112.560 106.390 114.620 ;
        RECT 106.710 113.240 106.850 114.620 ;
        RECT 107.510 114.085 109.390 114.455 ;
        RECT 106.650 112.920 106.910 113.240 ;
        RECT 106.190 112.240 106.450 112.560 ;
        RECT 114.470 112.240 114.730 112.560 ;
        RECT 106.190 110.540 106.450 110.860 ;
        RECT 106.250 105.760 106.390 110.540 ;
        RECT 109.870 109.860 110.130 110.180 ;
        RECT 107.510 108.645 109.390 109.015 ;
        RECT 106.190 105.440 106.450 105.760 ;
        RECT 105.730 104.760 105.990 105.080 ;
        RECT 107.510 103.205 109.390 103.575 ;
        RECT 109.930 102.440 110.070 109.860 ;
        RECT 109.010 102.300 110.070 102.440 ;
        RECT 109.010 92.720 109.150 102.300 ;
        RECT 114.530 92.720 114.670 112.240 ;
        RECT 114.920 108.305 115.200 108.675 ;
        RECT 114.990 107.460 115.130 108.305 ;
        RECT 114.930 107.140 115.190 107.460 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 48.220 92.240 48.500 92.720 ;
        RECT 46.910 92.100 48.500 92.240 ;
        RECT 42.700 90.720 42.980 92.100 ;
        RECT 48.220 90.720 48.500 92.100 ;
        RECT 53.740 90.720 54.020 92.720 ;
        RECT 59.260 90.720 59.540 92.720 ;
        RECT 64.780 90.720 65.060 92.720 ;
        RECT 70.300 90.720 70.580 92.720 ;
        RECT 75.820 90.720 76.100 92.720 ;
        RECT 81.340 90.720 81.620 92.720 ;
        RECT 86.860 90.720 87.140 92.720 ;
        RECT 92.380 90.720 92.660 92.720 ;
        RECT 97.900 90.720 98.180 92.720 ;
        RECT 103.420 90.720 103.700 92.720 ;
        RECT 108.940 90.720 109.220 92.720 ;
        RECT 114.460 90.720 114.740 92.720 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 32.460 203.865 34.440 204.195 ;
        RECT 62.460 203.865 64.440 204.195 ;
        RECT 92.460 203.865 94.440 204.195 ;
        RECT 17.460 201.145 19.440 201.475 ;
        RECT 47.460 201.145 49.440 201.475 ;
        RECT 77.460 201.145 79.440 201.475 ;
        RECT 107.460 201.145 109.440 201.475 ;
        RECT 32.460 198.425 34.440 198.755 ;
        RECT 62.460 198.425 64.440 198.755 ;
        RECT 92.460 198.425 94.440 198.755 ;
        RECT 17.460 195.705 19.440 196.035 ;
        RECT 47.460 195.705 49.440 196.035 ;
        RECT 77.460 195.705 79.440 196.035 ;
        RECT 107.460 195.705 109.440 196.035 ;
        RECT 67.975 195.010 68.305 195.015 ;
        RECT 67.720 195.000 68.305 195.010 ;
        RECT 67.720 194.700 68.530 195.000 ;
        RECT 67.720 194.690 68.305 194.700 ;
        RECT 67.975 194.685 68.305 194.690 ;
        RECT 32.460 192.985 34.440 193.315 ;
        RECT 62.460 192.985 64.440 193.315 ;
        RECT 92.460 192.985 94.440 193.315 ;
        RECT 17.460 190.265 19.440 190.595 ;
        RECT 47.460 190.265 49.440 190.595 ;
        RECT 77.460 190.265 79.440 190.595 ;
        RECT 107.460 190.265 109.440 190.595 ;
        RECT 32.460 187.545 34.440 187.875 ;
        RECT 62.460 187.545 64.440 187.875 ;
        RECT 92.460 187.545 94.440 187.875 ;
        RECT 17.460 184.825 19.440 185.155 ;
        RECT 47.460 184.825 49.440 185.155 ;
        RECT 77.460 184.825 79.440 185.155 ;
        RECT 107.460 184.825 109.440 185.155 ;
        RECT 32.460 182.105 34.440 182.435 ;
        RECT 62.460 182.105 64.440 182.435 ;
        RECT 92.460 182.105 94.440 182.435 ;
        RECT 17.460 179.385 19.440 179.715 ;
        RECT 47.460 179.385 49.440 179.715 ;
        RECT 77.460 179.385 79.440 179.715 ;
        RECT 107.460 179.385 109.440 179.715 ;
        RECT 35.315 177.320 35.645 177.335 ;
        RECT 39.455 177.330 39.785 177.335 ;
        RECT 36.440 177.320 36.820 177.330 ;
        RECT 35.315 177.020 36.820 177.320 ;
        RECT 35.315 177.005 35.645 177.020 ;
        RECT 36.440 177.010 36.820 177.020 ;
        RECT 39.200 177.320 39.785 177.330 ;
        RECT 39.200 177.020 40.010 177.320 ;
        RECT 39.200 177.010 39.785 177.020 ;
        RECT 39.455 177.005 39.785 177.010 ;
        RECT 32.460 176.665 34.440 176.995 ;
        RECT 62.460 176.665 64.440 176.995 ;
        RECT 92.460 176.665 94.440 176.995 ;
        RECT 17.460 173.945 19.440 174.275 ;
        RECT 47.460 173.945 49.440 174.275 ;
        RECT 77.460 173.945 79.440 174.275 ;
        RECT 107.460 173.945 109.440 174.275 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 68.895 171.890 69.225 171.895 ;
        RECT 68.640 171.880 69.225 171.890 ;
        RECT 68.640 171.580 69.450 171.880 ;
        RECT 68.640 171.570 69.225 171.580 ;
        RECT 68.895 171.565 69.225 171.570 ;
        RECT 32.460 171.225 34.440 171.555 ;
        RECT 62.460 171.225 64.440 171.555 ;
        RECT 92.460 171.225 94.440 171.555 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 55.760 169.840 56.140 169.850 ;
        RECT 75.795 169.840 76.125 169.855 ;
        RECT 87.755 169.840 88.085 169.855 ;
        RECT 55.760 169.540 88.085 169.840 ;
        RECT 55.760 169.530 56.140 169.540 ;
        RECT 75.795 169.525 76.125 169.540 ;
        RECT 87.755 169.525 88.085 169.540 ;
        RECT 41.295 169.170 41.625 169.175 ;
        RECT 41.040 169.160 41.625 169.170 ;
        RECT 41.040 168.860 41.850 169.160 ;
        RECT 41.040 168.850 41.625 168.860 ;
        RECT 41.295 168.845 41.625 168.850 ;
        RECT 17.460 168.505 19.440 168.835 ;
        RECT 47.460 168.505 49.440 168.835 ;
        RECT 77.460 168.505 79.440 168.835 ;
        RECT 107.460 168.505 109.440 168.835 ;
        RECT 113.515 168.480 113.845 168.495 ;
        RECT 116.970 168.480 118.970 168.630 ;
        RECT 113.515 168.180 118.970 168.480 ;
        RECT 113.515 168.165 113.845 168.180 ;
        RECT 116.970 168.030 118.970 168.180 ;
        RECT 32.460 165.785 34.440 166.115 ;
        RECT 62.460 165.785 64.440 166.115 ;
        RECT 92.460 165.785 94.440 166.115 ;
        RECT 17.460 163.065 19.440 163.395 ;
        RECT 47.460 163.065 49.440 163.395 ;
        RECT 77.460 163.065 79.440 163.395 ;
        RECT 107.460 163.065 109.440 163.395 ;
        RECT 32.460 160.345 34.440 160.675 ;
        RECT 62.460 160.345 64.440 160.675 ;
        RECT 92.460 160.345 94.440 160.675 ;
        RECT 92.355 159.640 92.685 159.655 ;
        RECT 96.495 159.640 96.825 159.655 ;
        RECT 92.355 159.340 96.825 159.640 ;
        RECT 92.355 159.325 92.685 159.340 ;
        RECT 96.495 159.325 96.825 159.340 ;
        RECT 37.615 158.960 37.945 158.975 ;
        RECT 44.515 158.960 44.845 158.975 ;
        RECT 37.615 158.660 44.845 158.960 ;
        RECT 37.615 158.645 37.945 158.660 ;
        RECT 44.515 158.645 44.845 158.660 ;
        RECT 46.815 158.960 47.145 158.975 ;
        RECT 66.135 158.960 66.465 158.975 ;
        RECT 46.815 158.660 66.465 158.960 ;
        RECT 46.815 158.645 47.145 158.660 ;
        RECT 66.135 158.645 66.465 158.660 ;
        RECT 69.355 158.290 69.685 158.295 ;
        RECT 69.355 158.280 69.940 158.290 ;
        RECT 69.355 157.980 70.140 158.280 ;
        RECT 69.355 157.970 69.940 157.980 ;
        RECT 69.355 157.965 69.685 157.970 ;
        RECT 17.460 157.625 19.440 157.955 ;
        RECT 47.460 157.625 49.440 157.955 ;
        RECT 77.460 157.625 79.440 157.955 ;
        RECT 107.460 157.625 109.440 157.955 ;
        RECT 32.555 157.600 32.885 157.615 ;
        RECT 41.295 157.600 41.625 157.615 ;
        RECT 32.555 157.300 41.625 157.600 ;
        RECT 32.555 157.285 32.885 157.300 ;
        RECT 41.295 157.285 41.625 157.300 ;
        RECT 28.415 156.920 28.745 156.935 ;
        RECT 53.715 156.920 54.045 156.935 ;
        RECT 28.415 156.620 54.045 156.920 ;
        RECT 28.415 156.605 28.745 156.620 ;
        RECT 53.715 156.605 54.045 156.620 ;
        RECT 66.800 156.920 67.180 156.930 ;
        RECT 70.275 156.920 70.605 156.935 ;
        RECT 66.800 156.620 70.605 156.920 ;
        RECT 66.800 156.610 67.180 156.620 ;
        RECT 70.275 156.605 70.605 156.620 ;
        RECT 28.875 156.240 29.205 156.255 ;
        RECT 28.875 155.940 46.900 156.240 ;
        RECT 28.875 155.925 29.205 155.940 ;
        RECT 32.460 154.905 34.440 155.235 ;
        RECT 46.600 154.890 46.900 155.940 ;
        RECT 62.460 154.905 64.440 155.235 ;
        RECT 92.460 154.905 94.440 155.235 ;
        RECT 55.555 154.890 55.885 154.895 ;
        RECT 46.560 154.880 46.940 154.890 ;
        RECT 55.555 154.880 56.140 154.890 ;
        RECT 46.560 154.580 56.140 154.880 ;
        RECT 46.560 154.570 46.940 154.580 ;
        RECT 55.555 154.570 56.140 154.580 ;
        RECT 55.555 154.565 55.885 154.570 ;
        RECT 29.795 154.200 30.125 154.215 ;
        RECT 33.475 154.200 33.805 154.215 ;
        RECT 59.695 154.200 60.025 154.215 ;
        RECT 87.755 154.200 88.085 154.215 ;
        RECT 94.195 154.200 94.525 154.215 ;
        RECT 29.795 153.900 94.525 154.200 ;
        RECT 29.795 153.885 30.125 153.900 ;
        RECT 33.475 153.885 33.805 153.900 ;
        RECT 59.695 153.885 60.025 153.900 ;
        RECT 87.755 153.885 88.085 153.900 ;
        RECT 94.195 153.885 94.525 153.900 ;
        RECT 31.635 153.520 31.965 153.535 ;
        RECT 33.015 153.520 33.345 153.535 ;
        RECT 31.635 153.220 33.345 153.520 ;
        RECT 31.635 153.205 31.965 153.220 ;
        RECT 33.015 153.205 33.345 153.220 ;
        RECT 61.280 153.520 61.660 153.530 ;
        RECT 61.995 153.520 62.325 153.535 ;
        RECT 61.280 153.220 62.325 153.520 ;
        RECT 61.280 153.210 61.660 153.220 ;
        RECT 61.995 153.205 62.325 153.220 ;
        RECT 66.595 152.840 66.925 152.855 ;
        RECT 67.515 152.840 67.845 152.855 ;
        RECT 66.595 152.540 67.845 152.840 ;
        RECT 66.595 152.525 66.925 152.540 ;
        RECT 67.515 152.525 67.845 152.540 ;
        RECT 17.460 152.185 19.440 152.515 ;
        RECT 47.460 152.185 49.440 152.515 ;
        RECT 77.460 152.185 79.440 152.515 ;
        RECT 107.460 152.185 109.440 152.515 ;
        RECT 72.575 151.480 72.905 151.495 ;
        RECT 90.515 151.480 90.845 151.495 ;
        RECT 98.795 151.480 99.125 151.495 ;
        RECT 101.095 151.480 101.425 151.495 ;
        RECT 72.575 151.180 101.425 151.480 ;
        RECT 72.575 151.165 72.905 151.180 ;
        RECT 90.515 151.165 90.845 151.180 ;
        RECT 98.795 151.165 99.125 151.180 ;
        RECT 101.095 151.165 101.425 151.180 ;
        RECT 31.175 150.800 31.505 150.815 ;
        RECT 33.935 150.800 34.265 150.815 ;
        RECT 58.315 150.800 58.645 150.815 ;
        RECT 70.275 150.800 70.605 150.815 ;
        RECT 31.175 150.500 70.605 150.800 ;
        RECT 31.175 150.485 31.505 150.500 ;
        RECT 33.935 150.485 34.265 150.500 ;
        RECT 58.315 150.485 58.645 150.500 ;
        RECT 70.275 150.485 70.605 150.500 ;
        RECT 92.355 150.800 92.685 150.815 ;
        RECT 92.355 150.500 95.660 150.800 ;
        RECT 92.355 150.485 92.685 150.500 ;
        RECT 95.360 150.135 95.660 150.500 ;
        RECT 95.360 149.820 95.905 150.135 ;
        RECT 95.575 149.805 95.905 149.820 ;
        RECT 32.460 149.465 34.440 149.795 ;
        RECT 62.460 149.465 64.440 149.795 ;
        RECT 92.460 149.465 94.440 149.795 ;
        RECT 66.135 148.760 66.465 148.775 ;
        RECT 67.720 148.760 68.100 148.770 ;
        RECT 69.815 148.760 70.145 148.775 ;
        RECT 66.135 148.460 70.145 148.760 ;
        RECT 66.135 148.445 66.465 148.460 ;
        RECT 67.720 148.450 68.100 148.460 ;
        RECT 69.815 148.445 70.145 148.460 ;
        RECT 90.975 148.760 91.305 148.775 ;
        RECT 97.875 148.760 98.205 148.775 ;
        RECT 90.975 148.460 98.205 148.760 ;
        RECT 90.975 148.445 91.305 148.460 ;
        RECT 97.875 148.445 98.205 148.460 ;
        RECT 67.055 148.090 67.385 148.095 ;
        RECT 66.800 148.080 67.385 148.090 ;
        RECT 66.600 147.780 67.385 148.080 ;
        RECT 66.800 147.770 67.385 147.780 ;
        RECT 67.055 147.765 67.385 147.770 ;
        RECT 17.460 146.745 19.440 147.075 ;
        RECT 47.460 146.745 49.440 147.075 ;
        RECT 77.460 146.745 79.440 147.075 ;
        RECT 107.460 146.745 109.440 147.075 ;
        RECT 32.460 144.025 34.440 144.355 ;
        RECT 62.460 144.025 64.440 144.355 ;
        RECT 92.460 144.025 94.440 144.355 ;
        RECT 17.460 141.305 19.440 141.635 ;
        RECT 47.460 141.305 49.440 141.635 ;
        RECT 77.460 141.305 79.440 141.635 ;
        RECT 107.460 141.305 109.440 141.635 ;
        RECT 32.460 138.585 34.440 138.915 ;
        RECT 62.460 138.585 64.440 138.915 ;
        RECT 92.460 138.585 94.440 138.915 ;
        RECT 38.995 138.570 39.325 138.575 ;
        RECT 69.355 138.570 69.685 138.575 ;
        RECT 38.995 138.560 39.580 138.570 ;
        RECT 69.355 138.560 69.940 138.570 ;
        RECT 116.970 138.560 118.970 138.710 ;
        RECT 38.995 138.260 39.780 138.560 ;
        RECT 69.130 138.260 69.940 138.560 ;
        RECT 38.995 138.250 39.580 138.260 ;
        RECT 69.355 138.250 69.940 138.260 ;
        RECT 105.020 138.260 118.970 138.560 ;
        RECT 38.995 138.245 39.325 138.250 ;
        RECT 69.355 138.245 69.685 138.250 ;
        RECT 36.440 137.880 36.820 137.890 ;
        RECT 37.615 137.880 37.945 137.895 ;
        RECT 36.440 137.580 37.945 137.880 ;
        RECT 36.440 137.570 36.820 137.580 ;
        RECT 37.615 137.565 37.945 137.580 ;
        RECT 61.280 137.880 61.660 137.890 ;
        RECT 105.020 137.880 105.320 138.260 ;
        RECT 116.970 138.110 118.970 138.260 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 61.280 137.580 105.320 137.880 ;
        RECT 61.280 137.570 61.660 137.580 ;
        RECT 17.460 135.865 19.440 136.195 ;
        RECT 47.460 135.865 49.440 136.195 ;
        RECT 77.460 135.865 79.440 136.195 ;
        RECT 107.460 135.865 109.440 136.195 ;
        RECT 45.435 134.480 45.765 134.495 ;
        RECT 49.115 134.480 49.445 134.495 ;
        RECT 67.975 134.480 68.305 134.495 ;
        RECT 45.435 134.180 68.305 134.480 ;
        RECT 45.435 134.165 45.765 134.180 ;
        RECT 49.115 134.165 49.445 134.180 ;
        RECT 67.975 134.165 68.305 134.180 ;
        RECT 32.460 133.145 34.440 133.475 ;
        RECT 62.460 133.145 64.440 133.475 ;
        RECT 92.460 133.145 94.440 133.475 ;
        RECT 41.295 131.770 41.625 131.775 ;
        RECT 68.895 131.770 69.225 131.775 ;
        RECT 41.040 131.760 41.625 131.770 ;
        RECT 68.640 131.760 69.225 131.770 ;
        RECT 40.840 131.460 41.625 131.760 ;
        RECT 68.440 131.460 69.225 131.760 ;
        RECT 41.040 131.450 41.625 131.460 ;
        RECT 68.640 131.450 69.225 131.460 ;
        RECT 41.295 131.445 41.625 131.450 ;
        RECT 68.895 131.445 69.225 131.450 ;
        RECT 17.460 130.425 19.440 130.755 ;
        RECT 47.460 130.425 49.440 130.755 ;
        RECT 77.460 130.425 79.440 130.755 ;
        RECT 107.460 130.425 109.440 130.755 ;
        RECT 32.460 127.705 34.440 128.035 ;
        RECT 62.460 127.705 64.440 128.035 ;
        RECT 92.460 127.705 94.440 128.035 ;
        RECT 46.560 127.680 46.940 127.690 ;
        RECT 47.735 127.680 48.065 127.695 ;
        RECT 46.560 127.380 57.020 127.680 ;
        RECT 46.560 127.370 46.940 127.380 ;
        RECT 47.735 127.365 48.065 127.380 ;
        RECT 56.720 127.000 57.020 127.380 ;
        RECT 83.615 127.000 83.945 127.015 ;
        RECT 56.720 126.700 83.945 127.000 ;
        RECT 83.615 126.685 83.945 126.700 ;
        RECT 46.560 125.640 46.940 125.650 ;
        RECT 32.800 125.340 46.940 125.640 ;
        RECT 17.460 124.985 19.440 125.315 ;
        RECT 32.800 124.975 33.100 125.340 ;
        RECT 46.560 125.330 46.940 125.340 ;
        RECT 47.460 124.985 49.440 125.315 ;
        RECT 77.460 124.985 79.440 125.315 ;
        RECT 107.460 124.985 109.440 125.315 ;
        RECT 32.555 124.660 33.100 124.975 ;
        RECT 32.555 124.645 32.885 124.660 ;
        RECT 32.460 122.265 34.440 122.595 ;
        RECT 62.460 122.265 64.440 122.595 ;
        RECT 92.460 122.265 94.440 122.595 ;
        RECT 83.615 120.880 83.945 120.895 ;
        RECT 87.295 120.880 87.625 120.895 ;
        RECT 83.615 120.580 87.625 120.880 ;
        RECT 83.615 120.565 83.945 120.580 ;
        RECT 87.295 120.565 87.625 120.580 ;
        RECT 17.460 119.545 19.440 119.875 ;
        RECT 47.460 119.545 49.440 119.875 ;
        RECT 77.460 119.545 79.440 119.875 ;
        RECT 107.460 119.545 109.440 119.875 ;
        RECT 32.460 116.825 34.440 117.155 ;
        RECT 62.460 116.825 64.440 117.155 ;
        RECT 92.460 116.825 94.440 117.155 ;
        RECT 17.460 114.105 19.440 114.435 ;
        RECT 47.460 114.105 49.440 114.435 ;
        RECT 77.460 114.105 79.440 114.435 ;
        RECT 107.460 114.105 109.440 114.435 ;
        RECT 32.460 111.385 34.440 111.715 ;
        RECT 62.460 111.385 64.440 111.715 ;
        RECT 92.460 111.385 94.440 111.715 ;
        RECT 17.460 108.665 19.440 108.995 ;
        RECT 47.460 108.665 49.440 108.995 ;
        RECT 77.460 108.665 79.440 108.995 ;
        RECT 107.460 108.665 109.440 108.995 ;
        RECT 114.895 108.640 115.225 108.655 ;
        RECT 116.970 108.640 118.970 108.790 ;
        RECT 114.895 108.340 118.970 108.640 ;
        RECT 114.895 108.325 115.225 108.340 ;
        RECT 116.970 108.190 118.970 108.340 ;
        RECT 32.460 105.945 34.440 106.275 ;
        RECT 62.460 105.945 64.440 106.275 ;
        RECT 92.460 105.945 94.440 106.275 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 17.460 103.225 19.440 103.555 ;
        RECT 47.460 103.225 49.440 103.555 ;
        RECT 77.460 103.225 79.440 103.555 ;
        RECT 107.460 103.225 109.440 103.555 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 17.450 103.150 19.450 204.270 ;
        RECT 32.450 103.150 34.450 204.270 ;
        RECT 36.465 177.005 36.795 177.335 ;
        RECT 39.225 177.005 39.555 177.335 ;
        RECT 36.480 137.895 36.780 177.005 ;
        RECT 39.240 138.575 39.540 177.005 ;
        RECT 41.065 168.845 41.395 169.175 ;
        RECT 39.225 138.245 39.555 138.575 ;
        RECT 36.465 137.565 36.795 137.895 ;
        RECT 41.080 131.775 41.380 168.845 ;
        RECT 46.585 154.565 46.915 154.895 ;
        RECT 41.065 131.445 41.395 131.775 ;
        RECT 46.600 127.695 46.900 154.565 ;
        RECT 46.585 127.365 46.915 127.695 ;
        RECT 46.600 125.655 46.900 127.365 ;
        RECT 46.585 125.325 46.915 125.655 ;
        RECT 47.450 103.150 49.450 204.270 ;
        RECT 55.785 169.525 56.115 169.855 ;
        RECT 55.800 154.895 56.100 169.525 ;
        RECT 55.785 154.565 56.115 154.895 ;
        RECT 61.305 153.205 61.635 153.535 ;
        RECT 61.320 137.895 61.620 153.205 ;
        RECT 61.305 137.565 61.635 137.895 ;
        RECT 62.450 103.150 64.450 204.270 ;
        RECT 67.745 194.685 68.075 195.015 ;
        RECT 66.825 156.605 67.155 156.935 ;
        RECT 66.840 148.095 67.140 156.605 ;
        RECT 67.760 148.775 68.060 194.685 ;
        RECT 68.665 171.565 68.995 171.895 ;
        RECT 67.745 148.445 68.075 148.775 ;
        RECT 66.825 147.765 67.155 148.095 ;
        RECT 68.680 131.775 68.980 171.565 ;
        RECT 69.585 157.965 69.915 158.295 ;
        RECT 69.600 138.575 69.900 157.965 ;
        RECT 69.585 138.245 69.915 138.575 ;
        RECT 68.665 131.445 68.995 131.775 ;
        RECT 77.450 103.150 79.450 204.270 ;
        RECT 92.450 103.150 94.450 204.270 ;
        RECT 107.450 103.150 109.450 204.270 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

