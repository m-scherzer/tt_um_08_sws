VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 18.310 193.515 18.480 193.705 ;
        RECT 20.150 193.560 20.310 193.670 ;
        RECT 20.610 193.515 20.780 193.705 ;
        RECT 24.750 193.515 24.920 193.705 ;
        RECT 30.270 193.515 30.440 193.705 ;
        RECT 30.730 193.515 30.900 193.705 ;
        RECT 34.410 193.515 34.580 193.705 ;
        RECT 35.385 193.565 35.505 193.675 ;
        RECT 37.170 193.515 37.340 193.705 ;
        RECT 42.690 193.515 42.860 193.705 ;
        RECT 44.070 193.515 44.240 193.705 ;
        RECT 45.450 193.515 45.620 193.705 ;
        RECT 46.830 193.515 47.000 193.705 ;
        RECT 47.345 193.565 47.465 193.675 ;
        RECT 51.430 193.515 51.600 193.705 ;
        RECT 52.810 193.515 52.980 193.705 ;
        RECT 54.650 193.515 54.820 193.705 ;
        RECT 60.170 193.515 60.340 193.705 ;
        RECT 63.390 193.515 63.560 193.705 ;
        RECT 64.770 193.515 64.940 193.705 ;
        RECT 65.285 193.565 65.405 193.675 ;
        RECT 66.610 193.515 66.780 193.705 ;
        RECT 67.530 193.560 67.690 193.670 ;
        RECT 73.050 193.515 73.220 193.705 ;
        RECT 74.025 193.565 74.145 193.675 ;
        RECT 75.810 193.515 75.980 193.705 ;
        RECT 79.675 193.515 79.845 193.705 ;
        RECT 80.465 193.565 80.585 193.675 ;
        RECT 85.930 193.515 86.100 193.705 ;
        RECT 88.230 193.515 88.400 193.705 ;
        RECT 89.610 193.515 89.780 193.705 ;
        RECT 90.530 193.560 90.690 193.670 ;
        RECT 96.050 193.515 96.220 193.705 ;
        RECT 96.510 193.515 96.680 193.705 ;
        RECT 98.810 193.515 98.980 193.705 ;
        RECT 99.730 193.515 99.900 193.705 ;
        RECT 101.165 193.565 101.285 193.675 ;
        RECT 110.310 193.515 110.480 193.705 ;
        RECT 110.825 193.565 110.945 193.675 ;
        RECT 112.150 193.515 112.320 193.705 ;
        RECT 18.170 192.705 19.540 193.515 ;
        RECT 20.480 192.605 21.830 193.515 ;
        RECT 21.860 192.645 22.290 193.430 ;
        RECT 22.310 192.705 25.060 193.515 ;
        RECT 25.070 192.705 30.580 193.515 ;
        RECT 30.590 192.735 31.960 193.515 ;
        RECT 31.970 192.705 34.720 193.515 ;
        RECT 34.740 192.645 35.170 193.430 ;
        RECT 35.650 192.705 37.480 193.515 ;
        RECT 37.490 192.705 43.000 193.515 ;
        RECT 43.020 192.605 44.370 193.515 ;
        RECT 44.390 192.705 45.760 193.515 ;
        RECT 45.770 192.735 47.140 193.515 ;
        RECT 47.620 192.645 48.050 193.430 ;
        RECT 48.070 192.705 51.740 193.515 ;
        RECT 51.760 192.605 53.110 193.515 ;
        RECT 53.130 192.705 54.960 193.515 ;
        RECT 54.970 192.705 60.480 193.515 ;
        RECT 60.500 192.645 60.930 193.430 ;
        RECT 60.950 192.705 63.700 193.515 ;
        RECT 63.720 192.605 65.070 193.515 ;
        RECT 65.560 192.605 66.910 193.515 ;
        RECT 67.850 192.705 73.360 193.515 ;
        RECT 73.380 192.645 73.810 193.430 ;
        RECT 74.290 192.705 76.120 193.515 ;
        RECT 76.360 192.835 80.260 193.515 ;
        RECT 79.330 192.605 80.260 192.835 ;
        RECT 80.730 192.705 86.240 193.515 ;
        RECT 86.260 192.645 86.690 193.430 ;
        RECT 86.710 192.705 88.540 193.515 ;
        RECT 88.550 192.735 89.920 193.515 ;
        RECT 90.850 192.705 96.360 193.515 ;
        RECT 96.380 192.605 97.730 193.515 ;
        RECT 97.750 192.705 99.120 193.515 ;
        RECT 99.140 192.645 99.570 193.430 ;
        RECT 99.590 192.735 100.960 193.515 ;
        RECT 101.430 192.835 110.620 193.515 ;
        RECT 101.430 192.605 102.350 192.835 ;
        RECT 105.180 192.615 106.110 192.835 ;
        RECT 111.090 192.705 112.460 193.515 ;
      LAYER nwell ;
        RECT 17.975 189.485 112.655 192.315 ;
      LAYER pwell ;
        RECT 18.170 188.285 19.540 189.095 ;
        RECT 23.125 188.965 24.045 189.195 ;
        RECT 20.580 188.285 24.045 188.965 ;
        RECT 24.150 188.965 25.070 189.195 ;
        RECT 27.900 188.965 28.830 189.185 ;
        RECT 24.150 188.285 33.340 188.965 ;
        RECT 33.350 188.285 34.720 189.095 ;
        RECT 34.740 188.370 35.170 189.155 ;
        RECT 36.480 189.085 37.400 189.195 ;
        RECT 36.480 188.965 38.815 189.085 ;
        RECT 43.480 188.965 44.400 189.185 ;
        RECT 36.480 188.285 45.760 188.965 ;
        RECT 46.230 188.285 47.600 189.065 ;
        RECT 52.120 188.965 53.050 189.185 ;
        RECT 55.880 188.965 57.220 189.195 ;
        RECT 47.610 188.285 57.220 188.965 ;
        RECT 57.730 188.285 60.480 189.095 ;
        RECT 60.500 188.370 60.930 189.155 ;
        RECT 60.950 188.965 61.870 189.195 ;
        RECT 64.700 188.965 65.630 189.185 ;
        RECT 60.950 188.285 70.140 188.965 ;
        RECT 70.150 188.285 73.820 189.095 ;
        RECT 74.200 189.085 75.120 189.195 ;
        RECT 74.200 188.965 76.535 189.085 ;
        RECT 81.200 188.965 82.120 189.185 ;
        RECT 74.200 188.285 83.480 188.965 ;
        RECT 83.490 188.285 84.860 189.095 ;
        RECT 84.880 188.285 86.230 189.195 ;
        RECT 86.260 188.370 86.690 189.155 ;
        RECT 91.220 188.965 92.150 189.185 ;
        RECT 94.980 188.965 95.900 189.195 ;
        RECT 86.710 188.285 95.900 188.965 ;
        RECT 95.910 188.965 96.830 189.195 ;
        RECT 99.660 188.965 100.590 189.185 ;
        RECT 95.910 188.285 105.100 188.965 ;
        RECT 105.120 188.285 106.470 189.195 ;
        RECT 107.410 188.285 111.080 189.095 ;
        RECT 111.090 188.285 112.460 189.095 ;
        RECT 18.310 188.075 18.480 188.285 ;
        RECT 20.150 188.120 20.310 188.240 ;
        RECT 20.610 188.075 20.780 188.285 ;
        RECT 22.910 188.120 23.070 188.230 ;
        RECT 23.370 188.075 23.540 188.265 ;
        RECT 28.155 188.075 28.325 188.265 ;
        RECT 33.030 188.095 33.200 188.285 ;
        RECT 34.410 188.095 34.580 188.285 ;
        RECT 35.790 188.130 35.950 188.240 ;
        RECT 37.630 188.075 37.800 188.265 ;
        RECT 45.450 188.095 45.620 188.285 ;
        RECT 45.965 188.125 46.085 188.235 ;
        RECT 47.290 188.075 47.460 188.285 ;
        RECT 47.750 188.095 47.920 188.285 ;
        RECT 48.265 188.125 48.385 188.235 ;
        RECT 49.590 188.075 49.760 188.265 ;
        RECT 52.810 188.075 52.980 188.265 ;
        RECT 56.490 188.075 56.660 188.265 ;
        RECT 57.465 188.125 57.585 188.235 ;
        RECT 57.870 188.075 58.040 188.265 ;
        RECT 18.170 187.265 19.540 188.075 ;
        RECT 20.480 187.165 21.830 188.075 ;
        RECT 21.860 187.205 22.290 187.990 ;
        RECT 23.240 187.165 24.590 188.075 ;
        RECT 24.840 187.395 28.740 188.075 ;
        RECT 27.810 187.165 28.740 187.395 ;
        RECT 28.750 187.395 37.940 188.075 ;
        RECT 38.320 187.395 47.600 188.075 ;
        RECT 28.750 187.165 29.670 187.395 ;
        RECT 32.500 187.175 33.430 187.395 ;
        RECT 38.320 187.275 40.655 187.395 ;
        RECT 38.320 187.165 39.240 187.275 ;
        RECT 45.320 187.175 46.240 187.395 ;
        RECT 47.620 187.205 48.050 187.990 ;
        RECT 48.540 187.165 49.890 188.075 ;
        RECT 49.910 187.165 53.020 188.075 ;
        RECT 53.225 187.395 56.690 188.075 ;
        RECT 53.225 187.165 54.145 187.395 ;
        RECT 56.810 187.265 58.180 188.075 ;
        RECT 58.330 188.045 58.500 188.265 ;
        RECT 60.170 188.095 60.340 188.285 ;
        RECT 61.550 188.075 61.720 188.265 ;
        RECT 69.830 188.095 70.000 188.285 ;
        RECT 71.670 188.075 71.840 188.265 ;
        RECT 73.050 188.075 73.220 188.265 ;
        RECT 73.510 188.095 73.680 188.285 ;
        RECT 74.025 188.125 74.145 188.235 ;
        RECT 83.170 188.095 83.340 188.285 ;
        RECT 83.630 188.075 83.800 188.265 ;
        RECT 84.550 188.095 84.720 188.285 ;
        RECT 85.010 188.095 85.180 188.285 ;
        RECT 86.850 188.095 87.020 188.285 ;
        RECT 87.495 188.075 87.665 188.265 ;
        RECT 89.150 188.075 89.320 188.265 ;
        RECT 90.530 188.075 90.700 188.265 ;
        RECT 91.045 188.125 91.165 188.235 ;
        RECT 92.830 188.075 93.000 188.265 ;
        RECT 93.290 188.075 93.460 188.265 ;
        RECT 94.725 188.125 94.845 188.235 ;
        RECT 98.535 188.075 98.705 188.265 ;
        RECT 103.135 188.075 103.305 188.265 ;
        RECT 103.925 188.125 104.045 188.235 ;
        RECT 104.790 188.095 104.960 188.285 ;
        RECT 105.250 188.095 105.420 188.285 ;
        RECT 105.710 188.075 105.880 188.265 ;
        RECT 106.170 188.075 106.340 188.265 ;
        RECT 107.090 188.130 107.250 188.240 ;
        RECT 110.770 188.075 110.940 188.285 ;
        RECT 112.150 188.075 112.320 188.285 ;
        RECT 60.455 188.045 61.400 188.075 ;
        RECT 58.330 187.845 61.400 188.045 ;
        RECT 58.190 187.365 61.400 187.845 ;
        RECT 58.190 187.165 59.120 187.365 ;
        RECT 60.455 187.165 61.400 187.365 ;
        RECT 61.410 187.295 62.780 188.075 ;
        RECT 62.790 187.395 71.980 188.075 ;
        RECT 62.790 187.165 63.710 187.395 ;
        RECT 66.540 187.175 67.470 187.395 ;
        RECT 72.000 187.165 73.350 188.075 ;
        RECT 73.380 187.205 73.810 187.990 ;
        RECT 74.660 187.395 83.940 188.075 ;
        RECT 84.180 187.395 88.080 188.075 ;
        RECT 74.660 187.275 76.995 187.395 ;
        RECT 74.660 187.165 75.580 187.275 ;
        RECT 81.660 187.175 82.580 187.395 ;
        RECT 87.150 187.165 88.080 187.395 ;
        RECT 88.090 187.265 89.460 188.075 ;
        RECT 89.480 187.165 90.830 188.075 ;
        RECT 91.310 187.265 93.140 188.075 ;
        RECT 93.150 187.295 94.520 188.075 ;
        RECT 95.220 187.395 99.120 188.075 ;
        RECT 98.190 187.165 99.120 187.395 ;
        RECT 99.140 187.205 99.570 187.990 ;
        RECT 99.820 187.395 103.720 188.075 ;
        RECT 102.790 187.165 103.720 187.395 ;
        RECT 104.190 187.265 106.020 188.075 ;
        RECT 106.030 187.295 107.400 188.075 ;
        RECT 107.410 187.265 111.080 188.075 ;
        RECT 111.090 187.265 112.460 188.075 ;
      LAYER nwell ;
        RECT 17.975 184.045 112.655 186.875 ;
      LAYER pwell ;
        RECT 18.170 182.845 19.540 183.655 ;
        RECT 19.560 182.845 20.910 183.755 ;
        RECT 25.440 183.525 26.370 183.745 ;
        RECT 29.200 183.525 30.120 183.755 ;
        RECT 33.790 183.525 34.720 183.755 ;
        RECT 20.930 182.845 30.120 183.525 ;
        RECT 30.820 182.845 34.720 183.525 ;
        RECT 34.740 182.930 35.170 183.715 ;
        RECT 35.650 182.845 37.020 183.625 ;
        RECT 37.500 182.845 38.850 183.755 ;
        RECT 42.070 183.525 43.000 183.755 ;
        RECT 46.210 183.525 47.140 183.755 ;
        RECT 39.100 182.845 43.000 183.525 ;
        RECT 43.240 182.845 47.140 183.525 ;
        RECT 48.270 183.525 50.480 183.755 ;
        RECT 53.200 183.525 54.130 183.745 ;
        RECT 48.270 182.845 58.640 183.525 ;
        RECT 58.650 182.845 60.020 183.625 ;
        RECT 60.500 182.930 60.930 183.715 ;
        RECT 60.950 183.555 61.895 183.755 ;
        RECT 63.230 183.555 64.160 183.755 ;
        RECT 60.950 183.075 64.160 183.555 ;
        RECT 60.950 182.875 64.020 183.075 ;
        RECT 60.950 182.845 61.895 182.875 ;
        RECT 18.310 182.635 18.480 182.845 ;
        RECT 20.150 182.680 20.310 182.790 ;
        RECT 20.610 182.635 20.780 182.845 ;
        RECT 21.070 182.655 21.240 182.845 ;
        RECT 22.450 182.635 22.620 182.825 ;
        RECT 26.590 182.680 26.750 182.790 ;
        RECT 27.325 182.635 27.495 182.825 ;
        RECT 30.325 182.685 30.445 182.795 ;
        RECT 34.135 182.655 34.305 182.845 ;
        RECT 35.385 182.685 35.505 182.795 ;
        RECT 35.790 182.655 35.960 182.845 ;
        RECT 37.225 182.685 37.345 182.795 ;
        RECT 37.630 182.655 37.800 182.845 ;
        RECT 39.930 182.635 40.100 182.825 ;
        RECT 41.770 182.635 41.940 182.825 ;
        RECT 42.415 182.655 42.585 182.845 ;
        RECT 46.555 182.655 46.725 182.845 ;
        RECT 47.290 182.635 47.460 182.825 ;
        RECT 47.750 182.690 47.910 182.800 ;
        RECT 49.590 182.635 49.760 182.825 ;
        RECT 55.110 182.635 55.280 182.825 ;
        RECT 55.570 182.635 55.740 182.825 ;
        RECT 57.875 182.635 58.045 182.825 ;
        RECT 58.330 182.655 58.500 182.845 ;
        RECT 59.710 182.655 59.880 182.845 ;
        RECT 60.225 182.685 60.345 182.795 ;
        RECT 62.470 182.635 62.640 182.825 ;
        RECT 62.985 182.685 63.105 182.795 ;
        RECT 63.850 182.655 64.020 182.875 ;
        RECT 64.170 182.845 66.460 183.755 ;
        RECT 66.780 183.525 67.710 183.755 ;
        RECT 66.780 182.845 68.615 183.525 ;
        RECT 68.870 182.845 71.980 183.755 ;
        RECT 71.990 182.845 73.340 183.755 ;
        RECT 74.300 182.845 75.650 183.755 ;
        RECT 78.870 183.525 79.800 183.755 ;
        RECT 75.900 182.845 79.800 183.525 ;
        RECT 80.270 182.845 81.640 183.625 ;
        RECT 81.650 182.845 83.020 183.625 ;
        RECT 83.490 182.845 86.240 183.655 ;
        RECT 86.260 182.930 86.690 183.715 ;
        RECT 86.710 183.525 87.630 183.755 ;
        RECT 90.460 183.525 91.390 183.745 ;
        RECT 99.110 183.525 100.040 183.755 ;
        RECT 103.250 183.525 104.180 183.755 ;
        RECT 86.710 182.845 95.900 183.525 ;
        RECT 96.140 182.845 100.040 183.525 ;
        RECT 100.280 182.845 104.180 183.525 ;
        RECT 104.200 182.845 105.550 183.755 ;
        RECT 106.030 182.845 107.400 183.625 ;
        RECT 107.410 182.845 111.080 183.655 ;
        RECT 111.090 182.845 112.460 183.655 ;
        RECT 65.690 182.635 65.860 182.825 ;
        RECT 66.145 182.655 66.315 182.845 ;
        RECT 68.450 182.825 68.615 182.845 ;
        RECT 67.990 182.635 68.160 182.825 ;
        RECT 68.450 182.655 68.620 182.825 ;
        RECT 68.910 182.655 69.080 182.845 ;
        RECT 73.055 182.825 73.225 182.845 ;
        RECT 69.370 182.635 69.540 182.825 ;
        RECT 73.050 182.655 73.225 182.825 ;
        RECT 73.970 182.795 74.130 182.800 ;
        RECT 73.970 182.690 74.145 182.795 ;
        RECT 74.025 182.685 74.145 182.690 ;
        RECT 74.430 182.655 74.600 182.845 ;
        RECT 73.050 182.635 73.220 182.655 ;
        RECT 75.810 182.635 75.980 182.825 ;
        RECT 79.215 182.655 79.385 182.845 ;
        RECT 79.675 182.635 79.845 182.825 ;
        RECT 80.410 182.795 80.580 182.845 ;
        RECT 80.005 182.685 80.125 182.795 ;
        RECT 80.410 182.685 80.585 182.795 ;
        RECT 80.410 182.655 80.580 182.685 ;
        RECT 82.710 182.655 82.880 182.845 ;
        RECT 83.225 182.685 83.345 182.795 ;
        RECT 84.090 182.635 84.260 182.825 ;
        RECT 85.930 182.655 86.100 182.845 ;
        RECT 89.610 182.635 89.780 182.825 ;
        RECT 95.590 182.655 95.760 182.845 ;
        RECT 98.810 182.635 98.980 182.825 ;
        RECT 99.455 182.655 99.625 182.845 ;
        RECT 100.650 182.635 100.820 182.825 ;
        RECT 103.595 182.655 103.765 182.845 ;
        RECT 105.250 182.655 105.420 182.845 ;
        RECT 105.765 182.685 105.885 182.795 ;
        RECT 106.170 182.655 106.340 182.845 ;
        RECT 109.850 182.635 110.020 182.825 ;
        RECT 110.770 182.655 110.940 182.845 ;
        RECT 112.150 182.635 112.320 182.845 ;
        RECT 18.170 181.825 19.540 182.635 ;
        RECT 20.470 181.855 21.840 182.635 ;
        RECT 21.860 181.765 22.290 182.550 ;
        RECT 22.420 181.955 25.885 182.635 ;
        RECT 24.965 181.725 25.885 181.955 ;
        RECT 26.910 181.955 30.810 182.635 ;
        RECT 31.050 181.955 40.240 182.635 ;
        RECT 26.910 181.725 27.840 181.955 ;
        RECT 31.050 181.725 31.970 181.955 ;
        RECT 34.800 181.735 35.730 181.955 ;
        RECT 40.250 181.825 42.080 182.635 ;
        RECT 42.090 181.825 47.600 182.635 ;
        RECT 47.620 181.765 48.050 182.550 ;
        RECT 48.070 181.825 49.900 182.635 ;
        RECT 49.910 181.825 55.420 182.635 ;
        RECT 55.430 181.955 57.720 182.635 ;
        RECT 56.800 181.725 57.720 181.955 ;
        RECT 57.730 181.725 60.650 182.635 ;
        RECT 60.950 181.955 62.780 182.635 ;
        RECT 60.950 181.725 62.295 181.955 ;
        RECT 63.250 181.825 66.000 182.635 ;
        RECT 66.010 181.955 68.300 182.635 ;
        RECT 66.010 181.725 66.930 181.955 ;
        RECT 68.310 181.825 69.680 182.635 ;
        RECT 69.690 181.825 73.360 182.635 ;
        RECT 73.380 181.765 73.810 182.550 ;
        RECT 74.290 181.825 76.120 182.635 ;
        RECT 76.360 181.955 80.260 182.635 ;
        RECT 79.330 181.725 80.260 181.955 ;
        RECT 80.730 181.825 84.400 182.635 ;
        RECT 84.410 181.825 89.920 182.635 ;
        RECT 89.930 181.955 99.120 182.635 ;
        RECT 89.930 181.725 90.850 181.955 ;
        RECT 93.680 181.735 94.610 181.955 ;
        RECT 99.140 181.765 99.570 182.550 ;
        RECT 99.590 181.855 100.960 182.635 ;
        RECT 100.970 181.955 110.160 182.635 ;
        RECT 100.970 181.725 101.890 181.955 ;
        RECT 104.720 181.735 105.650 181.955 ;
        RECT 111.090 181.825 112.460 182.635 ;
      LAYER nwell ;
        RECT 17.975 178.605 112.655 181.435 ;
      LAYER pwell ;
        RECT 18.170 177.405 19.540 178.215 ;
        RECT 20.010 178.085 20.930 178.315 ;
        RECT 23.760 178.085 24.690 178.305 ;
        RECT 20.010 177.405 29.200 178.085 ;
        RECT 29.210 177.405 30.580 178.185 ;
        RECT 33.790 178.085 34.720 178.315 ;
        RECT 30.820 177.405 34.720 178.085 ;
        RECT 34.740 177.490 35.170 178.275 ;
        RECT 35.200 177.405 36.550 178.315 ;
        RECT 37.030 177.405 38.400 178.185 ;
        RECT 38.410 177.405 39.780 178.185 ;
        RECT 39.790 177.405 43.460 178.215 ;
        RECT 43.480 177.405 44.830 178.315 ;
        RECT 45.220 178.205 46.140 178.315 ;
        RECT 45.220 178.085 47.555 178.205 ;
        RECT 52.220 178.085 53.140 178.305 ;
        RECT 45.220 177.405 54.500 178.085 ;
        RECT 54.970 177.405 56.800 178.215 ;
        RECT 59.550 178.085 60.480 178.315 ;
        RECT 56.810 177.405 60.480 178.085 ;
        RECT 60.500 177.490 60.930 178.275 ;
        RECT 60.950 177.405 62.780 178.085 ;
        RECT 63.250 177.405 66.920 178.215 ;
        RECT 66.940 177.405 68.290 178.315 ;
        RECT 68.320 177.405 69.670 178.315 ;
        RECT 69.690 177.405 72.300 178.315 ;
        RECT 72.460 177.405 73.810 178.315 ;
        RECT 73.830 178.085 74.750 178.315 ;
        RECT 77.580 178.085 78.510 178.305 ;
        RECT 73.830 177.405 83.020 178.085 ;
        RECT 83.030 177.405 84.400 178.215 ;
        RECT 84.420 177.405 85.770 178.315 ;
        RECT 86.260 177.490 86.690 178.275 ;
        RECT 86.720 177.405 88.070 178.315 ;
        RECT 88.090 177.405 89.460 178.185 ;
        RECT 93.590 178.085 94.520 178.315 ;
        RECT 90.620 177.405 94.520 178.085 ;
        RECT 95.000 177.405 96.350 178.315 ;
        RECT 96.830 177.405 102.340 178.215 ;
        RECT 102.360 177.405 103.710 178.315 ;
        RECT 103.730 177.405 105.560 178.215 ;
        RECT 105.570 177.405 106.940 178.185 ;
        RECT 107.410 177.405 111.080 178.215 ;
        RECT 111.090 177.405 112.460 178.215 ;
        RECT 18.310 177.195 18.480 177.405 ;
        RECT 19.745 177.245 19.865 177.355 ;
        RECT 21.530 177.195 21.700 177.385 ;
        RECT 23.830 177.195 24.000 177.385 ;
        RECT 27.695 177.195 27.865 177.385 ;
        RECT 28.890 177.215 29.060 177.405 ;
        RECT 30.270 177.215 30.440 177.405 ;
        RECT 34.135 177.215 34.305 177.405 ;
        RECT 36.250 177.215 36.420 177.405 ;
        RECT 36.765 177.245 36.885 177.355 ;
        RECT 37.170 177.215 37.340 177.405 ;
        RECT 37.630 177.195 37.800 177.385 ;
        RECT 38.090 177.195 38.260 177.385 ;
        RECT 39.470 177.215 39.640 177.405 ;
        RECT 43.150 177.215 43.320 177.405 ;
        RECT 44.530 177.215 44.700 177.405 ;
        RECT 51.615 177.195 51.785 177.385 ;
        RECT 52.350 177.195 52.520 177.385 ;
        RECT 54.190 177.215 54.360 177.405 ;
        RECT 54.705 177.245 54.825 177.355 ;
        RECT 56.490 177.215 56.660 177.405 ;
        RECT 56.950 177.195 57.120 177.405 ;
        RECT 58.790 177.195 58.960 177.385 ;
        RECT 59.250 177.195 59.420 177.385 ;
        RECT 61.090 177.215 61.260 177.405 ;
        RECT 62.985 177.245 63.105 177.355 ;
        RECT 66.610 177.215 66.780 177.405 ;
        RECT 67.990 177.215 68.160 177.405 ;
        RECT 68.450 177.215 68.620 177.405 ;
        RECT 69.835 177.215 70.005 177.405 ;
        RECT 72.590 177.195 72.760 177.385 ;
        RECT 73.105 177.245 73.225 177.355 ;
        RECT 73.510 177.215 73.680 177.405 ;
        RECT 74.025 177.245 74.145 177.355 ;
        RECT 79.490 177.195 79.660 177.385 ;
        RECT 79.950 177.195 80.120 177.385 ;
        RECT 81.385 177.245 81.505 177.355 ;
        RECT 82.710 177.215 82.880 177.405 ;
        RECT 84.090 177.215 84.260 177.405 ;
        RECT 85.470 177.215 85.640 177.405 ;
        RECT 85.985 177.245 86.105 177.355 ;
        RECT 86.850 177.215 87.020 177.405 ;
        RECT 88.230 177.215 88.400 177.405 ;
        RECT 90.070 177.250 90.230 177.360 ;
        RECT 90.530 177.195 90.700 177.385 ;
        RECT 91.910 177.195 92.080 177.385 ;
        RECT 93.935 177.215 94.105 177.405 ;
        RECT 94.725 177.245 94.845 177.355 ;
        RECT 96.050 177.215 96.220 177.405 ;
        RECT 96.565 177.245 96.685 177.355 ;
        RECT 97.430 177.195 97.600 177.385 ;
        RECT 97.890 177.195 98.060 177.385 ;
        RECT 99.785 177.245 99.905 177.355 ;
        RECT 102.030 177.215 102.200 177.405 ;
        RECT 102.490 177.215 102.660 177.405 ;
        RECT 105.250 177.215 105.420 177.405 ;
        RECT 105.710 177.215 105.880 177.405 ;
        RECT 107.145 177.245 107.265 177.355 ;
        RECT 108.930 177.195 109.100 177.385 ;
        RECT 110.770 177.195 110.940 177.405 ;
        RECT 112.150 177.195 112.320 177.405 ;
        RECT 18.170 176.385 19.540 177.195 ;
        RECT 20.010 176.385 21.840 177.195 ;
        RECT 21.860 176.325 22.290 177.110 ;
        RECT 22.310 176.385 24.140 177.195 ;
        RECT 24.380 176.515 28.280 177.195 ;
        RECT 27.350 176.285 28.280 176.515 ;
        RECT 28.660 176.515 37.940 177.195 ;
        RECT 37.950 176.515 47.230 177.195 ;
        RECT 28.660 176.395 30.995 176.515 ;
        RECT 28.660 176.285 29.580 176.395 ;
        RECT 35.660 176.295 36.580 176.515 ;
        RECT 39.310 176.295 40.230 176.515 ;
        RECT 44.895 176.395 47.230 176.515 ;
        RECT 46.310 176.285 47.230 176.395 ;
        RECT 47.620 176.325 48.050 177.110 ;
        RECT 48.300 176.515 52.200 177.195 ;
        RECT 51.270 176.285 52.200 176.515 ;
        RECT 52.210 176.415 53.580 177.195 ;
        RECT 53.590 176.385 57.260 177.195 ;
        RECT 57.270 176.515 59.100 177.195 ;
        RECT 59.110 176.965 60.680 177.195 ;
        RECT 62.770 177.155 63.690 177.195 ;
        RECT 62.770 176.965 63.700 177.155 ;
        RECT 59.110 176.605 63.700 176.965 ;
        RECT 59.110 176.515 63.690 176.605 ;
        RECT 57.270 176.285 58.615 176.515 ;
        RECT 60.690 176.285 63.690 176.515 ;
        RECT 63.710 176.515 72.900 177.195 ;
        RECT 63.710 176.285 64.630 176.515 ;
        RECT 67.460 176.295 68.390 176.515 ;
        RECT 73.380 176.325 73.810 177.110 ;
        RECT 74.290 176.385 79.800 177.195 ;
        RECT 79.810 176.415 81.180 177.195 ;
        RECT 81.650 176.515 90.840 177.195 ;
        RECT 81.650 176.285 82.570 176.515 ;
        RECT 85.400 176.295 86.330 176.515 ;
        RECT 90.850 176.385 92.220 177.195 ;
        RECT 92.230 176.385 97.740 177.195 ;
        RECT 97.760 176.285 99.110 177.195 ;
        RECT 99.140 176.325 99.570 177.110 ;
        RECT 100.050 176.515 109.240 177.195 ;
        RECT 100.050 176.285 100.970 176.515 ;
        RECT 103.800 176.295 104.730 176.515 ;
        RECT 109.250 176.385 111.080 177.195 ;
        RECT 111.090 176.385 112.460 177.195 ;
      LAYER nwell ;
        RECT 17.975 173.165 112.655 175.995 ;
      LAYER pwell ;
        RECT 18.170 171.965 19.540 172.775 ;
        RECT 20.010 171.965 22.760 172.775 ;
        RECT 25.425 172.645 26.345 172.875 ;
        RECT 22.880 171.965 26.345 172.645 ;
        RECT 26.910 171.965 30.580 172.775 ;
        RECT 33.790 172.645 34.720 172.875 ;
        RECT 30.820 171.965 34.720 172.645 ;
        RECT 34.740 172.050 35.170 172.835 ;
        RECT 35.650 171.965 38.400 172.775 ;
        RECT 38.420 171.965 39.770 172.875 ;
        RECT 40.710 171.965 44.380 172.775 ;
        RECT 44.390 171.965 45.760 172.745 ;
        RECT 45.770 172.645 46.700 172.875 ;
        RECT 45.770 171.965 49.670 172.645 ;
        RECT 49.920 171.965 51.270 172.875 ;
        RECT 51.290 171.965 54.960 172.775 ;
        RECT 54.970 171.965 60.480 172.775 ;
        RECT 60.500 172.050 60.930 172.835 ;
        RECT 61.165 172.195 63.920 172.875 ;
        RECT 61.650 171.965 63.920 172.195 ;
        RECT 64.170 171.965 66.920 172.775 ;
        RECT 66.930 171.965 69.670 172.645 ;
        RECT 69.690 171.965 72.430 172.645 ;
        RECT 72.910 171.965 75.520 172.875 ;
        RECT 75.680 171.965 77.030 172.875 ;
        RECT 77.050 172.645 77.970 172.875 ;
        RECT 80.800 172.645 81.730 172.865 ;
        RECT 77.050 171.965 86.240 172.645 ;
        RECT 86.260 172.050 86.690 172.835 ;
        RECT 86.720 171.965 88.070 172.875 ;
        RECT 88.090 172.645 89.010 172.875 ;
        RECT 91.840 172.645 92.770 172.865 ;
        RECT 88.090 171.965 97.280 172.645 ;
        RECT 97.760 171.965 99.110 172.875 ;
        RECT 99.590 172.645 100.510 172.875 ;
        RECT 103.340 172.645 104.270 172.865 ;
        RECT 99.590 171.965 108.780 172.645 ;
        RECT 108.790 171.965 110.160 172.745 ;
        RECT 111.090 171.965 112.460 172.775 ;
        RECT 18.310 171.755 18.480 171.965 ;
        RECT 19.745 171.805 19.865 171.915 ;
        RECT 20.150 171.800 20.310 171.910 ;
        RECT 20.610 171.755 20.780 171.945 ;
        RECT 22.450 171.755 22.620 171.965 ;
        RECT 22.910 171.775 23.080 171.965 ;
        RECT 26.645 171.805 26.765 171.915 ;
        RECT 30.270 171.775 30.440 171.965 ;
        RECT 34.135 171.775 34.305 171.965 ;
        RECT 34.865 171.755 35.035 171.945 ;
        RECT 35.335 171.755 35.505 171.945 ;
        RECT 38.090 171.775 38.260 171.965 ;
        RECT 39.065 171.805 39.185 171.915 ;
        RECT 39.470 171.775 39.640 171.965 ;
        RECT 40.390 171.810 40.550 171.920 ;
        RECT 42.690 171.755 42.860 171.945 ;
        RECT 43.155 171.755 43.325 171.945 ;
        RECT 44.070 171.775 44.240 171.965 ;
        RECT 45.450 171.775 45.620 171.965 ;
        RECT 46.185 171.775 46.355 171.965 ;
        RECT 47.290 171.800 47.450 171.910 ;
        RECT 48.215 171.755 48.385 171.945 ;
        RECT 50.970 171.775 51.140 171.965 ;
        RECT 53.270 171.755 53.440 171.945 ;
        RECT 54.650 171.775 54.820 171.965 ;
        RECT 56.030 171.755 56.200 171.945 ;
        RECT 56.950 171.800 57.110 171.910 ;
        RECT 57.410 171.755 57.580 171.945 ;
        RECT 59.250 171.775 59.420 171.945 ;
        RECT 60.170 171.775 60.340 171.965 ;
        RECT 63.850 171.945 63.920 171.965 ;
        RECT 59.350 171.755 59.420 171.775 ;
        RECT 63.390 171.755 63.560 171.945 ;
        RECT 63.850 171.755 64.020 171.945 ;
        RECT 66.610 171.775 66.780 171.965 ;
        RECT 67.070 171.775 67.240 171.965 ;
        RECT 69.830 171.775 70.000 171.965 ;
        RECT 71.210 171.775 71.380 171.945 ;
        RECT 71.725 171.805 71.845 171.915 ;
        RECT 71.210 171.755 71.280 171.775 ;
        RECT 72.130 171.755 72.300 171.945 ;
        RECT 72.645 171.805 72.765 171.915 ;
        RECT 73.055 171.775 73.225 171.965 ;
        RECT 73.970 171.755 74.140 171.945 ;
        RECT 75.810 171.775 75.980 171.965 ;
        RECT 85.930 171.775 86.100 171.965 ;
        RECT 87.035 171.755 87.205 171.945 ;
        RECT 87.770 171.755 87.940 171.965 ;
        RECT 94.855 171.755 95.025 171.945 ;
        RECT 96.510 171.755 96.680 171.945 ;
        RECT 96.970 171.775 97.140 171.965 ;
        RECT 97.485 171.805 97.605 171.915 ;
        RECT 97.890 171.755 98.060 171.965 ;
        RECT 98.810 171.800 98.970 171.910 ;
        RECT 99.325 171.805 99.445 171.915 ;
        RECT 100.190 171.800 100.350 171.910 ;
        RECT 104.055 171.755 104.225 171.945 ;
        RECT 105.065 171.755 105.235 171.945 ;
        RECT 108.470 171.775 108.640 171.965 ;
        RECT 108.985 171.805 109.105 171.915 ;
        RECT 109.850 171.775 110.020 171.965 ;
        RECT 110.770 171.755 110.940 171.945 ;
        RECT 112.150 171.755 112.320 171.965 ;
        RECT 18.170 170.945 19.540 171.755 ;
        RECT 20.480 170.845 21.830 171.755 ;
        RECT 21.860 170.885 22.290 171.670 ;
        RECT 22.310 171.075 31.500 171.755 ;
        RECT 26.820 170.855 27.750 171.075 ;
        RECT 30.580 170.845 31.500 171.075 ;
        RECT 31.705 170.845 35.180 171.755 ;
        RECT 35.190 170.845 38.665 171.755 ;
        RECT 39.330 170.945 43.000 171.755 ;
        RECT 43.010 170.845 46.485 171.755 ;
        RECT 47.620 170.885 48.050 171.670 ;
        RECT 48.070 170.845 51.545 171.755 ;
        RECT 51.750 170.945 53.580 171.755 ;
        RECT 53.600 171.075 56.340 171.755 ;
        RECT 57.270 171.075 59.100 171.755 ;
        RECT 57.755 170.845 59.100 171.075 ;
        RECT 59.350 171.525 61.620 171.755 ;
        RECT 59.350 170.845 62.105 171.525 ;
        RECT 62.330 170.945 63.700 171.755 ;
        RECT 63.710 171.525 65.280 171.755 ;
        RECT 67.370 171.715 68.290 171.755 ;
        RECT 67.370 171.525 68.300 171.715 ;
        RECT 69.010 171.525 71.280 171.755 ;
        RECT 63.710 171.165 68.300 171.525 ;
        RECT 63.710 171.075 68.290 171.165 ;
        RECT 65.290 170.845 68.290 171.075 ;
        RECT 68.525 170.845 71.280 171.525 ;
        RECT 71.990 170.975 73.360 171.755 ;
        RECT 73.380 170.885 73.810 171.670 ;
        RECT 73.830 171.075 83.110 171.755 ;
        RECT 83.720 171.075 87.620 171.755 ;
        RECT 87.740 171.075 91.205 171.755 ;
        RECT 91.540 171.075 95.440 171.755 ;
        RECT 75.190 170.855 76.110 171.075 ;
        RECT 80.775 170.955 83.110 171.075 ;
        RECT 82.190 170.845 83.110 170.955 ;
        RECT 86.690 170.845 87.620 171.075 ;
        RECT 90.285 170.845 91.205 171.075 ;
        RECT 94.510 170.845 95.440 171.075 ;
        RECT 95.450 170.975 96.820 171.755 ;
        RECT 96.830 170.975 98.200 171.755 ;
        RECT 99.140 170.885 99.570 171.670 ;
        RECT 100.740 171.075 104.640 171.755 ;
        RECT 103.710 170.845 104.640 171.075 ;
        RECT 104.650 171.075 108.550 171.755 ;
        RECT 104.650 170.845 105.580 171.075 ;
        RECT 109.250 170.945 111.080 171.755 ;
        RECT 111.090 170.945 112.460 171.755 ;
      LAYER nwell ;
        RECT 17.975 167.725 112.655 170.555 ;
      LAYER pwell ;
        RECT 18.170 166.525 19.540 167.335 ;
        RECT 20.010 166.525 21.840 167.335 ;
        RECT 21.860 166.525 23.210 167.435 ;
        RECT 23.230 166.525 24.600 167.305 ;
        RECT 24.610 167.205 25.540 167.435 ;
        RECT 24.610 166.525 28.510 167.205 ;
        RECT 28.750 166.525 30.120 167.305 ;
        RECT 31.245 166.525 34.720 167.435 ;
        RECT 34.740 166.610 35.170 167.395 ;
        RECT 35.190 166.525 38.665 167.435 ;
        RECT 38.880 166.525 40.230 167.435 ;
        RECT 40.445 166.525 43.920 167.435 ;
        RECT 44.025 167.205 44.945 167.435 ;
        RECT 44.025 166.525 47.490 167.205 ;
        RECT 47.805 166.525 51.280 167.435 ;
        RECT 52.210 166.525 55.880 167.335 ;
        RECT 55.890 167.205 57.235 167.435 ;
        RECT 55.890 166.525 57.720 167.205 ;
        RECT 57.730 166.525 60.450 167.435 ;
        RECT 60.500 166.610 60.930 167.395 ;
        RECT 62.085 166.755 64.840 167.435 ;
        RECT 62.570 166.525 64.840 166.755 ;
        RECT 65.090 166.525 67.810 167.435 ;
        RECT 67.860 166.525 69.210 167.435 ;
        RECT 70.170 166.525 81.180 167.435 ;
        RECT 84.390 167.205 85.320 167.435 ;
        RECT 81.420 166.525 85.320 167.205 ;
        RECT 86.260 166.610 86.690 167.395 ;
        RECT 86.905 166.525 90.380 167.435 ;
        RECT 90.585 166.525 94.060 167.435 ;
        RECT 94.265 166.525 97.740 167.435 ;
        RECT 98.210 166.525 100.960 167.335 ;
        RECT 104.170 167.205 105.100 167.435 ;
        RECT 101.200 166.525 105.100 167.205 ;
        RECT 105.570 166.525 106.940 167.305 ;
        RECT 107.410 166.525 111.080 167.335 ;
        RECT 111.090 166.525 112.460 167.335 ;
        RECT 18.310 166.315 18.480 166.525 ;
        RECT 19.745 166.365 19.865 166.475 ;
        RECT 21.530 166.315 21.700 166.525 ;
        RECT 21.990 166.335 22.160 166.525 ;
        RECT 24.290 166.335 24.460 166.525 ;
        RECT 25.025 166.335 25.195 166.525 ;
        RECT 28.890 166.335 29.060 166.525 ;
        RECT 30.730 166.370 30.890 166.480 ;
        RECT 31.190 166.315 31.360 166.505 ;
        RECT 32.570 166.315 32.740 166.505 ;
        RECT 34.405 166.335 34.575 166.525 ;
        RECT 35.335 166.335 35.505 166.525 ;
        RECT 36.435 166.315 36.605 166.505 ;
        RECT 39.010 166.335 39.180 166.525 ;
        RECT 43.605 166.335 43.775 166.525 ;
        RECT 46.370 166.315 46.540 166.505 ;
        RECT 47.290 166.335 47.460 166.525 ;
        RECT 49.130 166.315 49.300 166.505 ;
        RECT 49.590 166.315 49.760 166.505 ;
        RECT 50.965 166.335 51.135 166.525 ;
        RECT 51.890 166.370 52.050 166.480 ;
        RECT 54.375 166.315 54.545 166.505 ;
        RECT 55.570 166.335 55.740 166.525 ;
        RECT 56.030 166.315 56.200 166.505 ;
        RECT 57.410 166.315 57.580 166.525 ;
        RECT 57.870 166.335 58.040 166.525 ;
        RECT 64.770 166.505 64.840 166.525 ;
        RECT 59.250 166.315 59.420 166.505 ;
        RECT 61.550 166.370 61.710 166.480 ;
        RECT 63.390 166.315 63.560 166.505 ;
        RECT 64.770 166.315 64.940 166.505 ;
        RECT 65.230 166.475 65.400 166.525 ;
        RECT 65.230 166.365 65.405 166.475 ;
        RECT 65.230 166.335 65.400 166.365 ;
        RECT 67.990 166.335 68.160 166.525 ;
        RECT 68.905 166.315 69.075 166.505 ;
        RECT 69.830 166.370 69.990 166.480 ;
        RECT 72.775 166.315 72.945 166.505 ;
        RECT 73.970 166.315 74.140 166.505 ;
        RECT 80.865 166.335 81.035 166.525 ;
        RECT 83.225 166.365 83.345 166.475 ;
        RECT 84.735 166.335 84.905 166.525 ;
        RECT 85.930 166.370 86.090 166.480 ;
        RECT 90.065 166.335 90.235 166.525 ;
        RECT 92.830 166.315 93.000 166.505 ;
        RECT 93.745 166.335 93.915 166.525 ;
        RECT 94.210 166.315 94.380 166.505 ;
        RECT 94.675 166.315 94.845 166.505 ;
        RECT 97.425 166.335 97.595 166.525 ;
        RECT 97.945 166.365 98.065 166.475 ;
        RECT 98.810 166.360 98.970 166.470 ;
        RECT 99.785 166.365 99.905 166.475 ;
        RECT 100.650 166.335 100.820 166.525 ;
        RECT 104.515 166.335 104.685 166.525 ;
        RECT 105.305 166.365 105.425 166.475 ;
        RECT 105.710 166.335 105.880 166.525 ;
        RECT 107.145 166.365 107.265 166.475 ;
        RECT 108.930 166.315 109.100 166.505 ;
        RECT 110.770 166.315 110.940 166.525 ;
        RECT 112.150 166.315 112.320 166.525 ;
        RECT 18.170 165.505 19.540 166.315 ;
        RECT 20.010 165.505 21.840 166.315 ;
        RECT 21.860 165.445 22.290 166.230 ;
        RECT 22.310 165.635 31.500 166.315 ;
        RECT 22.310 165.405 23.230 165.635 ;
        RECT 26.060 165.415 26.990 165.635 ;
        RECT 31.510 165.505 32.880 166.315 ;
        RECT 33.120 165.635 37.020 166.315 ;
        RECT 36.090 165.405 37.020 165.635 ;
        RECT 37.400 165.635 46.680 166.315 ;
        RECT 37.400 165.515 39.735 165.635 ;
        RECT 37.400 165.405 38.320 165.515 ;
        RECT 44.400 165.415 45.320 165.635 ;
        RECT 47.620 165.445 48.050 166.230 ;
        RECT 48.070 165.535 49.440 166.315 ;
        RECT 49.460 165.405 50.810 166.315 ;
        RECT 51.060 165.635 54.960 166.315 ;
        RECT 54.030 165.405 54.960 165.635 ;
        RECT 55.890 165.535 57.260 166.315 ;
        RECT 57.270 165.635 59.100 166.315 ;
        RECT 59.110 165.635 60.940 166.315 ;
        RECT 60.960 165.635 63.700 166.315 ;
        RECT 57.755 165.405 59.100 165.635 ;
        RECT 59.595 165.405 60.940 165.635 ;
        RECT 63.710 165.535 65.080 166.315 ;
        RECT 65.745 165.405 69.220 166.315 ;
        RECT 69.460 165.635 73.360 166.315 ;
        RECT 72.430 165.405 73.360 165.635 ;
        RECT 73.380 165.445 73.810 166.230 ;
        RECT 73.830 165.635 82.935 166.315 ;
        RECT 83.860 165.635 93.140 166.315 ;
        RECT 83.860 165.515 86.195 165.635 ;
        RECT 83.860 165.405 84.780 165.515 ;
        RECT 90.860 165.415 91.780 165.635 ;
        RECT 93.150 165.505 94.520 166.315 ;
        RECT 94.530 165.405 98.005 166.315 ;
        RECT 99.140 165.445 99.570 166.230 ;
        RECT 100.050 165.635 109.240 166.315 ;
        RECT 100.050 165.405 100.970 165.635 ;
        RECT 103.800 165.415 104.730 165.635 ;
        RECT 109.250 165.505 111.080 166.315 ;
        RECT 111.090 165.505 112.460 166.315 ;
      LAYER nwell ;
        RECT 17.975 162.285 112.655 165.115 ;
      LAYER pwell ;
        RECT 18.170 161.085 19.540 161.895 ;
        RECT 19.560 161.085 20.910 161.995 ;
        RECT 20.930 161.085 22.300 161.865 ;
        RECT 22.310 161.765 23.230 161.995 ;
        RECT 26.060 161.765 26.990 161.985 ;
        RECT 22.310 161.085 31.500 161.765 ;
        RECT 31.970 161.085 34.720 161.895 ;
        RECT 34.740 161.170 35.170 161.955 ;
        RECT 35.190 161.085 37.020 161.895 ;
        RECT 37.115 161.085 46.220 161.765 ;
        RECT 46.230 161.085 49.390 161.995 ;
        RECT 49.450 161.765 50.370 161.995 ;
        RECT 53.200 161.765 54.130 161.985 ;
        RECT 49.450 161.085 58.640 161.765 ;
        RECT 58.650 161.085 60.480 161.895 ;
        RECT 60.500 161.170 60.930 161.955 ;
        RECT 61.410 161.085 63.240 161.895 ;
        RECT 63.250 161.765 64.595 161.995 ;
        RECT 63.250 161.085 65.080 161.765 ;
        RECT 65.090 161.085 67.840 161.895 ;
        RECT 67.850 161.085 69.220 161.865 ;
        RECT 69.230 161.085 70.600 161.895 ;
        RECT 70.610 161.085 74.085 161.995 ;
        RECT 74.290 161.765 75.220 161.995 ;
        RECT 81.630 161.765 82.560 161.995 ;
        RECT 74.290 161.085 78.190 161.765 ;
        RECT 78.660 161.085 82.560 161.765 ;
        RECT 83.500 161.085 84.850 161.995 ;
        RECT 84.870 161.085 86.240 161.865 ;
        RECT 86.260 161.170 86.690 161.955 ;
        RECT 90.830 161.765 91.760 161.995 ;
        RECT 87.860 161.085 91.760 161.765 ;
        RECT 91.770 161.085 93.140 161.865 ;
        RECT 93.150 161.085 94.520 161.895 ;
        RECT 94.530 161.085 98.005 161.995 ;
        RECT 98.670 161.085 100.500 161.895 ;
        RECT 103.710 161.765 104.640 161.995 ;
        RECT 100.740 161.085 104.640 161.765 ;
        RECT 104.660 161.085 106.010 161.995 ;
        RECT 106.950 161.085 108.780 161.765 ;
        RECT 108.790 161.085 110.160 161.865 ;
        RECT 111.090 161.085 112.460 161.895 ;
        RECT 18.310 160.875 18.480 161.085 ;
        RECT 19.745 160.925 19.865 161.035 ;
        RECT 20.610 160.895 20.780 161.085 ;
        RECT 21.070 160.895 21.240 161.085 ;
        RECT 21.530 160.875 21.700 161.065 ;
        RECT 22.455 160.875 22.625 161.065 ;
        RECT 29.535 160.875 29.705 161.065 ;
        RECT 31.190 160.895 31.360 161.085 ;
        RECT 31.705 160.925 31.825 161.035 ;
        RECT 34.410 160.895 34.580 161.085 ;
        RECT 36.710 160.895 36.880 161.085 ;
        RECT 40.845 160.875 41.015 161.065 ;
        RECT 41.365 160.925 41.485 161.035 ;
        RECT 43.150 160.875 43.320 161.065 ;
        RECT 45.910 160.895 46.080 161.085 ;
        RECT 47.015 160.875 47.185 161.065 ;
        RECT 48.215 160.875 48.385 161.065 ;
        RECT 49.130 160.895 49.300 161.085 ;
        RECT 51.895 160.875 52.065 161.065 ;
        RECT 57.865 160.875 58.035 161.065 ;
        RECT 58.330 160.895 58.500 161.085 ;
        RECT 59.250 160.875 59.420 161.065 ;
        RECT 60.170 160.895 60.340 161.085 ;
        RECT 61.090 161.035 61.260 161.065 ;
        RECT 61.090 160.925 61.265 161.035 ;
        RECT 61.090 160.875 61.260 160.925 ;
        RECT 62.930 160.875 63.100 161.085 ;
        RECT 64.770 160.875 64.940 161.085 ;
        RECT 66.610 160.875 66.780 161.065 ;
        RECT 67.530 160.895 67.700 161.085 ;
        RECT 68.910 160.895 69.080 161.085 ;
        RECT 69.370 160.875 69.540 161.065 ;
        RECT 69.835 160.875 70.005 161.065 ;
        RECT 70.290 160.895 70.460 161.085 ;
        RECT 70.755 160.895 70.925 161.085 ;
        RECT 74.705 160.895 74.875 161.085 ;
        RECT 74.890 160.875 75.060 161.065 ;
        RECT 75.350 160.875 75.520 161.065 ;
        RECT 81.975 160.895 82.145 161.085 ;
        RECT 83.170 160.930 83.330 161.040 ;
        RECT 83.630 160.895 83.800 161.085 ;
        RECT 85.930 160.875 86.100 161.085 ;
        RECT 87.310 160.930 87.470 161.040 ;
        RECT 91.175 160.895 91.345 161.085 ;
        RECT 92.830 160.895 93.000 161.085 ;
        RECT 94.210 160.895 94.380 161.085 ;
        RECT 94.675 160.895 94.845 161.085 ;
        RECT 95.130 160.875 95.300 161.065 ;
        RECT 95.595 160.875 95.765 161.065 ;
        RECT 98.405 160.925 98.525 161.035 ;
        RECT 100.190 160.895 100.360 161.085 ;
        RECT 101.110 160.875 101.280 161.065 ;
        RECT 104.055 160.895 104.225 161.085 ;
        RECT 104.790 160.895 104.960 161.085 ;
        RECT 106.630 160.930 106.790 161.040 ;
        RECT 108.470 160.895 108.640 161.085 ;
        RECT 108.930 160.895 109.100 161.085 ;
        RECT 110.770 160.875 110.940 161.065 ;
        RECT 112.150 160.875 112.320 161.085 ;
        RECT 18.170 160.065 19.540 160.875 ;
        RECT 20.010 160.065 21.840 160.875 ;
        RECT 21.860 160.005 22.290 160.790 ;
        RECT 22.310 159.965 25.785 160.875 ;
        RECT 26.220 160.195 30.120 160.875 ;
        RECT 29.190 159.965 30.120 160.195 ;
        RECT 30.150 159.965 41.160 160.875 ;
        RECT 41.630 160.065 43.460 160.875 ;
        RECT 43.700 160.195 47.600 160.875 ;
        RECT 46.670 159.965 47.600 160.195 ;
        RECT 47.620 160.005 48.050 160.790 ;
        RECT 48.070 159.965 51.545 160.875 ;
        RECT 51.750 159.965 55.225 160.875 ;
        RECT 55.570 159.965 58.180 160.875 ;
        RECT 58.190 160.095 59.560 160.875 ;
        RECT 59.570 160.195 61.400 160.875 ;
        RECT 61.410 160.195 63.240 160.875 ;
        RECT 63.250 160.195 65.080 160.875 ;
        RECT 65.090 160.195 66.920 160.875 ;
        RECT 59.570 159.965 60.915 160.195 ;
        RECT 61.410 159.965 62.755 160.195 ;
        RECT 63.250 159.965 64.595 160.195 ;
        RECT 65.090 159.965 66.435 160.195 ;
        RECT 66.930 160.065 69.680 160.875 ;
        RECT 69.690 159.965 73.165 160.875 ;
        RECT 73.380 160.005 73.810 160.790 ;
        RECT 73.840 159.965 75.190 160.875 ;
        RECT 75.210 160.095 76.580 160.875 ;
        RECT 76.960 160.195 86.240 160.875 ;
        RECT 86.335 160.195 95.440 160.875 ;
        RECT 76.960 160.075 79.295 160.195 ;
        RECT 76.960 159.965 77.880 160.075 ;
        RECT 83.960 159.975 84.880 160.195 ;
        RECT 95.450 159.965 98.925 160.875 ;
        RECT 99.140 160.005 99.570 160.790 ;
        RECT 99.590 160.065 101.420 160.875 ;
        RECT 101.800 160.195 111.080 160.875 ;
        RECT 101.800 160.075 104.135 160.195 ;
        RECT 101.800 159.965 102.720 160.075 ;
        RECT 108.800 159.975 109.720 160.195 ;
        RECT 111.090 160.065 112.460 160.875 ;
      LAYER nwell ;
        RECT 17.975 156.845 112.655 159.675 ;
      LAYER pwell ;
        RECT 18.170 155.645 19.540 156.455 ;
        RECT 20.020 155.645 21.370 156.555 ;
        RECT 21.390 156.325 22.320 156.555 ;
        RECT 25.530 156.325 26.450 156.555 ;
        RECT 29.280 156.325 30.210 156.545 ;
        RECT 21.390 155.645 25.290 156.325 ;
        RECT 25.530 155.645 34.720 156.325 ;
        RECT 34.740 155.730 35.170 156.515 ;
        RECT 35.190 156.325 36.110 156.555 ;
        RECT 38.940 156.325 39.870 156.545 ;
        RECT 35.190 155.645 44.380 156.325 ;
        RECT 45.310 155.645 48.785 156.555 ;
        RECT 49.185 155.645 52.660 156.555 ;
        RECT 52.810 155.645 55.420 156.555 ;
        RECT 55.430 155.645 57.260 156.455 ;
        RECT 57.280 155.645 58.630 156.555 ;
        RECT 58.650 156.325 59.995 156.555 ;
        RECT 58.650 155.645 60.480 156.325 ;
        RECT 60.500 155.730 60.930 156.515 ;
        RECT 60.960 155.645 63.700 156.325 ;
        RECT 63.710 155.645 65.080 156.455 ;
        RECT 65.090 155.645 67.700 156.555 ;
        RECT 68.335 156.325 69.680 156.555 ;
        RECT 67.850 155.645 69.680 156.325 ;
        RECT 69.690 155.645 73.165 156.555 ;
        RECT 73.740 156.445 74.660 156.555 ;
        RECT 73.740 156.325 76.075 156.445 ;
        RECT 80.740 156.325 81.660 156.545 ;
        RECT 73.740 155.645 83.020 156.325 ;
        RECT 83.490 155.645 86.240 156.455 ;
        RECT 86.260 155.730 86.690 156.515 ;
        RECT 87.170 155.645 88.535 156.325 ;
        RECT 89.010 155.645 92.485 156.555 ;
        RECT 93.345 155.645 96.820 156.555 ;
        RECT 96.830 155.645 100.305 156.555 ;
        RECT 100.970 155.645 102.800 156.455 ;
        RECT 102.950 155.645 105.560 156.555 ;
        RECT 105.570 155.645 111.080 156.455 ;
        RECT 111.090 155.645 112.460 156.455 ;
        RECT 18.310 155.435 18.480 155.645 ;
        RECT 19.745 155.485 19.865 155.595 ;
        RECT 20.150 155.480 20.310 155.590 ;
        RECT 21.070 155.455 21.240 155.645 ;
        RECT 21.530 155.435 21.700 155.625 ;
        RECT 21.805 155.455 21.975 155.645 ;
        RECT 22.505 155.485 22.625 155.595 ;
        RECT 22.910 155.435 23.080 155.625 ;
        RECT 24.290 155.435 24.460 155.625 ;
        RECT 31.375 155.435 31.545 155.625 ;
        RECT 34.410 155.455 34.580 155.645 ;
        RECT 40.850 155.435 41.020 155.625 ;
        RECT 41.310 155.435 41.480 155.625 ;
        RECT 43.610 155.435 43.780 155.625 ;
        RECT 44.070 155.455 44.240 155.645 ;
        RECT 44.990 155.490 45.150 155.600 ;
        RECT 45.455 155.455 45.625 155.645 ;
        RECT 47.285 155.435 47.455 155.625 ;
        RECT 49.590 155.435 49.760 155.625 ;
        RECT 52.345 155.455 52.515 155.645 ;
        RECT 55.105 155.625 55.275 155.645 ;
        RECT 55.105 155.455 55.280 155.625 ;
        RECT 56.950 155.455 57.120 155.645 ;
        RECT 57.410 155.455 57.580 155.645 ;
        RECT 60.170 155.455 60.340 155.645 ;
        RECT 63.390 155.455 63.560 155.645 ;
        RECT 55.110 155.435 55.280 155.455 ;
        RECT 64.770 155.435 64.940 155.645 ;
        RECT 65.235 155.455 65.405 155.645 ;
        RECT 65.690 155.480 65.850 155.590 ;
        RECT 66.150 155.435 66.320 155.625 ;
        RECT 67.990 155.455 68.160 155.645 ;
        RECT 68.910 155.435 69.080 155.625 ;
        RECT 69.835 155.455 70.005 155.645 ;
        RECT 73.050 155.435 73.220 155.625 ;
        RECT 74.025 155.485 74.145 155.595 ;
        RECT 74.430 155.435 74.600 155.625 ;
        RECT 77.650 155.480 77.810 155.590 ;
        RECT 79.030 155.435 79.200 155.625 ;
        RECT 79.545 155.485 79.665 155.595 ;
        RECT 82.250 155.435 82.420 155.625 ;
        RECT 82.710 155.455 82.880 155.645 ;
        RECT 83.225 155.485 83.345 155.595 ;
        RECT 85.930 155.455 86.100 155.645 ;
        RECT 86.905 155.485 87.025 155.595 ;
        RECT 87.770 155.435 87.940 155.625 ;
        RECT 88.235 155.435 88.405 155.625 ;
        RECT 88.690 155.455 88.860 155.625 ;
        RECT 89.155 155.455 89.325 155.645 ;
        RECT 91.965 155.485 92.085 155.595 ;
        RECT 92.375 155.435 92.545 155.625 ;
        RECT 92.885 155.485 93.005 155.595 ;
        RECT 96.105 155.485 96.225 155.595 ;
        RECT 96.505 155.455 96.675 155.645 ;
        RECT 96.975 155.455 97.145 155.645 ;
        RECT 102.490 155.625 102.660 155.645 ;
        RECT 98.810 155.435 98.980 155.625 ;
        RECT 100.705 155.485 100.825 155.595 ;
        RECT 102.030 155.435 102.200 155.625 ;
        RECT 102.490 155.455 102.665 155.625 ;
        RECT 105.245 155.595 105.415 155.645 ;
        RECT 105.245 155.485 105.425 155.595 ;
        RECT 105.245 155.455 105.415 155.485 ;
        RECT 102.495 155.435 102.665 155.455 ;
        RECT 105.710 155.435 105.880 155.625 ;
        RECT 107.145 155.485 107.265 155.595 ;
        RECT 110.770 155.435 110.940 155.645 ;
        RECT 112.150 155.435 112.320 155.645 ;
        RECT 18.170 154.625 19.540 155.435 ;
        RECT 20.480 154.525 21.830 155.435 ;
        RECT 21.860 154.565 22.290 155.350 ;
        RECT 22.780 154.525 24.130 155.435 ;
        RECT 24.260 154.755 27.725 155.435 ;
        RECT 28.060 154.755 31.960 155.435 ;
        RECT 32.055 154.755 41.160 155.435 ;
        RECT 26.805 154.525 27.725 154.755 ;
        RECT 31.030 154.525 31.960 154.755 ;
        RECT 41.170 154.655 42.540 155.435 ;
        RECT 42.550 154.625 43.920 155.435 ;
        RECT 44.125 154.525 47.600 155.435 ;
        RECT 47.620 154.565 48.050 155.350 ;
        RECT 48.070 154.625 49.900 155.435 ;
        RECT 49.910 154.625 55.420 155.435 ;
        RECT 55.800 154.755 65.080 155.435 ;
        RECT 55.800 154.635 58.135 154.755 ;
        RECT 55.800 154.525 56.720 154.635 ;
        RECT 62.800 154.535 63.720 154.755 ;
        RECT 66.010 154.525 68.730 155.435 ;
        RECT 68.770 154.755 70.600 155.435 ;
        RECT 69.255 154.525 70.600 154.755 ;
        RECT 70.610 154.625 73.360 155.435 ;
        RECT 73.380 154.565 73.810 155.350 ;
        RECT 74.290 154.755 77.030 155.435 ;
        RECT 77.980 154.525 79.330 155.435 ;
        RECT 79.810 154.625 82.560 155.435 ;
        RECT 82.570 154.625 88.080 155.435 ;
        RECT 88.090 154.525 91.565 155.435 ;
        RECT 92.230 154.525 95.705 155.435 ;
        RECT 96.370 154.625 99.120 155.435 ;
        RECT 99.140 154.565 99.570 155.350 ;
        RECT 99.590 154.625 102.340 155.435 ;
        RECT 102.350 154.525 104.960 155.435 ;
        RECT 105.570 154.655 106.940 155.435 ;
        RECT 107.410 154.625 111.080 155.435 ;
        RECT 111.090 154.625 112.460 155.435 ;
      LAYER nwell ;
        RECT 17.975 151.405 112.655 154.235 ;
      LAYER pwell ;
        RECT 18.170 150.205 19.540 151.015 ;
        RECT 20.010 150.885 20.930 151.115 ;
        RECT 23.760 150.885 24.690 151.105 ;
        RECT 20.010 150.205 29.200 150.885 ;
        RECT 29.210 150.205 30.580 150.985 ;
        RECT 30.590 150.205 31.960 150.985 ;
        RECT 31.970 150.915 32.915 151.115 ;
        RECT 31.970 150.235 34.720 150.915 ;
        RECT 34.740 150.290 35.170 151.075 ;
        RECT 31.970 150.205 32.915 150.235 ;
        RECT 18.310 149.995 18.480 150.205 ;
        RECT 19.745 150.045 19.865 150.155 ;
        RECT 21.530 149.995 21.700 150.185 ;
        RECT 23.370 149.995 23.540 150.185 ;
        RECT 27.235 149.995 27.405 150.185 ;
        RECT 28.025 150.045 28.145 150.155 ;
        RECT 28.890 150.015 29.060 150.205 ;
        RECT 29.810 149.995 29.980 150.185 ;
        RECT 30.270 150.015 30.440 150.205 ;
        RECT 30.730 150.015 30.900 150.205 ;
        RECT 31.190 149.995 31.360 150.185 ;
        RECT 31.655 149.995 31.825 150.185 ;
        RECT 34.405 150.015 34.575 150.235 ;
        RECT 35.190 150.205 38.665 151.115 ;
        RECT 39.330 150.205 43.000 151.015 ;
        RECT 43.010 150.915 43.955 151.115 ;
        RECT 45.770 150.915 46.715 151.115 ;
        RECT 43.010 150.235 45.760 150.915 ;
        RECT 45.770 150.235 48.520 150.915 ;
        RECT 43.010 150.205 43.955 150.235 ;
        RECT 35.335 150.015 35.505 150.205 ;
        RECT 35.790 150.040 35.950 150.150 ;
        RECT 36.255 149.995 36.425 150.185 ;
        RECT 39.065 150.045 39.185 150.155 ;
        RECT 39.930 149.995 40.100 150.185 ;
        RECT 42.690 150.015 42.860 150.205 ;
        RECT 45.445 150.015 45.615 150.235 ;
        RECT 45.770 150.205 46.715 150.235 ;
        RECT 47.015 149.995 47.185 150.185 ;
        RECT 48.205 150.155 48.375 150.235 ;
        RECT 48.530 150.205 52.005 151.115 ;
        RECT 55.410 150.885 56.340 151.115 ;
        RECT 59.465 150.885 60.385 151.115 ;
        RECT 52.440 150.205 56.340 150.885 ;
        RECT 56.920 150.205 60.385 150.885 ;
        RECT 60.500 150.290 60.930 151.075 ;
        RECT 62.355 150.885 63.700 151.115 ;
        RECT 66.955 150.885 68.300 151.115 ;
        RECT 68.795 150.885 70.140 151.115 ;
        RECT 61.870 150.205 63.700 150.885 ;
        RECT 63.720 150.205 66.460 150.885 ;
        RECT 66.470 150.205 68.300 150.885 ;
        RECT 68.310 150.205 70.140 150.885 ;
        RECT 70.610 150.205 72.440 151.015 ;
        RECT 72.450 150.205 75.925 151.115 ;
        RECT 76.130 150.205 79.605 151.115 ;
        RECT 80.740 150.205 82.090 151.115 ;
        RECT 85.310 150.885 86.240 151.115 ;
        RECT 82.340 150.205 86.240 150.885 ;
        RECT 86.260 150.290 86.690 151.075 ;
        RECT 87.630 150.205 89.000 150.985 ;
        RECT 89.010 150.205 91.760 151.015 ;
        RECT 91.965 150.205 95.440 151.115 ;
        RECT 95.450 150.205 98.925 151.115 ;
        RECT 99.600 150.205 100.950 151.115 ;
        RECT 100.970 150.885 101.890 151.115 ;
        RECT 104.720 150.885 105.650 151.105 ;
        RECT 100.970 150.205 110.160 150.885 ;
        RECT 111.090 150.205 112.460 151.015 ;
        RECT 48.205 150.045 48.385 150.155 ;
        RECT 48.205 150.015 48.375 150.045 ;
        RECT 48.675 150.015 48.845 150.205 ;
        RECT 55.755 150.015 55.925 150.205 ;
        RECT 56.545 150.045 56.665 150.155 ;
        RECT 56.950 150.015 57.120 150.205 ;
        RECT 57.410 149.995 57.580 150.185 ;
        RECT 58.790 149.995 58.960 150.185 ;
        RECT 59.255 149.995 59.425 150.185 ;
        RECT 61.550 150.050 61.710 150.160 ;
        RECT 62.010 150.015 62.180 150.205 ;
        RECT 65.690 149.995 65.860 150.185 ;
        RECT 66.150 149.995 66.320 150.205 ;
        RECT 66.610 150.015 66.780 150.205 ;
        RECT 67.990 149.995 68.160 150.185 ;
        RECT 68.450 150.015 68.620 150.205 ;
        RECT 70.345 150.045 70.465 150.155 ;
        RECT 72.130 150.015 72.300 150.205 ;
        RECT 72.595 150.015 72.765 150.205 ;
        RECT 73.045 149.995 73.215 150.185 ;
        RECT 73.975 149.995 74.145 150.185 ;
        RECT 76.275 150.015 76.445 150.205 ;
        RECT 78.110 150.040 78.270 150.150 ;
        RECT 80.410 150.050 80.570 150.160 ;
        RECT 80.870 150.015 81.040 150.205 ;
        RECT 81.790 149.995 81.960 150.185 ;
        RECT 85.655 150.015 85.825 150.205 ;
        RECT 87.310 150.050 87.470 150.160 ;
        RECT 87.770 150.015 87.940 150.205 ;
        RECT 90.990 149.995 91.160 150.185 ;
        RECT 91.450 150.015 91.620 150.205 ;
        RECT 94.665 149.995 94.835 150.185 ;
        RECT 95.125 150.015 95.295 150.205 ;
        RECT 95.595 150.015 95.765 150.205 ;
        RECT 98.535 149.995 98.705 150.185 ;
        RECT 99.325 150.045 99.445 150.155 ;
        RECT 99.730 150.015 99.900 150.205 ;
        RECT 101.110 149.995 101.280 150.185 ;
        RECT 109.850 150.015 110.020 150.205 ;
        RECT 110.770 149.995 110.940 150.185 ;
        RECT 112.150 149.995 112.320 150.205 ;
        RECT 18.170 149.185 19.540 149.995 ;
        RECT 20.010 149.185 21.840 149.995 ;
        RECT 21.860 149.125 22.290 149.910 ;
        RECT 22.310 149.185 23.680 149.995 ;
        RECT 23.920 149.315 27.820 149.995 ;
        RECT 26.890 149.085 27.820 149.315 ;
        RECT 28.290 149.185 30.120 149.995 ;
        RECT 30.140 149.085 31.490 149.995 ;
        RECT 31.510 149.085 34.985 149.995 ;
        RECT 36.110 149.085 39.585 149.995 ;
        RECT 39.900 149.315 43.365 149.995 ;
        RECT 43.700 149.315 47.600 149.995 ;
        RECT 42.445 149.085 43.365 149.315 ;
        RECT 46.670 149.085 47.600 149.315 ;
        RECT 47.620 149.125 48.050 149.910 ;
        RECT 48.530 149.315 57.720 149.995 ;
        RECT 48.530 149.085 49.450 149.315 ;
        RECT 52.280 149.095 53.210 149.315 ;
        RECT 57.730 149.215 59.100 149.995 ;
        RECT 59.110 149.085 62.585 149.995 ;
        RECT 62.790 149.085 66.000 149.995 ;
        RECT 66.010 149.315 67.840 149.995 ;
        RECT 67.850 149.315 69.680 149.995 ;
        RECT 66.495 149.085 67.840 149.315 ;
        RECT 68.335 149.085 69.680 149.315 ;
        RECT 69.885 149.085 73.360 149.995 ;
        RECT 73.380 149.125 73.810 149.910 ;
        RECT 73.830 149.085 77.305 149.995 ;
        RECT 78.430 149.185 82.100 149.995 ;
        RECT 82.110 149.315 91.300 149.995 ;
        RECT 82.110 149.085 83.030 149.315 ;
        RECT 85.860 149.095 86.790 149.315 ;
        RECT 91.505 149.085 94.980 149.995 ;
        RECT 95.220 149.315 99.120 149.995 ;
        RECT 98.190 149.085 99.120 149.315 ;
        RECT 99.140 149.125 99.570 149.910 ;
        RECT 99.590 149.185 101.420 149.995 ;
        RECT 101.800 149.315 111.080 149.995 ;
        RECT 101.800 149.195 104.135 149.315 ;
        RECT 101.800 149.085 102.720 149.195 ;
        RECT 108.800 149.095 109.720 149.315 ;
        RECT 111.090 149.185 112.460 149.995 ;
      LAYER nwell ;
        RECT 17.975 145.965 112.655 148.795 ;
      LAYER pwell ;
        RECT 18.170 144.765 19.540 145.575 ;
        RECT 19.550 145.445 20.470 145.675 ;
        RECT 23.300 145.445 24.230 145.665 ;
        RECT 19.550 144.765 28.740 145.445 ;
        RECT 28.750 144.765 30.120 145.545 ;
        RECT 31.245 144.765 34.720 145.675 ;
        RECT 34.740 144.850 35.170 145.635 ;
        RECT 35.190 144.765 38.665 145.675 ;
        RECT 39.700 145.565 40.620 145.675 ;
        RECT 39.700 145.445 42.035 145.565 ;
        RECT 46.700 145.445 47.620 145.665 ;
        RECT 39.700 144.765 48.980 145.445 ;
        RECT 48.990 144.765 50.360 145.545 ;
        RECT 50.840 144.765 52.190 145.675 ;
        RECT 52.670 144.765 56.145 145.675 ;
        RECT 59.550 145.445 60.480 145.675 ;
        RECT 56.580 144.765 60.480 145.445 ;
        RECT 60.500 144.850 60.930 145.635 ;
        RECT 61.410 144.765 63.240 145.575 ;
        RECT 63.735 145.445 65.080 145.675 ;
        RECT 63.250 144.765 65.080 145.445 ;
        RECT 65.100 144.765 66.450 145.675 ;
        RECT 66.470 144.765 67.840 145.545 ;
        RECT 68.310 144.765 70.140 145.575 ;
        RECT 70.150 145.475 71.095 145.675 ;
        RECT 70.150 144.795 72.900 145.475 ;
        RECT 70.150 144.765 71.095 144.795 ;
        RECT 18.310 144.555 18.480 144.765 ;
        RECT 20.150 144.600 20.310 144.710 ;
        RECT 20.610 144.555 20.780 144.745 ;
        RECT 28.430 144.575 28.600 144.765 ;
        RECT 28.890 144.575 29.060 144.765 ;
        RECT 30.730 144.610 30.890 144.720 ;
        RECT 31.190 144.555 31.360 144.745 ;
        RECT 32.110 144.600 32.270 144.710 ;
        RECT 34.405 144.575 34.575 144.765 ;
        RECT 35.335 144.575 35.505 144.765 ;
        RECT 35.785 144.555 35.955 144.745 ;
        RECT 37.170 144.555 37.340 144.745 ;
        RECT 37.635 144.555 37.805 144.745 ;
        RECT 39.065 144.605 39.185 144.715 ;
        RECT 41.365 144.605 41.485 144.715 ;
        RECT 43.150 144.555 43.320 144.745 ;
        RECT 43.885 144.555 44.055 144.745 ;
        RECT 48.265 144.605 48.385 144.715 ;
        RECT 48.670 144.575 48.840 144.765 ;
        RECT 50.050 144.575 50.220 144.765 ;
        RECT 50.565 144.605 50.685 144.715 ;
        RECT 50.970 144.575 51.140 144.765 ;
        RECT 51.890 144.555 52.060 144.745 ;
        RECT 52.405 144.605 52.525 144.715 ;
        RECT 52.815 144.575 52.985 144.765 ;
        RECT 59.895 144.575 60.065 144.765 ;
        RECT 61.090 144.715 61.260 144.745 ;
        RECT 61.090 144.605 61.265 144.715 ;
        RECT 61.090 144.555 61.260 144.605 ;
        RECT 62.930 144.575 63.100 144.765 ;
        RECT 63.390 144.575 63.560 144.765 ;
        RECT 66.150 144.575 66.320 144.765 ;
        RECT 66.610 144.575 66.780 144.765 ;
        RECT 68.045 144.605 68.165 144.715 ;
        RECT 69.830 144.575 70.000 144.765 ;
        RECT 70.750 144.555 70.920 144.745 ;
        RECT 71.265 144.605 71.385 144.715 ;
        RECT 72.585 144.575 72.755 144.795 ;
        RECT 72.910 144.765 76.385 145.675 ;
        RECT 76.960 145.565 77.880 145.675 ;
        RECT 76.960 145.445 79.295 145.565 ;
        RECT 83.960 145.445 84.880 145.665 ;
        RECT 76.960 144.765 86.240 145.445 ;
        RECT 86.260 144.850 86.690 145.635 ;
        RECT 86.720 144.765 88.070 145.675 ;
        RECT 88.090 144.765 91.760 145.575 ;
        RECT 91.770 145.475 92.715 145.675 ;
        RECT 96.335 145.475 97.280 145.675 ;
        RECT 91.770 144.795 94.520 145.475 ;
        RECT 94.530 144.795 97.280 145.475 ;
        RECT 91.770 144.765 92.715 144.795 ;
        RECT 73.055 144.745 73.225 144.765 ;
        RECT 73.050 144.575 73.225 144.745 ;
        RECT 73.050 144.555 73.220 144.575 ;
        RECT 79.030 144.555 79.200 144.745 ;
        RECT 82.895 144.555 83.065 144.745 ;
        RECT 84.090 144.600 84.250 144.710 ;
        RECT 85.470 144.555 85.640 144.745 ;
        RECT 85.930 144.575 86.100 144.765 ;
        RECT 86.850 144.555 87.020 144.745 ;
        RECT 87.770 144.575 87.940 144.765 ;
        RECT 91.450 144.575 91.620 144.765 ;
        RECT 92.370 144.555 92.540 144.745 ;
        RECT 94.205 144.575 94.375 144.795 ;
        RECT 94.675 144.575 94.845 144.795 ;
        RECT 96.335 144.765 97.280 144.795 ;
        RECT 97.750 144.765 100.500 145.575 ;
        RECT 103.710 145.445 104.640 145.675 ;
        RECT 100.740 144.765 104.640 145.445 ;
        RECT 104.660 144.765 106.010 145.675 ;
        RECT 106.490 144.765 107.860 145.545 ;
        RECT 108.330 144.765 111.080 145.575 ;
        RECT 111.090 144.765 112.460 145.575 ;
        RECT 18.170 143.745 19.540 144.555 ;
        RECT 20.470 143.775 21.840 144.555 ;
        RECT 21.860 143.685 22.290 144.470 ;
        RECT 22.310 143.875 31.500 144.555 ;
        RECT 22.310 143.645 23.230 143.875 ;
        RECT 26.060 143.655 26.990 143.875 ;
        RECT 32.625 143.645 36.100 144.555 ;
        RECT 36.110 143.745 37.480 144.555 ;
        RECT 37.490 143.645 40.965 144.555 ;
        RECT 41.630 143.745 43.460 144.555 ;
        RECT 43.470 143.875 47.370 144.555 ;
        RECT 43.470 143.645 44.400 143.875 ;
        RECT 47.620 143.685 48.050 144.470 ;
        RECT 48.530 143.745 52.200 144.555 ;
        RECT 52.295 143.875 61.400 144.555 ;
        RECT 61.780 143.875 71.060 144.555 ;
        RECT 61.780 143.755 64.115 143.875 ;
        RECT 61.780 143.645 62.700 143.755 ;
        RECT 68.780 143.655 69.700 143.875 ;
        RECT 71.530 143.745 73.360 144.555 ;
        RECT 73.380 143.685 73.810 144.470 ;
        RECT 73.830 143.745 79.340 144.555 ;
        RECT 79.580 143.875 83.480 144.555 ;
        RECT 82.550 143.645 83.480 143.875 ;
        RECT 84.410 143.775 85.780 144.555 ;
        RECT 85.790 143.745 87.160 144.555 ;
        RECT 87.170 143.745 92.680 144.555 ;
        RECT 92.690 144.525 93.635 144.555 ;
        RECT 95.125 144.525 95.295 144.745 ;
        RECT 95.595 144.555 95.765 144.745 ;
        RECT 97.485 144.605 97.605 144.715 ;
        RECT 100.190 144.575 100.360 144.765 ;
        RECT 104.055 144.575 104.225 144.765 ;
        RECT 104.790 144.555 104.960 144.765 ;
        RECT 105.250 144.555 105.420 144.745 ;
        RECT 106.225 144.605 106.345 144.715 ;
        RECT 106.630 144.555 106.800 144.765 ;
        RECT 108.065 144.605 108.185 144.715 ;
        RECT 110.770 144.555 110.940 144.765 ;
        RECT 112.150 144.555 112.320 144.765 ;
        RECT 92.690 143.845 95.440 144.525 ;
        RECT 92.690 143.645 93.635 143.845 ;
        RECT 95.450 143.645 98.925 144.555 ;
        RECT 99.140 143.685 99.570 144.470 ;
        RECT 99.590 143.745 105.100 144.555 ;
        RECT 105.120 143.645 106.470 144.555 ;
        RECT 106.490 143.775 107.860 144.555 ;
        RECT 108.330 143.745 111.080 144.555 ;
        RECT 111.090 143.745 112.460 144.555 ;
      LAYER nwell ;
        RECT 17.975 140.525 112.655 143.355 ;
      LAYER pwell ;
        RECT 18.170 139.325 19.540 140.135 ;
        RECT 20.020 139.325 21.370 140.235 ;
        RECT 21.400 139.325 22.750 140.235 ;
        RECT 22.770 140.005 23.700 140.235 ;
        RECT 30.110 140.005 31.040 140.235 ;
        RECT 22.770 139.325 26.670 140.005 ;
        RECT 27.140 139.325 31.040 140.005 ;
        RECT 31.970 140.035 32.915 140.235 ;
        RECT 31.970 139.355 34.720 140.035 ;
        RECT 34.740 139.410 35.170 140.195 ;
        RECT 31.970 139.325 32.915 139.355 ;
        RECT 18.310 139.115 18.480 139.325 ;
        RECT 19.745 139.165 19.865 139.275 ;
        RECT 21.070 139.135 21.240 139.325 ;
        RECT 21.530 139.115 21.700 139.325 ;
        RECT 22.910 139.160 23.070 139.270 ;
        RECT 23.185 139.135 23.355 139.325 ;
        RECT 26.590 139.115 26.760 139.305 ;
        RECT 30.455 139.135 30.625 139.325 ;
        RECT 31.650 139.170 31.810 139.280 ;
        RECT 32.110 139.115 32.280 139.305 ;
        RECT 18.170 138.305 19.540 139.115 ;
        RECT 20.010 138.305 21.840 139.115 ;
        RECT 21.860 138.245 22.290 139.030 ;
        RECT 23.230 138.305 26.900 139.115 ;
        RECT 26.910 138.305 32.420 139.115 ;
        RECT 32.575 139.085 32.745 139.305 ;
        RECT 34.405 139.135 34.575 139.355 ;
        RECT 36.110 139.325 39.780 140.135 ;
        RECT 39.800 139.325 41.150 140.235 ;
        RECT 41.540 140.125 42.460 140.235 ;
        RECT 41.540 140.005 43.875 140.125 ;
        RECT 48.540 140.005 49.460 140.225 ;
        RECT 50.830 140.035 51.775 140.235 ;
        RECT 41.540 139.325 50.820 140.005 ;
        RECT 50.830 139.355 53.580 140.035 ;
        RECT 50.830 139.325 51.775 139.355 ;
        RECT 35.790 139.170 35.950 139.280 ;
        RECT 37.630 139.115 37.800 139.305 ;
        RECT 38.095 139.115 38.265 139.305 ;
        RECT 39.470 139.135 39.640 139.325 ;
        RECT 39.930 139.135 40.100 139.325 ;
        RECT 43.150 139.115 43.320 139.305 ;
        RECT 43.610 139.115 43.780 139.305 ;
        RECT 34.235 139.085 35.180 139.115 ;
        RECT 32.430 138.405 35.180 139.085 ;
        RECT 34.235 138.205 35.180 138.405 ;
        RECT 35.190 138.305 37.940 139.115 ;
        RECT 37.950 138.205 41.425 139.115 ;
        RECT 41.630 138.305 43.460 139.115 ;
        RECT 43.470 138.335 44.840 139.115 ;
        RECT 44.850 139.085 45.795 139.115 ;
        RECT 47.285 139.085 47.455 139.305 ;
        RECT 50.510 139.115 50.680 139.325 ;
        RECT 53.265 139.135 53.435 139.355 ;
        RECT 53.590 139.325 56.340 140.135 ;
        RECT 56.350 139.325 59.825 140.235 ;
        RECT 60.500 139.410 60.930 140.195 ;
        RECT 61.320 140.125 62.240 140.235 ;
        RECT 61.320 140.005 63.655 140.125 ;
        RECT 68.320 140.005 69.240 140.225 ;
        RECT 61.320 139.325 70.600 140.005 ;
        RECT 71.070 139.325 72.900 140.135 ;
        RECT 72.910 139.325 76.385 140.235 ;
        RECT 76.960 140.125 77.880 140.235 ;
        RECT 76.960 140.005 79.295 140.125 ;
        RECT 83.960 140.005 84.880 140.225 ;
        RECT 76.960 139.325 86.240 140.005 ;
        RECT 86.260 139.410 86.690 140.195 ;
        RECT 86.720 139.325 88.070 140.235 ;
        RECT 88.090 139.325 90.840 140.135 ;
        RECT 90.850 140.035 91.795 140.235 ;
        RECT 90.850 139.355 93.600 140.035 ;
        RECT 90.850 139.325 91.795 139.355 ;
        RECT 56.030 139.115 56.200 139.325 ;
        RECT 56.495 139.115 56.665 139.325 ;
        RECT 60.225 139.165 60.345 139.275 ;
        RECT 60.630 139.160 60.790 139.270 ;
        RECT 64.495 139.115 64.665 139.305 ;
        RECT 66.140 139.115 66.310 139.305 ;
        RECT 67.530 139.115 67.700 139.305 ;
        RECT 67.990 139.115 68.160 139.305 ;
        RECT 70.290 139.115 70.460 139.325 ;
        RECT 70.805 139.165 70.925 139.275 ;
        RECT 72.590 139.135 72.760 139.325 ;
        RECT 73.055 139.305 73.225 139.325 ;
        RECT 73.045 139.135 73.225 139.305 ;
        RECT 74.430 139.160 74.590 139.270 ;
        RECT 44.850 138.405 47.600 139.085 ;
        RECT 44.850 138.205 45.795 138.405 ;
        RECT 47.620 138.245 48.050 139.030 ;
        RECT 48.070 138.305 50.820 139.115 ;
        RECT 50.830 138.305 56.340 139.115 ;
        RECT 56.350 138.205 59.825 139.115 ;
        RECT 61.180 138.435 65.080 139.115 ;
        RECT 64.150 138.205 65.080 138.435 ;
        RECT 65.090 138.335 66.460 139.115 ;
        RECT 66.480 138.205 67.830 139.115 ;
        RECT 67.850 138.335 69.220 139.115 ;
        RECT 69.230 138.305 70.600 139.115 ;
        RECT 70.610 139.085 71.555 139.115 ;
        RECT 73.045 139.085 73.215 139.135 ;
        RECT 78.110 139.115 78.280 139.305 ;
        RECT 81.975 139.115 82.145 139.305 ;
        RECT 82.710 139.115 82.880 139.305 ;
        RECT 85.930 139.135 86.100 139.325 ;
        RECT 70.610 138.405 73.360 139.085 ;
        RECT 70.610 138.205 71.555 138.405 ;
        RECT 73.380 138.245 73.810 139.030 ;
        RECT 74.750 138.305 78.420 139.115 ;
        RECT 78.660 138.435 82.560 139.115 ;
        RECT 81.630 138.205 82.560 138.435 ;
        RECT 82.570 138.335 83.940 139.115 ;
        RECT 83.950 139.085 84.895 139.115 ;
        RECT 86.385 139.085 86.555 139.305 ;
        RECT 87.770 139.135 87.940 139.325 ;
        RECT 90.530 139.305 90.700 139.325 ;
        RECT 90.065 139.115 90.235 139.305 ;
        RECT 90.530 139.135 90.705 139.305 ;
        RECT 93.285 139.135 93.455 139.355 ;
        RECT 93.610 139.325 97.085 140.235 ;
        RECT 100.490 140.005 101.420 140.235 ;
        RECT 97.520 139.325 101.420 140.005 ;
        RECT 101.800 140.125 102.720 140.235 ;
        RECT 101.800 140.005 104.135 140.125 ;
        RECT 108.800 140.005 109.720 140.225 ;
        RECT 101.800 139.325 111.080 140.005 ;
        RECT 111.090 139.325 112.460 140.135 ;
        RECT 93.755 139.135 93.925 139.325 ;
        RECT 94.670 139.160 94.830 139.270 ;
        RECT 90.535 139.115 90.705 139.135 ;
        RECT 98.535 139.115 98.705 139.305 ;
        RECT 99.785 139.165 99.905 139.275 ;
        RECT 100.190 139.115 100.360 139.305 ;
        RECT 100.835 139.135 101.005 139.325 ;
        RECT 110.770 139.115 110.940 139.325 ;
        RECT 112.150 139.115 112.320 139.325 ;
        RECT 83.950 138.405 86.700 139.085 ;
        RECT 83.950 138.205 84.895 138.405 ;
        RECT 86.905 138.205 90.380 139.115 ;
        RECT 90.390 138.205 93.865 139.115 ;
        RECT 95.220 138.435 99.120 139.115 ;
        RECT 98.190 138.205 99.120 138.435 ;
        RECT 99.140 138.245 99.570 139.030 ;
        RECT 100.060 138.205 101.410 139.115 ;
        RECT 101.800 138.435 111.080 139.115 ;
        RECT 101.800 138.315 104.135 138.435 ;
        RECT 101.800 138.205 102.720 138.315 ;
        RECT 108.800 138.215 109.720 138.435 ;
        RECT 111.090 138.305 112.460 139.115 ;
      LAYER nwell ;
        RECT 17.975 135.085 112.655 137.915 ;
      LAYER pwell ;
        RECT 18.170 133.885 19.540 134.695 ;
        RECT 19.550 133.885 20.920 134.695 ;
        RECT 20.930 133.885 26.440 134.695 ;
        RECT 26.450 133.885 31.960 134.695 ;
        RECT 33.775 134.595 34.720 134.795 ;
        RECT 31.970 133.915 34.720 134.595 ;
        RECT 34.740 133.970 35.170 134.755 ;
        RECT 18.310 133.675 18.480 133.885 ;
        RECT 19.745 133.725 19.865 133.835 ;
        RECT 20.610 133.695 20.780 133.885 ;
        RECT 21.530 133.675 21.700 133.865 ;
        RECT 22.505 133.725 22.625 133.835 ;
        RECT 22.910 133.675 23.080 133.865 ;
        RECT 24.750 133.720 24.910 133.830 ;
        RECT 25.485 133.675 25.655 133.865 ;
        RECT 26.130 133.695 26.300 133.885 ;
        RECT 30.270 133.675 30.440 133.865 ;
        RECT 31.650 133.695 31.820 133.885 ;
        RECT 32.115 133.695 32.285 133.915 ;
        RECT 33.775 133.885 34.720 133.915 ;
        RECT 35.650 133.885 37.480 134.695 ;
        RECT 37.500 133.885 38.850 134.795 ;
        RECT 38.870 133.885 42.345 134.795 ;
        RECT 43.010 133.885 45.760 134.695 ;
        RECT 46.140 134.685 47.060 134.795 ;
        RECT 46.140 134.565 48.475 134.685 ;
        RECT 53.140 134.565 54.060 134.785 ;
        RECT 59.550 134.565 60.480 134.795 ;
        RECT 46.140 133.885 55.420 134.565 ;
        RECT 56.580 133.885 60.480 134.565 ;
        RECT 60.500 133.970 60.930 134.755 ;
        RECT 61.320 134.685 62.240 134.795 ;
        RECT 61.320 134.565 63.655 134.685 ;
        RECT 68.320 134.565 69.240 134.785 ;
        RECT 61.320 133.885 70.600 134.565 ;
        RECT 71.070 133.885 73.820 134.695 ;
        RECT 73.830 133.885 77.305 134.795 ;
        RECT 77.510 133.885 79.340 134.695 ;
        RECT 82.550 134.565 83.480 134.795 ;
        RECT 79.580 133.885 83.480 134.565 ;
        RECT 83.490 133.885 84.860 134.665 ;
        RECT 84.870 133.885 86.240 134.695 ;
        RECT 86.260 133.970 86.690 134.755 ;
        RECT 87.170 133.885 89.920 134.695 ;
        RECT 93.130 134.565 94.060 134.795 ;
        RECT 90.160 133.885 94.060 134.565 ;
        RECT 94.070 134.595 95.015 134.795 ;
        RECT 97.200 134.685 98.120 134.795 ;
        RECT 94.070 133.915 96.820 134.595 ;
        RECT 97.200 134.565 99.535 134.685 ;
        RECT 104.200 134.565 105.120 134.785 ;
        RECT 94.070 133.885 95.015 133.915 ;
        RECT 18.170 132.865 19.540 133.675 ;
        RECT 20.010 132.865 21.840 133.675 ;
        RECT 21.860 132.805 22.290 133.590 ;
        RECT 22.780 132.765 24.130 133.675 ;
        RECT 25.070 132.995 28.970 133.675 ;
        RECT 25.070 132.765 26.000 132.995 ;
        RECT 29.210 132.865 30.580 133.675 ;
        RECT 30.590 133.645 31.535 133.675 ;
        RECT 33.025 133.645 33.195 133.865 ;
        RECT 35.330 133.835 35.500 133.865 ;
        RECT 35.330 133.725 35.505 133.835 ;
        RECT 35.330 133.695 35.500 133.725 ;
        RECT 35.330 133.675 35.480 133.695 ;
        RECT 35.795 133.675 35.965 133.865 ;
        RECT 37.170 133.695 37.340 133.885 ;
        RECT 37.630 133.695 37.800 133.885 ;
        RECT 39.015 133.695 39.185 133.885 ;
        RECT 42.745 133.725 42.865 133.835 ;
        RECT 42.875 133.675 43.045 133.865 ;
        RECT 45.450 133.695 45.620 133.885 ;
        RECT 47.015 133.675 47.185 133.865 ;
        RECT 48.670 133.720 48.830 133.830 ;
        RECT 49.130 133.675 49.300 133.865 ;
        RECT 50.510 133.675 50.680 133.865 ;
        RECT 51.895 133.675 52.065 133.865 ;
        RECT 55.110 133.695 55.280 133.885 ;
        RECT 56.030 133.730 56.190 133.840 ;
        RECT 59.895 133.695 60.065 133.885 ;
        RECT 64.770 133.675 64.940 133.865 ;
        RECT 66.150 133.675 66.320 133.865 ;
        RECT 66.610 133.675 66.780 133.865 ;
        RECT 70.290 133.675 70.460 133.885 ;
        RECT 70.805 133.725 70.925 133.835 ;
        RECT 30.590 132.965 33.340 133.645 ;
        RECT 30.590 132.765 31.535 132.965 ;
        RECT 33.550 132.855 35.480 133.675 ;
        RECT 33.550 132.765 34.500 132.855 ;
        RECT 35.650 132.765 39.125 133.675 ;
        RECT 39.560 132.995 43.460 133.675 ;
        RECT 43.700 132.995 47.600 133.675 ;
        RECT 42.530 132.765 43.460 132.995 ;
        RECT 46.670 132.765 47.600 132.995 ;
        RECT 47.620 132.805 48.050 133.590 ;
        RECT 49.000 132.765 50.350 133.675 ;
        RECT 50.370 132.895 51.740 133.675 ;
        RECT 51.750 132.765 55.225 133.675 ;
        RECT 55.800 132.995 65.080 133.675 ;
        RECT 55.800 132.875 58.135 132.995 ;
        RECT 55.800 132.765 56.720 132.875 ;
        RECT 62.800 132.775 63.720 132.995 ;
        RECT 65.100 132.765 66.450 133.675 ;
        RECT 66.470 132.895 67.840 133.675 ;
        RECT 67.850 132.865 70.600 133.675 ;
        RECT 70.610 133.645 71.555 133.675 ;
        RECT 73.045 133.645 73.215 133.865 ;
        RECT 73.510 133.695 73.680 133.885 ;
        RECT 73.975 133.675 74.145 133.885 ;
        RECT 79.030 133.695 79.200 133.885 ;
        RECT 82.895 133.695 83.065 133.885 ;
        RECT 83.630 133.695 83.800 133.885 ;
        RECT 85.930 133.695 86.100 133.885 ;
        RECT 86.850 133.835 87.020 133.865 ;
        RECT 86.850 133.725 87.025 133.835 ;
        RECT 86.850 133.675 87.020 133.725 ;
        RECT 89.610 133.695 89.780 133.885 ;
        RECT 93.475 133.695 93.645 133.885 ;
        RECT 96.505 133.865 96.675 133.915 ;
        RECT 97.200 133.885 106.480 134.565 ;
        RECT 106.490 133.885 107.860 134.665 ;
        RECT 108.330 133.885 111.080 134.695 ;
        RECT 111.090 133.885 112.460 134.695 ;
        RECT 96.505 133.695 96.680 133.865 ;
        RECT 97.430 133.720 97.590 133.830 ;
        RECT 96.510 133.675 96.680 133.695 ;
        RECT 97.890 133.675 98.060 133.865 ;
        RECT 103.135 133.675 103.305 133.865 ;
        RECT 103.870 133.675 104.040 133.865 ;
        RECT 105.305 133.725 105.425 133.835 ;
        RECT 106.170 133.695 106.340 133.885 ;
        RECT 106.630 133.695 106.800 133.885 ;
        RECT 108.065 133.725 108.185 133.835 ;
        RECT 110.770 133.675 110.940 133.885 ;
        RECT 112.150 133.675 112.320 133.885 ;
        RECT 70.610 132.965 73.360 133.645 ;
        RECT 70.610 132.765 71.555 132.965 ;
        RECT 73.380 132.805 73.810 133.590 ;
        RECT 73.830 132.765 77.305 133.675 ;
        RECT 77.880 132.995 87.160 133.675 ;
        RECT 87.540 132.995 96.820 133.675 ;
        RECT 77.880 132.875 80.215 132.995 ;
        RECT 77.880 132.765 78.800 132.875 ;
        RECT 84.880 132.775 85.800 132.995 ;
        RECT 87.540 132.875 89.875 132.995 ;
        RECT 87.540 132.765 88.460 132.875 ;
        RECT 94.540 132.775 95.460 132.995 ;
        RECT 97.760 132.765 99.110 133.675 ;
        RECT 99.140 132.805 99.570 133.590 ;
        RECT 99.820 132.995 103.720 133.675 ;
        RECT 102.790 132.765 103.720 132.995 ;
        RECT 103.730 132.895 105.100 133.675 ;
        RECT 105.570 132.865 111.080 133.675 ;
        RECT 111.090 132.865 112.460 133.675 ;
      LAYER nwell ;
        RECT 17.975 129.645 112.655 132.475 ;
      LAYER pwell ;
        RECT 18.170 128.445 19.540 129.255 ;
        RECT 19.920 129.245 20.840 129.355 ;
        RECT 19.920 129.125 22.255 129.245 ;
        RECT 26.920 129.125 27.840 129.345 ;
        RECT 19.920 128.445 29.200 129.125 ;
        RECT 29.680 128.445 31.030 129.355 ;
        RECT 32.190 129.265 33.140 129.355 ;
        RECT 31.210 128.445 33.140 129.265 ;
        RECT 33.350 128.445 34.720 129.255 ;
        RECT 34.740 128.530 35.170 129.315 ;
        RECT 35.850 129.265 36.800 129.355 ;
        RECT 35.850 128.445 37.780 129.265 ;
        RECT 38.320 129.245 39.240 129.355 ;
        RECT 38.320 129.125 40.655 129.245 ;
        RECT 45.320 129.125 46.240 129.345 ;
        RECT 47.610 129.155 48.555 129.355 ;
        RECT 38.320 128.445 47.600 129.125 ;
        RECT 47.610 128.475 50.360 129.155 ;
        RECT 47.610 128.445 48.555 128.475 ;
        RECT 18.310 128.235 18.480 128.445 ;
        RECT 20.150 128.280 20.310 128.390 ;
        RECT 20.610 128.235 20.780 128.425 ;
        RECT 22.725 128.235 22.895 128.425 ;
        RECT 26.590 128.235 26.760 128.425 ;
        RECT 28.890 128.255 29.060 128.445 ;
        RECT 29.405 128.285 29.525 128.395 ;
        RECT 29.810 128.255 29.980 128.445 ;
        RECT 31.210 128.425 31.360 128.445 ;
        RECT 31.190 128.255 31.360 128.425 ;
        RECT 34.410 128.255 34.580 128.445 ;
        RECT 37.630 128.425 37.780 128.445 ;
        RECT 35.385 128.285 35.505 128.395 ;
        RECT 37.170 128.235 37.340 128.425 ;
        RECT 37.630 128.255 37.800 128.425 ;
        RECT 37.905 128.235 38.075 128.425 ;
        RECT 41.770 128.235 41.940 128.425 ;
        RECT 43.150 128.255 43.320 128.425 ;
        RECT 45.450 128.255 45.620 128.425 ;
        RECT 47.290 128.255 47.460 128.445 ;
        RECT 48.265 128.285 48.385 128.395 ;
        RECT 50.045 128.255 50.215 128.475 ;
        RECT 50.370 128.445 55.880 129.255 ;
        RECT 59.090 129.125 60.020 129.355 ;
        RECT 56.120 128.445 60.020 129.125 ;
        RECT 60.500 128.530 60.930 129.315 ;
        RECT 60.950 128.445 62.320 129.225 ;
        RECT 62.340 128.445 63.690 129.355 ;
        RECT 69.450 129.265 70.400 129.355 ;
        RECT 64.630 128.445 68.300 129.255 ;
        RECT 68.470 128.445 70.400 129.265 ;
        RECT 70.695 128.445 79.800 129.125 ;
        RECT 80.270 128.445 82.100 129.255 ;
        RECT 82.120 128.445 83.470 129.355 ;
        RECT 83.490 128.445 84.860 129.255 ;
        RECT 84.880 128.445 86.230 129.355 ;
        RECT 86.260 128.530 86.690 129.315 ;
        RECT 86.710 128.445 95.815 129.125 ;
        RECT 95.910 128.445 97.280 129.225 ;
        RECT 97.290 128.445 100.040 129.255 ;
        RECT 100.050 128.445 105.560 129.255 ;
        RECT 105.570 128.445 111.080 129.255 ;
        RECT 111.090 128.445 112.460 129.255 ;
        RECT 50.510 128.255 50.680 128.425 ;
        RECT 43.170 128.235 43.320 128.255 ;
        RECT 45.470 128.235 45.620 128.255 ;
        RECT 50.510 128.235 50.660 128.255 ;
        RECT 51.890 128.235 52.060 128.425 ;
        RECT 55.110 128.255 55.280 128.425 ;
        RECT 55.570 128.255 55.740 128.445 ;
        RECT 56.950 128.235 57.120 128.425 ;
        RECT 57.410 128.235 57.580 128.425 ;
        RECT 58.790 128.235 58.960 128.425 ;
        RECT 59.435 128.255 59.605 128.445 ;
        RECT 60.225 128.285 60.345 128.395 ;
        RECT 61.090 128.255 61.260 128.445 ;
        RECT 62.010 128.235 62.180 128.425 ;
        RECT 63.390 128.255 63.560 128.445 ;
        RECT 64.310 128.255 64.480 128.425 ;
        RECT 64.310 128.235 64.460 128.255 ;
        RECT 67.990 128.235 68.160 128.445 ;
        RECT 68.470 128.425 68.620 128.445 ;
        RECT 68.450 128.255 68.620 128.425 ;
        RECT 68.470 128.235 68.620 128.255 ;
        RECT 18.170 127.425 19.540 128.235 ;
        RECT 20.470 127.455 21.840 128.235 ;
        RECT 21.860 127.365 22.290 128.150 ;
        RECT 22.310 127.555 26.210 128.235 ;
        RECT 22.310 127.325 23.240 127.555 ;
        RECT 26.450 127.455 27.820 128.235 ;
        RECT 28.200 127.555 37.480 128.235 ;
        RECT 37.490 127.555 41.390 128.235 ;
        RECT 28.200 127.435 30.535 127.555 ;
        RECT 28.200 127.325 29.120 127.435 ;
        RECT 35.200 127.335 36.120 127.555 ;
        RECT 37.490 127.325 38.420 127.555 ;
        RECT 41.630 127.455 43.000 128.235 ;
        RECT 43.170 127.415 45.100 128.235 ;
        RECT 45.470 127.415 47.400 128.235 ;
        RECT 44.150 127.325 45.100 127.415 ;
        RECT 46.450 127.325 47.400 127.415 ;
        RECT 47.620 127.365 48.050 128.150 ;
        RECT 48.730 127.415 50.660 128.235 ;
        RECT 50.830 127.425 52.200 128.235 ;
        RECT 52.590 127.555 55.015 128.235 ;
        RECT 55.430 127.425 57.260 128.235 ;
        RECT 57.270 127.455 58.640 128.235 ;
        RECT 58.650 127.555 60.480 128.235 ;
        RECT 60.490 127.555 62.320 128.235 ;
        RECT 62.530 127.415 64.460 128.235 ;
        RECT 64.630 127.425 68.300 128.235 ;
        RECT 68.470 127.415 70.400 128.235 ;
        RECT 48.730 127.325 49.680 127.415 ;
        RECT 62.530 127.325 63.480 127.415 ;
        RECT 69.450 127.325 70.400 127.415 ;
        RECT 70.610 128.205 71.555 128.235 ;
        RECT 73.045 128.205 73.215 128.425 ;
        RECT 74.025 128.285 74.145 128.395 ;
        RECT 77.835 128.235 78.005 128.425 ;
        RECT 79.490 128.255 79.660 128.445 ;
        RECT 80.005 128.285 80.125 128.395 ;
        RECT 80.870 128.235 81.040 128.425 ;
        RECT 81.790 128.255 81.960 128.445 ;
        RECT 82.250 128.235 82.420 128.425 ;
        RECT 82.765 128.285 82.885 128.395 ;
        RECT 83.170 128.235 83.340 128.445 ;
        RECT 84.550 128.255 84.720 128.445 ;
        RECT 85.010 128.255 85.180 128.445 ;
        RECT 86.850 128.255 87.020 128.445 ;
        RECT 93.290 128.280 93.450 128.390 ;
        RECT 95.590 128.255 95.760 128.425 ;
        RECT 96.510 128.280 96.670 128.390 ;
        RECT 96.970 128.255 97.140 128.445 ;
        RECT 98.810 128.255 98.980 128.425 ;
        RECT 99.730 128.395 99.900 128.445 ;
        RECT 99.730 128.285 99.905 128.395 ;
        RECT 99.730 128.255 99.900 128.285 ;
        RECT 95.590 128.235 95.740 128.255 ;
        RECT 98.810 128.235 98.960 128.255 ;
        RECT 100.190 128.235 100.360 128.425 ;
        RECT 105.250 128.255 105.420 128.445 ;
        RECT 110.770 128.235 110.940 128.445 ;
        RECT 112.150 128.235 112.320 128.445 ;
        RECT 70.610 127.525 73.360 128.205 ;
        RECT 70.610 127.325 71.555 127.525 ;
        RECT 73.380 127.365 73.810 128.150 ;
        RECT 74.520 127.555 78.420 128.235 ;
        RECT 77.490 127.325 78.420 127.555 ;
        RECT 79.090 127.425 81.180 128.235 ;
        RECT 81.200 127.325 82.550 128.235 ;
        RECT 83.030 127.555 92.310 128.235 ;
        RECT 84.390 127.335 85.310 127.555 ;
        RECT 89.975 127.435 92.310 127.555 ;
        RECT 91.390 127.325 92.310 127.435 ;
        RECT 93.810 127.415 95.740 128.235 ;
        RECT 97.030 127.415 98.960 128.235 ;
        RECT 93.810 127.325 94.760 127.415 ;
        RECT 97.030 127.325 97.980 127.415 ;
        RECT 99.140 127.365 99.570 128.150 ;
        RECT 100.060 127.325 101.410 128.235 ;
        RECT 101.800 127.555 111.080 128.235 ;
        RECT 101.800 127.435 104.135 127.555 ;
        RECT 101.800 127.325 102.720 127.435 ;
        RECT 108.800 127.335 109.720 127.555 ;
        RECT 111.090 127.425 112.460 128.235 ;
      LAYER nwell ;
        RECT 17.975 124.205 112.655 127.035 ;
      LAYER pwell ;
        RECT 18.170 123.005 19.540 123.815 ;
        RECT 19.920 123.805 20.840 123.915 ;
        RECT 19.920 123.685 22.255 123.805 ;
        RECT 26.920 123.685 27.840 123.905 ;
        RECT 30.810 123.825 31.760 123.915 ;
        RECT 19.920 123.005 29.200 123.685 ;
        RECT 29.830 123.005 31.760 123.825 ;
        RECT 32.170 123.825 33.120 123.915 ;
        RECT 32.170 123.005 34.100 123.825 ;
        RECT 34.740 123.090 35.170 123.875 ;
        RECT 35.275 123.005 44.380 123.685 ;
        RECT 44.850 123.005 46.220 123.785 ;
        RECT 46.230 123.005 55.335 123.685 ;
        RECT 55.430 123.005 56.800 123.815 ;
        RECT 56.820 123.005 59.560 123.685 ;
        RECT 60.500 123.090 60.930 123.875 ;
        RECT 60.950 123.005 62.780 123.815 ;
        RECT 62.790 123.005 65.530 123.685 ;
        RECT 65.550 123.005 67.380 123.815 ;
        RECT 67.400 123.005 68.750 123.915 ;
        RECT 69.910 123.825 70.860 123.915 ;
        RECT 72.210 123.825 73.160 123.915 ;
        RECT 68.930 123.005 70.860 123.825 ;
        RECT 71.230 123.005 73.160 123.825 ;
        RECT 74.200 123.805 75.120 123.915 ;
        RECT 74.200 123.685 76.535 123.805 ;
        RECT 81.200 123.685 82.120 123.905 ;
        RECT 74.200 123.005 83.480 123.685 ;
        RECT 83.490 123.005 84.860 123.815 ;
        RECT 84.880 123.005 86.230 123.915 ;
        RECT 86.260 123.090 86.690 123.875 ;
        RECT 88.290 123.825 89.240 123.915 ;
        RECT 94.730 123.825 95.680 123.915 ;
        RECT 97.030 123.825 97.980 123.915 ;
        RECT 86.710 123.005 88.080 123.785 ;
        RECT 88.290 123.005 90.220 123.825 ;
        RECT 90.850 123.005 94.520 123.815 ;
        RECT 94.730 123.005 96.660 123.825 ;
        RECT 97.030 123.005 98.960 123.825 ;
        RECT 102.330 123.685 103.260 123.915 ;
        RECT 99.360 123.005 103.260 123.685 ;
        RECT 104.190 123.005 105.560 123.785 ;
        RECT 106.030 123.005 107.400 123.785 ;
        RECT 107.410 123.005 111.080 123.815 ;
        RECT 111.090 123.005 112.460 123.815 ;
        RECT 18.310 122.795 18.480 123.005 ;
        RECT 20.150 122.840 20.310 122.950 ;
        RECT 21.530 122.795 21.700 122.985 ;
        RECT 28.890 122.815 29.060 123.005 ;
        RECT 29.830 122.985 29.980 123.005 ;
        RECT 33.950 122.985 34.100 123.005 ;
        RECT 29.405 122.845 29.525 122.955 ;
        RECT 29.810 122.815 29.980 122.985 ;
        RECT 31.650 122.795 31.820 122.985 ;
        RECT 32.385 122.795 32.555 122.985 ;
        RECT 33.950 122.815 34.120 122.985 ;
        RECT 34.465 122.845 34.585 122.955 ;
        RECT 37.170 122.795 37.340 122.985 ;
        RECT 38.090 122.840 38.250 122.950 ;
        RECT 38.550 122.795 38.720 122.985 ;
        RECT 40.850 122.815 41.020 122.985 ;
        RECT 41.310 122.815 41.480 122.985 ;
        RECT 41.330 122.795 41.480 122.815 ;
        RECT 43.885 122.795 44.055 122.985 ;
        RECT 44.070 122.815 44.240 123.005 ;
        RECT 44.585 122.845 44.705 122.955 ;
        RECT 44.990 122.815 45.160 123.005 ;
        RECT 46.370 122.815 46.540 123.005 ;
        RECT 48.670 122.840 48.830 122.950 ;
        RECT 49.130 122.795 49.300 122.985 ;
        RECT 50.510 122.815 50.680 122.985 ;
        RECT 50.530 122.795 50.680 122.815 ;
        RECT 56.215 122.795 56.385 122.985 ;
        RECT 56.490 122.815 56.660 123.005 ;
        RECT 59.250 122.985 59.420 123.005 ;
        RECT 59.245 122.815 59.420 122.985 ;
        RECT 59.765 122.845 59.885 122.955 ;
        RECT 60.170 122.850 60.330 122.960 ;
        RECT 62.470 122.815 62.640 123.005 ;
        RECT 62.930 122.815 63.100 123.005 ;
        RECT 59.245 122.795 59.415 122.815 ;
        RECT 63.390 122.795 63.560 122.985 ;
        RECT 63.850 122.795 64.020 122.985 ;
        RECT 67.070 122.815 67.240 123.005 ;
        RECT 67.530 122.815 67.700 123.005 ;
        RECT 68.930 122.985 69.080 123.005 ;
        RECT 71.230 122.985 71.380 123.005 ;
        RECT 68.910 122.815 69.080 122.985 ;
        RECT 71.210 122.815 71.380 122.985 ;
        RECT 73.565 122.845 73.685 122.955 ;
        RECT 74.025 122.845 74.145 122.955 ;
        RECT 75.350 122.795 75.520 122.985 ;
        RECT 75.865 122.845 75.985 122.955 ;
        RECT 78.570 122.795 78.740 122.985 ;
        RECT 79.030 122.795 79.200 122.985 ;
        RECT 80.465 122.845 80.585 122.955 ;
        RECT 83.170 122.795 83.340 123.005 ;
        RECT 84.550 122.815 84.720 123.005 ;
        RECT 85.010 122.815 85.180 123.005 ;
        RECT 87.035 122.795 87.205 122.985 ;
        RECT 87.770 122.815 87.940 123.005 ;
        RECT 90.070 122.985 90.220 123.005 ;
        RECT 88.045 122.795 88.215 122.985 ;
        RECT 90.070 122.815 90.240 122.985 ;
        RECT 90.585 122.845 90.705 122.955 ;
        RECT 91.910 122.815 92.080 122.985 ;
        RECT 94.210 122.815 94.380 123.005 ;
        RECT 96.510 122.985 96.660 123.005 ;
        RECT 98.810 122.985 98.960 123.005 ;
        RECT 96.510 122.815 96.680 122.985 ;
        RECT 91.930 122.795 92.080 122.815 ;
        RECT 97.615 122.795 97.785 122.985 ;
        RECT 98.810 122.815 98.980 122.985 ;
        RECT 100.190 122.840 100.350 122.950 ;
        RECT 102.675 122.815 102.845 123.005 ;
        RECT 103.870 122.850 104.030 122.960 ;
        RECT 104.055 122.795 104.225 122.985 ;
        RECT 104.330 122.815 104.500 123.005 ;
        RECT 104.790 122.795 104.960 122.985 ;
        RECT 106.170 122.955 106.340 123.005 ;
        RECT 105.765 122.845 105.885 122.955 ;
        RECT 106.170 122.845 106.345 122.955 ;
        RECT 106.170 122.815 106.340 122.845 ;
        RECT 106.630 122.795 106.800 122.985 ;
        RECT 108.065 122.845 108.185 122.955 ;
        RECT 110.770 122.795 110.940 123.005 ;
        RECT 112.150 122.795 112.320 123.005 ;
        RECT 18.170 121.985 19.540 122.795 ;
        RECT 20.480 121.885 21.830 122.795 ;
        RECT 21.860 121.925 22.290 122.710 ;
        RECT 22.680 122.115 31.960 122.795 ;
        RECT 31.970 122.115 35.870 122.795 ;
        RECT 22.680 121.995 25.015 122.115 ;
        RECT 22.680 121.885 23.600 121.995 ;
        RECT 29.680 121.895 30.600 122.115 ;
        RECT 31.970 121.885 32.900 122.115 ;
        RECT 36.110 122.015 37.480 122.795 ;
        RECT 38.420 121.885 39.770 122.795 ;
        RECT 39.790 122.115 40.745 122.795 ;
        RECT 41.330 121.975 43.260 122.795 ;
        RECT 42.310 121.885 43.260 121.975 ;
        RECT 43.470 122.115 47.370 122.795 ;
        RECT 43.470 121.885 44.400 122.115 ;
        RECT 47.620 121.925 48.050 122.710 ;
        RECT 49.000 121.885 50.350 122.795 ;
        RECT 50.530 121.975 52.460 122.795 ;
        RECT 52.900 122.115 56.800 122.795 ;
        RECT 51.510 121.885 52.460 121.975 ;
        RECT 55.870 121.885 56.800 122.115 ;
        RECT 56.950 121.885 59.560 122.795 ;
        RECT 60.030 121.985 63.700 122.795 ;
        RECT 63.710 122.115 72.990 122.795 ;
        RECT 65.070 121.895 65.990 122.115 ;
        RECT 70.655 121.995 72.990 122.115 ;
        RECT 72.070 121.885 72.990 121.995 ;
        RECT 73.380 121.925 73.810 122.710 ;
        RECT 74.290 122.015 75.660 122.795 ;
        RECT 76.130 121.985 78.880 122.795 ;
        RECT 78.890 122.015 80.260 122.795 ;
        RECT 80.730 121.985 83.480 122.795 ;
        RECT 83.720 122.115 87.620 122.795 ;
        RECT 86.690 121.885 87.620 122.115 ;
        RECT 87.630 122.115 91.530 122.795 ;
        RECT 87.630 121.885 88.560 122.115 ;
        RECT 91.930 121.975 93.860 122.795 ;
        RECT 94.300 122.115 98.200 122.795 ;
        RECT 92.910 121.885 93.860 121.975 ;
        RECT 97.270 121.885 98.200 122.115 ;
        RECT 99.140 121.925 99.570 122.710 ;
        RECT 100.740 122.115 104.640 122.795 ;
        RECT 103.710 121.885 104.640 122.115 ;
        RECT 104.660 121.885 106.010 122.795 ;
        RECT 106.490 122.015 107.860 122.795 ;
        RECT 108.330 121.985 111.080 122.795 ;
        RECT 111.090 121.985 112.460 122.795 ;
      LAYER nwell ;
        RECT 17.975 118.765 112.655 121.595 ;
      LAYER pwell ;
        RECT 18.170 117.565 19.540 118.375 ;
        RECT 19.550 117.565 20.920 118.375 ;
        RECT 24.130 118.245 25.060 118.475 ;
        RECT 21.160 117.565 25.060 118.245 ;
        RECT 25.440 118.365 26.360 118.475 ;
        RECT 25.440 118.245 27.775 118.365 ;
        RECT 32.440 118.245 33.360 118.465 ;
        RECT 25.440 117.565 34.720 118.245 ;
        RECT 34.740 117.650 35.170 118.435 ;
        RECT 35.660 117.565 37.010 118.475 ;
        RECT 37.030 118.245 37.960 118.475 ;
        RECT 41.540 118.365 42.460 118.475 ;
        RECT 41.540 118.245 43.875 118.365 ;
        RECT 48.540 118.245 49.460 118.465 ;
        RECT 51.200 118.365 52.120 118.475 ;
        RECT 51.200 118.245 53.535 118.365 ;
        RECT 58.200 118.245 59.120 118.465 ;
        RECT 37.030 117.565 40.930 118.245 ;
        RECT 41.540 117.565 50.820 118.245 ;
        RECT 51.200 117.565 60.480 118.245 ;
        RECT 60.500 117.650 60.930 118.435 ;
        RECT 63.620 118.365 64.540 118.475 ;
        RECT 60.950 117.565 62.320 118.345 ;
        RECT 63.620 118.245 65.955 118.365 ;
        RECT 70.620 118.245 71.540 118.465 ;
        RECT 72.910 118.245 73.840 118.475 ;
        RECT 63.620 117.565 72.900 118.245 ;
        RECT 72.910 117.565 76.810 118.245 ;
        RECT 77.050 117.565 78.420 118.375 ;
        RECT 78.430 118.245 79.360 118.475 ;
        RECT 78.430 117.565 82.330 118.245 ;
        RECT 82.570 117.565 86.240 118.375 ;
        RECT 86.260 117.650 86.690 118.435 ;
        RECT 86.710 117.565 88.080 118.375 ;
        RECT 88.100 117.565 89.450 118.475 ;
        RECT 89.840 118.365 90.760 118.475 ;
        RECT 89.840 118.245 92.175 118.365 ;
        RECT 96.840 118.245 97.760 118.465 ;
        RECT 89.840 117.565 99.120 118.245 ;
        RECT 100.060 117.565 101.410 118.475 ;
        RECT 101.800 118.365 102.720 118.475 ;
        RECT 101.800 118.245 104.135 118.365 ;
        RECT 108.800 118.245 109.720 118.465 ;
        RECT 101.800 117.565 111.080 118.245 ;
        RECT 111.090 117.565 112.460 118.375 ;
        RECT 18.310 117.355 18.480 117.565 ;
        RECT 19.745 117.405 19.865 117.515 ;
        RECT 20.610 117.375 20.780 117.565 ;
        RECT 21.530 117.355 21.700 117.545 ;
        RECT 22.910 117.400 23.070 117.510 ;
        RECT 23.370 117.355 23.540 117.545 ;
        RECT 24.475 117.375 24.645 117.565 ;
        RECT 25.210 117.400 25.370 117.510 ;
        RECT 25.670 117.355 25.840 117.545 ;
        RECT 27.050 117.355 27.220 117.545 ;
        RECT 28.430 117.355 28.600 117.545 ;
        RECT 34.410 117.375 34.580 117.565 ;
        RECT 35.385 117.405 35.505 117.515 ;
        RECT 36.710 117.375 36.880 117.565 ;
        RECT 37.445 117.375 37.615 117.565 ;
        RECT 47.290 117.355 47.460 117.545 ;
        RECT 48.670 117.400 48.830 117.510 ;
        RECT 50.510 117.375 50.680 117.565 ;
        RECT 52.535 117.355 52.705 117.545 ;
        RECT 60.170 117.375 60.340 117.565 ;
        RECT 62.010 117.375 62.180 117.565 ;
        RECT 62.470 117.355 62.640 117.545 ;
        RECT 62.930 117.515 63.090 117.520 ;
        RECT 62.930 117.410 63.105 117.515 ;
        RECT 62.985 117.405 63.105 117.410 ;
        RECT 65.690 117.355 65.860 117.545 ;
        RECT 66.150 117.355 66.320 117.545 ;
        RECT 70.935 117.355 71.105 117.545 ;
        RECT 72.590 117.355 72.760 117.565 ;
        RECT 73.105 117.405 73.225 117.515 ;
        RECT 73.325 117.375 73.495 117.565 ;
        RECT 74.430 117.400 74.590 117.510 ;
        RECT 78.110 117.375 78.280 117.565 ;
        RECT 78.845 117.375 79.015 117.565 ;
        RECT 84.090 117.355 84.260 117.545 ;
        RECT 85.930 117.375 86.100 117.565 ;
        RECT 87.770 117.375 87.940 117.565 ;
        RECT 88.230 117.375 88.400 117.565 ;
        RECT 93.750 117.355 93.920 117.545 ;
        RECT 94.670 117.400 94.830 117.510 ;
        RECT 98.535 117.355 98.705 117.545 ;
        RECT 98.810 117.375 98.980 117.565 ;
        RECT 99.730 117.410 99.890 117.520 ;
        RECT 100.190 117.375 100.360 117.565 ;
        RECT 108.930 117.355 109.100 117.545 ;
        RECT 110.770 117.355 110.940 117.565 ;
        RECT 112.150 117.355 112.320 117.565 ;
        RECT 18.170 116.545 19.540 117.355 ;
        RECT 20.010 116.545 21.840 117.355 ;
        RECT 21.860 116.485 22.290 117.270 ;
        RECT 23.240 116.445 24.590 117.355 ;
        RECT 25.530 116.575 26.900 117.355 ;
        RECT 26.920 116.445 28.270 117.355 ;
        RECT 28.290 116.675 37.570 117.355 ;
        RECT 29.650 116.455 30.570 116.675 ;
        RECT 35.235 116.555 37.570 116.675 ;
        RECT 36.650 116.445 37.570 116.555 ;
        RECT 38.320 116.675 47.600 117.355 ;
        RECT 38.320 116.555 40.655 116.675 ;
        RECT 38.320 116.445 39.240 116.555 ;
        RECT 45.320 116.455 46.240 116.675 ;
        RECT 47.620 116.485 48.050 117.270 ;
        RECT 49.220 116.675 53.120 117.355 ;
        RECT 52.190 116.445 53.120 116.675 ;
        RECT 53.500 116.675 62.780 117.355 ;
        RECT 53.500 116.555 55.835 116.675 ;
        RECT 53.500 116.445 54.420 116.555 ;
        RECT 60.500 116.455 61.420 116.675 ;
        RECT 63.250 116.545 66.000 117.355 ;
        RECT 66.020 116.445 67.370 117.355 ;
        RECT 67.620 116.675 71.520 117.355 ;
        RECT 70.590 116.445 71.520 116.675 ;
        RECT 71.530 116.575 72.900 117.355 ;
        RECT 73.380 116.485 73.810 117.270 ;
        RECT 75.120 116.675 84.400 117.355 ;
        RECT 84.780 116.675 94.060 117.355 ;
        RECT 95.220 116.675 99.120 117.355 ;
        RECT 75.120 116.555 77.455 116.675 ;
        RECT 75.120 116.445 76.040 116.555 ;
        RECT 82.120 116.455 83.040 116.675 ;
        RECT 84.780 116.555 87.115 116.675 ;
        RECT 84.780 116.445 85.700 116.555 ;
        RECT 91.780 116.455 92.700 116.675 ;
        RECT 98.190 116.445 99.120 116.675 ;
        RECT 99.140 116.485 99.570 117.270 ;
        RECT 99.960 116.675 109.240 117.355 ;
        RECT 99.960 116.555 102.295 116.675 ;
        RECT 99.960 116.445 100.880 116.555 ;
        RECT 106.960 116.455 107.880 116.675 ;
        RECT 109.250 116.545 111.080 117.355 ;
        RECT 111.090 116.545 112.460 117.355 ;
      LAYER nwell ;
        RECT 17.975 113.325 112.655 116.155 ;
      LAYER pwell ;
        RECT 18.170 112.125 19.540 112.935 ;
        RECT 19.750 112.805 21.960 113.035 ;
        RECT 24.680 112.805 25.610 113.025 ;
        RECT 19.750 112.125 30.120 112.805 ;
        RECT 30.130 112.125 31.960 112.935 ;
        RECT 31.970 112.125 33.340 112.905 ;
        RECT 33.360 112.125 34.710 113.035 ;
        RECT 34.740 112.210 35.170 112.995 ;
        RECT 35.650 112.125 37.020 112.905 ;
        RECT 37.030 112.125 40.700 112.935 ;
        RECT 40.720 112.125 42.070 113.035 ;
        RECT 45.290 112.805 46.220 113.035 ;
        RECT 42.320 112.125 46.220 112.805 ;
        RECT 46.230 112.125 47.600 112.905 ;
        RECT 48.070 112.125 50.820 112.935 ;
        RECT 50.830 112.125 56.340 112.935 ;
        RECT 56.360 112.125 57.710 113.035 ;
        RECT 58.190 112.125 59.560 112.905 ;
        RECT 60.500 112.210 60.930 112.995 ;
        RECT 61.410 112.125 63.240 112.935 ;
        RECT 63.250 112.125 68.760 112.935 ;
        RECT 68.780 112.125 70.130 113.035 ;
        RECT 70.610 112.125 72.440 112.935 ;
        RECT 72.450 112.125 77.960 112.935 ;
        RECT 77.980 112.125 79.330 113.035 ;
        RECT 79.810 112.125 81.180 112.905 ;
        RECT 81.200 112.125 82.550 113.035 ;
        RECT 82.570 112.125 86.240 112.935 ;
        RECT 86.260 112.210 86.690 112.995 ;
        RECT 86.710 112.125 88.540 112.935 ;
        RECT 88.550 112.125 89.920 112.905 ;
        RECT 90.850 112.125 96.360 112.935 ;
        RECT 96.370 112.125 97.740 112.905 ;
        RECT 98.210 112.125 100.040 112.935 ;
        RECT 100.050 112.125 105.560 112.935 ;
        RECT 105.570 112.125 111.080 112.935 ;
        RECT 111.090 112.125 112.460 112.935 ;
        RECT 18.310 111.915 18.480 112.125 ;
        RECT 19.745 111.965 19.865 112.075 ;
        RECT 21.530 111.915 21.700 112.105 ;
        RECT 27.510 111.915 27.680 112.105 ;
        RECT 28.890 111.915 29.060 112.105 ;
        RECT 29.405 111.965 29.525 112.075 ;
        RECT 29.810 111.915 29.980 112.125 ;
        RECT 31.650 111.935 31.820 112.125 ;
        RECT 32.110 111.935 32.280 112.125 ;
        RECT 33.490 111.935 33.660 112.125 ;
        RECT 35.385 111.965 35.505 112.075 ;
        RECT 36.710 111.935 36.880 112.125 ;
        RECT 40.390 111.935 40.560 112.125 ;
        RECT 40.850 111.935 41.020 112.125 ;
        RECT 41.310 111.915 41.480 112.105 ;
        RECT 42.230 111.960 42.390 112.070 ;
        RECT 43.610 111.915 43.780 112.105 ;
        RECT 44.990 111.915 45.160 112.105 ;
        RECT 45.450 111.915 45.620 112.105 ;
        RECT 45.635 111.935 45.805 112.125 ;
        RECT 47.290 111.935 47.460 112.125 ;
        RECT 47.805 111.965 47.925 112.075 ;
        RECT 50.510 111.915 50.680 112.125 ;
        RECT 51.890 111.915 52.060 112.105 ;
        RECT 52.405 111.965 52.525 112.075 ;
        RECT 54.190 111.915 54.360 112.105 ;
        RECT 56.030 111.935 56.200 112.125 ;
        RECT 56.490 111.935 56.660 112.125 ;
        RECT 56.945 111.915 57.115 112.105 ;
        RECT 57.925 111.965 58.045 112.075 ;
        RECT 58.330 111.935 58.500 112.125 ;
        RECT 60.170 111.970 60.330 112.080 ;
        RECT 61.145 111.965 61.265 112.075 ;
        RECT 62.930 111.935 63.100 112.125 ;
        RECT 67.530 111.915 67.700 112.105 ;
        RECT 68.450 111.935 68.620 112.125 ;
        RECT 68.910 111.915 69.080 112.105 ;
        RECT 69.830 111.935 70.000 112.125 ;
        RECT 70.290 112.075 70.460 112.105 ;
        RECT 70.290 111.965 70.465 112.075 ;
        RECT 70.290 111.915 70.460 111.965 ;
        RECT 70.755 111.915 70.925 112.105 ;
        RECT 72.130 111.935 72.300 112.125 ;
        RECT 77.190 111.915 77.360 112.105 ;
        RECT 77.650 111.915 77.820 112.125 ;
        RECT 78.110 111.935 78.280 112.125 ;
        RECT 79.085 111.965 79.205 112.075 ;
        RECT 79.545 111.965 79.665 112.075 ;
        RECT 79.950 111.935 80.120 112.125 ;
        RECT 81.330 111.935 81.500 112.125 ;
        RECT 82.710 111.915 82.880 112.105 ;
        RECT 83.170 111.915 83.340 112.105 ;
        RECT 85.930 111.915 86.100 112.125 ;
        RECT 86.390 111.915 86.560 112.105 ;
        RECT 88.230 111.935 88.400 112.125 ;
        RECT 88.690 111.915 88.860 112.125 ;
        RECT 89.150 111.915 89.320 112.105 ;
        RECT 90.530 111.970 90.690 112.080 ;
        RECT 90.990 111.960 91.150 112.070 ;
        RECT 92.370 111.915 92.540 112.105 ;
        RECT 93.290 111.960 93.450 112.070 ;
        RECT 93.750 111.915 93.920 112.105 ;
        RECT 96.050 111.935 96.220 112.125 ;
        RECT 97.430 111.915 97.600 112.125 ;
        RECT 97.890 112.075 98.060 112.105 ;
        RECT 99.730 112.075 99.900 112.125 ;
        RECT 97.890 111.965 98.065 112.075 ;
        RECT 99.730 111.965 99.905 112.075 ;
        RECT 97.890 111.915 98.060 111.965 ;
        RECT 99.730 111.935 99.900 111.965 ;
        RECT 100.190 111.915 100.360 112.105 ;
        RECT 101.625 111.965 101.745 112.075 ;
        RECT 104.330 111.915 104.500 112.105 ;
        RECT 104.790 111.915 104.960 112.105 ;
        RECT 105.250 111.935 105.420 112.125 ;
        RECT 110.770 112.105 110.940 112.125 ;
        RECT 106.170 111.915 106.340 112.105 ;
        RECT 107.550 111.915 107.720 112.105 ;
        RECT 109.390 111.960 109.550 112.070 ;
        RECT 110.760 111.935 110.940 112.105 ;
        RECT 110.760 111.915 110.930 111.935 ;
        RECT 112.150 111.915 112.320 112.125 ;
        RECT 18.170 111.105 19.540 111.915 ;
        RECT 20.010 111.105 21.840 111.915 ;
        RECT 21.860 111.045 22.290 111.830 ;
        RECT 22.310 111.105 27.820 111.915 ;
        RECT 27.830 111.135 29.200 111.915 ;
        RECT 29.670 111.135 31.040 111.915 ;
        RECT 31.250 111.235 41.620 111.915 ;
        RECT 31.250 111.005 33.460 111.235 ;
        RECT 36.180 111.015 37.110 111.235 ;
        RECT 42.550 111.135 43.920 111.915 ;
        RECT 43.930 111.135 45.300 111.915 ;
        RECT 45.310 111.135 46.680 111.915 ;
        RECT 47.620 111.045 48.050 111.830 ;
        RECT 48.070 111.105 50.820 111.915 ;
        RECT 50.830 111.135 52.200 111.915 ;
        RECT 52.670 111.105 54.500 111.915 ;
        RECT 54.650 111.005 57.260 111.915 ;
        RECT 57.470 111.235 67.840 111.915 ;
        RECT 57.470 111.005 59.680 111.235 ;
        RECT 62.400 111.015 63.330 111.235 ;
        RECT 67.850 111.105 69.220 111.915 ;
        RECT 69.230 111.135 70.600 111.915 ;
        RECT 70.610 111.005 73.220 111.915 ;
        RECT 73.380 111.045 73.810 111.830 ;
        RECT 73.830 111.105 77.500 111.915 ;
        RECT 77.510 111.135 78.880 111.915 ;
        RECT 79.350 111.105 83.020 111.915 ;
        RECT 83.030 111.135 84.400 111.915 ;
        RECT 84.410 111.105 86.240 111.915 ;
        RECT 86.260 111.005 87.610 111.915 ;
        RECT 87.630 111.105 89.000 111.915 ;
        RECT 89.010 111.135 90.380 111.915 ;
        RECT 91.320 111.005 92.670 111.915 ;
        RECT 93.610 111.135 94.980 111.915 ;
        RECT 94.990 111.105 97.740 111.915 ;
        RECT 97.760 111.005 99.110 111.915 ;
        RECT 99.140 111.045 99.570 111.830 ;
        RECT 100.050 111.135 101.420 111.915 ;
        RECT 101.890 111.105 104.640 111.915 ;
        RECT 104.660 111.005 106.010 111.915 ;
        RECT 106.030 111.135 107.400 111.915 ;
        RECT 107.410 111.135 108.780 111.915 ;
        RECT 109.710 111.135 111.080 111.915 ;
        RECT 111.090 111.105 112.460 111.915 ;
      LAYER nwell ;
        RECT 17.975 107.885 112.655 110.715 ;
      LAYER pwell ;
        RECT 18.170 106.685 19.540 107.495 ;
        RECT 20.010 106.685 22.760 107.495 ;
        RECT 22.780 106.685 24.130 107.595 ;
        RECT 24.350 107.365 26.560 107.595 ;
        RECT 29.280 107.365 30.210 107.585 ;
        RECT 24.350 106.685 34.720 107.365 ;
        RECT 34.740 106.770 35.170 107.555 ;
        RECT 36.110 106.685 37.480 107.465 ;
        RECT 37.690 107.365 39.900 107.595 ;
        RECT 42.620 107.365 43.550 107.585 ;
        RECT 49.190 107.365 51.400 107.595 ;
        RECT 54.120 107.365 55.050 107.585 ;
        RECT 37.690 106.685 48.060 107.365 ;
        RECT 49.190 106.685 59.560 107.365 ;
        RECT 60.500 106.770 60.930 107.555 ;
        RECT 60.950 106.685 62.320 107.465 ;
        RECT 63.250 106.685 64.620 107.465 ;
        RECT 64.830 107.365 67.040 107.595 ;
        RECT 69.760 107.365 70.690 107.585 ;
        RECT 75.870 107.365 78.080 107.595 ;
        RECT 80.800 107.365 81.730 107.585 ;
        RECT 64.830 106.685 75.200 107.365 ;
        RECT 75.870 106.685 86.240 107.365 ;
        RECT 86.260 106.770 86.690 107.555 ;
        RECT 86.910 107.365 89.120 107.595 ;
        RECT 91.840 107.365 92.770 107.585 ;
        RECT 86.910 106.685 97.280 107.365 ;
        RECT 97.290 106.685 98.660 107.465 ;
        RECT 98.680 106.685 100.030 107.595 ;
        RECT 100.710 107.365 102.920 107.595 ;
        RECT 105.640 107.365 106.570 107.585 ;
        RECT 100.710 106.685 111.080 107.365 ;
        RECT 111.090 106.685 112.460 107.495 ;
        RECT 18.310 106.475 18.480 106.685 ;
        RECT 19.745 106.525 19.865 106.635 ;
        RECT 21.530 106.475 21.700 106.665 ;
        RECT 22.450 106.495 22.620 106.685 ;
        RECT 23.370 106.475 23.540 106.665 ;
        RECT 23.830 106.475 24.000 106.685 ;
        RECT 25.210 106.475 25.380 106.665 ;
        RECT 34.410 106.495 34.580 106.685 ;
        RECT 35.790 106.530 35.950 106.640 ;
        RECT 36.710 106.475 36.880 106.665 ;
        RECT 37.170 106.475 37.340 106.685 ;
        RECT 47.750 106.495 47.920 106.685 ;
        RECT 48.670 106.530 48.830 106.640 ;
        RECT 49.130 106.475 49.300 106.665 ;
        RECT 50.510 106.475 50.680 106.665 ;
        RECT 51.890 106.475 52.060 106.665 ;
        RECT 52.350 106.475 52.520 106.665 ;
        RECT 53.730 106.475 53.900 106.665 ;
        RECT 59.250 106.495 59.420 106.685 ;
        RECT 60.170 106.530 60.330 106.640 ;
        RECT 61.090 106.495 61.260 106.685 ;
        RECT 62.930 106.530 63.090 106.640 ;
        RECT 63.390 106.495 63.560 106.685 ;
        RECT 65.230 106.475 65.400 106.665 ;
        RECT 65.745 106.525 65.865 106.635 ;
        RECT 68.450 106.475 68.620 106.665 ;
        RECT 69.830 106.475 70.000 106.665 ;
        RECT 71.210 106.475 71.380 106.665 ;
        RECT 71.725 106.525 71.845 106.635 ;
        RECT 72.130 106.475 72.300 106.665 ;
        RECT 74.890 106.495 75.060 106.685 ;
        RECT 75.405 106.525 75.525 106.635 ;
        RECT 84.090 106.475 84.260 106.665 ;
        RECT 85.930 106.495 86.100 106.685 ;
        RECT 94.670 106.475 94.840 106.665 ;
        RECT 96.970 106.495 97.140 106.685 ;
        RECT 97.430 106.475 97.600 106.665 ;
        RECT 97.890 106.475 98.060 106.665 ;
        RECT 98.350 106.495 98.520 106.685 ;
        RECT 99.730 106.495 99.900 106.685 ;
        RECT 100.245 106.525 100.365 106.635 ;
        RECT 109.850 106.475 110.020 106.665 ;
        RECT 110.770 106.495 110.940 106.685 ;
        RECT 112.150 106.475 112.320 106.685 ;
        RECT 18.170 105.665 19.540 106.475 ;
        RECT 20.010 105.665 21.840 106.475 ;
        RECT 21.860 105.605 22.290 106.390 ;
        RECT 22.310 105.665 23.680 106.475 ;
        RECT 23.700 105.565 25.050 106.475 ;
        RECT 25.080 105.565 26.430 106.475 ;
        RECT 26.650 105.795 37.020 106.475 ;
        RECT 37.030 105.795 47.400 106.475 ;
        RECT 26.650 105.565 28.860 105.795 ;
        RECT 31.580 105.575 32.510 105.795 ;
        RECT 41.540 105.575 42.470 105.795 ;
        RECT 45.190 105.565 47.400 105.795 ;
        RECT 47.620 105.605 48.050 106.390 ;
        RECT 48.070 105.665 49.440 106.475 ;
        RECT 49.460 105.565 50.810 106.475 ;
        RECT 50.830 105.665 52.200 106.475 ;
        RECT 52.220 105.565 53.570 106.475 ;
        RECT 53.590 105.695 54.960 106.475 ;
        RECT 55.170 105.795 65.540 106.475 ;
        RECT 55.170 105.565 57.380 105.795 ;
        RECT 60.100 105.575 61.030 105.795 ;
        RECT 66.010 105.665 68.760 106.475 ;
        RECT 68.780 105.565 70.130 106.475 ;
        RECT 70.160 105.565 71.510 106.475 ;
        RECT 71.990 105.695 73.360 106.475 ;
        RECT 73.380 105.605 73.810 106.390 ;
        RECT 74.030 105.795 84.400 106.475 ;
        RECT 84.610 105.795 94.980 106.475 ;
        RECT 74.030 105.565 76.240 105.795 ;
        RECT 78.960 105.575 79.890 105.795 ;
        RECT 84.610 105.565 86.820 105.795 ;
        RECT 89.540 105.575 90.470 105.795 ;
        RECT 94.990 105.665 97.740 106.475 ;
        RECT 97.760 105.565 99.110 106.475 ;
        RECT 99.140 105.605 99.570 106.390 ;
        RECT 99.790 105.795 110.160 106.475 ;
        RECT 99.790 105.565 102.000 105.795 ;
        RECT 104.720 105.575 105.650 105.795 ;
        RECT 111.090 105.665 112.460 106.475 ;
      LAYER nwell ;
        RECT 17.975 102.445 112.655 105.275 ;
      LAYER pwell ;
        RECT 18.170 101.245 19.540 102.055 ;
        RECT 20.010 101.245 21.840 102.055 ;
        RECT 21.860 101.330 22.290 102.115 ;
        RECT 22.510 101.925 24.720 102.155 ;
        RECT 27.440 101.925 28.370 102.145 ;
        RECT 22.510 101.245 32.880 101.925 ;
        RECT 32.890 101.245 34.720 102.055 ;
        RECT 34.740 101.330 35.170 102.115 ;
        RECT 35.650 101.245 38.400 102.055 ;
        RECT 38.420 101.245 39.770 102.155 ;
        RECT 39.790 101.245 41.160 102.055 ;
        RECT 41.180 101.245 42.530 102.155 ;
        RECT 42.550 101.245 43.920 102.055 ;
        RECT 43.930 101.245 47.600 102.055 ;
        RECT 47.620 101.330 48.050 102.115 ;
        RECT 48.530 101.245 52.200 102.055 ;
        RECT 52.210 101.245 57.720 102.055 ;
        RECT 57.740 101.245 59.090 102.155 ;
        RECT 59.120 101.245 60.470 102.155 ;
        RECT 60.500 101.330 60.930 102.115 ;
        RECT 60.950 101.245 62.780 102.055 ;
        RECT 67.300 101.925 68.230 102.145 ;
        RECT 70.950 101.925 73.160 102.155 ;
        RECT 62.790 101.245 73.160 101.925 ;
        RECT 73.380 101.330 73.810 102.115 ;
        RECT 73.830 101.245 76.580 102.055 ;
        RECT 76.600 101.245 77.950 102.155 ;
        RECT 77.970 101.245 81.640 102.055 ;
        RECT 81.660 101.245 83.010 102.155 ;
        RECT 83.490 101.245 86.240 102.055 ;
        RECT 86.260 101.330 86.690 102.115 ;
        RECT 86.710 101.245 88.540 102.055 ;
        RECT 88.750 101.925 90.960 102.155 ;
        RECT 93.680 101.925 94.610 102.145 ;
        RECT 88.750 101.245 99.120 101.925 ;
        RECT 99.140 101.330 99.570 102.115 ;
        RECT 100.710 101.925 102.920 102.155 ;
        RECT 105.640 101.925 106.570 102.145 ;
        RECT 100.710 101.245 111.080 101.925 ;
        RECT 111.090 101.245 112.460 102.055 ;
        RECT 18.310 101.055 18.480 101.245 ;
        RECT 19.745 101.085 19.865 101.195 ;
        RECT 21.530 101.055 21.700 101.245 ;
        RECT 32.570 101.055 32.740 101.245 ;
        RECT 34.410 101.055 34.580 101.245 ;
        RECT 35.385 101.085 35.505 101.195 ;
        RECT 38.090 101.055 38.260 101.245 ;
        RECT 39.470 101.055 39.640 101.245 ;
        RECT 40.850 101.055 41.020 101.245 ;
        RECT 41.310 101.055 41.480 101.245 ;
        RECT 43.610 101.055 43.780 101.245 ;
        RECT 47.290 101.055 47.460 101.245 ;
        RECT 48.265 101.085 48.385 101.195 ;
        RECT 51.890 101.055 52.060 101.245 ;
        RECT 57.410 101.055 57.580 101.245 ;
        RECT 57.870 101.055 58.040 101.245 ;
        RECT 59.250 101.055 59.420 101.245 ;
        RECT 62.470 101.055 62.640 101.245 ;
        RECT 62.930 101.055 63.100 101.245 ;
        RECT 76.270 101.055 76.440 101.245 ;
        RECT 76.730 101.055 76.900 101.245 ;
        RECT 81.330 101.055 81.500 101.245 ;
        RECT 82.710 101.055 82.880 101.245 ;
        RECT 83.225 101.085 83.345 101.195 ;
        RECT 85.930 101.055 86.100 101.245 ;
        RECT 88.230 101.055 88.400 101.245 ;
        RECT 98.810 101.055 98.980 101.245 ;
        RECT 100.190 101.090 100.350 101.200 ;
        RECT 110.770 101.055 110.940 101.245 ;
        RECT 112.150 101.055 112.320 101.245 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 18.165 193.535 112.465 193.705 ;
        RECT 18.250 192.785 19.460 193.535 ;
        RECT 18.250 192.245 18.770 192.785 ;
        RECT 20.590 192.715 20.820 193.535 ;
        RECT 20.990 192.735 21.320 193.365 ;
        RECT 18.940 192.075 19.460 192.615 ;
        RECT 20.570 192.295 20.900 192.545 ;
        RECT 21.070 192.135 21.320 192.735 ;
        RECT 21.490 192.715 21.700 193.535 ;
        RECT 21.930 192.810 22.220 193.535 ;
        RECT 22.390 192.765 24.980 193.535 ;
        RECT 25.155 192.990 30.500 193.535 ;
        RECT 18.250 190.985 19.460 192.075 ;
        RECT 20.590 190.985 20.820 192.125 ;
        RECT 20.990 191.155 21.320 192.135 ;
        RECT 21.490 190.985 21.700 192.125 ;
        RECT 21.930 190.985 22.220 192.150 ;
        RECT 22.390 192.075 23.600 192.595 ;
        RECT 23.770 192.245 24.980 192.765 ;
        RECT 22.390 190.985 24.980 192.075 ;
        RECT 26.745 191.420 27.095 192.670 ;
        RECT 28.575 192.160 28.915 192.990 ;
        RECT 30.760 192.985 30.930 193.365 ;
        RECT 31.110 193.155 31.440 193.535 ;
        RECT 30.760 192.815 31.425 192.985 ;
        RECT 31.620 192.860 31.880 193.365 ;
        RECT 30.690 192.265 31.020 192.635 ;
        RECT 31.255 192.560 31.425 192.815 ;
        RECT 31.255 192.230 31.540 192.560 ;
        RECT 31.255 192.085 31.425 192.230 ;
        RECT 30.760 191.915 31.425 192.085 ;
        RECT 31.710 192.060 31.880 192.860 ;
        RECT 32.050 192.765 34.640 193.535 ;
        RECT 34.810 192.810 35.100 193.535 ;
        RECT 35.730 192.765 37.400 193.535 ;
        RECT 37.575 192.990 42.920 193.535 ;
        RECT 25.155 190.985 30.500 191.420 ;
        RECT 30.760 191.155 30.930 191.915 ;
        RECT 31.110 190.985 31.440 191.745 ;
        RECT 31.610 191.155 31.880 192.060 ;
        RECT 32.050 192.075 33.260 192.595 ;
        RECT 33.430 192.245 34.640 192.765 ;
        RECT 32.050 190.985 34.640 192.075 ;
        RECT 34.810 190.985 35.100 192.150 ;
        RECT 35.730 192.075 36.480 192.595 ;
        RECT 36.650 192.245 37.400 192.765 ;
        RECT 35.730 190.985 37.400 192.075 ;
        RECT 39.165 191.420 39.515 192.670 ;
        RECT 40.995 192.160 41.335 192.990 ;
        RECT 43.150 192.715 43.360 193.535 ;
        RECT 43.530 192.735 43.860 193.365 ;
        RECT 43.530 192.135 43.780 192.735 ;
        RECT 44.030 192.715 44.260 193.535 ;
        RECT 44.470 192.785 45.680 193.535 ;
        RECT 43.950 192.295 44.280 192.545 ;
        RECT 37.575 190.985 42.920 191.420 ;
        RECT 43.150 190.985 43.360 192.125 ;
        RECT 43.530 191.155 43.860 192.135 ;
        RECT 44.030 190.985 44.260 192.125 ;
        RECT 44.470 192.075 44.990 192.615 ;
        RECT 45.160 192.245 45.680 192.785 ;
        RECT 45.850 192.860 46.110 193.365 ;
        RECT 46.290 193.155 46.620 193.535 ;
        RECT 46.800 192.985 46.970 193.365 ;
        RECT 44.470 190.985 45.680 192.075 ;
        RECT 45.850 192.060 46.020 192.860 ;
        RECT 46.305 192.815 46.970 192.985 ;
        RECT 46.305 192.560 46.475 192.815 ;
        RECT 47.690 192.810 47.980 193.535 ;
        RECT 48.150 192.765 51.660 193.535 ;
        RECT 46.190 192.230 46.475 192.560 ;
        RECT 46.710 192.265 47.040 192.635 ;
        RECT 46.305 192.085 46.475 192.230 ;
        RECT 45.850 191.155 46.120 192.060 ;
        RECT 46.305 191.915 46.970 192.085 ;
        RECT 46.290 190.985 46.620 191.745 ;
        RECT 46.800 191.155 46.970 191.915 ;
        RECT 47.690 190.985 47.980 192.150 ;
        RECT 48.150 192.075 49.840 192.595 ;
        RECT 50.010 192.245 51.660 192.765 ;
        RECT 51.890 192.715 52.100 193.535 ;
        RECT 52.270 192.735 52.600 193.365 ;
        RECT 52.270 192.135 52.520 192.735 ;
        RECT 52.770 192.715 53.000 193.535 ;
        RECT 53.210 192.765 54.880 193.535 ;
        RECT 55.055 192.990 60.400 193.535 ;
        RECT 52.690 192.295 53.020 192.545 ;
        RECT 48.150 190.985 51.660 192.075 ;
        RECT 51.890 190.985 52.100 192.125 ;
        RECT 52.270 191.155 52.600 192.135 ;
        RECT 52.770 190.985 53.000 192.125 ;
        RECT 53.210 192.075 53.960 192.595 ;
        RECT 54.130 192.245 54.880 192.765 ;
        RECT 53.210 190.985 54.880 192.075 ;
        RECT 56.645 191.420 56.995 192.670 ;
        RECT 58.475 192.160 58.815 192.990 ;
        RECT 60.570 192.810 60.860 193.535 ;
        RECT 61.030 192.765 63.620 193.535 ;
        RECT 55.055 190.985 60.400 191.420 ;
        RECT 60.570 190.985 60.860 192.150 ;
        RECT 61.030 192.075 62.240 192.595 ;
        RECT 62.410 192.245 63.620 192.765 ;
        RECT 63.850 192.715 64.060 193.535 ;
        RECT 64.230 192.735 64.560 193.365 ;
        RECT 64.230 192.135 64.480 192.735 ;
        RECT 64.730 192.715 64.960 193.535 ;
        RECT 65.690 192.715 65.900 193.535 ;
        RECT 66.070 192.735 66.400 193.365 ;
        RECT 64.650 192.295 64.980 192.545 ;
        RECT 66.070 192.135 66.320 192.735 ;
        RECT 66.570 192.715 66.800 193.535 ;
        RECT 67.935 192.990 73.280 193.535 ;
        RECT 66.490 192.295 66.820 192.545 ;
        RECT 61.030 190.985 63.620 192.075 ;
        RECT 63.850 190.985 64.060 192.125 ;
        RECT 64.230 191.155 64.560 192.135 ;
        RECT 64.730 190.985 64.960 192.125 ;
        RECT 65.690 190.985 65.900 192.125 ;
        RECT 66.070 191.155 66.400 192.135 ;
        RECT 66.570 190.985 66.800 192.125 ;
        RECT 69.525 191.420 69.875 192.670 ;
        RECT 71.355 192.160 71.695 192.990 ;
        RECT 73.450 192.810 73.740 193.535 ;
        RECT 74.370 192.765 76.040 193.535 ;
        RECT 67.935 190.985 73.280 191.420 ;
        RECT 73.450 190.985 73.740 192.150 ;
        RECT 74.370 192.075 75.120 192.595 ;
        RECT 75.290 192.245 76.040 192.765 ;
        RECT 76.485 192.725 76.730 193.330 ;
        RECT 76.950 193.000 77.460 193.535 ;
        RECT 76.210 192.555 77.440 192.725 ;
        RECT 74.370 190.985 76.040 192.075 ;
        RECT 76.210 191.745 76.550 192.555 ;
        RECT 76.720 191.990 77.470 192.180 ;
        RECT 76.210 191.335 76.725 191.745 ;
        RECT 76.960 190.985 77.130 191.745 ;
        RECT 77.300 191.325 77.470 191.990 ;
        RECT 77.640 192.005 77.830 193.365 ;
        RECT 78.000 192.515 78.275 193.365 ;
        RECT 78.465 193.000 78.995 193.365 ;
        RECT 79.420 193.135 79.750 193.535 ;
        RECT 78.820 192.965 78.995 193.000 ;
        RECT 78.000 192.345 78.280 192.515 ;
        RECT 78.000 192.205 78.275 192.345 ;
        RECT 78.480 192.005 78.650 192.805 ;
        RECT 77.640 191.835 78.650 192.005 ;
        RECT 78.820 192.795 79.750 192.965 ;
        RECT 79.920 192.795 80.175 193.365 ;
        RECT 80.815 192.990 86.160 193.535 ;
        RECT 78.820 191.665 78.990 192.795 ;
        RECT 79.580 192.625 79.750 192.795 ;
        RECT 77.865 191.495 78.990 191.665 ;
        RECT 79.160 192.295 79.355 192.625 ;
        RECT 79.580 192.295 79.835 192.625 ;
        RECT 79.160 191.325 79.330 192.295 ;
        RECT 80.005 192.125 80.175 192.795 ;
        RECT 77.300 191.155 79.330 191.325 ;
        RECT 79.500 190.985 79.670 192.125 ;
        RECT 79.840 191.155 80.175 192.125 ;
        RECT 82.405 191.420 82.755 192.670 ;
        RECT 84.235 192.160 84.575 192.990 ;
        RECT 86.330 192.810 86.620 193.535 ;
        RECT 86.790 192.765 88.460 193.535 ;
        RECT 80.815 190.985 86.160 191.420 ;
        RECT 86.330 190.985 86.620 192.150 ;
        RECT 86.790 192.075 87.540 192.595 ;
        RECT 87.710 192.245 88.460 192.765 ;
        RECT 88.630 192.860 88.890 193.365 ;
        RECT 89.070 193.155 89.400 193.535 ;
        RECT 89.580 192.985 89.750 193.365 ;
        RECT 90.935 192.990 96.280 193.535 ;
        RECT 86.790 190.985 88.460 192.075 ;
        RECT 88.630 192.060 88.800 192.860 ;
        RECT 89.085 192.815 89.750 192.985 ;
        RECT 89.085 192.560 89.255 192.815 ;
        RECT 88.970 192.230 89.255 192.560 ;
        RECT 89.490 192.265 89.820 192.635 ;
        RECT 89.085 192.085 89.255 192.230 ;
        RECT 88.630 191.155 88.900 192.060 ;
        RECT 89.085 191.915 89.750 192.085 ;
        RECT 89.070 190.985 89.400 191.745 ;
        RECT 89.580 191.155 89.750 191.915 ;
        RECT 92.525 191.420 92.875 192.670 ;
        RECT 94.355 192.160 94.695 192.990 ;
        RECT 96.490 192.715 96.720 193.535 ;
        RECT 96.890 192.735 97.220 193.365 ;
        RECT 96.470 192.295 96.800 192.545 ;
        RECT 96.970 192.135 97.220 192.735 ;
        RECT 97.390 192.715 97.600 193.535 ;
        RECT 97.830 192.785 99.040 193.535 ;
        RECT 99.210 192.810 99.500 193.535 ;
        RECT 99.760 192.985 99.930 193.365 ;
        RECT 100.110 193.155 100.440 193.535 ;
        RECT 99.760 192.815 100.425 192.985 ;
        RECT 100.620 192.860 100.880 193.365 ;
        RECT 90.935 190.985 96.280 191.420 ;
        RECT 96.490 190.985 96.720 192.125 ;
        RECT 96.890 191.155 97.220 192.135 ;
        RECT 97.390 190.985 97.600 192.125 ;
        RECT 97.830 192.075 98.350 192.615 ;
        RECT 98.520 192.245 99.040 192.785 ;
        RECT 99.690 192.265 100.020 192.635 ;
        RECT 100.255 192.560 100.425 192.815 ;
        RECT 100.255 192.230 100.540 192.560 ;
        RECT 97.830 190.985 99.040 192.075 ;
        RECT 99.210 190.985 99.500 192.150 ;
        RECT 100.255 192.085 100.425 192.230 ;
        RECT 99.760 191.915 100.425 192.085 ;
        RECT 100.710 192.060 100.880 192.860 ;
        RECT 99.760 191.155 99.930 191.915 ;
        RECT 100.110 190.985 100.440 191.745 ;
        RECT 100.610 191.155 100.880 192.060 ;
        RECT 101.515 192.825 101.770 193.355 ;
        RECT 101.940 193.075 102.245 193.535 ;
        RECT 102.490 193.155 103.560 193.325 ;
        RECT 101.515 192.175 101.725 192.825 ;
        RECT 102.490 192.800 102.810 193.155 ;
        RECT 102.485 192.625 102.810 192.800 ;
        RECT 101.895 192.325 102.810 192.625 ;
        RECT 102.980 192.585 103.220 192.985 ;
        RECT 103.390 192.925 103.560 193.155 ;
        RECT 103.730 193.095 103.920 193.535 ;
        RECT 104.090 193.085 105.040 193.365 ;
        RECT 105.260 193.175 105.610 193.345 ;
        RECT 103.390 192.755 103.920 192.925 ;
        RECT 101.895 192.295 102.635 192.325 ;
        RECT 101.515 191.295 101.770 192.175 ;
        RECT 101.940 190.985 102.245 192.125 ;
        RECT 102.465 191.705 102.635 192.295 ;
        RECT 102.980 192.215 103.520 192.585 ;
        RECT 103.700 192.475 103.920 192.755 ;
        RECT 104.090 192.305 104.260 193.085 ;
        RECT 103.855 192.135 104.260 192.305 ;
        RECT 104.430 192.295 104.780 192.915 ;
        RECT 103.855 192.045 104.025 192.135 ;
        RECT 104.950 192.125 105.160 192.915 ;
        RECT 102.805 191.875 104.025 192.045 ;
        RECT 104.485 191.965 105.160 192.125 ;
        RECT 102.465 191.535 103.265 191.705 ;
        RECT 102.585 190.985 102.915 191.365 ;
        RECT 103.095 191.245 103.265 191.535 ;
        RECT 103.855 191.495 104.025 191.875 ;
        RECT 104.195 191.955 105.160 191.965 ;
        RECT 105.350 192.785 105.610 193.175 ;
        RECT 105.820 193.075 106.150 193.535 ;
        RECT 107.025 193.145 107.880 193.315 ;
        RECT 108.085 193.145 108.580 193.315 ;
        RECT 108.750 193.175 109.080 193.535 ;
        RECT 105.350 192.095 105.520 192.785 ;
        RECT 105.690 192.435 105.860 192.615 ;
        RECT 106.030 192.605 106.820 192.855 ;
        RECT 107.025 192.435 107.195 193.145 ;
        RECT 107.365 192.635 107.720 192.855 ;
        RECT 105.690 192.265 107.380 192.435 ;
        RECT 104.195 191.665 104.655 191.955 ;
        RECT 105.350 191.925 106.850 192.095 ;
        RECT 105.350 191.785 105.520 191.925 ;
        RECT 104.960 191.615 105.520 191.785 ;
        RECT 103.435 190.985 103.685 191.445 ;
        RECT 103.855 191.155 104.725 191.495 ;
        RECT 104.960 191.155 105.130 191.615 ;
        RECT 105.965 191.585 107.040 191.755 ;
        RECT 105.300 190.985 105.670 191.445 ;
        RECT 105.965 191.245 106.135 191.585 ;
        RECT 106.305 190.985 106.635 191.415 ;
        RECT 106.870 191.245 107.040 191.585 ;
        RECT 107.210 191.485 107.380 192.265 ;
        RECT 107.550 192.045 107.720 192.635 ;
        RECT 107.890 192.235 108.240 192.855 ;
        RECT 107.550 191.655 108.015 192.045 ;
        RECT 108.410 191.785 108.580 193.145 ;
        RECT 108.750 191.955 109.210 193.005 ;
        RECT 108.185 191.615 108.580 191.785 ;
        RECT 108.185 191.485 108.355 191.615 ;
        RECT 107.210 191.155 107.890 191.485 ;
        RECT 108.105 191.155 108.355 191.485 ;
        RECT 108.525 190.985 108.775 191.445 ;
        RECT 108.945 191.170 109.270 191.955 ;
        RECT 109.440 191.155 109.610 193.275 ;
        RECT 109.780 193.155 110.110 193.535 ;
        RECT 110.280 192.985 110.535 193.275 ;
        RECT 109.785 192.815 110.535 192.985 ;
        RECT 109.785 191.825 110.015 192.815 ;
        RECT 111.170 192.785 112.380 193.535 ;
        RECT 110.185 191.995 110.535 192.645 ;
        RECT 111.170 192.075 111.690 192.615 ;
        RECT 111.860 192.245 112.380 192.785 ;
        RECT 109.785 191.655 110.535 191.825 ;
        RECT 109.780 190.985 110.110 191.485 ;
        RECT 110.280 191.155 110.535 191.655 ;
        RECT 111.170 190.985 112.380 192.075 ;
        RECT 18.165 190.815 112.465 190.985 ;
        RECT 18.250 189.725 19.460 190.815 ;
        RECT 20.665 190.185 20.950 190.645 ;
        RECT 21.120 190.355 21.390 190.815 ;
        RECT 20.665 189.965 21.620 190.185 ;
        RECT 18.250 189.015 18.770 189.555 ;
        RECT 18.940 189.185 19.460 189.725 ;
        RECT 20.550 189.235 21.240 189.795 ;
        RECT 21.410 189.065 21.620 189.965 ;
        RECT 18.250 188.265 19.460 189.015 ;
        RECT 20.665 188.895 21.620 189.065 ;
        RECT 21.790 189.795 22.190 190.645 ;
        RECT 22.380 190.185 22.660 190.645 ;
        RECT 23.180 190.355 23.505 190.815 ;
        RECT 22.380 189.965 23.505 190.185 ;
        RECT 21.790 189.235 22.885 189.795 ;
        RECT 23.055 189.505 23.505 189.965 ;
        RECT 23.675 189.675 24.060 190.645 ;
        RECT 20.665 188.435 20.950 188.895 ;
        RECT 21.120 188.265 21.390 188.725 ;
        RECT 21.790 188.435 22.190 189.235 ;
        RECT 23.055 189.175 23.610 189.505 ;
        RECT 23.055 189.065 23.505 189.175 ;
        RECT 22.380 188.895 23.505 189.065 ;
        RECT 23.780 189.005 24.060 189.675 ;
        RECT 22.380 188.435 22.660 188.895 ;
        RECT 23.180 188.265 23.505 188.725 ;
        RECT 23.675 188.435 24.060 189.005 ;
        RECT 24.235 189.625 24.490 190.505 ;
        RECT 24.660 189.675 24.965 190.815 ;
        RECT 25.305 190.435 25.635 190.815 ;
        RECT 25.815 190.265 25.985 190.555 ;
        RECT 26.155 190.355 26.405 190.815 ;
        RECT 25.185 190.095 25.985 190.265 ;
        RECT 26.575 190.305 27.445 190.645 ;
        RECT 24.235 188.975 24.445 189.625 ;
        RECT 25.185 189.505 25.355 190.095 ;
        RECT 26.575 189.925 26.745 190.305 ;
        RECT 27.680 190.185 27.850 190.645 ;
        RECT 28.020 190.355 28.390 190.815 ;
        RECT 28.685 190.215 28.855 190.555 ;
        RECT 29.025 190.385 29.355 190.815 ;
        RECT 29.590 190.215 29.760 190.555 ;
        RECT 25.525 189.755 26.745 189.925 ;
        RECT 26.915 189.845 27.375 190.135 ;
        RECT 27.680 190.015 28.240 190.185 ;
        RECT 28.685 190.045 29.760 190.215 ;
        RECT 29.930 190.315 30.610 190.645 ;
        RECT 30.825 190.315 31.075 190.645 ;
        RECT 31.245 190.355 31.495 190.815 ;
        RECT 28.070 189.875 28.240 190.015 ;
        RECT 26.915 189.835 27.880 189.845 ;
        RECT 26.575 189.665 26.745 189.755 ;
        RECT 27.205 189.675 27.880 189.835 ;
        RECT 24.615 189.475 25.355 189.505 ;
        RECT 24.615 189.175 25.530 189.475 ;
        RECT 25.205 189.000 25.530 189.175 ;
        RECT 24.235 188.445 24.490 188.975 ;
        RECT 24.660 188.265 24.965 188.725 ;
        RECT 25.210 188.645 25.530 189.000 ;
        RECT 25.700 189.215 26.240 189.585 ;
        RECT 26.575 189.495 26.980 189.665 ;
        RECT 25.700 188.815 25.940 189.215 ;
        RECT 26.420 189.045 26.640 189.325 ;
        RECT 26.110 188.875 26.640 189.045 ;
        RECT 26.110 188.645 26.280 188.875 ;
        RECT 26.810 188.715 26.980 189.495 ;
        RECT 27.150 188.885 27.500 189.505 ;
        RECT 27.670 188.885 27.880 189.675 ;
        RECT 28.070 189.705 29.570 189.875 ;
        RECT 28.070 189.015 28.240 189.705 ;
        RECT 29.930 189.535 30.100 190.315 ;
        RECT 30.905 190.185 31.075 190.315 ;
        RECT 28.410 189.365 30.100 189.535 ;
        RECT 30.270 189.755 30.735 190.145 ;
        RECT 30.905 190.015 31.300 190.185 ;
        RECT 28.410 189.185 28.580 189.365 ;
        RECT 25.210 188.475 26.280 188.645 ;
        RECT 26.450 188.265 26.640 188.705 ;
        RECT 26.810 188.435 27.760 188.715 ;
        RECT 28.070 188.625 28.330 189.015 ;
        RECT 28.750 188.945 29.540 189.195 ;
        RECT 27.980 188.455 28.330 188.625 ;
        RECT 28.540 188.265 28.870 188.725 ;
        RECT 29.745 188.655 29.915 189.365 ;
        RECT 30.270 189.165 30.440 189.755 ;
        RECT 30.085 188.945 30.440 189.165 ;
        RECT 30.610 188.945 30.960 189.565 ;
        RECT 31.130 188.655 31.300 190.015 ;
        RECT 31.665 189.845 31.990 190.630 ;
        RECT 31.470 188.795 31.930 189.845 ;
        RECT 29.745 188.485 30.600 188.655 ;
        RECT 30.805 188.485 31.300 188.655 ;
        RECT 31.470 188.265 31.800 188.625 ;
        RECT 32.160 188.525 32.330 190.645 ;
        RECT 32.500 190.315 32.830 190.815 ;
        RECT 33.000 190.145 33.255 190.645 ;
        RECT 32.505 189.975 33.255 190.145 ;
        RECT 32.505 188.985 32.735 189.975 ;
        RECT 32.905 189.155 33.255 189.805 ;
        RECT 33.430 189.725 34.640 190.815 ;
        RECT 33.430 189.185 33.950 189.725 ;
        RECT 34.810 189.650 35.100 190.815 ;
        RECT 36.565 189.835 36.820 190.505 ;
        RECT 37.000 190.015 37.285 190.815 ;
        RECT 37.465 190.095 37.795 190.605 ;
        RECT 34.120 189.015 34.640 189.555 ;
        RECT 32.505 188.815 33.255 188.985 ;
        RECT 32.500 188.265 32.830 188.645 ;
        RECT 33.000 188.525 33.255 188.815 ;
        RECT 33.430 188.265 34.640 189.015 ;
        RECT 34.810 188.265 35.100 188.990 ;
        RECT 36.565 188.975 36.745 189.835 ;
        RECT 37.465 189.505 37.715 190.095 ;
        RECT 38.065 189.945 38.235 190.555 ;
        RECT 38.405 190.125 38.735 190.815 ;
        RECT 38.965 190.265 39.205 190.555 ;
        RECT 39.405 190.435 39.825 190.815 ;
        RECT 40.005 190.345 40.635 190.595 ;
        RECT 41.105 190.435 41.435 190.815 ;
        RECT 40.005 190.265 40.175 190.345 ;
        RECT 41.605 190.265 41.775 190.555 ;
        RECT 41.955 190.435 42.335 190.815 ;
        RECT 42.575 190.430 43.405 190.600 ;
        RECT 38.965 190.095 40.175 190.265 ;
        RECT 36.915 189.175 37.715 189.505 ;
        RECT 36.565 188.775 36.820 188.975 ;
        RECT 36.480 188.605 36.820 188.775 ;
        RECT 36.565 188.445 36.820 188.605 ;
        RECT 37.000 188.265 37.285 188.725 ;
        RECT 37.465 188.525 37.715 189.175 ;
        RECT 37.915 189.925 38.235 189.945 ;
        RECT 37.915 189.755 39.835 189.925 ;
        RECT 37.915 188.860 38.105 189.755 ;
        RECT 40.005 189.585 40.175 190.095 ;
        RECT 40.345 189.835 40.865 190.145 ;
        RECT 38.275 189.415 40.175 189.585 ;
        RECT 38.275 189.355 38.605 189.415 ;
        RECT 38.755 189.185 39.085 189.245 ;
        RECT 38.425 188.915 39.085 189.185 ;
        RECT 37.915 188.530 38.235 188.860 ;
        RECT 38.415 188.265 39.075 188.745 ;
        RECT 39.275 188.655 39.445 189.415 ;
        RECT 40.345 189.245 40.525 189.655 ;
        RECT 39.615 189.075 39.945 189.195 ;
        RECT 40.695 189.075 40.865 189.835 ;
        RECT 39.615 188.905 40.865 189.075 ;
        RECT 41.035 190.015 42.405 190.265 ;
        RECT 41.035 189.245 41.225 190.015 ;
        RECT 42.155 189.755 42.405 190.015 ;
        RECT 41.395 189.585 41.645 189.745 ;
        RECT 42.575 189.585 42.745 190.430 ;
        RECT 43.640 190.145 43.810 190.645 ;
        RECT 43.980 190.315 44.310 190.815 ;
        RECT 42.915 189.755 43.415 190.135 ;
        RECT 43.640 189.975 44.335 190.145 ;
        RECT 41.395 189.415 42.745 189.585 ;
        RECT 42.325 189.375 42.745 189.415 ;
        RECT 41.035 188.905 41.455 189.245 ;
        RECT 41.745 188.915 42.155 189.245 ;
        RECT 39.275 188.485 40.125 188.655 ;
        RECT 40.685 188.265 41.005 188.725 ;
        RECT 41.205 188.475 41.455 188.905 ;
        RECT 41.745 188.265 42.155 188.705 ;
        RECT 42.325 188.645 42.495 189.375 ;
        RECT 42.665 188.825 43.015 189.195 ;
        RECT 43.195 188.885 43.415 189.755 ;
        RECT 43.585 189.185 43.995 189.805 ;
        RECT 44.165 189.005 44.335 189.975 ;
        RECT 43.640 188.815 44.335 189.005 ;
        RECT 42.325 188.445 43.340 188.645 ;
        RECT 43.640 188.485 43.810 188.815 ;
        RECT 43.980 188.265 44.310 188.645 ;
        RECT 44.525 188.525 44.750 190.645 ;
        RECT 44.920 190.315 45.250 190.815 ;
        RECT 45.420 190.145 45.590 190.645 ;
        RECT 44.925 189.975 45.590 190.145 ;
        RECT 44.925 188.985 45.155 189.975 ;
        RECT 45.325 189.155 45.675 189.805 ;
        RECT 46.310 189.740 46.580 190.645 ;
        RECT 46.750 190.055 47.080 190.815 ;
        RECT 47.260 189.885 47.430 190.645 ;
        RECT 47.695 190.145 47.950 190.645 ;
        RECT 48.120 190.315 48.450 190.815 ;
        RECT 47.695 189.975 48.445 190.145 ;
        RECT 44.925 188.815 45.590 188.985 ;
        RECT 44.920 188.265 45.250 188.645 ;
        RECT 45.420 188.525 45.590 188.815 ;
        RECT 46.310 188.940 46.480 189.740 ;
        RECT 46.765 189.715 47.430 189.885 ;
        RECT 46.765 189.570 46.935 189.715 ;
        RECT 46.650 189.240 46.935 189.570 ;
        RECT 46.765 188.985 46.935 189.240 ;
        RECT 47.170 189.165 47.500 189.535 ;
        RECT 47.695 189.155 48.045 189.805 ;
        RECT 48.215 188.985 48.445 189.975 ;
        RECT 46.310 188.435 46.570 188.940 ;
        RECT 46.765 188.815 47.430 188.985 ;
        RECT 46.750 188.265 47.080 188.645 ;
        RECT 47.260 188.435 47.430 188.815 ;
        RECT 47.695 188.815 48.445 188.985 ;
        RECT 47.695 188.525 47.950 188.815 ;
        RECT 48.120 188.265 48.450 188.645 ;
        RECT 48.620 188.525 48.790 190.645 ;
        RECT 48.960 189.845 49.285 190.630 ;
        RECT 49.455 190.355 49.705 190.815 ;
        RECT 49.875 190.315 50.125 190.645 ;
        RECT 50.340 190.315 51.020 190.645 ;
        RECT 49.875 190.185 50.045 190.315 ;
        RECT 49.650 190.015 50.045 190.185 ;
        RECT 49.020 188.795 49.480 189.845 ;
        RECT 49.650 188.655 49.820 190.015 ;
        RECT 50.215 189.755 50.680 190.145 ;
        RECT 49.990 188.945 50.340 189.565 ;
        RECT 50.510 189.165 50.680 189.755 ;
        RECT 50.850 189.535 51.020 190.315 ;
        RECT 51.190 190.215 51.360 190.555 ;
        RECT 51.595 190.385 51.925 190.815 ;
        RECT 52.095 190.215 52.265 190.555 ;
        RECT 52.560 190.355 52.930 190.815 ;
        RECT 51.190 190.045 52.265 190.215 ;
        RECT 53.100 190.185 53.270 190.645 ;
        RECT 53.505 190.305 54.375 190.645 ;
        RECT 54.545 190.355 54.795 190.815 ;
        RECT 52.710 190.015 53.270 190.185 ;
        RECT 52.710 189.875 52.880 190.015 ;
        RECT 51.380 189.705 52.880 189.875 ;
        RECT 53.575 189.845 54.035 190.135 ;
        RECT 50.850 189.365 52.540 189.535 ;
        RECT 50.510 188.945 50.865 189.165 ;
        RECT 51.035 188.655 51.205 189.365 ;
        RECT 51.410 188.945 52.200 189.195 ;
        RECT 52.370 189.185 52.540 189.365 ;
        RECT 52.710 189.015 52.880 189.705 ;
        RECT 49.150 188.265 49.480 188.625 ;
        RECT 49.650 188.485 50.145 188.655 ;
        RECT 50.350 188.485 51.205 188.655 ;
        RECT 52.080 188.265 52.410 188.725 ;
        RECT 52.620 188.625 52.880 189.015 ;
        RECT 53.070 189.835 54.035 189.845 ;
        RECT 54.205 189.925 54.375 190.305 ;
        RECT 54.965 190.265 55.135 190.555 ;
        RECT 55.315 190.435 55.645 190.815 ;
        RECT 54.965 190.095 55.765 190.265 ;
        RECT 53.070 189.675 53.745 189.835 ;
        RECT 54.205 189.755 55.425 189.925 ;
        RECT 53.070 188.885 53.280 189.675 ;
        RECT 54.205 189.665 54.375 189.755 ;
        RECT 53.450 188.885 53.800 189.505 ;
        RECT 53.970 189.495 54.375 189.665 ;
        RECT 53.970 188.715 54.140 189.495 ;
        RECT 54.310 189.045 54.530 189.325 ;
        RECT 54.710 189.215 55.250 189.585 ;
        RECT 55.595 189.505 55.765 190.095 ;
        RECT 55.985 189.675 56.290 190.815 ;
        RECT 56.460 189.625 56.710 190.505 ;
        RECT 56.880 189.675 57.130 190.815 ;
        RECT 57.810 189.725 60.400 190.815 ;
        RECT 55.595 189.475 56.335 189.505 ;
        RECT 54.310 188.875 54.840 189.045 ;
        RECT 52.620 188.455 52.970 188.625 ;
        RECT 53.190 188.435 54.140 188.715 ;
        RECT 54.310 188.265 54.500 188.705 ;
        RECT 54.670 188.645 54.840 188.875 ;
        RECT 55.010 188.815 55.250 189.215 ;
        RECT 55.420 189.175 56.335 189.475 ;
        RECT 55.420 189.000 55.745 189.175 ;
        RECT 55.420 188.645 55.740 189.000 ;
        RECT 56.505 188.975 56.710 189.625 ;
        RECT 57.810 189.205 59.020 189.725 ;
        RECT 60.570 189.650 60.860 190.815 ;
        RECT 61.035 189.625 61.290 190.505 ;
        RECT 61.460 189.675 61.765 190.815 ;
        RECT 62.105 190.435 62.435 190.815 ;
        RECT 62.615 190.265 62.785 190.555 ;
        RECT 62.955 190.355 63.205 190.815 ;
        RECT 61.985 190.095 62.785 190.265 ;
        RECT 63.375 190.305 64.245 190.645 ;
        RECT 59.190 189.035 60.400 189.555 ;
        RECT 54.670 188.475 55.740 188.645 ;
        RECT 55.985 188.265 56.290 188.725 ;
        RECT 56.460 188.445 56.710 188.975 ;
        RECT 56.880 188.265 57.130 189.020 ;
        RECT 57.810 188.265 60.400 189.035 ;
        RECT 60.570 188.265 60.860 188.990 ;
        RECT 61.035 188.975 61.245 189.625 ;
        RECT 61.985 189.505 62.155 190.095 ;
        RECT 63.375 189.925 63.545 190.305 ;
        RECT 64.480 190.185 64.650 190.645 ;
        RECT 64.820 190.355 65.190 190.815 ;
        RECT 65.485 190.215 65.655 190.555 ;
        RECT 65.825 190.385 66.155 190.815 ;
        RECT 66.390 190.215 66.560 190.555 ;
        RECT 62.325 189.755 63.545 189.925 ;
        RECT 63.715 189.845 64.175 190.135 ;
        RECT 64.480 190.015 65.040 190.185 ;
        RECT 65.485 190.045 66.560 190.215 ;
        RECT 66.730 190.315 67.410 190.645 ;
        RECT 67.625 190.315 67.875 190.645 ;
        RECT 68.045 190.355 68.295 190.815 ;
        RECT 64.870 189.875 65.040 190.015 ;
        RECT 63.715 189.835 64.680 189.845 ;
        RECT 63.375 189.665 63.545 189.755 ;
        RECT 64.005 189.675 64.680 189.835 ;
        RECT 61.415 189.475 62.155 189.505 ;
        RECT 61.415 189.175 62.330 189.475 ;
        RECT 62.005 189.000 62.330 189.175 ;
        RECT 61.035 188.445 61.290 188.975 ;
        RECT 61.460 188.265 61.765 188.725 ;
        RECT 62.010 188.645 62.330 189.000 ;
        RECT 62.500 189.215 63.040 189.585 ;
        RECT 63.375 189.495 63.780 189.665 ;
        RECT 62.500 188.815 62.740 189.215 ;
        RECT 63.220 189.045 63.440 189.325 ;
        RECT 62.910 188.875 63.440 189.045 ;
        RECT 62.910 188.645 63.080 188.875 ;
        RECT 63.610 188.715 63.780 189.495 ;
        RECT 63.950 188.885 64.300 189.505 ;
        RECT 64.470 188.885 64.680 189.675 ;
        RECT 64.870 189.705 66.370 189.875 ;
        RECT 64.870 189.015 65.040 189.705 ;
        RECT 66.730 189.535 66.900 190.315 ;
        RECT 67.705 190.185 67.875 190.315 ;
        RECT 65.210 189.365 66.900 189.535 ;
        RECT 67.070 189.755 67.535 190.145 ;
        RECT 67.705 190.015 68.100 190.185 ;
        RECT 65.210 189.185 65.380 189.365 ;
        RECT 62.010 188.475 63.080 188.645 ;
        RECT 63.250 188.265 63.440 188.705 ;
        RECT 63.610 188.435 64.560 188.715 ;
        RECT 64.870 188.625 65.130 189.015 ;
        RECT 65.550 188.945 66.340 189.195 ;
        RECT 64.780 188.455 65.130 188.625 ;
        RECT 65.340 188.265 65.670 188.725 ;
        RECT 66.545 188.655 66.715 189.365 ;
        RECT 67.070 189.165 67.240 189.755 ;
        RECT 66.885 188.945 67.240 189.165 ;
        RECT 67.410 188.945 67.760 189.565 ;
        RECT 67.930 188.655 68.100 190.015 ;
        RECT 68.465 189.845 68.790 190.630 ;
        RECT 68.270 188.795 68.730 189.845 ;
        RECT 66.545 188.485 67.400 188.655 ;
        RECT 67.605 188.485 68.100 188.655 ;
        RECT 68.270 188.265 68.600 188.625 ;
        RECT 68.960 188.525 69.130 190.645 ;
        RECT 69.300 190.315 69.630 190.815 ;
        RECT 69.800 190.145 70.055 190.645 ;
        RECT 69.305 189.975 70.055 190.145 ;
        RECT 69.305 188.985 69.535 189.975 ;
        RECT 69.705 189.155 70.055 189.805 ;
        RECT 70.230 189.725 73.740 190.815 ;
        RECT 74.285 189.835 74.540 190.505 ;
        RECT 74.720 190.015 75.005 190.815 ;
        RECT 75.185 190.095 75.515 190.605 ;
        RECT 70.230 189.205 71.920 189.725 ;
        RECT 72.090 189.035 73.740 189.555 ;
        RECT 69.305 188.815 70.055 188.985 ;
        RECT 69.300 188.265 69.630 188.645 ;
        RECT 69.800 188.525 70.055 188.815 ;
        RECT 70.230 188.265 73.740 189.035 ;
        RECT 74.285 188.975 74.465 189.835 ;
        RECT 75.185 189.505 75.435 190.095 ;
        RECT 75.785 189.945 75.955 190.555 ;
        RECT 76.125 190.125 76.455 190.815 ;
        RECT 76.685 190.265 76.925 190.555 ;
        RECT 77.125 190.435 77.545 190.815 ;
        RECT 77.725 190.345 78.355 190.595 ;
        RECT 78.825 190.435 79.155 190.815 ;
        RECT 77.725 190.265 77.895 190.345 ;
        RECT 79.325 190.265 79.495 190.555 ;
        RECT 79.675 190.435 80.055 190.815 ;
        RECT 80.295 190.430 81.125 190.600 ;
        RECT 76.685 190.095 77.895 190.265 ;
        RECT 74.635 189.175 75.435 189.505 ;
        RECT 74.285 188.775 74.540 188.975 ;
        RECT 74.200 188.605 74.540 188.775 ;
        RECT 74.285 188.445 74.540 188.605 ;
        RECT 74.720 188.265 75.005 188.725 ;
        RECT 75.185 188.525 75.435 189.175 ;
        RECT 75.635 189.925 75.955 189.945 ;
        RECT 75.635 189.755 77.555 189.925 ;
        RECT 75.635 188.860 75.825 189.755 ;
        RECT 77.725 189.585 77.895 190.095 ;
        RECT 78.065 189.835 78.585 190.145 ;
        RECT 75.995 189.415 77.895 189.585 ;
        RECT 75.995 189.355 76.325 189.415 ;
        RECT 76.475 189.185 76.805 189.245 ;
        RECT 76.145 188.915 76.805 189.185 ;
        RECT 75.635 188.530 75.955 188.860 ;
        RECT 76.135 188.265 76.795 188.745 ;
        RECT 76.995 188.655 77.165 189.415 ;
        RECT 78.065 189.245 78.245 189.655 ;
        RECT 77.335 189.075 77.665 189.195 ;
        RECT 78.415 189.075 78.585 189.835 ;
        RECT 77.335 188.905 78.585 189.075 ;
        RECT 78.755 190.015 80.125 190.265 ;
        RECT 78.755 189.245 78.945 190.015 ;
        RECT 79.875 189.755 80.125 190.015 ;
        RECT 79.115 189.585 79.365 189.745 ;
        RECT 80.295 189.585 80.465 190.430 ;
        RECT 81.360 190.145 81.530 190.645 ;
        RECT 81.700 190.315 82.030 190.815 ;
        RECT 80.635 189.755 81.135 190.135 ;
        RECT 81.360 189.975 82.055 190.145 ;
        RECT 79.115 189.415 80.465 189.585 ;
        RECT 80.045 189.375 80.465 189.415 ;
        RECT 78.755 188.905 79.175 189.245 ;
        RECT 79.465 188.915 79.875 189.245 ;
        RECT 76.995 188.485 77.845 188.655 ;
        RECT 78.405 188.265 78.725 188.725 ;
        RECT 78.925 188.475 79.175 188.905 ;
        RECT 79.465 188.265 79.875 188.705 ;
        RECT 80.045 188.645 80.215 189.375 ;
        RECT 80.385 188.825 80.735 189.195 ;
        RECT 80.915 188.885 81.135 189.755 ;
        RECT 81.305 189.185 81.715 189.805 ;
        RECT 81.885 189.005 82.055 189.975 ;
        RECT 81.360 188.815 82.055 189.005 ;
        RECT 80.045 188.445 81.060 188.645 ;
        RECT 81.360 188.485 81.530 188.815 ;
        RECT 81.700 188.265 82.030 188.645 ;
        RECT 82.245 188.525 82.470 190.645 ;
        RECT 82.640 190.315 82.970 190.815 ;
        RECT 83.140 190.145 83.310 190.645 ;
        RECT 82.645 189.975 83.310 190.145 ;
        RECT 82.645 188.985 82.875 189.975 ;
        RECT 83.045 189.155 83.395 189.805 ;
        RECT 83.570 189.725 84.780 190.815 ;
        RECT 83.570 189.185 84.090 189.725 ;
        RECT 84.990 189.675 85.220 190.815 ;
        RECT 85.390 189.665 85.720 190.645 ;
        RECT 85.890 189.675 86.100 190.815 ;
        RECT 84.260 189.015 84.780 189.555 ;
        RECT 84.970 189.255 85.300 189.505 ;
        RECT 82.645 188.815 83.310 188.985 ;
        RECT 82.640 188.265 82.970 188.645 ;
        RECT 83.140 188.525 83.310 188.815 ;
        RECT 83.570 188.265 84.780 189.015 ;
        RECT 84.990 188.265 85.220 189.085 ;
        RECT 85.470 189.065 85.720 189.665 ;
        RECT 86.330 189.650 86.620 190.815 ;
        RECT 86.795 190.145 87.050 190.645 ;
        RECT 87.220 190.315 87.550 190.815 ;
        RECT 86.795 189.975 87.545 190.145 ;
        RECT 86.795 189.155 87.145 189.805 ;
        RECT 85.390 188.435 85.720 189.065 ;
        RECT 85.890 188.265 86.100 189.085 ;
        RECT 86.330 188.265 86.620 188.990 ;
        RECT 87.315 188.985 87.545 189.975 ;
        RECT 86.795 188.815 87.545 188.985 ;
        RECT 86.795 188.525 87.050 188.815 ;
        RECT 87.220 188.265 87.550 188.645 ;
        RECT 87.720 188.525 87.890 190.645 ;
        RECT 88.060 189.845 88.385 190.630 ;
        RECT 88.555 190.355 88.805 190.815 ;
        RECT 88.975 190.315 89.225 190.645 ;
        RECT 89.440 190.315 90.120 190.645 ;
        RECT 88.975 190.185 89.145 190.315 ;
        RECT 88.750 190.015 89.145 190.185 ;
        RECT 88.120 188.795 88.580 189.845 ;
        RECT 88.750 188.655 88.920 190.015 ;
        RECT 89.315 189.755 89.780 190.145 ;
        RECT 89.090 188.945 89.440 189.565 ;
        RECT 89.610 189.165 89.780 189.755 ;
        RECT 89.950 189.535 90.120 190.315 ;
        RECT 90.290 190.215 90.460 190.555 ;
        RECT 90.695 190.385 91.025 190.815 ;
        RECT 91.195 190.215 91.365 190.555 ;
        RECT 91.660 190.355 92.030 190.815 ;
        RECT 90.290 190.045 91.365 190.215 ;
        RECT 92.200 190.185 92.370 190.645 ;
        RECT 92.605 190.305 93.475 190.645 ;
        RECT 93.645 190.355 93.895 190.815 ;
        RECT 91.810 190.015 92.370 190.185 ;
        RECT 91.810 189.875 91.980 190.015 ;
        RECT 90.480 189.705 91.980 189.875 ;
        RECT 92.675 189.845 93.135 190.135 ;
        RECT 89.950 189.365 91.640 189.535 ;
        RECT 89.610 188.945 89.965 189.165 ;
        RECT 90.135 188.655 90.305 189.365 ;
        RECT 90.510 188.945 91.300 189.195 ;
        RECT 91.470 189.185 91.640 189.365 ;
        RECT 91.810 189.015 91.980 189.705 ;
        RECT 88.250 188.265 88.580 188.625 ;
        RECT 88.750 188.485 89.245 188.655 ;
        RECT 89.450 188.485 90.305 188.655 ;
        RECT 91.180 188.265 91.510 188.725 ;
        RECT 91.720 188.625 91.980 189.015 ;
        RECT 92.170 189.835 93.135 189.845 ;
        RECT 93.305 189.925 93.475 190.305 ;
        RECT 94.065 190.265 94.235 190.555 ;
        RECT 94.415 190.435 94.745 190.815 ;
        RECT 94.065 190.095 94.865 190.265 ;
        RECT 92.170 189.675 92.845 189.835 ;
        RECT 93.305 189.755 94.525 189.925 ;
        RECT 92.170 188.885 92.380 189.675 ;
        RECT 93.305 189.665 93.475 189.755 ;
        RECT 92.550 188.885 92.900 189.505 ;
        RECT 93.070 189.495 93.475 189.665 ;
        RECT 93.070 188.715 93.240 189.495 ;
        RECT 93.410 189.045 93.630 189.325 ;
        RECT 93.810 189.215 94.350 189.585 ;
        RECT 94.695 189.505 94.865 190.095 ;
        RECT 95.085 189.675 95.390 190.815 ;
        RECT 95.560 189.625 95.815 190.505 ;
        RECT 94.695 189.475 95.435 189.505 ;
        RECT 93.410 188.875 93.940 189.045 ;
        RECT 91.720 188.455 92.070 188.625 ;
        RECT 92.290 188.435 93.240 188.715 ;
        RECT 93.410 188.265 93.600 188.705 ;
        RECT 93.770 188.645 93.940 188.875 ;
        RECT 94.110 188.815 94.350 189.215 ;
        RECT 94.520 189.175 95.435 189.475 ;
        RECT 94.520 189.000 94.845 189.175 ;
        RECT 94.520 188.645 94.840 189.000 ;
        RECT 95.605 188.975 95.815 189.625 ;
        RECT 93.770 188.475 94.840 188.645 ;
        RECT 95.085 188.265 95.390 188.725 ;
        RECT 95.560 188.445 95.815 188.975 ;
        RECT 95.995 189.625 96.250 190.505 ;
        RECT 96.420 189.675 96.725 190.815 ;
        RECT 97.065 190.435 97.395 190.815 ;
        RECT 97.575 190.265 97.745 190.555 ;
        RECT 97.915 190.355 98.165 190.815 ;
        RECT 96.945 190.095 97.745 190.265 ;
        RECT 98.335 190.305 99.205 190.645 ;
        RECT 95.995 188.975 96.205 189.625 ;
        RECT 96.945 189.505 97.115 190.095 ;
        RECT 98.335 189.925 98.505 190.305 ;
        RECT 99.440 190.185 99.610 190.645 ;
        RECT 99.780 190.355 100.150 190.815 ;
        RECT 100.445 190.215 100.615 190.555 ;
        RECT 100.785 190.385 101.115 190.815 ;
        RECT 101.350 190.215 101.520 190.555 ;
        RECT 97.285 189.755 98.505 189.925 ;
        RECT 98.675 189.845 99.135 190.135 ;
        RECT 99.440 190.015 100.000 190.185 ;
        RECT 100.445 190.045 101.520 190.215 ;
        RECT 101.690 190.315 102.370 190.645 ;
        RECT 102.585 190.315 102.835 190.645 ;
        RECT 103.005 190.355 103.255 190.815 ;
        RECT 99.830 189.875 100.000 190.015 ;
        RECT 98.675 189.835 99.640 189.845 ;
        RECT 98.335 189.665 98.505 189.755 ;
        RECT 98.965 189.675 99.640 189.835 ;
        RECT 96.375 189.475 97.115 189.505 ;
        RECT 96.375 189.175 97.290 189.475 ;
        RECT 96.965 189.000 97.290 189.175 ;
        RECT 95.995 188.445 96.250 188.975 ;
        RECT 96.420 188.265 96.725 188.725 ;
        RECT 96.970 188.645 97.290 189.000 ;
        RECT 97.460 189.215 98.000 189.585 ;
        RECT 98.335 189.495 98.740 189.665 ;
        RECT 97.460 188.815 97.700 189.215 ;
        RECT 98.180 189.045 98.400 189.325 ;
        RECT 97.870 188.875 98.400 189.045 ;
        RECT 97.870 188.645 98.040 188.875 ;
        RECT 98.570 188.715 98.740 189.495 ;
        RECT 98.910 188.885 99.260 189.505 ;
        RECT 99.430 188.885 99.640 189.675 ;
        RECT 99.830 189.705 101.330 189.875 ;
        RECT 99.830 189.015 100.000 189.705 ;
        RECT 101.690 189.535 101.860 190.315 ;
        RECT 102.665 190.185 102.835 190.315 ;
        RECT 100.170 189.365 101.860 189.535 ;
        RECT 102.030 189.755 102.495 190.145 ;
        RECT 102.665 190.015 103.060 190.185 ;
        RECT 100.170 189.185 100.340 189.365 ;
        RECT 96.970 188.475 98.040 188.645 ;
        RECT 98.210 188.265 98.400 188.705 ;
        RECT 98.570 188.435 99.520 188.715 ;
        RECT 99.830 188.625 100.090 189.015 ;
        RECT 100.510 188.945 101.300 189.195 ;
        RECT 99.740 188.455 100.090 188.625 ;
        RECT 100.300 188.265 100.630 188.725 ;
        RECT 101.505 188.655 101.675 189.365 ;
        RECT 102.030 189.165 102.200 189.755 ;
        RECT 101.845 188.945 102.200 189.165 ;
        RECT 102.370 188.945 102.720 189.565 ;
        RECT 102.890 188.655 103.060 190.015 ;
        RECT 103.425 189.845 103.750 190.630 ;
        RECT 103.230 188.795 103.690 189.845 ;
        RECT 101.505 188.485 102.360 188.655 ;
        RECT 102.565 188.485 103.060 188.655 ;
        RECT 103.230 188.265 103.560 188.625 ;
        RECT 103.920 188.525 104.090 190.645 ;
        RECT 104.260 190.315 104.590 190.815 ;
        RECT 104.760 190.145 105.015 190.645 ;
        RECT 104.265 189.975 105.015 190.145 ;
        RECT 104.265 188.985 104.495 189.975 ;
        RECT 104.665 189.155 105.015 189.805 ;
        RECT 105.230 189.675 105.460 190.815 ;
        RECT 105.630 189.665 105.960 190.645 ;
        RECT 106.130 189.675 106.340 190.815 ;
        RECT 107.490 189.725 111.000 190.815 ;
        RECT 111.170 189.725 112.380 190.815 ;
        RECT 105.210 189.255 105.540 189.505 ;
        RECT 104.265 188.815 105.015 188.985 ;
        RECT 104.260 188.265 104.590 188.645 ;
        RECT 104.760 188.525 105.015 188.815 ;
        RECT 105.230 188.265 105.460 189.085 ;
        RECT 105.710 189.065 105.960 189.665 ;
        RECT 107.490 189.205 109.180 189.725 ;
        RECT 105.630 188.435 105.960 189.065 ;
        RECT 106.130 188.265 106.340 189.085 ;
        RECT 109.350 189.035 111.000 189.555 ;
        RECT 111.170 189.185 111.690 189.725 ;
        RECT 107.490 188.265 111.000 189.035 ;
        RECT 111.860 189.015 112.380 189.555 ;
        RECT 111.170 188.265 112.380 189.015 ;
        RECT 18.165 188.095 112.465 188.265 ;
        RECT 18.250 187.345 19.460 188.095 ;
        RECT 18.250 186.805 18.770 187.345 ;
        RECT 20.590 187.275 20.820 188.095 ;
        RECT 20.990 187.295 21.320 187.925 ;
        RECT 18.940 186.635 19.460 187.175 ;
        RECT 20.570 186.855 20.900 187.105 ;
        RECT 21.070 186.695 21.320 187.295 ;
        RECT 21.490 187.275 21.700 188.095 ;
        RECT 21.930 187.370 22.220 188.095 ;
        RECT 23.350 187.275 23.580 188.095 ;
        RECT 23.750 187.295 24.080 187.925 ;
        RECT 23.330 186.855 23.660 187.105 ;
        RECT 18.250 185.545 19.460 186.635 ;
        RECT 20.590 185.545 20.820 186.685 ;
        RECT 20.990 185.715 21.320 186.695 ;
        RECT 21.490 185.545 21.700 186.685 ;
        RECT 21.930 185.545 22.220 186.710 ;
        RECT 23.830 186.695 24.080 187.295 ;
        RECT 24.250 187.275 24.460 188.095 ;
        RECT 24.965 187.285 25.210 187.890 ;
        RECT 25.430 187.560 25.940 188.095 ;
        RECT 23.350 185.545 23.580 186.685 ;
        RECT 23.750 185.715 24.080 186.695 ;
        RECT 24.690 187.115 25.920 187.285 ;
        RECT 24.250 185.545 24.460 186.685 ;
        RECT 24.690 186.305 25.030 187.115 ;
        RECT 25.200 186.550 25.950 186.740 ;
        RECT 24.690 185.895 25.205 186.305 ;
        RECT 25.440 185.545 25.610 186.305 ;
        RECT 25.780 185.885 25.950 186.550 ;
        RECT 26.120 186.565 26.310 187.925 ;
        RECT 26.480 187.755 26.755 187.925 ;
        RECT 26.480 187.585 26.760 187.755 ;
        RECT 26.480 186.765 26.755 187.585 ;
        RECT 26.945 187.560 27.475 187.925 ;
        RECT 27.900 187.695 28.230 188.095 ;
        RECT 27.300 187.525 27.475 187.560 ;
        RECT 26.960 186.565 27.130 187.365 ;
        RECT 26.120 186.395 27.130 186.565 ;
        RECT 27.300 187.355 28.230 187.525 ;
        RECT 28.400 187.355 28.655 187.925 ;
        RECT 27.300 186.225 27.470 187.355 ;
        RECT 28.060 187.185 28.230 187.355 ;
        RECT 26.345 186.055 27.470 186.225 ;
        RECT 27.640 186.855 27.835 187.185 ;
        RECT 28.060 186.855 28.315 187.185 ;
        RECT 27.640 185.885 27.810 186.855 ;
        RECT 28.485 186.685 28.655 187.355 ;
        RECT 25.780 185.715 27.810 185.885 ;
        RECT 27.980 185.545 28.150 186.685 ;
        RECT 28.320 185.715 28.655 186.685 ;
        RECT 28.835 187.385 29.090 187.915 ;
        RECT 29.260 187.635 29.565 188.095 ;
        RECT 29.810 187.715 30.880 187.885 ;
        RECT 28.835 186.735 29.045 187.385 ;
        RECT 29.810 187.360 30.130 187.715 ;
        RECT 29.805 187.185 30.130 187.360 ;
        RECT 29.215 186.885 30.130 187.185 ;
        RECT 30.300 187.145 30.540 187.545 ;
        RECT 30.710 187.485 30.880 187.715 ;
        RECT 31.050 187.655 31.240 188.095 ;
        RECT 31.410 187.645 32.360 187.925 ;
        RECT 32.580 187.735 32.930 187.905 ;
        RECT 30.710 187.315 31.240 187.485 ;
        RECT 29.215 186.855 29.955 186.885 ;
        RECT 28.835 185.855 29.090 186.735 ;
        RECT 29.260 185.545 29.565 186.685 ;
        RECT 29.785 186.265 29.955 186.855 ;
        RECT 30.300 186.775 30.840 187.145 ;
        RECT 31.020 187.035 31.240 187.315 ;
        RECT 31.410 186.865 31.580 187.645 ;
        RECT 31.175 186.695 31.580 186.865 ;
        RECT 31.750 186.855 32.100 187.475 ;
        RECT 31.175 186.605 31.345 186.695 ;
        RECT 32.270 186.685 32.480 187.475 ;
        RECT 30.125 186.435 31.345 186.605 ;
        RECT 31.805 186.525 32.480 186.685 ;
        RECT 29.785 186.095 30.585 186.265 ;
        RECT 29.905 185.545 30.235 185.925 ;
        RECT 30.415 185.805 30.585 186.095 ;
        RECT 31.175 186.055 31.345 186.435 ;
        RECT 31.515 186.515 32.480 186.525 ;
        RECT 32.670 187.345 32.930 187.735 ;
        RECT 33.140 187.635 33.470 188.095 ;
        RECT 34.345 187.705 35.200 187.875 ;
        RECT 35.405 187.705 35.900 187.875 ;
        RECT 36.070 187.735 36.400 188.095 ;
        RECT 32.670 186.655 32.840 187.345 ;
        RECT 33.010 186.995 33.180 187.175 ;
        RECT 33.350 187.165 34.140 187.415 ;
        RECT 34.345 186.995 34.515 187.705 ;
        RECT 34.685 187.195 35.040 187.415 ;
        RECT 33.010 186.825 34.700 186.995 ;
        RECT 31.515 186.225 31.975 186.515 ;
        RECT 32.670 186.485 34.170 186.655 ;
        RECT 32.670 186.345 32.840 186.485 ;
        RECT 32.280 186.175 32.840 186.345 ;
        RECT 30.755 185.545 31.005 186.005 ;
        RECT 31.175 185.715 32.045 186.055 ;
        RECT 32.280 185.715 32.450 186.175 ;
        RECT 33.285 186.145 34.360 186.315 ;
        RECT 32.620 185.545 32.990 186.005 ;
        RECT 33.285 185.805 33.455 186.145 ;
        RECT 33.625 185.545 33.955 185.975 ;
        RECT 34.190 185.805 34.360 186.145 ;
        RECT 34.530 186.045 34.700 186.825 ;
        RECT 34.870 186.605 35.040 187.195 ;
        RECT 35.210 186.795 35.560 187.415 ;
        RECT 34.870 186.215 35.335 186.605 ;
        RECT 35.730 186.345 35.900 187.705 ;
        RECT 36.070 186.515 36.530 187.565 ;
        RECT 35.505 186.175 35.900 186.345 ;
        RECT 35.505 186.045 35.675 186.175 ;
        RECT 34.530 185.715 35.210 186.045 ;
        RECT 35.425 185.715 35.675 186.045 ;
        RECT 35.845 185.545 36.095 186.005 ;
        RECT 36.265 185.730 36.590 186.515 ;
        RECT 36.760 185.715 36.930 187.835 ;
        RECT 37.100 187.715 37.430 188.095 ;
        RECT 37.600 187.545 37.855 187.835 ;
        RECT 37.105 187.375 37.855 187.545 ;
        RECT 38.405 187.385 38.660 187.915 ;
        RECT 38.840 187.635 39.125 188.095 ;
        RECT 37.105 186.385 37.335 187.375 ;
        RECT 37.505 186.555 37.855 187.205 ;
        RECT 38.405 186.525 38.585 187.385 ;
        RECT 39.305 187.185 39.555 187.835 ;
        RECT 38.755 186.855 39.555 187.185 ;
        RECT 37.105 186.215 37.855 186.385 ;
        RECT 37.100 185.545 37.430 186.045 ;
        RECT 37.600 185.715 37.855 186.215 ;
        RECT 38.405 186.055 38.660 186.525 ;
        RECT 38.320 185.885 38.660 186.055 ;
        RECT 38.405 185.855 38.660 185.885 ;
        RECT 38.840 185.545 39.125 186.345 ;
        RECT 39.305 186.265 39.555 186.855 ;
        RECT 39.755 187.500 40.075 187.830 ;
        RECT 40.255 187.615 40.915 188.095 ;
        RECT 41.115 187.705 41.965 187.875 ;
        RECT 39.755 186.605 39.945 187.500 ;
        RECT 40.265 187.175 40.925 187.445 ;
        RECT 40.595 187.115 40.925 187.175 ;
        RECT 40.115 186.945 40.445 187.005 ;
        RECT 41.115 186.945 41.285 187.705 ;
        RECT 42.525 187.635 42.845 188.095 ;
        RECT 43.045 187.455 43.295 187.885 ;
        RECT 43.585 187.655 43.995 188.095 ;
        RECT 44.165 187.715 45.180 187.915 ;
        RECT 41.455 187.285 42.705 187.455 ;
        RECT 41.455 187.165 41.785 187.285 ;
        RECT 40.115 186.775 42.015 186.945 ;
        RECT 39.755 186.435 41.675 186.605 ;
        RECT 39.755 186.415 40.075 186.435 ;
        RECT 39.305 185.755 39.635 186.265 ;
        RECT 39.905 185.805 40.075 186.415 ;
        RECT 41.845 186.265 42.015 186.775 ;
        RECT 42.185 186.705 42.365 187.115 ;
        RECT 42.535 186.525 42.705 187.285 ;
        RECT 40.245 185.545 40.575 186.235 ;
        RECT 40.805 186.095 42.015 186.265 ;
        RECT 42.185 186.215 42.705 186.525 ;
        RECT 42.875 187.115 43.295 187.455 ;
        RECT 43.585 187.115 43.995 187.445 ;
        RECT 42.875 186.345 43.065 187.115 ;
        RECT 44.165 186.985 44.335 187.715 ;
        RECT 45.480 187.545 45.650 187.875 ;
        RECT 45.820 187.715 46.150 188.095 ;
        RECT 44.505 187.165 44.855 187.535 ;
        RECT 44.165 186.945 44.585 186.985 ;
        RECT 43.235 186.775 44.585 186.945 ;
        RECT 43.235 186.615 43.485 186.775 ;
        RECT 43.995 186.345 44.245 186.605 ;
        RECT 42.875 186.095 44.245 186.345 ;
        RECT 40.805 185.805 41.045 186.095 ;
        RECT 41.845 186.015 42.015 186.095 ;
        RECT 41.245 185.545 41.665 185.925 ;
        RECT 41.845 185.765 42.475 186.015 ;
        RECT 42.945 185.545 43.275 185.925 ;
        RECT 43.445 185.805 43.615 186.095 ;
        RECT 44.415 185.930 44.585 186.775 ;
        RECT 45.035 186.605 45.255 187.475 ;
        RECT 45.480 187.355 46.175 187.545 ;
        RECT 44.755 186.225 45.255 186.605 ;
        RECT 45.425 186.555 45.835 187.175 ;
        RECT 46.005 186.385 46.175 187.355 ;
        RECT 45.480 186.215 46.175 186.385 ;
        RECT 43.795 185.545 44.175 185.925 ;
        RECT 44.415 185.760 45.245 185.930 ;
        RECT 45.480 185.715 45.650 186.215 ;
        RECT 45.820 185.545 46.150 186.045 ;
        RECT 46.365 185.715 46.590 187.835 ;
        RECT 46.760 187.715 47.090 188.095 ;
        RECT 47.260 187.545 47.430 187.835 ;
        RECT 46.765 187.375 47.430 187.545 ;
        RECT 46.765 186.385 46.995 187.375 ;
        RECT 47.690 187.370 47.980 188.095 ;
        RECT 48.670 187.275 48.880 188.095 ;
        RECT 49.050 187.295 49.380 187.925 ;
        RECT 47.165 186.555 47.515 187.205 ;
        RECT 46.765 186.215 47.430 186.385 ;
        RECT 46.760 185.545 47.090 186.045 ;
        RECT 47.260 185.715 47.430 186.215 ;
        RECT 47.690 185.545 47.980 186.710 ;
        RECT 49.050 186.695 49.300 187.295 ;
        RECT 49.550 187.275 49.780 188.095 ;
        RECT 49.990 187.355 50.310 187.835 ;
        RECT 50.480 187.525 50.710 187.925 ;
        RECT 50.880 187.705 51.230 188.095 ;
        RECT 50.480 187.445 50.990 187.525 ;
        RECT 51.400 187.445 51.730 187.925 ;
        RECT 50.480 187.355 51.730 187.445 ;
        RECT 49.470 186.855 49.800 187.105 ;
        RECT 48.670 185.545 48.880 186.685 ;
        RECT 49.050 185.715 49.380 186.695 ;
        RECT 49.550 185.545 49.780 186.685 ;
        RECT 49.990 186.425 50.160 187.355 ;
        RECT 50.820 187.275 51.730 187.355 ;
        RECT 51.900 187.275 52.070 188.095 ;
        RECT 52.575 187.355 53.040 187.900 ;
        RECT 50.330 186.765 50.500 187.185 ;
        RECT 50.730 186.935 51.330 187.105 ;
        RECT 50.330 186.595 50.990 186.765 ;
        RECT 49.990 186.225 50.650 186.425 ;
        RECT 50.820 186.395 50.990 186.595 ;
        RECT 51.160 186.735 51.330 186.935 ;
        RECT 51.500 186.905 52.195 187.105 ;
        RECT 52.455 186.735 52.700 187.185 ;
        RECT 51.160 186.565 52.700 186.735 ;
        RECT 52.870 186.395 53.040 187.355 ;
        RECT 50.820 186.225 53.040 186.395 ;
        RECT 53.210 187.355 53.595 187.925 ;
        RECT 53.765 187.635 54.090 188.095 ;
        RECT 54.610 187.465 54.890 187.925 ;
        RECT 53.210 186.685 53.490 187.355 ;
        RECT 53.765 187.295 54.890 187.465 ;
        RECT 53.765 187.185 54.215 187.295 ;
        RECT 53.660 186.855 54.215 187.185 ;
        RECT 55.080 187.125 55.480 187.925 ;
        RECT 55.880 187.635 56.150 188.095 ;
        RECT 56.320 187.465 56.605 187.925 ;
        RECT 50.480 186.055 50.650 186.225 ;
        RECT 50.010 185.545 50.310 186.055 ;
        RECT 50.480 185.885 50.860 186.055 ;
        RECT 51.440 185.545 52.070 186.055 ;
        RECT 52.240 185.715 52.570 186.225 ;
        RECT 52.740 185.545 53.040 186.055 ;
        RECT 53.210 185.715 53.595 186.685 ;
        RECT 53.765 186.395 54.215 186.855 ;
        RECT 54.385 186.565 55.480 187.125 ;
        RECT 53.765 186.175 54.890 186.395 ;
        RECT 53.765 185.545 54.090 186.005 ;
        RECT 54.610 185.715 54.890 186.175 ;
        RECT 55.080 185.715 55.480 186.565 ;
        RECT 55.650 187.295 56.605 187.465 ;
        RECT 56.890 187.345 58.100 188.095 ;
        RECT 55.650 186.395 55.860 187.295 ;
        RECT 56.030 186.565 56.720 187.125 ;
        RECT 56.890 186.635 57.410 187.175 ;
        RECT 57.580 186.805 58.100 187.345 ;
        RECT 58.270 187.275 58.530 188.095 ;
        RECT 58.700 187.275 59.030 187.695 ;
        RECT 59.210 187.525 59.470 187.925 ;
        RECT 59.640 187.695 59.970 188.095 ;
        RECT 60.140 187.525 60.310 187.875 ;
        RECT 60.480 187.695 60.855 188.095 ;
        RECT 59.210 187.355 60.875 187.525 ;
        RECT 61.045 187.420 61.320 187.765 ;
        RECT 58.780 187.185 59.030 187.275 ;
        RECT 60.705 187.185 60.875 187.355 ;
        RECT 58.275 186.855 58.610 187.105 ;
        RECT 58.780 186.855 59.495 187.185 ;
        RECT 59.710 186.855 60.535 187.185 ;
        RECT 60.705 186.855 60.980 187.185 ;
        RECT 55.650 186.175 56.605 186.395 ;
        RECT 55.880 185.545 56.150 186.005 ;
        RECT 56.320 185.715 56.605 186.175 ;
        RECT 56.890 185.545 58.100 186.635 ;
        RECT 58.270 185.545 58.530 186.685 ;
        RECT 58.780 186.295 58.950 186.855 ;
        RECT 59.210 186.395 59.540 186.685 ;
        RECT 59.710 186.565 59.955 186.855 ;
        RECT 60.705 186.685 60.875 186.855 ;
        RECT 61.150 186.685 61.320 187.420 ;
        RECT 61.580 187.545 61.750 187.925 ;
        RECT 61.930 187.715 62.260 188.095 ;
        RECT 61.580 187.375 62.245 187.545 ;
        RECT 62.440 187.420 62.700 187.925 ;
        RECT 61.510 186.825 61.840 187.195 ;
        RECT 62.075 187.120 62.245 187.375 ;
        RECT 60.215 186.515 60.875 186.685 ;
        RECT 60.215 186.395 60.385 186.515 ;
        RECT 59.210 186.225 60.385 186.395 ;
        RECT 58.770 185.725 60.385 186.055 ;
        RECT 60.555 185.545 60.835 186.345 ;
        RECT 61.045 185.715 61.320 186.685 ;
        RECT 62.075 186.790 62.360 187.120 ;
        RECT 62.075 186.645 62.245 186.790 ;
        RECT 61.580 186.475 62.245 186.645 ;
        RECT 62.530 186.620 62.700 187.420 ;
        RECT 61.580 185.715 61.750 186.475 ;
        RECT 61.930 185.545 62.260 186.305 ;
        RECT 62.430 185.715 62.700 186.620 ;
        RECT 62.875 187.385 63.130 187.915 ;
        RECT 63.300 187.635 63.605 188.095 ;
        RECT 63.850 187.715 64.920 187.885 ;
        RECT 62.875 186.735 63.085 187.385 ;
        RECT 63.850 187.360 64.170 187.715 ;
        RECT 63.845 187.185 64.170 187.360 ;
        RECT 63.255 186.885 64.170 187.185 ;
        RECT 64.340 187.145 64.580 187.545 ;
        RECT 64.750 187.485 64.920 187.715 ;
        RECT 65.090 187.655 65.280 188.095 ;
        RECT 65.450 187.645 66.400 187.925 ;
        RECT 66.620 187.735 66.970 187.905 ;
        RECT 64.750 187.315 65.280 187.485 ;
        RECT 63.255 186.855 63.995 186.885 ;
        RECT 62.875 185.855 63.130 186.735 ;
        RECT 63.300 185.545 63.605 186.685 ;
        RECT 63.825 186.265 63.995 186.855 ;
        RECT 64.340 186.775 64.880 187.145 ;
        RECT 65.060 187.035 65.280 187.315 ;
        RECT 65.450 186.865 65.620 187.645 ;
        RECT 65.215 186.695 65.620 186.865 ;
        RECT 65.790 186.855 66.140 187.475 ;
        RECT 65.215 186.605 65.385 186.695 ;
        RECT 66.310 186.685 66.520 187.475 ;
        RECT 64.165 186.435 65.385 186.605 ;
        RECT 65.845 186.525 66.520 186.685 ;
        RECT 63.825 186.095 64.625 186.265 ;
        RECT 63.945 185.545 64.275 185.925 ;
        RECT 64.455 185.805 64.625 186.095 ;
        RECT 65.215 186.055 65.385 186.435 ;
        RECT 65.555 186.515 66.520 186.525 ;
        RECT 66.710 187.345 66.970 187.735 ;
        RECT 67.180 187.635 67.510 188.095 ;
        RECT 68.385 187.705 69.240 187.875 ;
        RECT 69.445 187.705 69.940 187.875 ;
        RECT 70.110 187.735 70.440 188.095 ;
        RECT 66.710 186.655 66.880 187.345 ;
        RECT 67.050 186.995 67.220 187.175 ;
        RECT 67.390 187.165 68.180 187.415 ;
        RECT 68.385 186.995 68.555 187.705 ;
        RECT 68.725 187.195 69.080 187.415 ;
        RECT 67.050 186.825 68.740 186.995 ;
        RECT 65.555 186.225 66.015 186.515 ;
        RECT 66.710 186.485 68.210 186.655 ;
        RECT 66.710 186.345 66.880 186.485 ;
        RECT 66.320 186.175 66.880 186.345 ;
        RECT 64.795 185.545 65.045 186.005 ;
        RECT 65.215 185.715 66.085 186.055 ;
        RECT 66.320 185.715 66.490 186.175 ;
        RECT 67.325 186.145 68.400 186.315 ;
        RECT 66.660 185.545 67.030 186.005 ;
        RECT 67.325 185.805 67.495 186.145 ;
        RECT 67.665 185.545 67.995 185.975 ;
        RECT 68.230 185.805 68.400 186.145 ;
        RECT 68.570 186.045 68.740 186.825 ;
        RECT 68.910 186.605 69.080 187.195 ;
        RECT 69.250 186.795 69.600 187.415 ;
        RECT 68.910 186.215 69.375 186.605 ;
        RECT 69.770 186.345 69.940 187.705 ;
        RECT 70.110 186.515 70.570 187.565 ;
        RECT 69.545 186.175 69.940 186.345 ;
        RECT 69.545 186.045 69.715 186.175 ;
        RECT 68.570 185.715 69.250 186.045 ;
        RECT 69.465 185.715 69.715 186.045 ;
        RECT 69.885 185.545 70.135 186.005 ;
        RECT 70.305 185.730 70.630 186.515 ;
        RECT 70.800 185.715 70.970 187.835 ;
        RECT 71.140 187.715 71.470 188.095 ;
        RECT 71.640 187.545 71.895 187.835 ;
        RECT 71.145 187.375 71.895 187.545 ;
        RECT 71.145 186.385 71.375 187.375 ;
        RECT 72.130 187.275 72.340 188.095 ;
        RECT 72.510 187.295 72.840 187.925 ;
        RECT 71.545 186.555 71.895 187.205 ;
        RECT 72.510 186.695 72.760 187.295 ;
        RECT 73.010 187.275 73.240 188.095 ;
        RECT 73.450 187.370 73.740 188.095 ;
        RECT 74.745 187.385 75.000 187.915 ;
        RECT 75.180 187.635 75.465 188.095 ;
        RECT 72.930 186.855 73.260 187.105 ;
        RECT 71.145 186.215 71.895 186.385 ;
        RECT 71.140 185.545 71.470 186.045 ;
        RECT 71.640 185.715 71.895 186.215 ;
        RECT 72.130 185.545 72.340 186.685 ;
        RECT 72.510 185.715 72.840 186.695 ;
        RECT 73.010 185.545 73.240 186.685 ;
        RECT 73.450 185.545 73.740 186.710 ;
        RECT 74.745 186.525 74.925 187.385 ;
        RECT 75.645 187.185 75.895 187.835 ;
        RECT 75.095 186.855 75.895 187.185 ;
        RECT 74.745 186.055 75.000 186.525 ;
        RECT 74.660 185.885 75.000 186.055 ;
        RECT 74.745 185.855 75.000 185.885 ;
        RECT 75.180 185.545 75.465 186.345 ;
        RECT 75.645 186.265 75.895 186.855 ;
        RECT 76.095 187.500 76.415 187.830 ;
        RECT 76.595 187.615 77.255 188.095 ;
        RECT 77.455 187.705 78.305 187.875 ;
        RECT 76.095 186.605 76.285 187.500 ;
        RECT 76.605 187.175 77.265 187.445 ;
        RECT 76.935 187.115 77.265 187.175 ;
        RECT 76.455 186.945 76.785 187.005 ;
        RECT 77.455 186.945 77.625 187.705 ;
        RECT 78.865 187.635 79.185 188.095 ;
        RECT 79.385 187.455 79.635 187.885 ;
        RECT 79.925 187.655 80.335 188.095 ;
        RECT 80.505 187.715 81.520 187.915 ;
        RECT 77.795 187.285 79.045 187.455 ;
        RECT 77.795 187.165 78.125 187.285 ;
        RECT 76.455 186.775 78.355 186.945 ;
        RECT 76.095 186.435 78.015 186.605 ;
        RECT 76.095 186.415 76.415 186.435 ;
        RECT 75.645 185.755 75.975 186.265 ;
        RECT 76.245 185.805 76.415 186.415 ;
        RECT 78.185 186.265 78.355 186.775 ;
        RECT 78.525 186.705 78.705 187.115 ;
        RECT 78.875 186.525 79.045 187.285 ;
        RECT 76.585 185.545 76.915 186.235 ;
        RECT 77.145 186.095 78.355 186.265 ;
        RECT 78.525 186.215 79.045 186.525 ;
        RECT 79.215 187.115 79.635 187.455 ;
        RECT 79.925 187.115 80.335 187.445 ;
        RECT 79.215 186.345 79.405 187.115 ;
        RECT 80.505 186.985 80.675 187.715 ;
        RECT 81.820 187.545 81.990 187.875 ;
        RECT 82.160 187.715 82.490 188.095 ;
        RECT 80.845 187.165 81.195 187.535 ;
        RECT 80.505 186.945 80.925 186.985 ;
        RECT 79.575 186.775 80.925 186.945 ;
        RECT 79.575 186.615 79.825 186.775 ;
        RECT 80.335 186.345 80.585 186.605 ;
        RECT 79.215 186.095 80.585 186.345 ;
        RECT 77.145 185.805 77.385 186.095 ;
        RECT 78.185 186.015 78.355 186.095 ;
        RECT 77.585 185.545 78.005 185.925 ;
        RECT 78.185 185.765 78.815 186.015 ;
        RECT 79.285 185.545 79.615 185.925 ;
        RECT 79.785 185.805 79.955 186.095 ;
        RECT 80.755 185.930 80.925 186.775 ;
        RECT 81.375 186.605 81.595 187.475 ;
        RECT 81.820 187.355 82.515 187.545 ;
        RECT 81.095 186.225 81.595 186.605 ;
        RECT 81.765 186.555 82.175 187.175 ;
        RECT 82.345 186.385 82.515 187.355 ;
        RECT 81.820 186.215 82.515 186.385 ;
        RECT 80.135 185.545 80.515 185.925 ;
        RECT 80.755 185.760 81.585 185.930 ;
        RECT 81.820 185.715 81.990 186.215 ;
        RECT 82.160 185.545 82.490 186.045 ;
        RECT 82.705 185.715 82.930 187.835 ;
        RECT 83.100 187.715 83.430 188.095 ;
        RECT 83.600 187.545 83.770 187.835 ;
        RECT 83.105 187.375 83.770 187.545 ;
        RECT 83.105 186.385 83.335 187.375 ;
        RECT 84.305 187.285 84.550 187.890 ;
        RECT 84.770 187.560 85.280 188.095 ;
        RECT 83.505 186.555 83.855 187.205 ;
        RECT 84.030 187.115 85.260 187.285 ;
        RECT 83.105 186.215 83.770 186.385 ;
        RECT 83.100 185.545 83.430 186.045 ;
        RECT 83.600 185.715 83.770 186.215 ;
        RECT 84.030 186.305 84.370 187.115 ;
        RECT 84.540 186.550 85.290 186.740 ;
        RECT 84.030 185.895 84.545 186.305 ;
        RECT 84.780 185.545 84.950 186.305 ;
        RECT 85.120 185.885 85.290 186.550 ;
        RECT 85.460 186.565 85.650 187.925 ;
        RECT 85.820 187.415 86.095 187.925 ;
        RECT 86.285 187.560 86.815 187.925 ;
        RECT 87.240 187.695 87.570 188.095 ;
        RECT 86.640 187.525 86.815 187.560 ;
        RECT 85.820 187.245 86.100 187.415 ;
        RECT 85.820 186.765 86.095 187.245 ;
        RECT 86.300 186.565 86.470 187.365 ;
        RECT 85.460 186.395 86.470 186.565 ;
        RECT 86.640 187.355 87.570 187.525 ;
        RECT 87.740 187.355 87.995 187.925 ;
        RECT 86.640 186.225 86.810 187.355 ;
        RECT 87.400 187.185 87.570 187.355 ;
        RECT 85.685 186.055 86.810 186.225 ;
        RECT 86.980 186.855 87.175 187.185 ;
        RECT 87.400 186.855 87.655 187.185 ;
        RECT 86.980 185.885 87.150 186.855 ;
        RECT 87.825 186.685 87.995 187.355 ;
        RECT 88.170 187.345 89.380 188.095 ;
        RECT 85.120 185.715 87.150 185.885 ;
        RECT 87.320 185.545 87.490 186.685 ;
        RECT 87.660 185.715 87.995 186.685 ;
        RECT 88.170 186.635 88.690 187.175 ;
        RECT 88.860 186.805 89.380 187.345 ;
        RECT 89.610 187.275 89.820 188.095 ;
        RECT 89.990 187.295 90.320 187.925 ;
        RECT 89.990 186.695 90.240 187.295 ;
        RECT 90.490 187.275 90.720 188.095 ;
        RECT 91.390 187.325 93.060 188.095 ;
        RECT 93.320 187.545 93.490 187.925 ;
        RECT 93.670 187.715 94.000 188.095 ;
        RECT 93.320 187.375 93.985 187.545 ;
        RECT 94.180 187.420 94.440 187.925 ;
        RECT 90.410 186.855 90.740 187.105 ;
        RECT 88.170 185.545 89.380 186.635 ;
        RECT 89.610 185.545 89.820 186.685 ;
        RECT 89.990 185.715 90.320 186.695 ;
        RECT 90.490 185.545 90.720 186.685 ;
        RECT 91.390 186.635 92.140 187.155 ;
        RECT 92.310 186.805 93.060 187.325 ;
        RECT 93.250 186.825 93.580 187.195 ;
        RECT 93.815 187.120 93.985 187.375 ;
        RECT 93.815 186.790 94.100 187.120 ;
        RECT 93.815 186.645 93.985 186.790 ;
        RECT 91.390 185.545 93.060 186.635 ;
        RECT 93.320 186.475 93.985 186.645 ;
        RECT 94.270 186.620 94.440 187.420 ;
        RECT 95.345 187.285 95.590 187.890 ;
        RECT 95.810 187.560 96.320 188.095 ;
        RECT 93.320 185.715 93.490 186.475 ;
        RECT 93.670 185.545 94.000 186.305 ;
        RECT 94.170 185.715 94.440 186.620 ;
        RECT 95.070 187.115 96.300 187.285 ;
        RECT 95.070 186.305 95.410 187.115 ;
        RECT 95.580 186.550 96.330 186.740 ;
        RECT 95.070 185.895 95.585 186.305 ;
        RECT 95.820 185.545 95.990 186.305 ;
        RECT 96.160 185.885 96.330 186.550 ;
        RECT 96.500 186.565 96.690 187.925 ;
        RECT 96.860 187.415 97.135 187.925 ;
        RECT 97.325 187.560 97.855 187.925 ;
        RECT 98.280 187.695 98.610 188.095 ;
        RECT 97.680 187.525 97.855 187.560 ;
        RECT 96.860 187.245 97.140 187.415 ;
        RECT 96.860 186.765 97.135 187.245 ;
        RECT 97.340 186.565 97.510 187.365 ;
        RECT 96.500 186.395 97.510 186.565 ;
        RECT 97.680 187.355 98.610 187.525 ;
        RECT 98.780 187.355 99.035 187.925 ;
        RECT 99.210 187.370 99.500 188.095 ;
        RECT 97.680 186.225 97.850 187.355 ;
        RECT 98.440 187.185 98.610 187.355 ;
        RECT 96.725 186.055 97.850 186.225 ;
        RECT 98.020 186.855 98.215 187.185 ;
        RECT 98.440 186.855 98.695 187.185 ;
        RECT 98.020 185.885 98.190 186.855 ;
        RECT 98.865 186.685 99.035 187.355 ;
        RECT 99.945 187.285 100.190 187.890 ;
        RECT 100.410 187.560 100.920 188.095 ;
        RECT 99.670 187.115 100.900 187.285 ;
        RECT 96.160 185.715 98.190 185.885 ;
        RECT 98.360 185.545 98.530 186.685 ;
        RECT 98.700 185.715 99.035 186.685 ;
        RECT 99.210 185.545 99.500 186.710 ;
        RECT 99.670 186.305 100.010 187.115 ;
        RECT 100.180 186.550 100.930 186.740 ;
        RECT 99.670 185.895 100.185 186.305 ;
        RECT 100.420 185.545 100.590 186.305 ;
        RECT 100.760 185.885 100.930 186.550 ;
        RECT 101.100 186.565 101.290 187.925 ;
        RECT 101.460 187.075 101.735 187.925 ;
        RECT 101.925 187.560 102.455 187.925 ;
        RECT 102.880 187.695 103.210 188.095 ;
        RECT 102.280 187.525 102.455 187.560 ;
        RECT 101.460 186.905 101.740 187.075 ;
        RECT 101.460 186.765 101.735 186.905 ;
        RECT 101.940 186.565 102.110 187.365 ;
        RECT 101.100 186.395 102.110 186.565 ;
        RECT 102.280 187.355 103.210 187.525 ;
        RECT 103.380 187.355 103.635 187.925 ;
        RECT 102.280 186.225 102.450 187.355 ;
        RECT 103.040 187.185 103.210 187.355 ;
        RECT 101.325 186.055 102.450 186.225 ;
        RECT 102.620 186.855 102.815 187.185 ;
        RECT 103.040 186.855 103.295 187.185 ;
        RECT 102.620 185.885 102.790 186.855 ;
        RECT 103.465 186.685 103.635 187.355 ;
        RECT 104.270 187.325 105.940 188.095 ;
        RECT 106.200 187.545 106.370 187.925 ;
        RECT 106.550 187.715 106.880 188.095 ;
        RECT 106.200 187.375 106.865 187.545 ;
        RECT 107.060 187.420 107.320 187.925 ;
        RECT 100.760 185.715 102.790 185.885 ;
        RECT 102.960 185.545 103.130 186.685 ;
        RECT 103.300 185.715 103.635 186.685 ;
        RECT 104.270 186.635 105.020 187.155 ;
        RECT 105.190 186.805 105.940 187.325 ;
        RECT 106.130 186.825 106.460 187.195 ;
        RECT 106.695 187.120 106.865 187.375 ;
        RECT 106.695 186.790 106.980 187.120 ;
        RECT 106.695 186.645 106.865 186.790 ;
        RECT 104.270 185.545 105.940 186.635 ;
        RECT 106.200 186.475 106.865 186.645 ;
        RECT 107.150 186.620 107.320 187.420 ;
        RECT 107.490 187.325 111.000 188.095 ;
        RECT 111.170 187.345 112.380 188.095 ;
        RECT 106.200 185.715 106.370 186.475 ;
        RECT 106.550 185.545 106.880 186.305 ;
        RECT 107.050 185.715 107.320 186.620 ;
        RECT 107.490 186.635 109.180 187.155 ;
        RECT 109.350 186.805 111.000 187.325 ;
        RECT 111.170 186.635 111.690 187.175 ;
        RECT 111.860 186.805 112.380 187.345 ;
        RECT 107.490 185.545 111.000 186.635 ;
        RECT 111.170 185.545 112.380 186.635 ;
        RECT 18.165 185.375 112.465 185.545 ;
        RECT 18.250 184.285 19.460 185.375 ;
        RECT 18.250 183.575 18.770 184.115 ;
        RECT 18.940 183.745 19.460 184.285 ;
        RECT 19.690 184.235 19.900 185.375 ;
        RECT 20.070 184.225 20.400 185.205 ;
        RECT 20.570 184.235 20.800 185.375 ;
        RECT 21.015 184.705 21.270 185.205 ;
        RECT 21.440 184.875 21.770 185.375 ;
        RECT 21.015 184.535 21.765 184.705 ;
        RECT 18.250 182.825 19.460 183.575 ;
        RECT 19.690 182.825 19.900 183.645 ;
        RECT 20.070 183.625 20.320 184.225 ;
        RECT 20.490 183.815 20.820 184.065 ;
        RECT 21.015 183.715 21.365 184.365 ;
        RECT 20.070 182.995 20.400 183.625 ;
        RECT 20.570 182.825 20.800 183.645 ;
        RECT 21.535 183.545 21.765 184.535 ;
        RECT 21.015 183.375 21.765 183.545 ;
        RECT 21.015 183.085 21.270 183.375 ;
        RECT 21.440 182.825 21.770 183.205 ;
        RECT 21.940 183.085 22.110 185.205 ;
        RECT 22.280 184.405 22.605 185.190 ;
        RECT 22.775 184.915 23.025 185.375 ;
        RECT 23.195 184.875 23.445 185.205 ;
        RECT 23.660 184.875 24.340 185.205 ;
        RECT 23.195 184.745 23.365 184.875 ;
        RECT 22.970 184.575 23.365 184.745 ;
        RECT 22.340 183.355 22.800 184.405 ;
        RECT 22.970 183.215 23.140 184.575 ;
        RECT 23.535 184.315 24.000 184.705 ;
        RECT 23.310 183.505 23.660 184.125 ;
        RECT 23.830 183.725 24.000 184.315 ;
        RECT 24.170 184.095 24.340 184.875 ;
        RECT 24.510 184.775 24.680 185.115 ;
        RECT 24.915 184.945 25.245 185.375 ;
        RECT 25.415 184.775 25.585 185.115 ;
        RECT 25.880 184.915 26.250 185.375 ;
        RECT 24.510 184.605 25.585 184.775 ;
        RECT 26.420 184.745 26.590 185.205 ;
        RECT 26.825 184.865 27.695 185.205 ;
        RECT 27.865 184.915 28.115 185.375 ;
        RECT 26.030 184.575 26.590 184.745 ;
        RECT 26.030 184.435 26.200 184.575 ;
        RECT 24.700 184.265 26.200 184.435 ;
        RECT 26.895 184.405 27.355 184.695 ;
        RECT 24.170 183.925 25.860 184.095 ;
        RECT 23.830 183.505 24.185 183.725 ;
        RECT 24.355 183.215 24.525 183.925 ;
        RECT 24.730 183.505 25.520 183.755 ;
        RECT 25.690 183.745 25.860 183.925 ;
        RECT 26.030 183.575 26.200 184.265 ;
        RECT 22.470 182.825 22.800 183.185 ;
        RECT 22.970 183.045 23.465 183.215 ;
        RECT 23.670 183.045 24.525 183.215 ;
        RECT 25.400 182.825 25.730 183.285 ;
        RECT 25.940 183.185 26.200 183.575 ;
        RECT 26.390 184.395 27.355 184.405 ;
        RECT 27.525 184.485 27.695 184.865 ;
        RECT 28.285 184.825 28.455 185.115 ;
        RECT 28.635 184.995 28.965 185.375 ;
        RECT 28.285 184.655 29.085 184.825 ;
        RECT 26.390 184.235 27.065 184.395 ;
        RECT 27.525 184.315 28.745 184.485 ;
        RECT 26.390 183.445 26.600 184.235 ;
        RECT 27.525 184.225 27.695 184.315 ;
        RECT 26.770 183.445 27.120 184.065 ;
        RECT 27.290 184.055 27.695 184.225 ;
        RECT 27.290 183.275 27.460 184.055 ;
        RECT 27.630 183.605 27.850 183.885 ;
        RECT 28.030 183.775 28.570 184.145 ;
        RECT 28.915 184.065 29.085 184.655 ;
        RECT 29.305 184.235 29.610 185.375 ;
        RECT 29.780 184.185 30.035 185.065 ;
        RECT 28.915 184.035 29.655 184.065 ;
        RECT 27.630 183.435 28.160 183.605 ;
        RECT 25.940 183.015 26.290 183.185 ;
        RECT 26.510 182.995 27.460 183.275 ;
        RECT 27.630 182.825 27.820 183.265 ;
        RECT 27.990 183.205 28.160 183.435 ;
        RECT 28.330 183.375 28.570 183.775 ;
        RECT 28.740 183.735 29.655 184.035 ;
        RECT 28.740 183.560 29.065 183.735 ;
        RECT 28.740 183.205 29.060 183.560 ;
        RECT 29.825 183.535 30.035 184.185 ;
        RECT 30.670 184.615 31.185 185.025 ;
        RECT 31.420 184.615 31.590 185.375 ;
        RECT 31.760 185.035 33.790 185.205 ;
        RECT 30.670 183.805 31.010 184.615 ;
        RECT 31.760 184.370 31.930 185.035 ;
        RECT 32.325 184.695 33.450 184.865 ;
        RECT 31.180 184.180 31.930 184.370 ;
        RECT 32.100 184.355 33.110 184.525 ;
        RECT 30.670 183.635 31.900 183.805 ;
        RECT 27.990 183.035 29.060 183.205 ;
        RECT 29.305 182.825 29.610 183.285 ;
        RECT 29.780 183.005 30.035 183.535 ;
        RECT 30.945 183.030 31.190 183.635 ;
        RECT 31.410 182.825 31.920 183.360 ;
        RECT 32.100 182.995 32.290 184.355 ;
        RECT 32.460 183.675 32.735 184.155 ;
        RECT 32.460 183.505 32.740 183.675 ;
        RECT 32.940 183.555 33.110 184.355 ;
        RECT 33.280 183.565 33.450 184.695 ;
        RECT 33.620 184.065 33.790 185.035 ;
        RECT 33.960 184.235 34.130 185.375 ;
        RECT 34.300 184.235 34.635 185.205 ;
        RECT 33.620 183.735 33.815 184.065 ;
        RECT 34.040 183.735 34.295 184.065 ;
        RECT 34.040 183.565 34.210 183.735 ;
        RECT 34.465 183.565 34.635 184.235 ;
        RECT 34.810 184.210 35.100 185.375 ;
        RECT 35.820 184.445 35.990 185.205 ;
        RECT 36.170 184.615 36.500 185.375 ;
        RECT 35.820 184.275 36.485 184.445 ;
        RECT 36.670 184.300 36.940 185.205 ;
        RECT 36.315 184.130 36.485 184.275 ;
        RECT 35.750 183.725 36.080 184.095 ;
        RECT 36.315 183.800 36.600 184.130 ;
        RECT 32.460 182.995 32.735 183.505 ;
        RECT 33.280 183.395 34.210 183.565 ;
        RECT 33.280 183.360 33.455 183.395 ;
        RECT 32.925 182.995 33.455 183.360 ;
        RECT 33.880 182.825 34.210 183.225 ;
        RECT 34.380 182.995 34.635 183.565 ;
        RECT 34.810 182.825 35.100 183.550 ;
        RECT 36.315 183.545 36.485 183.800 ;
        RECT 35.820 183.375 36.485 183.545 ;
        RECT 36.770 183.500 36.940 184.300 ;
        RECT 37.610 184.235 37.840 185.375 ;
        RECT 38.010 184.225 38.340 185.205 ;
        RECT 38.510 184.235 38.720 185.375 ;
        RECT 38.950 184.615 39.465 185.025 ;
        RECT 39.700 184.615 39.870 185.375 ;
        RECT 40.040 185.035 42.070 185.205 ;
        RECT 37.590 183.815 37.920 184.065 ;
        RECT 35.820 182.995 35.990 183.375 ;
        RECT 36.170 182.825 36.500 183.205 ;
        RECT 36.680 182.995 36.940 183.500 ;
        RECT 37.610 182.825 37.840 183.645 ;
        RECT 38.090 183.625 38.340 184.225 ;
        RECT 38.950 183.805 39.290 184.615 ;
        RECT 40.040 184.370 40.210 185.035 ;
        RECT 40.605 184.695 41.730 184.865 ;
        RECT 39.460 184.180 40.210 184.370 ;
        RECT 40.380 184.355 41.390 184.525 ;
        RECT 38.010 182.995 38.340 183.625 ;
        RECT 38.510 182.825 38.720 183.645 ;
        RECT 38.950 183.635 40.180 183.805 ;
        RECT 39.225 183.030 39.470 183.635 ;
        RECT 39.690 182.825 40.200 183.360 ;
        RECT 40.380 182.995 40.570 184.355 ;
        RECT 40.740 184.015 41.015 184.155 ;
        RECT 40.740 183.845 41.020 184.015 ;
        RECT 40.740 182.995 41.015 183.845 ;
        RECT 41.220 183.555 41.390 184.355 ;
        RECT 41.560 183.565 41.730 184.695 ;
        RECT 41.900 184.065 42.070 185.035 ;
        RECT 42.240 184.235 42.410 185.375 ;
        RECT 42.580 184.235 42.915 185.205 ;
        RECT 41.900 183.735 42.095 184.065 ;
        RECT 42.320 183.735 42.575 184.065 ;
        RECT 42.320 183.565 42.490 183.735 ;
        RECT 42.745 183.565 42.915 184.235 ;
        RECT 43.090 184.615 43.605 185.025 ;
        RECT 43.840 184.615 44.010 185.375 ;
        RECT 44.180 185.035 46.210 185.205 ;
        RECT 43.090 183.805 43.430 184.615 ;
        RECT 44.180 184.370 44.350 185.035 ;
        RECT 44.745 184.695 45.870 184.865 ;
        RECT 43.600 184.180 44.350 184.370 ;
        RECT 44.520 184.355 45.530 184.525 ;
        RECT 43.090 183.635 44.320 183.805 ;
        RECT 41.560 183.395 42.490 183.565 ;
        RECT 41.560 183.360 41.735 183.395 ;
        RECT 41.205 182.995 41.735 183.360 ;
        RECT 42.160 182.825 42.490 183.225 ;
        RECT 42.660 182.995 42.915 183.565 ;
        RECT 43.365 183.030 43.610 183.635 ;
        RECT 43.830 182.825 44.340 183.360 ;
        RECT 44.520 182.995 44.710 184.355 ;
        RECT 44.880 183.335 45.155 184.155 ;
        RECT 45.360 183.555 45.530 184.355 ;
        RECT 45.700 183.565 45.870 184.695 ;
        RECT 46.040 184.065 46.210 185.035 ;
        RECT 46.380 184.235 46.550 185.375 ;
        RECT 46.720 184.235 47.055 185.205 ;
        RECT 48.460 184.535 48.630 185.375 ;
        RECT 48.840 184.365 49.090 185.205 ;
        RECT 49.300 184.535 49.470 185.375 ;
        RECT 49.640 184.365 49.930 185.205 ;
        RECT 46.040 183.735 46.235 184.065 ;
        RECT 46.460 183.735 46.715 184.065 ;
        RECT 46.460 183.565 46.630 183.735 ;
        RECT 46.885 183.565 47.055 184.235 ;
        RECT 45.700 183.395 46.630 183.565 ;
        RECT 45.700 183.360 45.875 183.395 ;
        RECT 44.880 183.165 45.160 183.335 ;
        RECT 44.880 182.995 45.155 183.165 ;
        RECT 45.345 182.995 45.875 183.360 ;
        RECT 46.300 182.825 46.630 183.225 ;
        RECT 46.800 182.995 47.055 183.565 ;
        RECT 48.205 184.195 49.930 184.365 ;
        RECT 50.140 184.315 50.310 185.375 ;
        RECT 50.605 184.995 50.935 185.375 ;
        RECT 51.115 184.825 51.285 185.115 ;
        RECT 51.455 184.915 51.705 185.375 ;
        RECT 50.485 184.655 51.285 184.825 ;
        RECT 51.875 184.865 52.745 185.205 ;
        RECT 48.205 183.645 48.615 184.195 ;
        RECT 50.485 184.035 50.655 184.655 ;
        RECT 51.875 184.485 52.045 184.865 ;
        RECT 52.980 184.745 53.150 185.205 ;
        RECT 53.320 184.915 53.690 185.375 ;
        RECT 53.985 184.775 54.155 185.115 ;
        RECT 54.325 184.945 54.655 185.375 ;
        RECT 54.890 184.775 55.060 185.115 ;
        RECT 50.825 184.315 52.045 184.485 ;
        RECT 52.215 184.405 52.675 184.695 ;
        RECT 52.980 184.575 53.540 184.745 ;
        RECT 53.985 184.605 55.060 184.775 ;
        RECT 55.230 184.875 55.910 185.205 ;
        RECT 56.125 184.875 56.375 185.205 ;
        RECT 56.545 184.915 56.795 185.375 ;
        RECT 53.370 184.435 53.540 184.575 ;
        RECT 52.215 184.395 53.180 184.405 ;
        RECT 51.875 184.225 52.045 184.315 ;
        RECT 52.505 184.235 53.180 184.395 ;
        RECT 50.485 184.025 50.830 184.035 ;
        RECT 48.800 183.815 50.830 184.025 ;
        RECT 48.205 183.475 49.970 183.645 ;
        RECT 48.460 182.825 48.630 183.295 ;
        RECT 48.800 182.995 49.130 183.475 ;
        RECT 49.300 182.825 49.470 183.295 ;
        RECT 49.640 182.995 49.970 183.475 ;
        RECT 50.140 182.825 50.310 183.635 ;
        RECT 50.505 183.560 50.830 183.815 ;
        RECT 50.510 183.205 50.830 183.560 ;
        RECT 51.000 183.775 51.540 184.145 ;
        RECT 51.875 184.055 52.280 184.225 ;
        RECT 51.000 183.375 51.240 183.775 ;
        RECT 51.720 183.605 51.940 183.885 ;
        RECT 51.410 183.435 51.940 183.605 ;
        RECT 51.410 183.205 51.580 183.435 ;
        RECT 52.110 183.275 52.280 184.055 ;
        RECT 52.450 183.445 52.800 184.065 ;
        RECT 52.970 183.445 53.180 184.235 ;
        RECT 53.370 184.265 54.870 184.435 ;
        RECT 53.370 183.575 53.540 184.265 ;
        RECT 55.230 184.095 55.400 184.875 ;
        RECT 56.205 184.745 56.375 184.875 ;
        RECT 53.710 183.925 55.400 184.095 ;
        RECT 55.570 184.315 56.035 184.705 ;
        RECT 56.205 184.575 56.600 184.745 ;
        RECT 53.710 183.745 53.880 183.925 ;
        RECT 50.510 183.035 51.580 183.205 ;
        RECT 51.750 182.825 51.940 183.265 ;
        RECT 52.110 182.995 53.060 183.275 ;
        RECT 53.370 183.185 53.630 183.575 ;
        RECT 54.050 183.505 54.840 183.755 ;
        RECT 53.280 183.015 53.630 183.185 ;
        RECT 53.840 182.825 54.170 183.285 ;
        RECT 55.045 183.215 55.215 183.925 ;
        RECT 55.570 183.725 55.740 184.315 ;
        RECT 55.385 183.505 55.740 183.725 ;
        RECT 55.910 183.505 56.260 184.125 ;
        RECT 56.430 183.215 56.600 184.575 ;
        RECT 56.965 184.405 57.290 185.190 ;
        RECT 56.770 183.355 57.230 184.405 ;
        RECT 55.045 183.045 55.900 183.215 ;
        RECT 56.105 183.045 56.600 183.215 ;
        RECT 56.770 182.825 57.100 183.185 ;
        RECT 57.460 183.085 57.630 185.205 ;
        RECT 57.800 184.875 58.130 185.375 ;
        RECT 58.300 184.705 58.555 185.205 ;
        RECT 57.805 184.535 58.555 184.705 ;
        RECT 57.805 183.545 58.035 184.535 ;
        RECT 58.205 183.715 58.555 184.365 ;
        RECT 58.730 184.300 59.000 185.205 ;
        RECT 59.170 184.615 59.500 185.375 ;
        RECT 59.680 184.445 59.850 185.205 ;
        RECT 57.805 183.375 58.555 183.545 ;
        RECT 57.800 182.825 58.130 183.205 ;
        RECT 58.300 183.085 58.555 183.375 ;
        RECT 58.730 183.500 58.900 184.300 ;
        RECT 59.185 184.275 59.850 184.445 ;
        RECT 59.185 184.130 59.355 184.275 ;
        RECT 60.570 184.210 60.860 185.375 ;
        RECT 61.030 184.235 61.305 185.205 ;
        RECT 61.515 184.575 61.795 185.375 ;
        RECT 61.965 184.865 63.580 185.195 ;
        RECT 61.965 184.525 63.140 184.695 ;
        RECT 61.965 184.405 62.135 184.525 ;
        RECT 61.475 184.235 62.135 184.405 ;
        RECT 59.070 183.800 59.355 184.130 ;
        RECT 59.185 183.545 59.355 183.800 ;
        RECT 59.590 183.725 59.920 184.095 ;
        RECT 58.730 182.995 58.990 183.500 ;
        RECT 59.185 183.375 59.850 183.545 ;
        RECT 59.170 182.825 59.500 183.205 ;
        RECT 59.680 182.995 59.850 183.375 ;
        RECT 60.570 182.825 60.860 183.550 ;
        RECT 61.030 183.500 61.200 184.235 ;
        RECT 61.475 184.065 61.645 184.235 ;
        RECT 62.395 184.065 62.640 184.355 ;
        RECT 62.810 184.235 63.140 184.525 ;
        RECT 63.400 184.065 63.570 184.625 ;
        RECT 63.820 184.235 64.080 185.375 ;
        RECT 64.270 184.575 64.550 185.375 ;
        RECT 64.750 184.405 65.080 185.205 ;
        RECT 65.280 184.575 65.450 185.375 ;
        RECT 65.620 184.405 65.950 185.205 ;
        RECT 61.370 183.735 61.645 184.065 ;
        RECT 61.815 183.735 62.640 184.065 ;
        RECT 62.855 183.735 63.570 184.065 ;
        RECT 63.740 183.815 64.075 184.065 ;
        RECT 64.250 183.735 64.490 184.405 ;
        RECT 64.670 184.235 65.950 184.405 ;
        RECT 66.120 184.235 66.380 185.375 ;
        RECT 66.585 184.585 67.120 185.205 ;
        RECT 61.475 183.565 61.645 183.735 ;
        RECT 63.320 183.645 63.570 183.735 ;
        RECT 61.030 183.155 61.305 183.500 ;
        RECT 61.475 183.395 63.140 183.565 ;
        RECT 61.495 182.825 61.870 183.225 ;
        RECT 62.040 183.045 62.210 183.395 ;
        RECT 62.380 182.825 62.710 183.225 ;
        RECT 62.880 182.995 63.140 183.395 ;
        RECT 63.320 183.225 63.650 183.645 ;
        RECT 63.820 182.825 64.080 183.645 ;
        RECT 64.670 183.565 64.840 184.235 ;
        RECT 65.010 183.735 65.320 184.065 ;
        RECT 65.490 183.735 65.870 184.065 ;
        RECT 66.070 183.735 66.355 184.065 ;
        RECT 65.115 183.565 65.320 183.735 ;
        RECT 64.250 182.995 64.945 183.565 ;
        RECT 65.115 183.040 65.465 183.565 ;
        RECT 65.655 183.040 65.870 183.735 ;
        RECT 66.585 183.565 66.900 184.585 ;
        RECT 67.290 184.575 67.620 185.375 ;
        RECT 68.850 184.865 69.150 185.375 ;
        RECT 69.320 184.695 69.650 185.205 ;
        RECT 69.820 184.865 70.450 185.375 ;
        RECT 71.030 184.865 71.410 185.035 ;
        RECT 71.580 184.865 71.880 185.375 ;
        RECT 71.240 184.695 71.410 184.865 ;
        RECT 68.105 184.405 68.495 184.580 ;
        RECT 67.070 184.235 68.495 184.405 ;
        RECT 68.850 184.525 71.070 184.695 ;
        RECT 67.070 183.735 67.240 184.235 ;
        RECT 66.040 182.825 66.375 183.565 ;
        RECT 66.585 182.995 67.200 183.565 ;
        RECT 67.490 183.505 67.755 184.065 ;
        RECT 67.925 183.335 68.095 184.235 ;
        RECT 68.265 183.505 68.620 184.065 ;
        RECT 68.850 183.565 69.020 184.525 ;
        RECT 69.190 184.185 70.730 184.355 ;
        RECT 69.190 183.735 69.435 184.185 ;
        RECT 69.695 183.815 70.390 184.015 ;
        RECT 70.560 183.985 70.730 184.185 ;
        RECT 70.900 184.325 71.070 184.525 ;
        RECT 71.240 184.495 71.900 184.695 ;
        RECT 70.900 184.155 71.560 184.325 ;
        RECT 70.560 183.815 71.160 183.985 ;
        RECT 71.390 183.735 71.560 184.155 ;
        RECT 67.370 182.825 67.585 183.335 ;
        RECT 67.815 183.005 68.095 183.335 ;
        RECT 68.275 182.825 68.515 183.335 ;
        RECT 68.850 183.020 69.315 183.565 ;
        RECT 69.820 182.825 69.990 183.645 ;
        RECT 70.160 183.565 71.070 183.645 ;
        RECT 71.730 183.565 71.900 184.495 ;
        RECT 72.070 184.235 72.330 185.375 ;
        RECT 72.500 184.225 72.830 185.205 ;
        RECT 73.000 184.235 73.280 185.375 ;
        RECT 74.410 184.235 74.640 185.375 ;
        RECT 74.810 184.225 75.140 185.205 ;
        RECT 75.310 184.235 75.520 185.375 ;
        RECT 75.750 184.615 76.265 185.025 ;
        RECT 76.500 184.615 76.670 185.375 ;
        RECT 76.840 185.035 78.870 185.205 ;
        RECT 72.090 183.815 72.425 184.065 ;
        RECT 72.595 183.625 72.765 184.225 ;
        RECT 72.935 183.795 73.270 184.065 ;
        RECT 74.390 183.815 74.720 184.065 ;
        RECT 70.160 183.475 71.410 183.565 ;
        RECT 70.160 182.995 70.490 183.475 ;
        RECT 70.900 183.395 71.410 183.475 ;
        RECT 70.660 182.825 71.010 183.215 ;
        RECT 71.180 182.995 71.410 183.395 ;
        RECT 71.580 183.085 71.900 183.565 ;
        RECT 72.070 182.995 72.765 183.625 ;
        RECT 72.970 182.825 73.280 183.625 ;
        RECT 74.410 182.825 74.640 183.645 ;
        RECT 74.890 183.625 75.140 184.225 ;
        RECT 75.750 183.805 76.090 184.615 ;
        RECT 76.840 184.370 77.010 185.035 ;
        RECT 77.405 184.695 78.530 184.865 ;
        RECT 76.260 184.180 77.010 184.370 ;
        RECT 77.180 184.355 78.190 184.525 ;
        RECT 74.810 182.995 75.140 183.625 ;
        RECT 75.310 182.825 75.520 183.645 ;
        RECT 75.750 183.635 76.980 183.805 ;
        RECT 76.025 183.030 76.270 183.635 ;
        RECT 76.490 182.825 77.000 183.360 ;
        RECT 77.180 182.995 77.370 184.355 ;
        RECT 77.540 183.335 77.815 184.155 ;
        RECT 78.020 183.555 78.190 184.355 ;
        RECT 78.360 183.565 78.530 184.695 ;
        RECT 78.700 184.065 78.870 185.035 ;
        RECT 79.040 184.235 79.210 185.375 ;
        RECT 79.380 184.235 79.715 185.205 ;
        RECT 80.440 184.445 80.610 185.205 ;
        RECT 80.790 184.615 81.120 185.375 ;
        RECT 80.440 184.275 81.105 184.445 ;
        RECT 81.290 184.300 81.560 185.205 ;
        RECT 78.700 183.735 78.895 184.065 ;
        RECT 79.120 183.735 79.375 184.065 ;
        RECT 79.120 183.565 79.290 183.735 ;
        RECT 79.545 183.565 79.715 184.235 ;
        RECT 80.935 184.130 81.105 184.275 ;
        RECT 80.370 183.725 80.700 184.095 ;
        RECT 80.935 183.800 81.220 184.130 ;
        RECT 78.360 183.395 79.290 183.565 ;
        RECT 78.360 183.360 78.535 183.395 ;
        RECT 77.540 183.165 77.820 183.335 ;
        RECT 77.540 182.995 77.815 183.165 ;
        RECT 78.005 182.995 78.535 183.360 ;
        RECT 78.960 182.825 79.290 183.225 ;
        RECT 79.460 182.995 79.715 183.565 ;
        RECT 80.935 183.545 81.105 183.800 ;
        RECT 80.440 183.375 81.105 183.545 ;
        RECT 81.390 183.500 81.560 184.300 ;
        RECT 80.440 182.995 80.610 183.375 ;
        RECT 80.790 182.825 81.120 183.205 ;
        RECT 81.300 182.995 81.560 183.500 ;
        RECT 81.730 184.300 82.000 185.205 ;
        RECT 82.170 184.615 82.500 185.375 ;
        RECT 82.680 184.445 82.850 185.205 ;
        RECT 81.730 183.500 81.900 184.300 ;
        RECT 82.185 184.275 82.850 184.445 ;
        RECT 83.570 184.285 86.160 185.375 ;
        RECT 82.185 184.130 82.355 184.275 ;
        RECT 82.070 183.800 82.355 184.130 ;
        RECT 82.185 183.545 82.355 183.800 ;
        RECT 82.590 183.725 82.920 184.095 ;
        RECT 83.570 183.765 84.780 184.285 ;
        RECT 86.330 184.210 86.620 185.375 ;
        RECT 86.795 184.185 87.050 185.065 ;
        RECT 87.220 184.235 87.525 185.375 ;
        RECT 87.865 184.995 88.195 185.375 ;
        RECT 88.375 184.825 88.545 185.115 ;
        RECT 88.715 184.915 88.965 185.375 ;
        RECT 87.745 184.655 88.545 184.825 ;
        RECT 89.135 184.865 90.005 185.205 ;
        RECT 84.950 183.595 86.160 184.115 ;
        RECT 81.730 182.995 81.990 183.500 ;
        RECT 82.185 183.375 82.850 183.545 ;
        RECT 82.170 182.825 82.500 183.205 ;
        RECT 82.680 182.995 82.850 183.375 ;
        RECT 83.570 182.825 86.160 183.595 ;
        RECT 86.330 182.825 86.620 183.550 ;
        RECT 86.795 183.535 87.005 184.185 ;
        RECT 87.745 184.065 87.915 184.655 ;
        RECT 89.135 184.485 89.305 184.865 ;
        RECT 90.240 184.745 90.410 185.205 ;
        RECT 90.580 184.915 90.950 185.375 ;
        RECT 91.245 184.775 91.415 185.115 ;
        RECT 91.585 184.945 91.915 185.375 ;
        RECT 92.150 184.775 92.320 185.115 ;
        RECT 88.085 184.315 89.305 184.485 ;
        RECT 89.475 184.405 89.935 184.695 ;
        RECT 90.240 184.575 90.800 184.745 ;
        RECT 91.245 184.605 92.320 184.775 ;
        RECT 92.490 184.875 93.170 185.205 ;
        RECT 93.385 184.875 93.635 185.205 ;
        RECT 93.805 184.915 94.055 185.375 ;
        RECT 90.630 184.435 90.800 184.575 ;
        RECT 89.475 184.395 90.440 184.405 ;
        RECT 89.135 184.225 89.305 184.315 ;
        RECT 89.765 184.235 90.440 184.395 ;
        RECT 87.175 184.035 87.915 184.065 ;
        RECT 87.175 183.735 88.090 184.035 ;
        RECT 87.765 183.560 88.090 183.735 ;
        RECT 86.795 183.005 87.050 183.535 ;
        RECT 87.220 182.825 87.525 183.285 ;
        RECT 87.770 183.205 88.090 183.560 ;
        RECT 88.260 183.775 88.800 184.145 ;
        RECT 89.135 184.055 89.540 184.225 ;
        RECT 88.260 183.375 88.500 183.775 ;
        RECT 88.980 183.605 89.200 183.885 ;
        RECT 88.670 183.435 89.200 183.605 ;
        RECT 88.670 183.205 88.840 183.435 ;
        RECT 89.370 183.275 89.540 184.055 ;
        RECT 89.710 183.445 90.060 184.065 ;
        RECT 90.230 183.445 90.440 184.235 ;
        RECT 90.630 184.265 92.130 184.435 ;
        RECT 90.630 183.575 90.800 184.265 ;
        RECT 92.490 184.095 92.660 184.875 ;
        RECT 93.465 184.745 93.635 184.875 ;
        RECT 90.970 183.925 92.660 184.095 ;
        RECT 92.830 184.315 93.295 184.705 ;
        RECT 93.465 184.575 93.860 184.745 ;
        RECT 90.970 183.745 91.140 183.925 ;
        RECT 87.770 183.035 88.840 183.205 ;
        RECT 89.010 182.825 89.200 183.265 ;
        RECT 89.370 182.995 90.320 183.275 ;
        RECT 90.630 183.185 90.890 183.575 ;
        RECT 91.310 183.505 92.100 183.755 ;
        RECT 90.540 183.015 90.890 183.185 ;
        RECT 91.100 182.825 91.430 183.285 ;
        RECT 92.305 183.215 92.475 183.925 ;
        RECT 92.830 183.725 93.000 184.315 ;
        RECT 92.645 183.505 93.000 183.725 ;
        RECT 93.170 183.505 93.520 184.125 ;
        RECT 93.690 183.215 93.860 184.575 ;
        RECT 94.225 184.405 94.550 185.190 ;
        RECT 94.030 183.355 94.490 184.405 ;
        RECT 92.305 183.045 93.160 183.215 ;
        RECT 93.365 183.045 93.860 183.215 ;
        RECT 94.030 182.825 94.360 183.185 ;
        RECT 94.720 183.085 94.890 185.205 ;
        RECT 95.060 184.875 95.390 185.375 ;
        RECT 95.560 184.705 95.815 185.205 ;
        RECT 95.065 184.535 95.815 184.705 ;
        RECT 95.990 184.615 96.505 185.025 ;
        RECT 96.740 184.615 96.910 185.375 ;
        RECT 97.080 185.035 99.110 185.205 ;
        RECT 95.065 183.545 95.295 184.535 ;
        RECT 95.465 183.715 95.815 184.365 ;
        RECT 95.990 183.805 96.330 184.615 ;
        RECT 97.080 184.370 97.250 185.035 ;
        RECT 97.645 184.695 98.770 184.865 ;
        RECT 96.500 184.180 97.250 184.370 ;
        RECT 97.420 184.355 98.430 184.525 ;
        RECT 95.990 183.635 97.220 183.805 ;
        RECT 95.065 183.375 95.815 183.545 ;
        RECT 95.060 182.825 95.390 183.205 ;
        RECT 95.560 183.085 95.815 183.375 ;
        RECT 96.265 183.030 96.510 183.635 ;
        RECT 96.730 182.825 97.240 183.360 ;
        RECT 97.420 182.995 97.610 184.355 ;
        RECT 97.780 183.675 98.055 184.155 ;
        RECT 97.780 183.505 98.060 183.675 ;
        RECT 98.260 183.555 98.430 184.355 ;
        RECT 98.600 183.565 98.770 184.695 ;
        RECT 98.940 184.065 99.110 185.035 ;
        RECT 99.280 184.235 99.450 185.375 ;
        RECT 99.620 184.235 99.955 185.205 ;
        RECT 98.940 183.735 99.135 184.065 ;
        RECT 99.360 183.735 99.615 184.065 ;
        RECT 99.360 183.565 99.530 183.735 ;
        RECT 99.785 183.565 99.955 184.235 ;
        RECT 100.130 184.615 100.645 185.025 ;
        RECT 100.880 184.615 101.050 185.375 ;
        RECT 101.220 185.035 103.250 185.205 ;
        RECT 100.130 183.805 100.470 184.615 ;
        RECT 101.220 184.370 101.390 185.035 ;
        RECT 101.785 184.695 102.910 184.865 ;
        RECT 100.640 184.180 101.390 184.370 ;
        RECT 101.560 184.355 102.570 184.525 ;
        RECT 100.130 183.635 101.360 183.805 ;
        RECT 97.780 182.995 98.055 183.505 ;
        RECT 98.600 183.395 99.530 183.565 ;
        RECT 98.600 183.360 98.775 183.395 ;
        RECT 98.245 182.995 98.775 183.360 ;
        RECT 99.200 182.825 99.530 183.225 ;
        RECT 99.700 182.995 99.955 183.565 ;
        RECT 100.405 183.030 100.650 183.635 ;
        RECT 100.870 182.825 101.380 183.360 ;
        RECT 101.560 182.995 101.750 184.355 ;
        RECT 101.920 184.015 102.195 184.155 ;
        RECT 101.920 183.845 102.200 184.015 ;
        RECT 101.920 182.995 102.195 183.845 ;
        RECT 102.400 183.555 102.570 184.355 ;
        RECT 102.740 183.565 102.910 184.695 ;
        RECT 103.080 184.065 103.250 185.035 ;
        RECT 103.420 184.235 103.590 185.375 ;
        RECT 103.760 184.235 104.095 185.205 ;
        RECT 104.330 184.235 104.540 185.375 ;
        RECT 103.080 183.735 103.275 184.065 ;
        RECT 103.500 183.735 103.755 184.065 ;
        RECT 103.500 183.565 103.670 183.735 ;
        RECT 103.925 183.565 104.095 184.235 ;
        RECT 104.710 184.225 105.040 185.205 ;
        RECT 105.210 184.235 105.440 185.375 ;
        RECT 106.200 184.445 106.370 185.205 ;
        RECT 106.550 184.615 106.880 185.375 ;
        RECT 106.200 184.275 106.865 184.445 ;
        RECT 107.050 184.300 107.320 185.205 ;
        RECT 102.740 183.395 103.670 183.565 ;
        RECT 102.740 183.360 102.915 183.395 ;
        RECT 102.385 182.995 102.915 183.360 ;
        RECT 103.340 182.825 103.670 183.225 ;
        RECT 103.840 182.995 104.095 183.565 ;
        RECT 104.330 182.825 104.540 183.645 ;
        RECT 104.710 183.625 104.960 184.225 ;
        RECT 106.695 184.130 106.865 184.275 ;
        RECT 105.130 183.815 105.460 184.065 ;
        RECT 106.130 183.725 106.460 184.095 ;
        RECT 106.695 183.800 106.980 184.130 ;
        RECT 104.710 182.995 105.040 183.625 ;
        RECT 105.210 182.825 105.440 183.645 ;
        RECT 106.695 183.545 106.865 183.800 ;
        RECT 106.200 183.375 106.865 183.545 ;
        RECT 107.150 183.500 107.320 184.300 ;
        RECT 107.490 184.285 111.000 185.375 ;
        RECT 111.170 184.285 112.380 185.375 ;
        RECT 107.490 183.765 109.180 184.285 ;
        RECT 109.350 183.595 111.000 184.115 ;
        RECT 111.170 183.745 111.690 184.285 ;
        RECT 106.200 182.995 106.370 183.375 ;
        RECT 106.550 182.825 106.880 183.205 ;
        RECT 107.060 182.995 107.320 183.500 ;
        RECT 107.490 182.825 111.000 183.595 ;
        RECT 111.860 183.575 112.380 184.115 ;
        RECT 111.170 182.825 112.380 183.575 ;
        RECT 18.165 182.655 112.465 182.825 ;
        RECT 18.250 181.905 19.460 182.655 ;
        RECT 20.640 182.105 20.810 182.485 ;
        RECT 20.990 182.275 21.320 182.655 ;
        RECT 20.640 181.935 21.305 182.105 ;
        RECT 21.500 181.980 21.760 182.485 ;
        RECT 18.250 181.365 18.770 181.905 ;
        RECT 18.940 181.195 19.460 181.735 ;
        RECT 20.570 181.385 20.900 181.755 ;
        RECT 21.135 181.680 21.305 181.935 ;
        RECT 21.135 181.350 21.420 181.680 ;
        RECT 21.135 181.205 21.305 181.350 ;
        RECT 18.250 180.105 19.460 181.195 ;
        RECT 20.640 181.035 21.305 181.205 ;
        RECT 21.590 181.180 21.760 181.980 ;
        RECT 21.930 181.930 22.220 182.655 ;
        RECT 22.505 182.025 22.790 182.485 ;
        RECT 22.960 182.195 23.230 182.655 ;
        RECT 22.505 181.855 23.460 182.025 ;
        RECT 20.640 180.275 20.810 181.035 ;
        RECT 20.990 180.105 21.320 180.865 ;
        RECT 21.490 180.275 21.760 181.180 ;
        RECT 21.930 180.105 22.220 181.270 ;
        RECT 22.390 181.125 23.080 181.685 ;
        RECT 23.250 180.955 23.460 181.855 ;
        RECT 22.505 180.735 23.460 180.955 ;
        RECT 23.630 181.685 24.030 182.485 ;
        RECT 24.220 182.025 24.500 182.485 ;
        RECT 25.020 182.195 25.345 182.655 ;
        RECT 24.220 181.855 25.345 182.025 ;
        RECT 25.515 181.915 25.900 182.485 ;
        RECT 24.895 181.745 25.345 181.855 ;
        RECT 23.630 181.125 24.725 181.685 ;
        RECT 24.895 181.415 25.450 181.745 ;
        RECT 22.505 180.275 22.790 180.735 ;
        RECT 22.960 180.105 23.230 180.565 ;
        RECT 23.630 180.275 24.030 181.125 ;
        RECT 24.895 180.955 25.345 181.415 ;
        RECT 25.620 181.245 25.900 181.915 ;
        RECT 24.220 180.735 25.345 180.955 ;
        RECT 24.220 180.275 24.500 180.735 ;
        RECT 25.020 180.105 25.345 180.565 ;
        RECT 25.515 180.275 25.900 181.245 ;
        RECT 26.995 181.915 27.250 182.485 ;
        RECT 27.420 182.255 27.750 182.655 ;
        RECT 28.175 182.120 28.705 182.485 ;
        RECT 28.175 182.085 28.350 182.120 ;
        RECT 27.420 181.915 28.350 182.085 ;
        RECT 26.995 181.245 27.165 181.915 ;
        RECT 27.420 181.745 27.590 181.915 ;
        RECT 27.335 181.415 27.590 181.745 ;
        RECT 27.815 181.415 28.010 181.745 ;
        RECT 26.995 180.275 27.330 181.245 ;
        RECT 27.500 180.105 27.670 181.245 ;
        RECT 27.840 180.445 28.010 181.415 ;
        RECT 28.180 180.785 28.350 181.915 ;
        RECT 28.520 181.125 28.690 181.925 ;
        RECT 28.895 181.635 29.170 182.485 ;
        RECT 28.890 181.465 29.170 181.635 ;
        RECT 28.895 181.325 29.170 181.465 ;
        RECT 29.340 181.125 29.530 182.485 ;
        RECT 29.710 182.120 30.220 182.655 ;
        RECT 30.440 181.845 30.685 182.450 ;
        RECT 31.135 181.945 31.390 182.475 ;
        RECT 31.560 182.195 31.865 182.655 ;
        RECT 32.110 182.275 33.180 182.445 ;
        RECT 29.730 181.675 30.960 181.845 ;
        RECT 28.520 180.955 29.530 181.125 ;
        RECT 29.700 181.110 30.450 181.300 ;
        RECT 28.180 180.615 29.305 180.785 ;
        RECT 29.700 180.445 29.870 181.110 ;
        RECT 30.620 180.865 30.960 181.675 ;
        RECT 27.840 180.275 29.870 180.445 ;
        RECT 30.040 180.105 30.210 180.865 ;
        RECT 30.445 180.455 30.960 180.865 ;
        RECT 31.135 181.295 31.345 181.945 ;
        RECT 32.110 181.920 32.430 182.275 ;
        RECT 32.105 181.745 32.430 181.920 ;
        RECT 31.515 181.445 32.430 181.745 ;
        RECT 32.600 181.705 32.840 182.105 ;
        RECT 33.010 182.045 33.180 182.275 ;
        RECT 33.350 182.215 33.540 182.655 ;
        RECT 33.710 182.205 34.660 182.485 ;
        RECT 34.880 182.295 35.230 182.465 ;
        RECT 33.010 181.875 33.540 182.045 ;
        RECT 31.515 181.415 32.255 181.445 ;
        RECT 31.135 180.415 31.390 181.295 ;
        RECT 31.560 180.105 31.865 181.245 ;
        RECT 32.085 180.825 32.255 181.415 ;
        RECT 32.600 181.335 33.140 181.705 ;
        RECT 33.320 181.595 33.540 181.875 ;
        RECT 33.710 181.425 33.880 182.205 ;
        RECT 33.475 181.255 33.880 181.425 ;
        RECT 34.050 181.415 34.400 182.035 ;
        RECT 33.475 181.165 33.645 181.255 ;
        RECT 34.570 181.245 34.780 182.035 ;
        RECT 32.425 180.995 33.645 181.165 ;
        RECT 34.105 181.085 34.780 181.245 ;
        RECT 32.085 180.655 32.885 180.825 ;
        RECT 32.205 180.105 32.535 180.485 ;
        RECT 32.715 180.365 32.885 180.655 ;
        RECT 33.475 180.615 33.645 180.995 ;
        RECT 33.815 181.075 34.780 181.085 ;
        RECT 34.970 181.905 35.230 182.295 ;
        RECT 35.440 182.195 35.770 182.655 ;
        RECT 36.645 182.265 37.500 182.435 ;
        RECT 37.705 182.265 38.200 182.435 ;
        RECT 38.370 182.295 38.700 182.655 ;
        RECT 34.970 181.215 35.140 181.905 ;
        RECT 35.310 181.555 35.480 181.735 ;
        RECT 35.650 181.725 36.440 181.975 ;
        RECT 36.645 181.555 36.815 182.265 ;
        RECT 36.985 181.755 37.340 181.975 ;
        RECT 35.310 181.385 37.000 181.555 ;
        RECT 33.815 180.785 34.275 181.075 ;
        RECT 34.970 181.045 36.470 181.215 ;
        RECT 34.970 180.905 35.140 181.045 ;
        RECT 34.580 180.735 35.140 180.905 ;
        RECT 33.055 180.105 33.305 180.565 ;
        RECT 33.475 180.275 34.345 180.615 ;
        RECT 34.580 180.275 34.750 180.735 ;
        RECT 35.585 180.705 36.660 180.875 ;
        RECT 34.920 180.105 35.290 180.565 ;
        RECT 35.585 180.365 35.755 180.705 ;
        RECT 35.925 180.105 36.255 180.535 ;
        RECT 36.490 180.365 36.660 180.705 ;
        RECT 36.830 180.605 37.000 181.385 ;
        RECT 37.170 181.165 37.340 181.755 ;
        RECT 37.510 181.355 37.860 181.975 ;
        RECT 37.170 180.775 37.635 181.165 ;
        RECT 38.030 180.905 38.200 182.265 ;
        RECT 38.370 181.075 38.830 182.125 ;
        RECT 37.805 180.735 38.200 180.905 ;
        RECT 37.805 180.605 37.975 180.735 ;
        RECT 36.830 180.275 37.510 180.605 ;
        RECT 37.725 180.275 37.975 180.605 ;
        RECT 38.145 180.105 38.395 180.565 ;
        RECT 38.565 180.290 38.890 181.075 ;
        RECT 39.060 180.275 39.230 182.395 ;
        RECT 39.400 182.275 39.730 182.655 ;
        RECT 39.900 182.105 40.155 182.395 ;
        RECT 39.405 181.935 40.155 182.105 ;
        RECT 39.405 180.945 39.635 181.935 ;
        RECT 40.330 181.885 42.000 182.655 ;
        RECT 42.175 182.110 47.520 182.655 ;
        RECT 39.805 181.115 40.155 181.765 ;
        RECT 40.330 181.195 41.080 181.715 ;
        RECT 41.250 181.365 42.000 181.885 ;
        RECT 39.405 180.775 40.155 180.945 ;
        RECT 39.400 180.105 39.730 180.605 ;
        RECT 39.900 180.275 40.155 180.775 ;
        RECT 40.330 180.105 42.000 181.195 ;
        RECT 43.765 180.540 44.115 181.790 ;
        RECT 45.595 181.280 45.935 182.110 ;
        RECT 47.690 181.930 47.980 182.655 ;
        RECT 48.150 181.885 49.820 182.655 ;
        RECT 49.995 182.110 55.340 182.655 ;
        RECT 55.510 182.275 56.400 182.445 ;
        RECT 42.175 180.105 47.520 180.540 ;
        RECT 47.690 180.105 47.980 181.270 ;
        RECT 48.150 181.195 48.900 181.715 ;
        RECT 49.070 181.365 49.820 181.885 ;
        RECT 48.150 180.105 49.820 181.195 ;
        RECT 51.585 180.540 51.935 181.790 ;
        RECT 53.415 181.280 53.755 182.110 ;
        RECT 55.510 181.720 56.060 182.105 ;
        RECT 56.230 181.550 56.400 182.275 ;
        RECT 55.510 181.480 56.400 181.550 ;
        RECT 56.570 181.975 56.790 182.435 ;
        RECT 56.960 182.115 57.210 182.655 ;
        RECT 57.380 182.005 57.640 182.485 ;
        RECT 56.570 181.950 56.820 181.975 ;
        RECT 56.570 181.525 56.900 181.950 ;
        RECT 55.510 181.455 56.405 181.480 ;
        RECT 55.510 181.440 56.415 181.455 ;
        RECT 55.510 181.425 56.420 181.440 ;
        RECT 55.510 181.420 56.430 181.425 ;
        RECT 55.510 181.410 56.435 181.420 ;
        RECT 55.510 181.400 56.440 181.410 ;
        RECT 55.510 181.395 56.450 181.400 ;
        RECT 55.510 181.385 56.460 181.395 ;
        RECT 55.510 181.380 56.470 181.385 ;
        RECT 55.510 180.930 55.770 181.380 ;
        RECT 56.135 181.375 56.470 181.380 ;
        RECT 56.135 181.370 56.485 181.375 ;
        RECT 56.135 181.360 56.500 181.370 ;
        RECT 56.135 181.355 56.525 181.360 ;
        RECT 57.070 181.355 57.300 181.750 ;
        RECT 56.135 181.350 57.300 181.355 ;
        RECT 56.165 181.315 57.300 181.350 ;
        RECT 56.200 181.290 57.300 181.315 ;
        RECT 56.230 181.260 57.300 181.290 ;
        RECT 56.250 181.230 57.300 181.260 ;
        RECT 56.270 181.200 57.300 181.230 ;
        RECT 56.340 181.190 57.300 181.200 ;
        RECT 56.365 181.180 57.300 181.190 ;
        RECT 56.385 181.165 57.300 181.180 ;
        RECT 56.405 181.150 57.300 181.165 ;
        RECT 56.410 181.140 57.195 181.150 ;
        RECT 56.425 181.105 57.195 181.140 ;
        RECT 55.940 180.785 56.270 181.030 ;
        RECT 56.440 180.855 57.195 181.105 ;
        RECT 57.470 180.975 57.640 182.005 ;
        RECT 55.940 180.760 56.125 180.785 ;
        RECT 55.510 180.660 56.125 180.760 ;
        RECT 49.995 180.105 55.340 180.540 ;
        RECT 55.510 180.105 56.115 180.660 ;
        RECT 56.290 180.275 56.770 180.615 ;
        RECT 56.940 180.105 57.195 180.650 ;
        RECT 57.365 180.275 57.640 180.975 ;
        RECT 57.820 181.930 58.150 182.440 ;
        RECT 58.320 182.255 58.650 182.655 ;
        RECT 59.700 182.085 60.030 182.425 ;
        RECT 60.200 182.255 60.530 182.655 ;
        RECT 57.820 181.165 58.010 181.930 ;
        RECT 58.320 181.915 60.685 182.085 ;
        RECT 58.320 181.745 58.490 181.915 ;
        RECT 58.180 181.415 58.490 181.745 ;
        RECT 58.660 181.415 58.965 181.745 ;
        RECT 57.820 180.315 58.150 181.165 ;
        RECT 58.320 180.105 58.570 181.245 ;
        RECT 58.750 181.085 58.965 181.415 ;
        RECT 59.140 181.085 59.425 181.745 ;
        RECT 59.620 181.085 59.885 181.745 ;
        RECT 60.100 181.085 60.345 181.745 ;
        RECT 60.515 180.915 60.685 181.915 ;
        RECT 61.035 181.815 61.295 182.655 ;
        RECT 61.470 181.910 61.725 182.485 ;
        RECT 61.895 182.275 62.225 182.655 ;
        RECT 62.440 182.105 62.610 182.485 ;
        RECT 61.895 181.935 62.610 182.105 ;
        RECT 58.760 180.745 60.050 180.915 ;
        RECT 58.760 180.325 59.010 180.745 ;
        RECT 59.240 180.105 59.570 180.575 ;
        RECT 59.800 180.325 60.050 180.745 ;
        RECT 60.230 180.745 60.685 180.915 ;
        RECT 60.230 180.315 60.560 180.745 ;
        RECT 61.035 180.105 61.295 181.255 ;
        RECT 61.470 181.180 61.640 181.910 ;
        RECT 61.895 181.745 62.065 181.935 ;
        RECT 63.330 181.885 65.920 182.655 ;
        RECT 61.810 181.415 62.065 181.745 ;
        RECT 61.895 181.205 62.065 181.415 ;
        RECT 62.345 181.385 62.700 181.755 ;
        RECT 61.470 180.275 61.725 181.180 ;
        RECT 61.895 181.035 62.610 181.205 ;
        RECT 61.895 180.105 62.225 180.865 ;
        RECT 62.440 180.275 62.610 181.035 ;
        RECT 63.330 181.195 64.540 181.715 ;
        RECT 64.710 181.365 65.920 181.885 ;
        RECT 66.090 182.005 66.350 182.485 ;
        RECT 66.520 182.115 66.770 182.655 ;
        RECT 63.330 180.105 65.920 181.195 ;
        RECT 66.090 180.975 66.260 182.005 ;
        RECT 66.940 181.975 67.160 182.435 ;
        RECT 66.910 181.950 67.160 181.975 ;
        RECT 66.430 181.355 66.660 181.750 ;
        RECT 66.830 181.525 67.160 181.950 ;
        RECT 67.330 182.275 68.220 182.445 ;
        RECT 67.330 181.550 67.500 182.275 ;
        RECT 67.670 181.720 68.220 182.105 ;
        RECT 68.390 181.905 69.600 182.655 ;
        RECT 67.330 181.480 68.220 181.550 ;
        RECT 67.325 181.455 68.220 181.480 ;
        RECT 67.315 181.440 68.220 181.455 ;
        RECT 67.310 181.425 68.220 181.440 ;
        RECT 67.300 181.420 68.220 181.425 ;
        RECT 67.295 181.410 68.220 181.420 ;
        RECT 67.290 181.400 68.220 181.410 ;
        RECT 67.280 181.395 68.220 181.400 ;
        RECT 67.270 181.385 68.220 181.395 ;
        RECT 67.260 181.380 68.220 181.385 ;
        RECT 67.260 181.375 67.595 181.380 ;
        RECT 67.245 181.370 67.595 181.375 ;
        RECT 67.230 181.360 67.595 181.370 ;
        RECT 67.205 181.355 67.595 181.360 ;
        RECT 66.430 181.350 67.595 181.355 ;
        RECT 66.430 181.315 67.565 181.350 ;
        RECT 66.430 181.290 67.530 181.315 ;
        RECT 66.430 181.260 67.500 181.290 ;
        RECT 66.430 181.230 67.480 181.260 ;
        RECT 66.430 181.200 67.460 181.230 ;
        RECT 66.430 181.190 67.390 181.200 ;
        RECT 66.430 181.180 67.365 181.190 ;
        RECT 66.430 181.165 67.345 181.180 ;
        RECT 66.430 181.150 67.325 181.165 ;
        RECT 66.535 181.140 67.320 181.150 ;
        RECT 66.535 181.105 67.305 181.140 ;
        RECT 66.090 180.275 66.365 180.975 ;
        RECT 66.535 180.855 67.290 181.105 ;
        RECT 67.460 180.785 67.790 181.030 ;
        RECT 67.960 180.930 68.220 181.380 ;
        RECT 68.390 181.195 68.910 181.735 ;
        RECT 69.080 181.365 69.600 181.905 ;
        RECT 69.770 181.885 73.280 182.655 ;
        RECT 73.450 181.930 73.740 182.655 ;
        RECT 74.370 181.885 76.040 182.655 ;
        RECT 69.770 181.195 71.460 181.715 ;
        RECT 71.630 181.365 73.280 181.885 ;
        RECT 67.605 180.760 67.790 180.785 ;
        RECT 67.605 180.660 68.220 180.760 ;
        RECT 66.535 180.105 66.790 180.650 ;
        RECT 66.960 180.275 67.440 180.615 ;
        RECT 67.615 180.105 68.220 180.660 ;
        RECT 68.390 180.105 69.600 181.195 ;
        RECT 69.770 180.105 73.280 181.195 ;
        RECT 73.450 180.105 73.740 181.270 ;
        RECT 74.370 181.195 75.120 181.715 ;
        RECT 75.290 181.365 76.040 181.885 ;
        RECT 76.485 181.845 76.730 182.450 ;
        RECT 76.950 182.120 77.460 182.655 ;
        RECT 76.210 181.675 77.440 181.845 ;
        RECT 74.370 180.105 76.040 181.195 ;
        RECT 76.210 180.865 76.550 181.675 ;
        RECT 76.720 181.110 77.470 181.300 ;
        RECT 76.210 180.455 76.725 180.865 ;
        RECT 76.960 180.105 77.130 180.865 ;
        RECT 77.300 180.445 77.470 181.110 ;
        RECT 77.640 181.125 77.830 182.485 ;
        RECT 78.000 181.635 78.275 182.485 ;
        RECT 78.465 182.120 78.995 182.485 ;
        RECT 79.420 182.255 79.750 182.655 ;
        RECT 78.820 182.085 78.995 182.120 ;
        RECT 78.000 181.465 78.280 181.635 ;
        RECT 78.000 181.325 78.275 181.465 ;
        RECT 78.480 181.125 78.650 181.925 ;
        RECT 77.640 180.955 78.650 181.125 ;
        RECT 78.820 181.915 79.750 182.085 ;
        RECT 79.920 181.915 80.175 182.485 ;
        RECT 78.820 180.785 78.990 181.915 ;
        RECT 79.580 181.745 79.750 181.915 ;
        RECT 77.865 180.615 78.990 180.785 ;
        RECT 79.160 181.415 79.355 181.745 ;
        RECT 79.580 181.415 79.835 181.745 ;
        RECT 79.160 180.445 79.330 181.415 ;
        RECT 80.005 181.245 80.175 181.915 ;
        RECT 80.810 181.885 84.320 182.655 ;
        RECT 84.495 182.110 89.840 182.655 ;
        RECT 77.300 180.275 79.330 180.445 ;
        RECT 79.500 180.105 79.670 181.245 ;
        RECT 79.840 180.275 80.175 181.245 ;
        RECT 80.810 181.195 82.500 181.715 ;
        RECT 82.670 181.365 84.320 181.885 ;
        RECT 80.810 180.105 84.320 181.195 ;
        RECT 86.085 180.540 86.435 181.790 ;
        RECT 87.915 181.280 88.255 182.110 ;
        RECT 90.015 181.945 90.270 182.475 ;
        RECT 90.440 182.195 90.745 182.655 ;
        RECT 90.990 182.275 92.060 182.445 ;
        RECT 90.015 181.295 90.225 181.945 ;
        RECT 90.990 181.920 91.310 182.275 ;
        RECT 90.985 181.745 91.310 181.920 ;
        RECT 90.395 181.445 91.310 181.745 ;
        RECT 91.480 181.705 91.720 182.105 ;
        RECT 91.890 182.045 92.060 182.275 ;
        RECT 92.230 182.215 92.420 182.655 ;
        RECT 92.590 182.205 93.540 182.485 ;
        RECT 93.760 182.295 94.110 182.465 ;
        RECT 91.890 181.875 92.420 182.045 ;
        RECT 90.395 181.415 91.135 181.445 ;
        RECT 84.495 180.105 89.840 180.540 ;
        RECT 90.015 180.415 90.270 181.295 ;
        RECT 90.440 180.105 90.745 181.245 ;
        RECT 90.965 180.825 91.135 181.415 ;
        RECT 91.480 181.335 92.020 181.705 ;
        RECT 92.200 181.595 92.420 181.875 ;
        RECT 92.590 181.425 92.760 182.205 ;
        RECT 92.355 181.255 92.760 181.425 ;
        RECT 92.930 181.415 93.280 182.035 ;
        RECT 92.355 181.165 92.525 181.255 ;
        RECT 93.450 181.245 93.660 182.035 ;
        RECT 91.305 180.995 92.525 181.165 ;
        RECT 92.985 181.085 93.660 181.245 ;
        RECT 90.965 180.655 91.765 180.825 ;
        RECT 91.085 180.105 91.415 180.485 ;
        RECT 91.595 180.365 91.765 180.655 ;
        RECT 92.355 180.615 92.525 180.995 ;
        RECT 92.695 181.075 93.660 181.085 ;
        RECT 93.850 181.905 94.110 182.295 ;
        RECT 94.320 182.195 94.650 182.655 ;
        RECT 95.525 182.265 96.380 182.435 ;
        RECT 96.585 182.265 97.080 182.435 ;
        RECT 97.250 182.295 97.580 182.655 ;
        RECT 93.850 181.215 94.020 181.905 ;
        RECT 94.190 181.555 94.360 181.735 ;
        RECT 94.530 181.725 95.320 181.975 ;
        RECT 95.525 181.555 95.695 182.265 ;
        RECT 95.865 181.755 96.220 181.975 ;
        RECT 94.190 181.385 95.880 181.555 ;
        RECT 92.695 180.785 93.155 181.075 ;
        RECT 93.850 181.045 95.350 181.215 ;
        RECT 93.850 180.905 94.020 181.045 ;
        RECT 93.460 180.735 94.020 180.905 ;
        RECT 91.935 180.105 92.185 180.565 ;
        RECT 92.355 180.275 93.225 180.615 ;
        RECT 93.460 180.275 93.630 180.735 ;
        RECT 94.465 180.705 95.540 180.875 ;
        RECT 93.800 180.105 94.170 180.565 ;
        RECT 94.465 180.365 94.635 180.705 ;
        RECT 94.805 180.105 95.135 180.535 ;
        RECT 95.370 180.365 95.540 180.705 ;
        RECT 95.710 180.605 95.880 181.385 ;
        RECT 96.050 181.165 96.220 181.755 ;
        RECT 96.390 181.355 96.740 181.975 ;
        RECT 96.050 180.775 96.515 181.165 ;
        RECT 96.910 180.905 97.080 182.265 ;
        RECT 97.250 181.075 97.710 182.125 ;
        RECT 96.685 180.735 97.080 180.905 ;
        RECT 96.685 180.605 96.855 180.735 ;
        RECT 95.710 180.275 96.390 180.605 ;
        RECT 96.605 180.275 96.855 180.605 ;
        RECT 97.025 180.105 97.275 180.565 ;
        RECT 97.445 180.290 97.770 181.075 ;
        RECT 97.940 180.275 98.110 182.395 ;
        RECT 98.280 182.275 98.610 182.655 ;
        RECT 98.780 182.105 99.035 182.395 ;
        RECT 98.285 181.935 99.035 182.105 ;
        RECT 98.285 180.945 98.515 181.935 ;
        RECT 99.210 181.930 99.500 182.655 ;
        RECT 99.670 181.980 99.930 182.485 ;
        RECT 100.110 182.275 100.440 182.655 ;
        RECT 100.620 182.105 100.790 182.485 ;
        RECT 98.685 181.115 99.035 181.765 ;
        RECT 98.285 180.775 99.035 180.945 ;
        RECT 98.280 180.105 98.610 180.605 ;
        RECT 98.780 180.275 99.035 180.775 ;
        RECT 99.210 180.105 99.500 181.270 ;
        RECT 99.670 181.180 99.840 181.980 ;
        RECT 100.125 181.935 100.790 182.105 ;
        RECT 101.055 181.945 101.310 182.475 ;
        RECT 101.480 182.195 101.785 182.655 ;
        RECT 102.030 182.275 103.100 182.445 ;
        RECT 100.125 181.680 100.295 181.935 ;
        RECT 100.010 181.350 100.295 181.680 ;
        RECT 100.530 181.385 100.860 181.755 ;
        RECT 100.125 181.205 100.295 181.350 ;
        RECT 101.055 181.295 101.265 181.945 ;
        RECT 102.030 181.920 102.350 182.275 ;
        RECT 102.025 181.745 102.350 181.920 ;
        RECT 101.435 181.445 102.350 181.745 ;
        RECT 102.520 181.705 102.760 182.105 ;
        RECT 102.930 182.045 103.100 182.275 ;
        RECT 103.270 182.215 103.460 182.655 ;
        RECT 103.630 182.205 104.580 182.485 ;
        RECT 104.800 182.295 105.150 182.465 ;
        RECT 102.930 181.875 103.460 182.045 ;
        RECT 101.435 181.415 102.175 181.445 ;
        RECT 99.670 180.275 99.940 181.180 ;
        RECT 100.125 181.035 100.790 181.205 ;
        RECT 100.110 180.105 100.440 180.865 ;
        RECT 100.620 180.275 100.790 181.035 ;
        RECT 101.055 180.415 101.310 181.295 ;
        RECT 101.480 180.105 101.785 181.245 ;
        RECT 102.005 180.825 102.175 181.415 ;
        RECT 102.520 181.335 103.060 181.705 ;
        RECT 103.240 181.595 103.460 181.875 ;
        RECT 103.630 181.425 103.800 182.205 ;
        RECT 103.395 181.255 103.800 181.425 ;
        RECT 103.970 181.415 104.320 182.035 ;
        RECT 103.395 181.165 103.565 181.255 ;
        RECT 104.490 181.245 104.700 182.035 ;
        RECT 102.345 180.995 103.565 181.165 ;
        RECT 104.025 181.085 104.700 181.245 ;
        RECT 102.005 180.655 102.805 180.825 ;
        RECT 102.125 180.105 102.455 180.485 ;
        RECT 102.635 180.365 102.805 180.655 ;
        RECT 103.395 180.615 103.565 180.995 ;
        RECT 103.735 181.075 104.700 181.085 ;
        RECT 104.890 181.905 105.150 182.295 ;
        RECT 105.360 182.195 105.690 182.655 ;
        RECT 106.565 182.265 107.420 182.435 ;
        RECT 107.625 182.265 108.120 182.435 ;
        RECT 108.290 182.295 108.620 182.655 ;
        RECT 104.890 181.215 105.060 181.905 ;
        RECT 105.230 181.555 105.400 181.735 ;
        RECT 105.570 181.725 106.360 181.975 ;
        RECT 106.565 181.555 106.735 182.265 ;
        RECT 106.905 181.755 107.260 181.975 ;
        RECT 105.230 181.385 106.920 181.555 ;
        RECT 103.735 180.785 104.195 181.075 ;
        RECT 104.890 181.045 106.390 181.215 ;
        RECT 104.890 180.905 105.060 181.045 ;
        RECT 104.500 180.735 105.060 180.905 ;
        RECT 102.975 180.105 103.225 180.565 ;
        RECT 103.395 180.275 104.265 180.615 ;
        RECT 104.500 180.275 104.670 180.735 ;
        RECT 105.505 180.705 106.580 180.875 ;
        RECT 104.840 180.105 105.210 180.565 ;
        RECT 105.505 180.365 105.675 180.705 ;
        RECT 105.845 180.105 106.175 180.535 ;
        RECT 106.410 180.365 106.580 180.705 ;
        RECT 106.750 180.605 106.920 181.385 ;
        RECT 107.090 181.165 107.260 181.755 ;
        RECT 107.430 181.355 107.780 181.975 ;
        RECT 107.090 180.775 107.555 181.165 ;
        RECT 107.950 180.905 108.120 182.265 ;
        RECT 108.290 181.075 108.750 182.125 ;
        RECT 107.725 180.735 108.120 180.905 ;
        RECT 107.725 180.605 107.895 180.735 ;
        RECT 106.750 180.275 107.430 180.605 ;
        RECT 107.645 180.275 107.895 180.605 ;
        RECT 108.065 180.105 108.315 180.565 ;
        RECT 108.485 180.290 108.810 181.075 ;
        RECT 108.980 180.275 109.150 182.395 ;
        RECT 109.320 182.275 109.650 182.655 ;
        RECT 109.820 182.105 110.075 182.395 ;
        RECT 109.325 181.935 110.075 182.105 ;
        RECT 109.325 180.945 109.555 181.935 ;
        RECT 111.170 181.905 112.380 182.655 ;
        RECT 109.725 181.115 110.075 181.765 ;
        RECT 111.170 181.195 111.690 181.735 ;
        RECT 111.860 181.365 112.380 181.905 ;
        RECT 109.325 180.775 110.075 180.945 ;
        RECT 109.320 180.105 109.650 180.605 ;
        RECT 109.820 180.275 110.075 180.775 ;
        RECT 111.170 180.105 112.380 181.195 ;
        RECT 18.165 179.935 112.465 180.105 ;
        RECT 18.250 178.845 19.460 179.935 ;
        RECT 18.250 178.135 18.770 178.675 ;
        RECT 18.940 178.305 19.460 178.845 ;
        RECT 20.095 178.745 20.350 179.625 ;
        RECT 20.520 178.795 20.825 179.935 ;
        RECT 21.165 179.555 21.495 179.935 ;
        RECT 21.675 179.385 21.845 179.675 ;
        RECT 22.015 179.475 22.265 179.935 ;
        RECT 21.045 179.215 21.845 179.385 ;
        RECT 22.435 179.425 23.305 179.765 ;
        RECT 18.250 177.385 19.460 178.135 ;
        RECT 20.095 178.095 20.305 178.745 ;
        RECT 21.045 178.625 21.215 179.215 ;
        RECT 22.435 179.045 22.605 179.425 ;
        RECT 23.540 179.305 23.710 179.765 ;
        RECT 23.880 179.475 24.250 179.935 ;
        RECT 24.545 179.335 24.715 179.675 ;
        RECT 24.885 179.505 25.215 179.935 ;
        RECT 25.450 179.335 25.620 179.675 ;
        RECT 21.385 178.875 22.605 179.045 ;
        RECT 22.775 178.965 23.235 179.255 ;
        RECT 23.540 179.135 24.100 179.305 ;
        RECT 24.545 179.165 25.620 179.335 ;
        RECT 25.790 179.435 26.470 179.765 ;
        RECT 26.685 179.435 26.935 179.765 ;
        RECT 27.105 179.475 27.355 179.935 ;
        RECT 23.930 178.995 24.100 179.135 ;
        RECT 22.775 178.955 23.740 178.965 ;
        RECT 22.435 178.785 22.605 178.875 ;
        RECT 23.065 178.795 23.740 178.955 ;
        RECT 20.475 178.595 21.215 178.625 ;
        RECT 20.475 178.295 21.390 178.595 ;
        RECT 21.065 178.120 21.390 178.295 ;
        RECT 20.095 177.565 20.350 178.095 ;
        RECT 20.520 177.385 20.825 177.845 ;
        RECT 21.070 177.765 21.390 178.120 ;
        RECT 21.560 178.335 22.100 178.705 ;
        RECT 22.435 178.615 22.840 178.785 ;
        RECT 21.560 177.935 21.800 178.335 ;
        RECT 22.280 178.165 22.500 178.445 ;
        RECT 21.970 177.995 22.500 178.165 ;
        RECT 21.970 177.765 22.140 177.995 ;
        RECT 22.670 177.835 22.840 178.615 ;
        RECT 23.010 178.005 23.360 178.625 ;
        RECT 23.530 178.005 23.740 178.795 ;
        RECT 23.930 178.825 25.430 178.995 ;
        RECT 23.930 178.135 24.100 178.825 ;
        RECT 25.790 178.655 25.960 179.435 ;
        RECT 26.765 179.305 26.935 179.435 ;
        RECT 24.270 178.485 25.960 178.655 ;
        RECT 26.130 178.875 26.595 179.265 ;
        RECT 26.765 179.135 27.160 179.305 ;
        RECT 24.270 178.305 24.440 178.485 ;
        RECT 21.070 177.595 22.140 177.765 ;
        RECT 22.310 177.385 22.500 177.825 ;
        RECT 22.670 177.555 23.620 177.835 ;
        RECT 23.930 177.745 24.190 178.135 ;
        RECT 24.610 178.065 25.400 178.315 ;
        RECT 23.840 177.575 24.190 177.745 ;
        RECT 24.400 177.385 24.730 177.845 ;
        RECT 25.605 177.775 25.775 178.485 ;
        RECT 26.130 178.285 26.300 178.875 ;
        RECT 25.945 178.065 26.300 178.285 ;
        RECT 26.470 178.065 26.820 178.685 ;
        RECT 26.990 177.775 27.160 179.135 ;
        RECT 27.525 178.965 27.850 179.750 ;
        RECT 27.330 177.915 27.790 178.965 ;
        RECT 25.605 177.605 26.460 177.775 ;
        RECT 26.665 177.605 27.160 177.775 ;
        RECT 27.330 177.385 27.660 177.745 ;
        RECT 28.020 177.645 28.190 179.765 ;
        RECT 28.360 179.435 28.690 179.935 ;
        RECT 28.860 179.265 29.115 179.765 ;
        RECT 28.365 179.095 29.115 179.265 ;
        RECT 28.365 178.105 28.595 179.095 ;
        RECT 28.765 178.275 29.115 178.925 ;
        RECT 29.290 178.860 29.560 179.765 ;
        RECT 29.730 179.175 30.060 179.935 ;
        RECT 30.240 179.005 30.410 179.765 ;
        RECT 28.365 177.935 29.115 178.105 ;
        RECT 28.360 177.385 28.690 177.765 ;
        RECT 28.860 177.645 29.115 177.935 ;
        RECT 29.290 178.060 29.460 178.860 ;
        RECT 29.745 178.835 30.410 179.005 ;
        RECT 30.670 179.175 31.185 179.585 ;
        RECT 31.420 179.175 31.590 179.935 ;
        RECT 31.760 179.595 33.790 179.765 ;
        RECT 29.745 178.690 29.915 178.835 ;
        RECT 29.630 178.360 29.915 178.690 ;
        RECT 29.745 178.105 29.915 178.360 ;
        RECT 30.150 178.285 30.480 178.655 ;
        RECT 30.670 178.365 31.010 179.175 ;
        RECT 31.760 178.930 31.930 179.595 ;
        RECT 32.325 179.255 33.450 179.425 ;
        RECT 31.180 178.740 31.930 178.930 ;
        RECT 32.100 178.915 33.110 179.085 ;
        RECT 30.670 178.195 31.900 178.365 ;
        RECT 29.290 177.555 29.550 178.060 ;
        RECT 29.745 177.935 30.410 178.105 ;
        RECT 29.730 177.385 30.060 177.765 ;
        RECT 30.240 177.555 30.410 177.935 ;
        RECT 30.945 177.590 31.190 178.195 ;
        RECT 31.410 177.385 31.920 177.920 ;
        RECT 32.100 177.555 32.290 178.915 ;
        RECT 32.460 177.895 32.735 178.715 ;
        RECT 32.940 178.115 33.110 178.915 ;
        RECT 33.280 178.125 33.450 179.255 ;
        RECT 33.620 178.625 33.790 179.595 ;
        RECT 33.960 178.795 34.130 179.935 ;
        RECT 34.300 178.795 34.635 179.765 ;
        RECT 33.620 178.295 33.815 178.625 ;
        RECT 34.040 178.295 34.295 178.625 ;
        RECT 34.040 178.125 34.210 178.295 ;
        RECT 34.465 178.125 34.635 178.795 ;
        RECT 34.810 178.770 35.100 179.935 ;
        RECT 35.330 178.795 35.540 179.935 ;
        RECT 35.710 178.785 36.040 179.765 ;
        RECT 36.210 178.795 36.440 179.935 ;
        RECT 37.200 179.005 37.370 179.765 ;
        RECT 37.550 179.175 37.880 179.935 ;
        RECT 37.200 178.835 37.865 179.005 ;
        RECT 38.050 178.860 38.320 179.765 ;
        RECT 33.280 177.955 34.210 178.125 ;
        RECT 33.280 177.920 33.455 177.955 ;
        RECT 32.460 177.725 32.740 177.895 ;
        RECT 32.460 177.555 32.735 177.725 ;
        RECT 32.925 177.555 33.455 177.920 ;
        RECT 33.880 177.385 34.210 177.785 ;
        RECT 34.380 177.555 34.635 178.125 ;
        RECT 34.810 177.385 35.100 178.110 ;
        RECT 35.330 177.385 35.540 178.205 ;
        RECT 35.710 178.185 35.960 178.785 ;
        RECT 37.695 178.690 37.865 178.835 ;
        RECT 36.130 178.375 36.460 178.625 ;
        RECT 37.130 178.285 37.460 178.655 ;
        RECT 37.695 178.360 37.980 178.690 ;
        RECT 35.710 177.555 36.040 178.185 ;
        RECT 36.210 177.385 36.440 178.205 ;
        RECT 37.695 178.105 37.865 178.360 ;
        RECT 37.200 177.935 37.865 178.105 ;
        RECT 38.150 178.060 38.320 178.860 ;
        RECT 37.200 177.555 37.370 177.935 ;
        RECT 37.550 177.385 37.880 177.765 ;
        RECT 38.060 177.555 38.320 178.060 ;
        RECT 38.490 178.860 38.760 179.765 ;
        RECT 38.930 179.175 39.260 179.935 ;
        RECT 39.440 179.005 39.610 179.765 ;
        RECT 38.490 178.060 38.660 178.860 ;
        RECT 38.945 178.835 39.610 179.005 ;
        RECT 39.870 178.845 43.380 179.935 ;
        RECT 38.945 178.690 39.115 178.835 ;
        RECT 38.830 178.360 39.115 178.690 ;
        RECT 38.945 178.105 39.115 178.360 ;
        RECT 39.350 178.285 39.680 178.655 ;
        RECT 39.870 178.325 41.560 178.845 ;
        RECT 43.610 178.795 43.820 179.935 ;
        RECT 43.990 178.785 44.320 179.765 ;
        RECT 44.490 178.795 44.720 179.935 ;
        RECT 45.305 178.955 45.560 179.625 ;
        RECT 45.740 179.135 46.025 179.935 ;
        RECT 46.205 179.215 46.535 179.725 ;
        RECT 41.730 178.155 43.380 178.675 ;
        RECT 38.490 177.555 38.750 178.060 ;
        RECT 38.945 177.935 39.610 178.105 ;
        RECT 38.930 177.385 39.260 177.765 ;
        RECT 39.440 177.555 39.610 177.935 ;
        RECT 39.870 177.385 43.380 178.155 ;
        RECT 43.610 177.385 43.820 178.205 ;
        RECT 43.990 178.185 44.240 178.785 ;
        RECT 44.410 178.375 44.740 178.625 ;
        RECT 43.990 177.555 44.320 178.185 ;
        RECT 44.490 177.385 44.720 178.205 ;
        RECT 45.305 178.095 45.485 178.955 ;
        RECT 46.205 178.625 46.455 179.215 ;
        RECT 46.805 179.065 46.975 179.675 ;
        RECT 47.145 179.245 47.475 179.935 ;
        RECT 47.705 179.385 47.945 179.675 ;
        RECT 48.145 179.555 48.565 179.935 ;
        RECT 48.745 179.465 49.375 179.715 ;
        RECT 49.845 179.555 50.175 179.935 ;
        RECT 48.745 179.385 48.915 179.465 ;
        RECT 50.345 179.385 50.515 179.675 ;
        RECT 50.695 179.555 51.075 179.935 ;
        RECT 51.315 179.550 52.145 179.720 ;
        RECT 47.705 179.215 48.915 179.385 ;
        RECT 45.655 178.295 46.455 178.625 ;
        RECT 45.305 177.895 45.560 178.095 ;
        RECT 45.220 177.725 45.560 177.895 ;
        RECT 45.305 177.565 45.560 177.725 ;
        RECT 45.740 177.385 46.025 177.845 ;
        RECT 46.205 177.645 46.455 178.295 ;
        RECT 46.655 179.045 46.975 179.065 ;
        RECT 46.655 178.875 48.575 179.045 ;
        RECT 46.655 177.980 46.845 178.875 ;
        RECT 48.745 178.705 48.915 179.215 ;
        RECT 49.085 178.955 49.605 179.265 ;
        RECT 47.015 178.535 48.915 178.705 ;
        RECT 47.015 178.475 47.345 178.535 ;
        RECT 47.495 178.305 47.825 178.365 ;
        RECT 47.165 178.035 47.825 178.305 ;
        RECT 46.655 177.650 46.975 177.980 ;
        RECT 47.155 177.385 47.815 177.865 ;
        RECT 48.015 177.775 48.185 178.535 ;
        RECT 49.085 178.365 49.265 178.775 ;
        RECT 48.355 178.195 48.685 178.315 ;
        RECT 49.435 178.195 49.605 178.955 ;
        RECT 48.355 178.025 49.605 178.195 ;
        RECT 49.775 179.135 51.145 179.385 ;
        RECT 49.775 178.365 49.965 179.135 ;
        RECT 50.895 178.875 51.145 179.135 ;
        RECT 50.135 178.705 50.385 178.865 ;
        RECT 51.315 178.705 51.485 179.550 ;
        RECT 52.380 179.265 52.550 179.765 ;
        RECT 52.720 179.435 53.050 179.935 ;
        RECT 51.655 178.875 52.155 179.255 ;
        RECT 52.380 179.095 53.075 179.265 ;
        RECT 50.135 178.535 51.485 178.705 ;
        RECT 51.065 178.495 51.485 178.535 ;
        RECT 49.775 178.025 50.195 178.365 ;
        RECT 50.485 178.035 50.895 178.365 ;
        RECT 48.015 177.605 48.865 177.775 ;
        RECT 49.425 177.385 49.745 177.845 ;
        RECT 49.945 177.595 50.195 178.025 ;
        RECT 50.485 177.385 50.895 177.825 ;
        RECT 51.065 177.765 51.235 178.495 ;
        RECT 51.405 177.945 51.755 178.315 ;
        RECT 51.935 178.005 52.155 178.875 ;
        RECT 52.325 178.305 52.735 178.925 ;
        RECT 52.905 178.125 53.075 179.095 ;
        RECT 52.380 177.935 53.075 178.125 ;
        RECT 51.065 177.565 52.080 177.765 ;
        RECT 52.380 177.605 52.550 177.935 ;
        RECT 52.720 177.385 53.050 177.765 ;
        RECT 53.265 177.645 53.490 179.765 ;
        RECT 53.660 179.435 53.990 179.935 ;
        RECT 54.160 179.265 54.330 179.765 ;
        RECT 53.665 179.095 54.330 179.265 ;
        RECT 53.665 178.105 53.895 179.095 ;
        RECT 54.065 178.275 54.415 178.925 ;
        RECT 55.050 178.845 56.720 179.935 ;
        RECT 56.975 179.315 57.150 179.765 ;
        RECT 57.320 179.495 57.650 179.935 ;
        RECT 57.955 179.345 58.125 179.765 ;
        RECT 58.360 179.525 59.030 179.935 ;
        RECT 59.245 179.345 59.415 179.765 ;
        RECT 59.615 179.525 59.945 179.935 ;
        RECT 56.975 179.145 57.605 179.315 ;
        RECT 55.050 178.325 55.800 178.845 ;
        RECT 55.970 178.155 56.720 178.675 ;
        RECT 56.890 178.295 57.255 178.975 ;
        RECT 57.435 178.625 57.605 179.145 ;
        RECT 57.955 179.175 59.970 179.345 ;
        RECT 57.435 178.295 57.785 178.625 ;
        RECT 53.665 177.935 54.330 178.105 ;
        RECT 53.660 177.385 53.990 177.765 ;
        RECT 54.160 177.645 54.330 177.935 ;
        RECT 55.050 177.385 56.720 178.155 ;
        RECT 57.435 178.125 57.605 178.295 ;
        RECT 56.975 177.955 57.605 178.125 ;
        RECT 56.975 177.555 57.150 177.955 ;
        RECT 57.955 177.885 58.125 179.175 ;
        RECT 57.320 177.385 57.650 177.765 ;
        RECT 57.895 177.555 58.125 177.885 ;
        RECT 58.325 177.720 58.605 178.995 ;
        RECT 58.830 177.895 59.100 178.995 ;
        RECT 59.290 177.965 59.630 178.995 ;
        RECT 59.800 178.625 59.970 179.175 ;
        RECT 60.140 178.795 60.400 179.765 ;
        RECT 59.800 178.295 60.060 178.625 ;
        RECT 60.230 178.105 60.400 178.795 ;
        RECT 60.570 178.770 60.860 179.935 ;
        RECT 61.030 178.965 61.300 179.735 ;
        RECT 61.470 179.155 61.800 179.935 ;
        RECT 62.005 179.330 62.190 179.735 ;
        RECT 62.360 179.510 62.695 179.935 ;
        RECT 62.005 179.155 62.670 179.330 ;
        RECT 61.030 178.795 62.160 178.965 ;
        RECT 58.790 177.725 59.100 177.895 ;
        RECT 58.830 177.720 59.100 177.725 ;
        RECT 59.560 177.385 59.890 177.765 ;
        RECT 60.060 177.640 60.400 178.105 ;
        RECT 60.060 177.595 60.395 177.640 ;
        RECT 60.570 177.385 60.860 178.110 ;
        RECT 61.030 177.885 61.200 178.795 ;
        RECT 61.370 178.045 61.730 178.625 ;
        RECT 61.910 178.295 62.160 178.795 ;
        RECT 62.330 178.125 62.670 179.155 ;
        RECT 63.330 178.845 66.840 179.935 ;
        RECT 63.330 178.325 65.020 178.845 ;
        RECT 67.070 178.795 67.280 179.935 ;
        RECT 67.450 178.785 67.780 179.765 ;
        RECT 67.950 178.795 68.180 179.935 ;
        RECT 68.430 178.795 68.660 179.935 ;
        RECT 68.830 178.785 69.160 179.765 ;
        RECT 69.330 178.795 69.540 179.935 ;
        RECT 69.780 178.955 70.110 179.765 ;
        RECT 70.280 179.135 70.520 179.935 ;
        RECT 69.780 178.785 70.495 178.955 ;
        RECT 65.190 178.155 66.840 178.675 ;
        RECT 61.985 177.955 62.670 178.125 ;
        RECT 61.030 177.555 61.290 177.885 ;
        RECT 61.500 177.385 61.775 177.865 ;
        RECT 61.985 177.555 62.190 177.955 ;
        RECT 62.360 177.385 62.695 177.785 ;
        RECT 63.330 177.385 66.840 178.155 ;
        RECT 67.070 177.385 67.280 178.205 ;
        RECT 67.450 178.185 67.700 178.785 ;
        RECT 67.870 178.375 68.200 178.625 ;
        RECT 68.410 178.375 68.740 178.625 ;
        RECT 67.450 177.555 67.780 178.185 ;
        RECT 67.950 177.385 68.180 178.205 ;
        RECT 68.430 177.385 68.660 178.205 ;
        RECT 68.910 178.185 69.160 178.785 ;
        RECT 69.775 178.375 70.155 178.615 ;
        RECT 70.325 178.545 70.495 178.785 ;
        RECT 70.700 178.915 70.870 179.765 ;
        RECT 71.040 179.135 71.370 179.935 ;
        RECT 71.540 178.915 71.710 179.765 ;
        RECT 70.700 178.745 71.710 178.915 ;
        RECT 71.880 178.785 72.210 179.935 ;
        RECT 72.590 178.795 72.800 179.935 ;
        RECT 72.970 178.785 73.300 179.765 ;
        RECT 73.470 178.795 73.700 179.935 ;
        RECT 70.325 178.375 70.825 178.545 ;
        RECT 70.325 178.205 70.495 178.375 ;
        RECT 71.215 178.205 71.710 178.745 ;
        RECT 68.830 177.555 69.160 178.185 ;
        RECT 69.330 177.385 69.540 178.205 ;
        RECT 69.860 178.035 70.495 178.205 ;
        RECT 70.700 178.035 71.710 178.205 ;
        RECT 69.860 177.555 70.030 178.035 ;
        RECT 70.210 177.385 70.450 177.865 ;
        RECT 70.700 177.555 70.870 178.035 ;
        RECT 71.040 177.385 71.370 177.865 ;
        RECT 71.540 177.555 71.710 178.035 ;
        RECT 71.880 177.385 72.210 178.185 ;
        RECT 72.590 177.385 72.800 178.205 ;
        RECT 72.970 178.185 73.220 178.785 ;
        RECT 73.915 178.745 74.170 179.625 ;
        RECT 74.340 178.795 74.645 179.935 ;
        RECT 74.985 179.555 75.315 179.935 ;
        RECT 75.495 179.385 75.665 179.675 ;
        RECT 75.835 179.475 76.085 179.935 ;
        RECT 74.865 179.215 75.665 179.385 ;
        RECT 76.255 179.425 77.125 179.765 ;
        RECT 73.390 178.375 73.720 178.625 ;
        RECT 72.970 177.555 73.300 178.185 ;
        RECT 73.470 177.385 73.700 178.205 ;
        RECT 73.915 178.095 74.125 178.745 ;
        RECT 74.865 178.625 75.035 179.215 ;
        RECT 76.255 179.045 76.425 179.425 ;
        RECT 77.360 179.305 77.530 179.765 ;
        RECT 77.700 179.475 78.070 179.935 ;
        RECT 78.365 179.335 78.535 179.675 ;
        RECT 78.705 179.505 79.035 179.935 ;
        RECT 79.270 179.335 79.440 179.675 ;
        RECT 75.205 178.875 76.425 179.045 ;
        RECT 76.595 178.965 77.055 179.255 ;
        RECT 77.360 179.135 77.920 179.305 ;
        RECT 78.365 179.165 79.440 179.335 ;
        RECT 79.610 179.435 80.290 179.765 ;
        RECT 80.505 179.435 80.755 179.765 ;
        RECT 80.925 179.475 81.175 179.935 ;
        RECT 77.750 178.995 77.920 179.135 ;
        RECT 76.595 178.955 77.560 178.965 ;
        RECT 76.255 178.785 76.425 178.875 ;
        RECT 76.885 178.795 77.560 178.955 ;
        RECT 74.295 178.595 75.035 178.625 ;
        RECT 74.295 178.295 75.210 178.595 ;
        RECT 74.885 178.120 75.210 178.295 ;
        RECT 73.915 177.565 74.170 178.095 ;
        RECT 74.340 177.385 74.645 177.845 ;
        RECT 74.890 177.765 75.210 178.120 ;
        RECT 75.380 178.335 75.920 178.705 ;
        RECT 76.255 178.615 76.660 178.785 ;
        RECT 75.380 177.935 75.620 178.335 ;
        RECT 76.100 178.165 76.320 178.445 ;
        RECT 75.790 177.995 76.320 178.165 ;
        RECT 75.790 177.765 75.960 177.995 ;
        RECT 76.490 177.835 76.660 178.615 ;
        RECT 76.830 178.005 77.180 178.625 ;
        RECT 77.350 178.005 77.560 178.795 ;
        RECT 77.750 178.825 79.250 178.995 ;
        RECT 77.750 178.135 77.920 178.825 ;
        RECT 79.610 178.655 79.780 179.435 ;
        RECT 80.585 179.305 80.755 179.435 ;
        RECT 78.090 178.485 79.780 178.655 ;
        RECT 79.950 178.875 80.415 179.265 ;
        RECT 80.585 179.135 80.980 179.305 ;
        RECT 78.090 178.305 78.260 178.485 ;
        RECT 74.890 177.595 75.960 177.765 ;
        RECT 76.130 177.385 76.320 177.825 ;
        RECT 76.490 177.555 77.440 177.835 ;
        RECT 77.750 177.745 78.010 178.135 ;
        RECT 78.430 178.065 79.220 178.315 ;
        RECT 77.660 177.575 78.010 177.745 ;
        RECT 78.220 177.385 78.550 177.845 ;
        RECT 79.425 177.775 79.595 178.485 ;
        RECT 79.950 178.285 80.120 178.875 ;
        RECT 79.765 178.065 80.120 178.285 ;
        RECT 80.290 178.065 80.640 178.685 ;
        RECT 80.810 177.775 80.980 179.135 ;
        RECT 81.345 178.965 81.670 179.750 ;
        RECT 81.150 177.915 81.610 178.965 ;
        RECT 79.425 177.605 80.280 177.775 ;
        RECT 80.485 177.605 80.980 177.775 ;
        RECT 81.150 177.385 81.480 177.745 ;
        RECT 81.840 177.645 82.010 179.765 ;
        RECT 82.180 179.435 82.510 179.935 ;
        RECT 82.680 179.265 82.935 179.765 ;
        RECT 82.185 179.095 82.935 179.265 ;
        RECT 82.185 178.105 82.415 179.095 ;
        RECT 82.585 178.275 82.935 178.925 ;
        RECT 83.110 178.845 84.320 179.935 ;
        RECT 83.110 178.305 83.630 178.845 ;
        RECT 84.550 178.795 84.760 179.935 ;
        RECT 84.930 178.785 85.260 179.765 ;
        RECT 85.430 178.795 85.660 179.935 ;
        RECT 83.800 178.135 84.320 178.675 ;
        RECT 82.185 177.935 82.935 178.105 ;
        RECT 82.180 177.385 82.510 177.765 ;
        RECT 82.680 177.645 82.935 177.935 ;
        RECT 83.110 177.385 84.320 178.135 ;
        RECT 84.550 177.385 84.760 178.205 ;
        RECT 84.930 178.185 85.180 178.785 ;
        RECT 86.330 178.770 86.620 179.935 ;
        RECT 86.830 178.795 87.060 179.935 ;
        RECT 87.230 178.785 87.560 179.765 ;
        RECT 87.730 178.795 87.940 179.935 ;
        RECT 88.260 179.005 88.430 179.765 ;
        RECT 88.610 179.175 88.940 179.935 ;
        RECT 88.260 178.835 88.925 179.005 ;
        RECT 89.110 178.860 89.380 179.765 ;
        RECT 85.350 178.375 85.680 178.625 ;
        RECT 86.810 178.375 87.140 178.625 ;
        RECT 84.930 177.555 85.260 178.185 ;
        RECT 85.430 177.385 85.660 178.205 ;
        RECT 86.330 177.385 86.620 178.110 ;
        RECT 86.830 177.385 87.060 178.205 ;
        RECT 87.310 178.185 87.560 178.785 ;
        RECT 88.755 178.690 88.925 178.835 ;
        RECT 88.190 178.285 88.520 178.655 ;
        RECT 88.755 178.360 89.040 178.690 ;
        RECT 87.230 177.555 87.560 178.185 ;
        RECT 87.730 177.385 87.940 178.205 ;
        RECT 88.755 178.105 88.925 178.360 ;
        RECT 88.260 177.935 88.925 178.105 ;
        RECT 89.210 178.060 89.380 178.860 ;
        RECT 90.470 179.175 90.985 179.585 ;
        RECT 91.220 179.175 91.390 179.935 ;
        RECT 91.560 179.595 93.590 179.765 ;
        RECT 90.470 178.365 90.810 179.175 ;
        RECT 91.560 178.930 91.730 179.595 ;
        RECT 92.125 179.255 93.250 179.425 ;
        RECT 90.980 178.740 91.730 178.930 ;
        RECT 91.900 178.915 92.910 179.085 ;
        RECT 90.470 178.195 91.700 178.365 ;
        RECT 88.260 177.555 88.430 177.935 ;
        RECT 88.610 177.385 88.940 177.765 ;
        RECT 89.120 177.555 89.380 178.060 ;
        RECT 90.745 177.590 90.990 178.195 ;
        RECT 91.210 177.385 91.720 177.920 ;
        RECT 91.900 177.555 92.090 178.915 ;
        RECT 92.260 177.895 92.535 178.715 ;
        RECT 92.740 178.115 92.910 178.915 ;
        RECT 93.080 178.125 93.250 179.255 ;
        RECT 93.420 178.625 93.590 179.595 ;
        RECT 93.760 178.795 93.930 179.935 ;
        RECT 94.100 178.795 94.435 179.765 ;
        RECT 95.130 178.795 95.340 179.935 ;
        RECT 93.420 178.295 93.615 178.625 ;
        RECT 93.840 178.295 94.095 178.625 ;
        RECT 93.840 178.125 94.010 178.295 ;
        RECT 94.265 178.125 94.435 178.795 ;
        RECT 95.510 178.785 95.840 179.765 ;
        RECT 96.010 178.795 96.240 179.935 ;
        RECT 96.915 179.500 102.260 179.935 ;
        RECT 93.080 177.955 94.010 178.125 ;
        RECT 93.080 177.920 93.255 177.955 ;
        RECT 92.260 177.725 92.540 177.895 ;
        RECT 92.260 177.555 92.535 177.725 ;
        RECT 92.725 177.555 93.255 177.920 ;
        RECT 93.680 177.385 94.010 177.785 ;
        RECT 94.180 177.555 94.435 178.125 ;
        RECT 95.130 177.385 95.340 178.205 ;
        RECT 95.510 178.185 95.760 178.785 ;
        RECT 95.930 178.375 96.260 178.625 ;
        RECT 98.505 178.250 98.855 179.500 ;
        RECT 102.470 178.795 102.700 179.935 ;
        RECT 102.870 178.785 103.200 179.765 ;
        RECT 103.370 178.795 103.580 179.935 ;
        RECT 103.810 178.845 105.480 179.935 ;
        RECT 105.740 179.005 105.910 179.765 ;
        RECT 106.090 179.175 106.420 179.935 ;
        RECT 95.510 177.555 95.840 178.185 ;
        RECT 96.010 177.385 96.240 178.205 ;
        RECT 100.335 177.930 100.675 178.760 ;
        RECT 102.450 178.375 102.780 178.625 ;
        RECT 96.915 177.385 102.260 177.930 ;
        RECT 102.470 177.385 102.700 178.205 ;
        RECT 102.950 178.185 103.200 178.785 ;
        RECT 103.810 178.325 104.560 178.845 ;
        RECT 105.740 178.835 106.405 179.005 ;
        RECT 106.590 178.860 106.860 179.765 ;
        RECT 106.235 178.690 106.405 178.835 ;
        RECT 102.870 177.555 103.200 178.185 ;
        RECT 103.370 177.385 103.580 178.205 ;
        RECT 104.730 178.155 105.480 178.675 ;
        RECT 105.670 178.285 106.000 178.655 ;
        RECT 106.235 178.360 106.520 178.690 ;
        RECT 103.810 177.385 105.480 178.155 ;
        RECT 106.235 178.105 106.405 178.360 ;
        RECT 105.740 177.935 106.405 178.105 ;
        RECT 106.690 178.060 106.860 178.860 ;
        RECT 107.490 178.845 111.000 179.935 ;
        RECT 111.170 178.845 112.380 179.935 ;
        RECT 107.490 178.325 109.180 178.845 ;
        RECT 109.350 178.155 111.000 178.675 ;
        RECT 111.170 178.305 111.690 178.845 ;
        RECT 105.740 177.555 105.910 177.935 ;
        RECT 106.090 177.385 106.420 177.765 ;
        RECT 106.600 177.555 106.860 178.060 ;
        RECT 107.490 177.385 111.000 178.155 ;
        RECT 111.860 178.135 112.380 178.675 ;
        RECT 111.170 177.385 112.380 178.135 ;
        RECT 18.165 177.215 112.465 177.385 ;
        RECT 18.250 176.465 19.460 177.215 ;
        RECT 18.250 175.925 18.770 176.465 ;
        RECT 20.090 176.445 21.760 177.215 ;
        RECT 21.930 176.490 22.220 177.215 ;
        RECT 22.390 176.445 24.060 177.215 ;
        RECT 18.940 175.755 19.460 176.295 ;
        RECT 18.250 174.665 19.460 175.755 ;
        RECT 20.090 175.755 20.840 176.275 ;
        RECT 21.010 175.925 21.760 176.445 ;
        RECT 20.090 174.665 21.760 175.755 ;
        RECT 21.930 174.665 22.220 175.830 ;
        RECT 22.390 175.755 23.140 176.275 ;
        RECT 23.310 175.925 24.060 176.445 ;
        RECT 24.505 176.405 24.750 177.010 ;
        RECT 24.970 176.680 25.480 177.215 ;
        RECT 24.230 176.235 25.460 176.405 ;
        RECT 22.390 174.665 24.060 175.755 ;
        RECT 24.230 175.425 24.570 176.235 ;
        RECT 24.740 175.670 25.490 175.860 ;
        RECT 24.230 175.015 24.745 175.425 ;
        RECT 24.980 174.665 25.150 175.425 ;
        RECT 25.320 175.005 25.490 175.670 ;
        RECT 25.660 175.685 25.850 177.045 ;
        RECT 26.020 176.875 26.295 177.045 ;
        RECT 26.020 176.705 26.300 176.875 ;
        RECT 26.020 175.885 26.295 176.705 ;
        RECT 26.485 176.680 27.015 177.045 ;
        RECT 27.440 176.815 27.770 177.215 ;
        RECT 26.840 176.645 27.015 176.680 ;
        RECT 26.500 175.685 26.670 176.485 ;
        RECT 25.660 175.515 26.670 175.685 ;
        RECT 26.840 176.475 27.770 176.645 ;
        RECT 27.940 176.475 28.195 177.045 ;
        RECT 28.745 176.875 29.000 177.035 ;
        RECT 28.660 176.705 29.000 176.875 ;
        RECT 29.180 176.755 29.465 177.215 ;
        RECT 26.840 175.345 27.010 176.475 ;
        RECT 27.600 176.305 27.770 176.475 ;
        RECT 25.885 175.175 27.010 175.345 ;
        RECT 27.180 175.975 27.375 176.305 ;
        RECT 27.600 175.975 27.855 176.305 ;
        RECT 27.180 175.005 27.350 175.975 ;
        RECT 28.025 175.805 28.195 176.475 ;
        RECT 25.320 174.835 27.350 175.005 ;
        RECT 27.520 174.665 27.690 175.805 ;
        RECT 27.860 174.835 28.195 175.805 ;
        RECT 28.745 176.505 29.000 176.705 ;
        RECT 28.745 175.645 28.925 176.505 ;
        RECT 29.645 176.305 29.895 176.955 ;
        RECT 29.095 175.975 29.895 176.305 ;
        RECT 28.745 174.975 29.000 175.645 ;
        RECT 29.180 174.665 29.465 175.465 ;
        RECT 29.645 175.385 29.895 175.975 ;
        RECT 30.095 176.620 30.415 176.950 ;
        RECT 30.595 176.735 31.255 177.215 ;
        RECT 31.455 176.825 32.305 176.995 ;
        RECT 30.095 175.725 30.285 176.620 ;
        RECT 30.605 176.295 31.265 176.565 ;
        RECT 30.935 176.235 31.265 176.295 ;
        RECT 30.455 176.065 30.785 176.125 ;
        RECT 31.455 176.065 31.625 176.825 ;
        RECT 32.865 176.755 33.185 177.215 ;
        RECT 33.385 176.575 33.635 177.005 ;
        RECT 33.925 176.775 34.335 177.215 ;
        RECT 34.505 176.835 35.520 177.035 ;
        RECT 31.795 176.405 33.045 176.575 ;
        RECT 31.795 176.285 32.125 176.405 ;
        RECT 30.455 175.895 32.355 176.065 ;
        RECT 30.095 175.555 32.015 175.725 ;
        RECT 30.095 175.535 30.415 175.555 ;
        RECT 29.645 174.875 29.975 175.385 ;
        RECT 30.245 174.925 30.415 175.535 ;
        RECT 32.185 175.385 32.355 175.895 ;
        RECT 32.525 175.825 32.705 176.235 ;
        RECT 32.875 175.645 33.045 176.405 ;
        RECT 30.585 174.665 30.915 175.355 ;
        RECT 31.145 175.215 32.355 175.385 ;
        RECT 32.525 175.335 33.045 175.645 ;
        RECT 33.215 176.235 33.635 176.575 ;
        RECT 33.925 176.235 34.335 176.565 ;
        RECT 33.215 175.465 33.405 176.235 ;
        RECT 34.505 176.105 34.675 176.835 ;
        RECT 35.820 176.665 35.990 176.995 ;
        RECT 36.160 176.835 36.490 177.215 ;
        RECT 34.845 176.285 35.195 176.655 ;
        RECT 34.505 176.065 34.925 176.105 ;
        RECT 33.575 175.895 34.925 176.065 ;
        RECT 33.575 175.735 33.825 175.895 ;
        RECT 34.335 175.465 34.585 175.725 ;
        RECT 33.215 175.215 34.585 175.465 ;
        RECT 31.145 174.925 31.385 175.215 ;
        RECT 32.185 175.135 32.355 175.215 ;
        RECT 31.585 174.665 32.005 175.045 ;
        RECT 32.185 174.885 32.815 175.135 ;
        RECT 33.285 174.665 33.615 175.045 ;
        RECT 33.785 174.925 33.955 175.215 ;
        RECT 34.755 175.050 34.925 175.895 ;
        RECT 35.375 175.725 35.595 176.595 ;
        RECT 35.820 176.475 36.515 176.665 ;
        RECT 35.095 175.345 35.595 175.725 ;
        RECT 35.765 175.675 36.175 176.295 ;
        RECT 36.345 175.505 36.515 176.475 ;
        RECT 35.820 175.335 36.515 175.505 ;
        RECT 34.135 174.665 34.515 175.045 ;
        RECT 34.755 174.880 35.585 175.050 ;
        RECT 35.820 174.835 35.990 175.335 ;
        RECT 36.160 174.665 36.490 175.165 ;
        RECT 36.705 174.835 36.930 176.955 ;
        RECT 37.100 176.835 37.430 177.215 ;
        RECT 37.600 176.665 37.770 176.955 ;
        RECT 37.105 176.495 37.770 176.665 ;
        RECT 38.120 176.665 38.290 176.955 ;
        RECT 38.460 176.835 38.790 177.215 ;
        RECT 38.120 176.495 38.785 176.665 ;
        RECT 37.105 175.505 37.335 176.495 ;
        RECT 37.505 175.675 37.855 176.325 ;
        RECT 38.035 175.675 38.385 176.325 ;
        RECT 38.555 175.505 38.785 176.495 ;
        RECT 37.105 175.335 37.770 175.505 ;
        RECT 37.100 174.665 37.430 175.165 ;
        RECT 37.600 174.835 37.770 175.335 ;
        RECT 38.120 175.335 38.785 175.505 ;
        RECT 38.120 174.835 38.290 175.335 ;
        RECT 38.460 174.665 38.790 175.165 ;
        RECT 38.960 174.835 39.185 176.955 ;
        RECT 39.400 176.835 39.730 177.215 ;
        RECT 39.900 176.665 40.070 176.995 ;
        RECT 40.370 176.835 41.385 177.035 ;
        RECT 39.375 176.475 40.070 176.665 ;
        RECT 39.375 175.505 39.545 176.475 ;
        RECT 39.715 175.675 40.125 176.295 ;
        RECT 40.295 175.725 40.515 176.595 ;
        RECT 40.695 176.285 41.045 176.655 ;
        RECT 41.215 176.105 41.385 176.835 ;
        RECT 41.555 176.775 41.965 177.215 ;
        RECT 42.255 176.575 42.505 177.005 ;
        RECT 42.705 176.755 43.025 177.215 ;
        RECT 43.585 176.825 44.435 176.995 ;
        RECT 41.555 176.235 41.965 176.565 ;
        RECT 42.255 176.235 42.675 176.575 ;
        RECT 40.965 176.065 41.385 176.105 ;
        RECT 40.965 175.895 42.315 176.065 ;
        RECT 39.375 175.335 40.070 175.505 ;
        RECT 40.295 175.345 40.795 175.725 ;
        RECT 39.400 174.665 39.730 175.165 ;
        RECT 39.900 174.835 40.070 175.335 ;
        RECT 40.965 175.050 41.135 175.895 ;
        RECT 42.065 175.735 42.315 175.895 ;
        RECT 41.305 175.465 41.555 175.725 ;
        RECT 42.485 175.465 42.675 176.235 ;
        RECT 41.305 175.215 42.675 175.465 ;
        RECT 42.845 176.405 44.095 176.575 ;
        RECT 42.845 175.645 43.015 176.405 ;
        RECT 43.765 176.285 44.095 176.405 ;
        RECT 43.185 175.825 43.365 176.235 ;
        RECT 44.265 176.065 44.435 176.825 ;
        RECT 44.635 176.735 45.295 177.215 ;
        RECT 45.475 176.620 45.795 176.950 ;
        RECT 44.625 176.295 45.285 176.565 ;
        RECT 44.625 176.235 44.955 176.295 ;
        RECT 45.105 176.065 45.435 176.125 ;
        RECT 43.535 175.895 45.435 176.065 ;
        RECT 42.845 175.335 43.365 175.645 ;
        RECT 43.535 175.385 43.705 175.895 ;
        RECT 45.605 175.725 45.795 176.620 ;
        RECT 43.875 175.555 45.795 175.725 ;
        RECT 45.475 175.535 45.795 175.555 ;
        RECT 45.995 176.305 46.245 176.955 ;
        RECT 46.425 176.755 46.710 177.215 ;
        RECT 46.890 176.875 47.145 177.035 ;
        RECT 46.890 176.705 47.230 176.875 ;
        RECT 46.890 176.505 47.145 176.705 ;
        RECT 45.995 175.975 46.795 176.305 ;
        RECT 43.535 175.215 44.745 175.385 ;
        RECT 40.305 174.880 41.135 175.050 ;
        RECT 41.375 174.665 41.755 175.045 ;
        RECT 41.935 174.925 42.105 175.215 ;
        RECT 43.535 175.135 43.705 175.215 ;
        RECT 42.275 174.665 42.605 175.045 ;
        RECT 43.075 174.885 43.705 175.135 ;
        RECT 43.885 174.665 44.305 175.045 ;
        RECT 44.505 174.925 44.745 175.215 ;
        RECT 44.975 174.665 45.305 175.355 ;
        RECT 45.475 174.925 45.645 175.535 ;
        RECT 45.995 175.385 46.245 175.975 ;
        RECT 46.965 175.645 47.145 176.505 ;
        RECT 47.690 176.490 47.980 177.215 ;
        RECT 48.425 176.405 48.670 177.010 ;
        RECT 48.890 176.680 49.400 177.215 ;
        RECT 48.150 176.235 49.380 176.405 ;
        RECT 45.915 174.875 46.245 175.385 ;
        RECT 46.425 174.665 46.710 175.465 ;
        RECT 46.890 174.975 47.145 175.645 ;
        RECT 47.690 174.665 47.980 175.830 ;
        RECT 48.150 175.425 48.490 176.235 ;
        RECT 48.660 175.670 49.410 175.860 ;
        RECT 48.150 175.015 48.665 175.425 ;
        RECT 48.900 174.665 49.070 175.425 ;
        RECT 49.240 175.005 49.410 175.670 ;
        RECT 49.580 175.685 49.770 177.045 ;
        RECT 49.940 176.535 50.215 177.045 ;
        RECT 50.405 176.680 50.935 177.045 ;
        RECT 51.360 176.815 51.690 177.215 ;
        RECT 50.760 176.645 50.935 176.680 ;
        RECT 49.940 176.365 50.220 176.535 ;
        RECT 49.940 175.885 50.215 176.365 ;
        RECT 50.420 175.685 50.590 176.485 ;
        RECT 49.580 175.515 50.590 175.685 ;
        RECT 50.760 176.475 51.690 176.645 ;
        RECT 51.860 176.475 52.115 177.045 ;
        RECT 52.380 176.665 52.550 177.045 ;
        RECT 52.730 176.835 53.060 177.215 ;
        RECT 52.380 176.495 53.045 176.665 ;
        RECT 53.240 176.540 53.500 177.045 ;
        RECT 50.760 175.345 50.930 176.475 ;
        RECT 51.520 176.305 51.690 176.475 ;
        RECT 49.805 175.175 50.930 175.345 ;
        RECT 51.100 175.975 51.295 176.305 ;
        RECT 51.520 175.975 51.775 176.305 ;
        RECT 51.100 175.005 51.270 175.975 ;
        RECT 51.945 175.805 52.115 176.475 ;
        RECT 52.310 175.945 52.640 176.315 ;
        RECT 52.875 176.240 53.045 176.495 ;
        RECT 49.240 174.835 51.270 175.005 ;
        RECT 51.440 174.665 51.610 175.805 ;
        RECT 51.780 174.835 52.115 175.805 ;
        RECT 52.875 175.910 53.160 176.240 ;
        RECT 52.875 175.765 53.045 175.910 ;
        RECT 52.380 175.595 53.045 175.765 ;
        RECT 53.330 175.740 53.500 176.540 ;
        RECT 53.670 176.445 57.180 177.215 ;
        RECT 52.380 174.835 52.550 175.595 ;
        RECT 52.730 174.665 53.060 175.425 ;
        RECT 53.230 174.835 53.500 175.740 ;
        RECT 53.670 175.755 55.360 176.275 ;
        RECT 55.530 175.925 57.180 176.445 ;
        RECT 57.355 176.375 57.615 177.215 ;
        RECT 57.790 176.470 58.045 177.045 ;
        RECT 58.215 176.835 58.545 177.215 ;
        RECT 58.760 176.665 58.930 177.045 ;
        RECT 58.215 176.495 58.930 176.665 ;
        RECT 59.190 176.715 59.450 177.045 ;
        RECT 59.760 176.835 60.090 177.215 ;
        RECT 60.270 176.875 61.750 177.045 ;
        RECT 53.670 174.665 57.180 175.755 ;
        RECT 57.355 174.665 57.615 175.815 ;
        RECT 57.790 175.740 57.960 176.470 ;
        RECT 58.215 176.305 58.385 176.495 ;
        RECT 58.130 175.975 58.385 176.305 ;
        RECT 58.215 175.765 58.385 175.975 ;
        RECT 58.665 175.945 59.020 176.315 ;
        RECT 59.190 176.015 59.360 176.715 ;
        RECT 60.270 176.545 60.670 176.875 ;
        RECT 59.710 176.355 59.920 176.535 ;
        RECT 59.710 176.185 60.330 176.355 ;
        RECT 60.500 176.065 60.670 176.545 ;
        RECT 60.860 176.375 61.410 176.705 ;
        RECT 59.190 175.845 60.320 176.015 ;
        RECT 60.500 175.895 61.070 176.065 ;
        RECT 57.790 174.835 58.045 175.740 ;
        RECT 58.215 175.595 58.930 175.765 ;
        RECT 58.215 174.665 58.545 175.425 ;
        RECT 58.760 174.835 58.930 175.595 ;
        RECT 59.190 175.165 59.360 175.845 ;
        RECT 60.150 175.725 60.320 175.845 ;
        RECT 59.530 175.345 59.880 175.675 ;
        RECT 60.150 175.555 60.730 175.725 ;
        RECT 60.900 175.385 61.070 175.895 ;
        RECT 60.330 175.215 61.070 175.385 ;
        RECT 61.240 175.385 61.410 176.375 ;
        RECT 61.580 175.975 61.750 176.875 ;
        RECT 62.000 176.305 62.185 176.885 ;
        RECT 62.455 176.305 62.650 176.880 ;
        RECT 62.860 176.835 63.190 177.215 ;
        RECT 62.000 175.975 62.230 176.305 ;
        RECT 62.455 175.975 62.710 176.305 ;
        RECT 62.000 175.665 62.185 175.975 ;
        RECT 62.455 175.665 62.650 175.975 ;
        RECT 63.020 175.385 63.190 176.305 ;
        RECT 61.240 175.215 63.190 175.385 ;
        RECT 59.190 174.835 59.450 175.165 ;
        RECT 59.760 174.665 60.090 175.045 ;
        RECT 60.330 174.835 60.520 175.215 ;
        RECT 60.770 174.665 61.100 175.045 ;
        RECT 61.310 174.835 61.480 175.215 ;
        RECT 61.675 174.665 62.005 175.045 ;
        RECT 62.265 174.835 62.435 175.215 ;
        RECT 62.860 174.665 63.190 175.045 ;
        RECT 63.360 174.835 63.620 177.045 ;
        RECT 63.795 176.505 64.050 177.035 ;
        RECT 64.220 176.755 64.525 177.215 ;
        RECT 64.770 176.835 65.840 177.005 ;
        RECT 63.795 175.855 64.005 176.505 ;
        RECT 64.770 176.480 65.090 176.835 ;
        RECT 64.765 176.305 65.090 176.480 ;
        RECT 64.175 176.005 65.090 176.305 ;
        RECT 65.260 176.265 65.500 176.665 ;
        RECT 65.670 176.605 65.840 176.835 ;
        RECT 66.010 176.775 66.200 177.215 ;
        RECT 66.370 176.765 67.320 177.045 ;
        RECT 67.540 176.855 67.890 177.025 ;
        RECT 65.670 176.435 66.200 176.605 ;
        RECT 64.175 175.975 64.915 176.005 ;
        RECT 63.795 174.975 64.050 175.855 ;
        RECT 64.220 174.665 64.525 175.805 ;
        RECT 64.745 175.385 64.915 175.975 ;
        RECT 65.260 175.895 65.800 176.265 ;
        RECT 65.980 176.155 66.200 176.435 ;
        RECT 66.370 175.985 66.540 176.765 ;
        RECT 66.135 175.815 66.540 175.985 ;
        RECT 66.710 175.975 67.060 176.595 ;
        RECT 66.135 175.725 66.305 175.815 ;
        RECT 67.230 175.805 67.440 176.595 ;
        RECT 65.085 175.555 66.305 175.725 ;
        RECT 66.765 175.645 67.440 175.805 ;
        RECT 64.745 175.215 65.545 175.385 ;
        RECT 64.865 174.665 65.195 175.045 ;
        RECT 65.375 174.925 65.545 175.215 ;
        RECT 66.135 175.175 66.305 175.555 ;
        RECT 66.475 175.635 67.440 175.645 ;
        RECT 67.630 176.465 67.890 176.855 ;
        RECT 68.100 176.755 68.430 177.215 ;
        RECT 69.305 176.825 70.160 176.995 ;
        RECT 70.365 176.825 70.860 176.995 ;
        RECT 71.030 176.855 71.360 177.215 ;
        RECT 67.630 175.775 67.800 176.465 ;
        RECT 67.970 176.115 68.140 176.295 ;
        RECT 68.310 176.285 69.100 176.535 ;
        RECT 69.305 176.115 69.475 176.825 ;
        RECT 69.645 176.315 70.000 176.535 ;
        RECT 67.970 175.945 69.660 176.115 ;
        RECT 66.475 175.345 66.935 175.635 ;
        RECT 67.630 175.605 69.130 175.775 ;
        RECT 67.630 175.465 67.800 175.605 ;
        RECT 67.240 175.295 67.800 175.465 ;
        RECT 65.715 174.665 65.965 175.125 ;
        RECT 66.135 174.835 67.005 175.175 ;
        RECT 67.240 174.835 67.410 175.295 ;
        RECT 68.245 175.265 69.320 175.435 ;
        RECT 67.580 174.665 67.950 175.125 ;
        RECT 68.245 174.925 68.415 175.265 ;
        RECT 68.585 174.665 68.915 175.095 ;
        RECT 69.150 174.925 69.320 175.265 ;
        RECT 69.490 175.165 69.660 175.945 ;
        RECT 69.830 175.725 70.000 176.315 ;
        RECT 70.170 175.915 70.520 176.535 ;
        RECT 69.830 175.335 70.295 175.725 ;
        RECT 70.690 175.465 70.860 176.825 ;
        RECT 71.030 175.635 71.490 176.685 ;
        RECT 70.465 175.295 70.860 175.465 ;
        RECT 70.465 175.165 70.635 175.295 ;
        RECT 69.490 174.835 70.170 175.165 ;
        RECT 70.385 174.835 70.635 175.165 ;
        RECT 70.805 174.665 71.055 175.125 ;
        RECT 71.225 174.850 71.550 175.635 ;
        RECT 71.720 174.835 71.890 176.955 ;
        RECT 72.060 176.835 72.390 177.215 ;
        RECT 72.560 176.665 72.815 176.955 ;
        RECT 72.065 176.495 72.815 176.665 ;
        RECT 72.065 175.505 72.295 176.495 ;
        RECT 73.450 176.490 73.740 177.215 ;
        RECT 74.375 176.670 79.720 177.215 ;
        RECT 72.465 175.675 72.815 176.325 ;
        RECT 72.065 175.335 72.815 175.505 ;
        RECT 72.060 174.665 72.390 175.165 ;
        RECT 72.560 174.835 72.815 175.335 ;
        RECT 73.450 174.665 73.740 175.830 ;
        RECT 75.965 175.100 76.315 176.350 ;
        RECT 77.795 175.840 78.135 176.670 ;
        RECT 79.980 176.665 80.150 177.045 ;
        RECT 80.330 176.835 80.660 177.215 ;
        RECT 79.980 176.495 80.645 176.665 ;
        RECT 80.840 176.540 81.100 177.045 ;
        RECT 79.910 175.945 80.240 176.315 ;
        RECT 80.475 176.240 80.645 176.495 ;
        RECT 80.475 175.910 80.760 176.240 ;
        RECT 80.475 175.765 80.645 175.910 ;
        RECT 79.980 175.595 80.645 175.765 ;
        RECT 80.930 175.740 81.100 176.540 ;
        RECT 74.375 174.665 79.720 175.100 ;
        RECT 79.980 174.835 80.150 175.595 ;
        RECT 80.330 174.665 80.660 175.425 ;
        RECT 80.830 174.835 81.100 175.740 ;
        RECT 81.735 176.505 81.990 177.035 ;
        RECT 82.160 176.755 82.465 177.215 ;
        RECT 82.710 176.835 83.780 177.005 ;
        RECT 81.735 175.855 81.945 176.505 ;
        RECT 82.710 176.480 83.030 176.835 ;
        RECT 82.705 176.305 83.030 176.480 ;
        RECT 82.115 176.005 83.030 176.305 ;
        RECT 83.200 176.265 83.440 176.665 ;
        RECT 83.610 176.605 83.780 176.835 ;
        RECT 83.950 176.775 84.140 177.215 ;
        RECT 84.310 176.765 85.260 177.045 ;
        RECT 85.480 176.855 85.830 177.025 ;
        RECT 83.610 176.435 84.140 176.605 ;
        RECT 82.115 175.975 82.855 176.005 ;
        RECT 81.735 174.975 81.990 175.855 ;
        RECT 82.160 174.665 82.465 175.805 ;
        RECT 82.685 175.385 82.855 175.975 ;
        RECT 83.200 175.895 83.740 176.265 ;
        RECT 83.920 176.155 84.140 176.435 ;
        RECT 84.310 175.985 84.480 176.765 ;
        RECT 84.075 175.815 84.480 175.985 ;
        RECT 84.650 175.975 85.000 176.595 ;
        RECT 84.075 175.725 84.245 175.815 ;
        RECT 85.170 175.805 85.380 176.595 ;
        RECT 83.025 175.555 84.245 175.725 ;
        RECT 84.705 175.645 85.380 175.805 ;
        RECT 82.685 175.215 83.485 175.385 ;
        RECT 82.805 174.665 83.135 175.045 ;
        RECT 83.315 174.925 83.485 175.215 ;
        RECT 84.075 175.175 84.245 175.555 ;
        RECT 84.415 175.635 85.380 175.645 ;
        RECT 85.570 176.465 85.830 176.855 ;
        RECT 86.040 176.755 86.370 177.215 ;
        RECT 87.245 176.825 88.100 176.995 ;
        RECT 88.305 176.825 88.800 176.995 ;
        RECT 88.970 176.855 89.300 177.215 ;
        RECT 85.570 175.775 85.740 176.465 ;
        RECT 85.910 176.115 86.080 176.295 ;
        RECT 86.250 176.285 87.040 176.535 ;
        RECT 87.245 176.115 87.415 176.825 ;
        RECT 87.585 176.315 87.940 176.535 ;
        RECT 85.910 175.945 87.600 176.115 ;
        RECT 84.415 175.345 84.875 175.635 ;
        RECT 85.570 175.605 87.070 175.775 ;
        RECT 85.570 175.465 85.740 175.605 ;
        RECT 85.180 175.295 85.740 175.465 ;
        RECT 83.655 174.665 83.905 175.125 ;
        RECT 84.075 174.835 84.945 175.175 ;
        RECT 85.180 174.835 85.350 175.295 ;
        RECT 86.185 175.265 87.260 175.435 ;
        RECT 85.520 174.665 85.890 175.125 ;
        RECT 86.185 174.925 86.355 175.265 ;
        RECT 86.525 174.665 86.855 175.095 ;
        RECT 87.090 174.925 87.260 175.265 ;
        RECT 87.430 175.165 87.600 175.945 ;
        RECT 87.770 175.725 87.940 176.315 ;
        RECT 88.110 175.915 88.460 176.535 ;
        RECT 87.770 175.335 88.235 175.725 ;
        RECT 88.630 175.465 88.800 176.825 ;
        RECT 88.970 175.635 89.430 176.685 ;
        RECT 88.405 175.295 88.800 175.465 ;
        RECT 88.405 175.165 88.575 175.295 ;
        RECT 87.430 174.835 88.110 175.165 ;
        RECT 88.325 174.835 88.575 175.165 ;
        RECT 88.745 174.665 88.995 175.125 ;
        RECT 89.165 174.850 89.490 175.635 ;
        RECT 89.660 174.835 89.830 176.955 ;
        RECT 90.000 176.835 90.330 177.215 ;
        RECT 90.500 176.665 90.755 176.955 ;
        RECT 90.005 176.495 90.755 176.665 ;
        RECT 90.005 175.505 90.235 176.495 ;
        RECT 90.930 176.465 92.140 177.215 ;
        RECT 92.315 176.670 97.660 177.215 ;
        RECT 90.405 175.675 90.755 176.325 ;
        RECT 90.930 175.755 91.450 176.295 ;
        RECT 91.620 175.925 92.140 176.465 ;
        RECT 90.005 175.335 90.755 175.505 ;
        RECT 90.000 174.665 90.330 175.165 ;
        RECT 90.500 174.835 90.755 175.335 ;
        RECT 90.930 174.665 92.140 175.755 ;
        RECT 93.905 175.100 94.255 176.350 ;
        RECT 95.735 175.840 96.075 176.670 ;
        RECT 97.870 176.395 98.100 177.215 ;
        RECT 98.270 176.415 98.600 177.045 ;
        RECT 97.850 175.975 98.180 176.225 ;
        RECT 98.350 175.815 98.600 176.415 ;
        RECT 98.770 176.395 98.980 177.215 ;
        RECT 99.210 176.490 99.500 177.215 ;
        RECT 100.135 176.505 100.390 177.035 ;
        RECT 100.560 176.755 100.865 177.215 ;
        RECT 101.110 176.835 102.180 177.005 ;
        RECT 100.135 175.855 100.345 176.505 ;
        RECT 101.110 176.480 101.430 176.835 ;
        RECT 101.105 176.305 101.430 176.480 ;
        RECT 100.515 176.005 101.430 176.305 ;
        RECT 101.600 176.265 101.840 176.665 ;
        RECT 102.010 176.605 102.180 176.835 ;
        RECT 102.350 176.775 102.540 177.215 ;
        RECT 102.710 176.765 103.660 177.045 ;
        RECT 103.880 176.855 104.230 177.025 ;
        RECT 102.010 176.435 102.540 176.605 ;
        RECT 100.515 175.975 101.255 176.005 ;
        RECT 92.315 174.665 97.660 175.100 ;
        RECT 97.870 174.665 98.100 175.805 ;
        RECT 98.270 174.835 98.600 175.815 ;
        RECT 98.770 174.665 98.980 175.805 ;
        RECT 99.210 174.665 99.500 175.830 ;
        RECT 100.135 174.975 100.390 175.855 ;
        RECT 100.560 174.665 100.865 175.805 ;
        RECT 101.085 175.385 101.255 175.975 ;
        RECT 101.600 175.895 102.140 176.265 ;
        RECT 102.320 176.155 102.540 176.435 ;
        RECT 102.710 175.985 102.880 176.765 ;
        RECT 102.475 175.815 102.880 175.985 ;
        RECT 103.050 175.975 103.400 176.595 ;
        RECT 102.475 175.725 102.645 175.815 ;
        RECT 103.570 175.805 103.780 176.595 ;
        RECT 101.425 175.555 102.645 175.725 ;
        RECT 103.105 175.645 103.780 175.805 ;
        RECT 101.085 175.215 101.885 175.385 ;
        RECT 101.205 174.665 101.535 175.045 ;
        RECT 101.715 174.925 101.885 175.215 ;
        RECT 102.475 175.175 102.645 175.555 ;
        RECT 102.815 175.635 103.780 175.645 ;
        RECT 103.970 176.465 104.230 176.855 ;
        RECT 104.440 176.755 104.770 177.215 ;
        RECT 105.645 176.825 106.500 176.995 ;
        RECT 106.705 176.825 107.200 176.995 ;
        RECT 107.370 176.855 107.700 177.215 ;
        RECT 103.970 175.775 104.140 176.465 ;
        RECT 104.310 176.115 104.480 176.295 ;
        RECT 104.650 176.285 105.440 176.535 ;
        RECT 105.645 176.115 105.815 176.825 ;
        RECT 105.985 176.315 106.340 176.535 ;
        RECT 104.310 175.945 106.000 176.115 ;
        RECT 102.815 175.345 103.275 175.635 ;
        RECT 103.970 175.605 105.470 175.775 ;
        RECT 103.970 175.465 104.140 175.605 ;
        RECT 103.580 175.295 104.140 175.465 ;
        RECT 102.055 174.665 102.305 175.125 ;
        RECT 102.475 174.835 103.345 175.175 ;
        RECT 103.580 174.835 103.750 175.295 ;
        RECT 104.585 175.265 105.660 175.435 ;
        RECT 103.920 174.665 104.290 175.125 ;
        RECT 104.585 174.925 104.755 175.265 ;
        RECT 104.925 174.665 105.255 175.095 ;
        RECT 105.490 174.925 105.660 175.265 ;
        RECT 105.830 175.165 106.000 175.945 ;
        RECT 106.170 175.725 106.340 176.315 ;
        RECT 106.510 175.915 106.860 176.535 ;
        RECT 106.170 175.335 106.635 175.725 ;
        RECT 107.030 175.465 107.200 176.825 ;
        RECT 107.370 175.635 107.830 176.685 ;
        RECT 106.805 175.295 107.200 175.465 ;
        RECT 106.805 175.165 106.975 175.295 ;
        RECT 105.830 174.835 106.510 175.165 ;
        RECT 106.725 174.835 106.975 175.165 ;
        RECT 107.145 174.665 107.395 175.125 ;
        RECT 107.565 174.850 107.890 175.635 ;
        RECT 108.060 174.835 108.230 176.955 ;
        RECT 108.400 176.835 108.730 177.215 ;
        RECT 108.900 176.665 109.155 176.955 ;
        RECT 108.405 176.495 109.155 176.665 ;
        RECT 108.405 175.505 108.635 176.495 ;
        RECT 109.330 176.445 111.000 177.215 ;
        RECT 111.170 176.465 112.380 177.215 ;
        RECT 108.805 175.675 109.155 176.325 ;
        RECT 109.330 175.755 110.080 176.275 ;
        RECT 110.250 175.925 111.000 176.445 ;
        RECT 111.170 175.755 111.690 176.295 ;
        RECT 111.860 175.925 112.380 176.465 ;
        RECT 108.405 175.335 109.155 175.505 ;
        RECT 108.400 174.665 108.730 175.165 ;
        RECT 108.900 174.835 109.155 175.335 ;
        RECT 109.330 174.665 111.000 175.755 ;
        RECT 111.170 174.665 112.380 175.755 ;
        RECT 18.165 174.495 112.465 174.665 ;
        RECT 18.250 173.405 19.460 174.495 ;
        RECT 18.250 172.695 18.770 173.235 ;
        RECT 18.940 172.865 19.460 173.405 ;
        RECT 20.090 173.405 22.680 174.495 ;
        RECT 22.965 173.865 23.250 174.325 ;
        RECT 23.420 174.035 23.690 174.495 ;
        RECT 22.965 173.645 23.920 173.865 ;
        RECT 20.090 172.885 21.300 173.405 ;
        RECT 21.470 172.715 22.680 173.235 ;
        RECT 22.850 172.915 23.540 173.475 ;
        RECT 23.710 172.745 23.920 173.645 ;
        RECT 18.250 171.945 19.460 172.695 ;
        RECT 20.090 171.945 22.680 172.715 ;
        RECT 22.965 172.575 23.920 172.745 ;
        RECT 24.090 173.475 24.490 174.325 ;
        RECT 24.680 173.865 24.960 174.325 ;
        RECT 25.480 174.035 25.805 174.495 ;
        RECT 24.680 173.645 25.805 173.865 ;
        RECT 24.090 172.915 25.185 173.475 ;
        RECT 25.355 173.185 25.805 173.645 ;
        RECT 25.975 173.355 26.360 174.325 ;
        RECT 22.965 172.115 23.250 172.575 ;
        RECT 23.420 171.945 23.690 172.405 ;
        RECT 24.090 172.115 24.490 172.915 ;
        RECT 25.355 172.855 25.910 173.185 ;
        RECT 25.355 172.745 25.805 172.855 ;
        RECT 24.680 172.575 25.805 172.745 ;
        RECT 26.080 172.685 26.360 173.355 ;
        RECT 26.990 173.405 30.500 174.495 ;
        RECT 30.670 173.735 31.185 174.145 ;
        RECT 31.420 173.735 31.590 174.495 ;
        RECT 31.760 174.155 33.790 174.325 ;
        RECT 26.990 172.885 28.680 173.405 ;
        RECT 28.850 172.715 30.500 173.235 ;
        RECT 30.670 172.925 31.010 173.735 ;
        RECT 31.760 173.490 31.930 174.155 ;
        RECT 32.325 173.815 33.450 173.985 ;
        RECT 31.180 173.300 31.930 173.490 ;
        RECT 32.100 173.475 33.110 173.645 ;
        RECT 30.670 172.755 31.900 172.925 ;
        RECT 24.680 172.115 24.960 172.575 ;
        RECT 25.480 171.945 25.805 172.405 ;
        RECT 25.975 172.115 26.360 172.685 ;
        RECT 26.990 171.945 30.500 172.715 ;
        RECT 30.945 172.150 31.190 172.755 ;
        RECT 31.410 171.945 31.920 172.480 ;
        RECT 32.100 172.115 32.290 173.475 ;
        RECT 32.460 172.455 32.735 173.275 ;
        RECT 32.940 172.675 33.110 173.475 ;
        RECT 33.280 172.685 33.450 173.815 ;
        RECT 33.620 173.185 33.790 174.155 ;
        RECT 33.960 173.355 34.130 174.495 ;
        RECT 34.300 173.355 34.635 174.325 ;
        RECT 33.620 172.855 33.815 173.185 ;
        RECT 34.040 172.855 34.295 173.185 ;
        RECT 34.040 172.685 34.210 172.855 ;
        RECT 34.465 172.685 34.635 173.355 ;
        RECT 34.810 173.330 35.100 174.495 ;
        RECT 35.730 173.405 38.320 174.495 ;
        RECT 35.730 172.885 36.940 173.405 ;
        RECT 38.550 173.355 38.760 174.495 ;
        RECT 38.930 173.345 39.260 174.325 ;
        RECT 39.430 173.355 39.660 174.495 ;
        RECT 40.790 173.405 44.300 174.495 ;
        RECT 44.470 173.420 44.740 174.325 ;
        RECT 44.910 173.735 45.240 174.495 ;
        RECT 45.420 173.565 45.590 174.325 ;
        RECT 37.110 172.715 38.320 173.235 ;
        RECT 33.280 172.515 34.210 172.685 ;
        RECT 33.280 172.480 33.455 172.515 ;
        RECT 32.460 172.285 32.740 172.455 ;
        RECT 32.460 172.115 32.735 172.285 ;
        RECT 32.925 172.115 33.455 172.480 ;
        RECT 33.880 171.945 34.210 172.345 ;
        RECT 34.380 172.115 34.635 172.685 ;
        RECT 34.810 171.945 35.100 172.670 ;
        RECT 35.730 171.945 38.320 172.715 ;
        RECT 38.550 171.945 38.760 172.765 ;
        RECT 38.930 172.745 39.180 173.345 ;
        RECT 39.350 172.935 39.680 173.185 ;
        RECT 40.790 172.885 42.480 173.405 ;
        RECT 38.930 172.115 39.260 172.745 ;
        RECT 39.430 171.945 39.660 172.765 ;
        RECT 42.650 172.715 44.300 173.235 ;
        RECT 40.790 171.945 44.300 172.715 ;
        RECT 44.470 172.620 44.640 173.420 ;
        RECT 44.925 173.395 45.590 173.565 ;
        RECT 44.925 173.250 45.095 173.395 ;
        RECT 44.810 172.920 45.095 173.250 ;
        RECT 45.855 173.355 46.190 174.325 ;
        RECT 46.360 173.355 46.530 174.495 ;
        RECT 46.700 174.155 48.730 174.325 ;
        RECT 44.925 172.665 45.095 172.920 ;
        RECT 45.330 172.845 45.660 173.215 ;
        RECT 45.855 172.685 46.025 173.355 ;
        RECT 46.700 173.185 46.870 174.155 ;
        RECT 46.195 172.855 46.450 173.185 ;
        RECT 46.675 172.855 46.870 173.185 ;
        RECT 47.040 173.815 48.165 173.985 ;
        RECT 46.280 172.685 46.450 172.855 ;
        RECT 47.040 172.685 47.210 173.815 ;
        RECT 44.470 172.115 44.730 172.620 ;
        RECT 44.925 172.495 45.590 172.665 ;
        RECT 44.910 171.945 45.240 172.325 ;
        RECT 45.420 172.115 45.590 172.495 ;
        RECT 45.855 172.115 46.110 172.685 ;
        RECT 46.280 172.515 47.210 172.685 ;
        RECT 47.380 173.475 48.390 173.645 ;
        RECT 47.380 172.675 47.550 173.475 ;
        RECT 47.755 173.135 48.030 173.275 ;
        RECT 47.750 172.965 48.030 173.135 ;
        RECT 47.035 172.480 47.210 172.515 ;
        RECT 46.280 171.945 46.610 172.345 ;
        RECT 47.035 172.115 47.565 172.480 ;
        RECT 47.755 172.115 48.030 172.965 ;
        RECT 48.200 172.115 48.390 173.475 ;
        RECT 48.560 173.490 48.730 174.155 ;
        RECT 48.900 173.735 49.070 174.495 ;
        RECT 49.305 173.735 49.820 174.145 ;
        RECT 48.560 173.300 49.310 173.490 ;
        RECT 49.480 172.925 49.820 173.735 ;
        RECT 50.050 173.355 50.260 174.495 ;
        RECT 48.590 172.755 49.820 172.925 ;
        RECT 50.430 173.345 50.760 174.325 ;
        RECT 50.930 173.355 51.160 174.495 ;
        RECT 51.370 173.405 54.880 174.495 ;
        RECT 55.055 174.060 60.400 174.495 ;
        RECT 48.570 171.945 49.080 172.480 ;
        RECT 49.300 172.150 49.545 172.755 ;
        RECT 50.050 171.945 50.260 172.765 ;
        RECT 50.430 172.745 50.680 173.345 ;
        RECT 50.850 172.935 51.180 173.185 ;
        RECT 51.370 172.885 53.060 173.405 ;
        RECT 50.430 172.115 50.760 172.745 ;
        RECT 50.930 171.945 51.160 172.765 ;
        RECT 53.230 172.715 54.880 173.235 ;
        RECT 56.645 172.810 56.995 174.060 ;
        RECT 60.570 173.330 60.860 174.495 ;
        RECT 61.740 174.045 62.070 174.495 ;
        RECT 61.030 173.655 63.640 173.865 ;
        RECT 51.370 171.945 54.880 172.715 ;
        RECT 58.475 172.490 58.815 173.320 ;
        RECT 61.030 172.685 61.200 173.655 ;
        RECT 61.370 172.855 61.720 173.475 ;
        RECT 61.890 172.855 62.210 173.475 ;
        RECT 62.380 172.855 62.710 173.475 ;
        RECT 62.880 172.855 63.180 173.475 ;
        RECT 63.420 172.855 63.640 173.655 ;
        RECT 63.820 172.685 64.080 174.310 ;
        RECT 64.250 173.405 66.840 174.495 ;
        RECT 67.010 173.525 67.320 174.325 ;
        RECT 67.490 173.695 67.800 174.495 ;
        RECT 67.970 173.865 68.230 174.325 ;
        RECT 68.400 174.035 68.655 174.495 ;
        RECT 68.830 173.865 69.090 174.325 ;
        RECT 67.970 173.695 69.090 173.865 ;
        RECT 64.250 172.885 65.460 173.405 ;
        RECT 67.010 173.355 68.040 173.525 ;
        RECT 65.630 172.715 66.840 173.235 ;
        RECT 55.055 171.945 60.400 172.490 ;
        RECT 60.570 171.945 60.860 172.670 ;
        RECT 61.030 172.515 61.505 172.685 ;
        RECT 61.335 172.265 61.505 172.515 ;
        RECT 61.740 171.945 62.070 172.685 ;
        RECT 62.240 172.515 64.080 172.685 ;
        RECT 62.240 172.170 62.440 172.515 ;
        RECT 62.610 171.945 62.940 172.345 ;
        RECT 63.110 172.160 63.310 172.515 ;
        RECT 63.480 171.945 63.810 172.340 ;
        RECT 64.250 171.945 66.840 172.715 ;
        RECT 67.010 172.445 67.180 173.355 ;
        RECT 67.350 172.615 67.700 173.185 ;
        RECT 67.870 173.105 68.040 173.355 ;
        RECT 68.830 173.445 69.090 173.695 ;
        RECT 69.260 173.625 69.545 174.495 ;
        RECT 69.770 173.525 70.080 174.325 ;
        RECT 70.250 173.695 70.560 174.495 ;
        RECT 70.730 173.865 70.990 174.325 ;
        RECT 71.160 174.035 71.415 174.495 ;
        RECT 71.590 173.865 71.850 174.325 ;
        RECT 70.730 173.695 71.850 173.865 ;
        RECT 68.830 173.275 69.585 173.445 ;
        RECT 67.870 172.935 69.010 173.105 ;
        RECT 69.180 172.765 69.585 173.275 ;
        RECT 67.935 172.595 69.585 172.765 ;
        RECT 69.770 173.355 70.800 173.525 ;
        RECT 67.010 172.115 67.310 172.445 ;
        RECT 67.480 171.945 67.755 172.425 ;
        RECT 67.935 172.205 68.230 172.595 ;
        RECT 68.400 171.945 68.655 172.425 ;
        RECT 68.830 172.205 69.090 172.595 ;
        RECT 69.770 172.445 69.940 173.355 ;
        RECT 70.110 172.615 70.460 173.185 ;
        RECT 70.630 173.105 70.800 173.355 ;
        RECT 71.590 173.445 71.850 173.695 ;
        RECT 72.020 173.625 72.305 174.495 ;
        RECT 73.000 173.515 73.330 174.325 ;
        RECT 73.500 173.695 73.740 174.495 ;
        RECT 71.590 173.275 72.345 173.445 ;
        RECT 73.000 173.345 73.715 173.515 ;
        RECT 70.630 172.935 71.770 173.105 ;
        RECT 71.940 172.765 72.345 173.275 ;
        RECT 72.995 172.935 73.375 173.175 ;
        RECT 73.545 173.105 73.715 173.345 ;
        RECT 73.920 173.475 74.090 174.325 ;
        RECT 74.260 173.695 74.590 174.495 ;
        RECT 74.760 173.475 74.930 174.325 ;
        RECT 73.920 173.305 74.930 173.475 ;
        RECT 75.100 173.345 75.430 174.495 ;
        RECT 75.790 173.355 76.020 174.495 ;
        RECT 76.190 173.345 76.520 174.325 ;
        RECT 76.690 173.355 76.900 174.495 ;
        RECT 73.545 172.935 74.045 173.105 ;
        RECT 73.545 172.765 73.715 172.935 ;
        RECT 74.435 172.765 74.930 173.305 ;
        RECT 75.770 172.935 76.100 173.185 ;
        RECT 70.695 172.595 72.345 172.765 ;
        RECT 73.080 172.595 73.715 172.765 ;
        RECT 73.920 172.595 74.930 172.765 ;
        RECT 69.260 171.945 69.540 172.425 ;
        RECT 69.770 172.115 70.070 172.445 ;
        RECT 70.240 171.945 70.515 172.425 ;
        RECT 70.695 172.205 70.990 172.595 ;
        RECT 71.160 171.945 71.415 172.425 ;
        RECT 71.590 172.205 71.850 172.595 ;
        RECT 72.020 171.945 72.300 172.425 ;
        RECT 73.080 172.115 73.250 172.595 ;
        RECT 73.430 171.945 73.670 172.425 ;
        RECT 73.920 172.115 74.090 172.595 ;
        RECT 74.260 171.945 74.590 172.425 ;
        RECT 74.760 172.115 74.930 172.595 ;
        RECT 75.100 171.945 75.430 172.745 ;
        RECT 75.790 171.945 76.020 172.765 ;
        RECT 76.270 172.745 76.520 173.345 ;
        RECT 77.135 173.305 77.390 174.185 ;
        RECT 77.560 173.355 77.865 174.495 ;
        RECT 78.205 174.115 78.535 174.495 ;
        RECT 78.715 173.945 78.885 174.235 ;
        RECT 79.055 174.035 79.305 174.495 ;
        RECT 78.085 173.775 78.885 173.945 ;
        RECT 79.475 173.985 80.345 174.325 ;
        RECT 76.190 172.115 76.520 172.745 ;
        RECT 76.690 171.945 76.900 172.765 ;
        RECT 77.135 172.655 77.345 173.305 ;
        RECT 78.085 173.185 78.255 173.775 ;
        RECT 79.475 173.605 79.645 173.985 ;
        RECT 80.580 173.865 80.750 174.325 ;
        RECT 80.920 174.035 81.290 174.495 ;
        RECT 81.585 173.895 81.755 174.235 ;
        RECT 81.925 174.065 82.255 174.495 ;
        RECT 82.490 173.895 82.660 174.235 ;
        RECT 78.425 173.435 79.645 173.605 ;
        RECT 79.815 173.525 80.275 173.815 ;
        RECT 80.580 173.695 81.140 173.865 ;
        RECT 81.585 173.725 82.660 173.895 ;
        RECT 82.830 173.995 83.510 174.325 ;
        RECT 83.725 173.995 83.975 174.325 ;
        RECT 84.145 174.035 84.395 174.495 ;
        RECT 80.970 173.555 81.140 173.695 ;
        RECT 79.815 173.515 80.780 173.525 ;
        RECT 79.475 173.345 79.645 173.435 ;
        RECT 80.105 173.355 80.780 173.515 ;
        RECT 77.515 173.155 78.255 173.185 ;
        RECT 77.515 172.855 78.430 173.155 ;
        RECT 78.105 172.680 78.430 172.855 ;
        RECT 77.135 172.125 77.390 172.655 ;
        RECT 77.560 171.945 77.865 172.405 ;
        RECT 78.110 172.325 78.430 172.680 ;
        RECT 78.600 172.895 79.140 173.265 ;
        RECT 79.475 173.175 79.880 173.345 ;
        RECT 78.600 172.495 78.840 172.895 ;
        RECT 79.320 172.725 79.540 173.005 ;
        RECT 79.010 172.555 79.540 172.725 ;
        RECT 79.010 172.325 79.180 172.555 ;
        RECT 79.710 172.395 79.880 173.175 ;
        RECT 80.050 172.565 80.400 173.185 ;
        RECT 80.570 172.565 80.780 173.355 ;
        RECT 80.970 173.385 82.470 173.555 ;
        RECT 80.970 172.695 81.140 173.385 ;
        RECT 82.830 173.215 83.000 173.995 ;
        RECT 83.805 173.865 83.975 173.995 ;
        RECT 81.310 173.045 83.000 173.215 ;
        RECT 83.170 173.435 83.635 173.825 ;
        RECT 83.805 173.695 84.200 173.865 ;
        RECT 81.310 172.865 81.480 173.045 ;
        RECT 78.110 172.155 79.180 172.325 ;
        RECT 79.350 171.945 79.540 172.385 ;
        RECT 79.710 172.115 80.660 172.395 ;
        RECT 80.970 172.305 81.230 172.695 ;
        RECT 81.650 172.625 82.440 172.875 ;
        RECT 80.880 172.135 81.230 172.305 ;
        RECT 81.440 171.945 81.770 172.405 ;
        RECT 82.645 172.335 82.815 173.045 ;
        RECT 83.170 172.845 83.340 173.435 ;
        RECT 82.985 172.625 83.340 172.845 ;
        RECT 83.510 172.625 83.860 173.245 ;
        RECT 84.030 172.335 84.200 173.695 ;
        RECT 84.565 173.525 84.890 174.310 ;
        RECT 84.370 172.475 84.830 173.525 ;
        RECT 82.645 172.165 83.500 172.335 ;
        RECT 83.705 172.165 84.200 172.335 ;
        RECT 84.370 171.945 84.700 172.305 ;
        RECT 85.060 172.205 85.230 174.325 ;
        RECT 85.400 173.995 85.730 174.495 ;
        RECT 85.900 173.825 86.155 174.325 ;
        RECT 85.405 173.655 86.155 173.825 ;
        RECT 85.405 172.665 85.635 173.655 ;
        RECT 85.805 172.835 86.155 173.485 ;
        RECT 86.330 173.330 86.620 174.495 ;
        RECT 86.850 173.355 87.060 174.495 ;
        RECT 87.230 173.345 87.560 174.325 ;
        RECT 87.730 173.355 87.960 174.495 ;
        RECT 85.405 172.495 86.155 172.665 ;
        RECT 85.400 171.945 85.730 172.325 ;
        RECT 85.900 172.205 86.155 172.495 ;
        RECT 86.330 171.945 86.620 172.670 ;
        RECT 86.850 171.945 87.060 172.765 ;
        RECT 87.230 172.745 87.480 173.345 ;
        RECT 88.175 173.305 88.430 174.185 ;
        RECT 88.600 173.355 88.905 174.495 ;
        RECT 89.245 174.115 89.575 174.495 ;
        RECT 89.755 173.945 89.925 174.235 ;
        RECT 90.095 174.035 90.345 174.495 ;
        RECT 89.125 173.775 89.925 173.945 ;
        RECT 90.515 173.985 91.385 174.325 ;
        RECT 87.650 172.935 87.980 173.185 ;
        RECT 87.230 172.115 87.560 172.745 ;
        RECT 87.730 171.945 87.960 172.765 ;
        RECT 88.175 172.655 88.385 173.305 ;
        RECT 89.125 173.185 89.295 173.775 ;
        RECT 90.515 173.605 90.685 173.985 ;
        RECT 91.620 173.865 91.790 174.325 ;
        RECT 91.960 174.035 92.330 174.495 ;
        RECT 92.625 173.895 92.795 174.235 ;
        RECT 92.965 174.065 93.295 174.495 ;
        RECT 93.530 173.895 93.700 174.235 ;
        RECT 89.465 173.435 90.685 173.605 ;
        RECT 90.855 173.525 91.315 173.815 ;
        RECT 91.620 173.695 92.180 173.865 ;
        RECT 92.625 173.725 93.700 173.895 ;
        RECT 93.870 173.995 94.550 174.325 ;
        RECT 94.765 173.995 95.015 174.325 ;
        RECT 95.185 174.035 95.435 174.495 ;
        RECT 92.010 173.555 92.180 173.695 ;
        RECT 90.855 173.515 91.820 173.525 ;
        RECT 90.515 173.345 90.685 173.435 ;
        RECT 91.145 173.355 91.820 173.515 ;
        RECT 88.555 173.155 89.295 173.185 ;
        RECT 88.555 172.855 89.470 173.155 ;
        RECT 89.145 172.680 89.470 172.855 ;
        RECT 88.175 172.125 88.430 172.655 ;
        RECT 88.600 171.945 88.905 172.405 ;
        RECT 89.150 172.325 89.470 172.680 ;
        RECT 89.640 172.895 90.180 173.265 ;
        RECT 90.515 173.175 90.920 173.345 ;
        RECT 89.640 172.495 89.880 172.895 ;
        RECT 90.360 172.725 90.580 173.005 ;
        RECT 90.050 172.555 90.580 172.725 ;
        RECT 90.050 172.325 90.220 172.555 ;
        RECT 90.750 172.395 90.920 173.175 ;
        RECT 91.090 172.565 91.440 173.185 ;
        RECT 91.610 172.565 91.820 173.355 ;
        RECT 92.010 173.385 93.510 173.555 ;
        RECT 92.010 172.695 92.180 173.385 ;
        RECT 93.870 173.215 94.040 173.995 ;
        RECT 94.845 173.865 95.015 173.995 ;
        RECT 92.350 173.045 94.040 173.215 ;
        RECT 94.210 173.435 94.675 173.825 ;
        RECT 94.845 173.695 95.240 173.865 ;
        RECT 92.350 172.865 92.520 173.045 ;
        RECT 89.150 172.155 90.220 172.325 ;
        RECT 90.390 171.945 90.580 172.385 ;
        RECT 90.750 172.115 91.700 172.395 ;
        RECT 92.010 172.305 92.270 172.695 ;
        RECT 92.690 172.625 93.480 172.875 ;
        RECT 91.920 172.135 92.270 172.305 ;
        RECT 92.480 171.945 92.810 172.405 ;
        RECT 93.685 172.335 93.855 173.045 ;
        RECT 94.210 172.845 94.380 173.435 ;
        RECT 94.025 172.625 94.380 172.845 ;
        RECT 94.550 172.625 94.900 173.245 ;
        RECT 95.070 172.335 95.240 173.695 ;
        RECT 95.605 173.525 95.930 174.310 ;
        RECT 95.410 172.475 95.870 173.525 ;
        RECT 93.685 172.165 94.540 172.335 ;
        RECT 94.745 172.165 95.240 172.335 ;
        RECT 95.410 171.945 95.740 172.305 ;
        RECT 96.100 172.205 96.270 174.325 ;
        RECT 96.440 173.995 96.770 174.495 ;
        RECT 96.940 173.825 97.195 174.325 ;
        RECT 96.445 173.655 97.195 173.825 ;
        RECT 96.445 172.665 96.675 173.655 ;
        RECT 96.845 172.835 97.195 173.485 ;
        RECT 97.870 173.355 98.100 174.495 ;
        RECT 98.270 173.345 98.600 174.325 ;
        RECT 98.770 173.355 98.980 174.495 ;
        RECT 97.850 172.935 98.180 173.185 ;
        RECT 96.445 172.495 97.195 172.665 ;
        RECT 96.440 171.945 96.770 172.325 ;
        RECT 96.940 172.205 97.195 172.495 ;
        RECT 97.870 171.945 98.100 172.765 ;
        RECT 98.350 172.745 98.600 173.345 ;
        RECT 99.675 173.305 99.930 174.185 ;
        RECT 100.100 173.355 100.405 174.495 ;
        RECT 100.745 174.115 101.075 174.495 ;
        RECT 101.255 173.945 101.425 174.235 ;
        RECT 101.595 174.035 101.845 174.495 ;
        RECT 100.625 173.775 101.425 173.945 ;
        RECT 102.015 173.985 102.885 174.325 ;
        RECT 98.270 172.115 98.600 172.745 ;
        RECT 98.770 171.945 98.980 172.765 ;
        RECT 99.675 172.655 99.885 173.305 ;
        RECT 100.625 173.185 100.795 173.775 ;
        RECT 102.015 173.605 102.185 173.985 ;
        RECT 103.120 173.865 103.290 174.325 ;
        RECT 103.460 174.035 103.830 174.495 ;
        RECT 104.125 173.895 104.295 174.235 ;
        RECT 104.465 174.065 104.795 174.495 ;
        RECT 105.030 173.895 105.200 174.235 ;
        RECT 100.965 173.435 102.185 173.605 ;
        RECT 102.355 173.525 102.815 173.815 ;
        RECT 103.120 173.695 103.680 173.865 ;
        RECT 104.125 173.725 105.200 173.895 ;
        RECT 105.370 173.995 106.050 174.325 ;
        RECT 106.265 173.995 106.515 174.325 ;
        RECT 106.685 174.035 106.935 174.495 ;
        RECT 103.510 173.555 103.680 173.695 ;
        RECT 102.355 173.515 103.320 173.525 ;
        RECT 102.015 173.345 102.185 173.435 ;
        RECT 102.645 173.355 103.320 173.515 ;
        RECT 100.055 173.155 100.795 173.185 ;
        RECT 100.055 172.855 100.970 173.155 ;
        RECT 100.645 172.680 100.970 172.855 ;
        RECT 99.675 172.125 99.930 172.655 ;
        RECT 100.100 171.945 100.405 172.405 ;
        RECT 100.650 172.325 100.970 172.680 ;
        RECT 101.140 172.895 101.680 173.265 ;
        RECT 102.015 173.175 102.420 173.345 ;
        RECT 101.140 172.495 101.380 172.895 ;
        RECT 101.860 172.725 102.080 173.005 ;
        RECT 101.550 172.555 102.080 172.725 ;
        RECT 101.550 172.325 101.720 172.555 ;
        RECT 102.250 172.395 102.420 173.175 ;
        RECT 102.590 172.565 102.940 173.185 ;
        RECT 103.110 172.565 103.320 173.355 ;
        RECT 103.510 173.385 105.010 173.555 ;
        RECT 103.510 172.695 103.680 173.385 ;
        RECT 105.370 173.215 105.540 173.995 ;
        RECT 106.345 173.865 106.515 173.995 ;
        RECT 103.850 173.045 105.540 173.215 ;
        RECT 105.710 173.435 106.175 173.825 ;
        RECT 106.345 173.695 106.740 173.865 ;
        RECT 103.850 172.865 104.020 173.045 ;
        RECT 100.650 172.155 101.720 172.325 ;
        RECT 101.890 171.945 102.080 172.385 ;
        RECT 102.250 172.115 103.200 172.395 ;
        RECT 103.510 172.305 103.770 172.695 ;
        RECT 104.190 172.625 104.980 172.875 ;
        RECT 103.420 172.135 103.770 172.305 ;
        RECT 103.980 171.945 104.310 172.405 ;
        RECT 105.185 172.335 105.355 173.045 ;
        RECT 105.710 172.845 105.880 173.435 ;
        RECT 105.525 172.625 105.880 172.845 ;
        RECT 106.050 172.625 106.400 173.245 ;
        RECT 106.570 172.335 106.740 173.695 ;
        RECT 107.105 173.525 107.430 174.310 ;
        RECT 106.910 172.475 107.370 173.525 ;
        RECT 105.185 172.165 106.040 172.335 ;
        RECT 106.245 172.165 106.740 172.335 ;
        RECT 106.910 171.945 107.240 172.305 ;
        RECT 107.600 172.205 107.770 174.325 ;
        RECT 107.940 173.995 108.270 174.495 ;
        RECT 108.440 173.825 108.695 174.325 ;
        RECT 107.945 173.655 108.695 173.825 ;
        RECT 107.945 172.665 108.175 173.655 ;
        RECT 108.345 172.835 108.695 173.485 ;
        RECT 108.870 173.420 109.140 174.325 ;
        RECT 109.310 173.735 109.640 174.495 ;
        RECT 109.820 173.565 109.990 174.325 ;
        RECT 107.945 172.495 108.695 172.665 ;
        RECT 107.940 171.945 108.270 172.325 ;
        RECT 108.440 172.205 108.695 172.495 ;
        RECT 108.870 172.620 109.040 173.420 ;
        RECT 109.325 173.395 109.990 173.565 ;
        RECT 111.170 173.405 112.380 174.495 ;
        RECT 109.325 173.250 109.495 173.395 ;
        RECT 109.210 172.920 109.495 173.250 ;
        RECT 109.325 172.665 109.495 172.920 ;
        RECT 109.730 172.845 110.060 173.215 ;
        RECT 111.170 172.865 111.690 173.405 ;
        RECT 111.860 172.695 112.380 173.235 ;
        RECT 108.870 172.115 109.130 172.620 ;
        RECT 109.325 172.495 109.990 172.665 ;
        RECT 109.310 171.945 109.640 172.325 ;
        RECT 109.820 172.115 109.990 172.495 ;
        RECT 111.170 171.945 112.380 172.695 ;
        RECT 18.165 171.775 112.465 171.945 ;
        RECT 18.250 171.025 19.460 171.775 ;
        RECT 18.250 170.485 18.770 171.025 ;
        RECT 20.590 170.955 20.820 171.775 ;
        RECT 20.990 170.975 21.320 171.605 ;
        RECT 18.940 170.315 19.460 170.855 ;
        RECT 20.570 170.535 20.900 170.785 ;
        RECT 21.070 170.375 21.320 170.975 ;
        RECT 21.490 170.955 21.700 171.775 ;
        RECT 21.930 171.050 22.220 171.775 ;
        RECT 22.395 171.225 22.650 171.515 ;
        RECT 22.820 171.395 23.150 171.775 ;
        RECT 22.395 171.055 23.145 171.225 ;
        RECT 18.250 169.225 19.460 170.315 ;
        RECT 20.590 169.225 20.820 170.365 ;
        RECT 20.990 169.395 21.320 170.375 ;
        RECT 21.490 169.225 21.700 170.365 ;
        RECT 21.930 169.225 22.220 170.390 ;
        RECT 22.395 170.235 22.745 170.885 ;
        RECT 22.915 170.065 23.145 171.055 ;
        RECT 22.395 169.895 23.145 170.065 ;
        RECT 22.395 169.395 22.650 169.895 ;
        RECT 22.820 169.225 23.150 169.725 ;
        RECT 23.320 169.395 23.490 171.515 ;
        RECT 23.850 171.415 24.180 171.775 ;
        RECT 24.350 171.385 24.845 171.555 ;
        RECT 25.050 171.385 25.905 171.555 ;
        RECT 23.720 170.195 24.180 171.245 ;
        RECT 23.660 169.410 23.985 170.195 ;
        RECT 24.350 170.025 24.520 171.385 ;
        RECT 24.690 170.475 25.040 171.095 ;
        RECT 25.210 170.875 25.565 171.095 ;
        RECT 25.210 170.285 25.380 170.875 ;
        RECT 25.735 170.675 25.905 171.385 ;
        RECT 26.780 171.315 27.110 171.775 ;
        RECT 27.320 171.415 27.670 171.585 ;
        RECT 26.110 170.845 26.900 171.095 ;
        RECT 27.320 171.025 27.580 171.415 ;
        RECT 27.890 171.325 28.840 171.605 ;
        RECT 29.010 171.335 29.200 171.775 ;
        RECT 29.370 171.395 30.440 171.565 ;
        RECT 27.070 170.675 27.240 170.855 ;
        RECT 24.350 169.855 24.745 170.025 ;
        RECT 24.915 169.895 25.380 170.285 ;
        RECT 25.550 170.505 27.240 170.675 ;
        RECT 24.575 169.725 24.745 169.855 ;
        RECT 25.550 169.725 25.720 170.505 ;
        RECT 27.410 170.335 27.580 171.025 ;
        RECT 26.080 170.165 27.580 170.335 ;
        RECT 27.770 170.365 27.980 171.155 ;
        RECT 28.150 170.535 28.500 171.155 ;
        RECT 28.670 170.545 28.840 171.325 ;
        RECT 29.370 171.165 29.540 171.395 ;
        RECT 29.010 170.995 29.540 171.165 ;
        RECT 29.010 170.715 29.230 170.995 ;
        RECT 29.710 170.825 29.950 171.225 ;
        RECT 28.670 170.375 29.075 170.545 ;
        RECT 29.410 170.455 29.950 170.825 ;
        RECT 30.120 171.040 30.440 171.395 ;
        RECT 30.685 171.315 30.990 171.775 ;
        RECT 31.160 171.065 31.415 171.595 ;
        RECT 30.120 170.865 30.445 171.040 ;
        RECT 30.120 170.565 31.035 170.865 ;
        RECT 30.295 170.535 31.035 170.565 ;
        RECT 27.770 170.205 28.445 170.365 ;
        RECT 28.905 170.285 29.075 170.375 ;
        RECT 27.770 170.195 28.735 170.205 ;
        RECT 27.410 170.025 27.580 170.165 ;
        RECT 24.155 169.225 24.405 169.685 ;
        RECT 24.575 169.395 24.825 169.725 ;
        RECT 25.040 169.395 25.720 169.725 ;
        RECT 25.890 169.825 26.965 169.995 ;
        RECT 27.410 169.855 27.970 170.025 ;
        RECT 28.275 169.905 28.735 170.195 ;
        RECT 28.905 170.115 30.125 170.285 ;
        RECT 25.890 169.485 26.060 169.825 ;
        RECT 26.295 169.225 26.625 169.655 ;
        RECT 26.795 169.485 26.965 169.825 ;
        RECT 27.260 169.225 27.630 169.685 ;
        RECT 27.800 169.395 27.970 169.855 ;
        RECT 28.905 169.735 29.075 170.115 ;
        RECT 30.295 169.945 30.465 170.535 ;
        RECT 31.205 170.415 31.415 171.065 ;
        RECT 31.795 170.995 32.295 171.605 ;
        RECT 31.590 170.535 31.940 170.785 ;
        RECT 28.205 169.395 29.075 169.735 ;
        RECT 29.665 169.775 30.465 169.945 ;
        RECT 29.245 169.225 29.495 169.685 ;
        RECT 29.665 169.485 29.835 169.775 ;
        RECT 30.015 169.225 30.345 169.605 ;
        RECT 30.685 169.225 30.990 170.365 ;
        RECT 31.160 169.535 31.415 170.415 ;
        RECT 32.125 170.365 32.295 170.995 ;
        RECT 32.925 171.125 33.255 171.605 ;
        RECT 33.425 171.315 33.650 171.775 ;
        RECT 33.820 171.125 34.150 171.605 ;
        RECT 32.925 170.955 34.150 171.125 ;
        RECT 34.340 170.975 34.590 171.775 ;
        RECT 34.760 170.975 35.100 171.605 ;
        RECT 32.465 170.585 32.795 170.785 ;
        RECT 32.965 170.585 33.295 170.785 ;
        RECT 33.465 170.585 33.885 170.785 ;
        RECT 34.060 170.615 34.755 170.785 ;
        RECT 34.060 170.365 34.230 170.615 ;
        RECT 34.925 170.365 35.100 170.975 ;
        RECT 31.795 170.195 34.230 170.365 ;
        RECT 31.795 169.395 32.125 170.195 ;
        RECT 32.295 169.225 32.625 170.025 ;
        RECT 32.925 169.395 33.255 170.195 ;
        RECT 33.900 169.225 34.150 170.025 ;
        RECT 34.420 169.225 34.590 170.365 ;
        RECT 34.760 169.395 35.100 170.365 ;
        RECT 35.270 170.975 35.610 171.605 ;
        RECT 35.780 170.975 36.030 171.775 ;
        RECT 36.220 171.125 36.550 171.605 ;
        RECT 36.720 171.315 36.945 171.775 ;
        RECT 37.115 171.125 37.445 171.605 ;
        RECT 35.270 170.365 35.445 170.975 ;
        RECT 36.220 170.955 37.445 171.125 ;
        RECT 38.075 170.995 38.575 171.605 ;
        RECT 39.410 171.005 42.920 171.775 ;
        RECT 35.615 170.615 36.310 170.785 ;
        RECT 36.140 170.365 36.310 170.615 ;
        RECT 36.485 170.585 36.905 170.785 ;
        RECT 37.075 170.585 37.405 170.785 ;
        RECT 37.575 170.585 37.905 170.785 ;
        RECT 38.075 170.365 38.245 170.995 ;
        RECT 38.430 170.535 38.780 170.785 ;
        RECT 35.270 169.395 35.610 170.365 ;
        RECT 35.780 169.225 35.950 170.365 ;
        RECT 36.140 170.195 38.575 170.365 ;
        RECT 36.220 169.225 36.470 170.025 ;
        RECT 37.115 169.395 37.445 170.195 ;
        RECT 37.745 169.225 38.075 170.025 ;
        RECT 38.245 169.395 38.575 170.195 ;
        RECT 39.410 170.315 41.100 170.835 ;
        RECT 41.270 170.485 42.920 171.005 ;
        RECT 43.090 170.975 43.430 171.605 ;
        RECT 43.600 170.975 43.850 171.775 ;
        RECT 44.040 171.125 44.370 171.605 ;
        RECT 44.540 171.315 44.765 171.775 ;
        RECT 44.935 171.125 45.265 171.605 ;
        RECT 43.090 170.365 43.265 170.975 ;
        RECT 44.040 170.955 45.265 171.125 ;
        RECT 45.895 170.995 46.395 171.605 ;
        RECT 47.690 171.050 47.980 171.775 ;
        RECT 43.435 170.615 44.130 170.785 ;
        RECT 43.960 170.365 44.130 170.615 ;
        RECT 44.305 170.585 44.725 170.785 ;
        RECT 44.895 170.585 45.225 170.785 ;
        RECT 45.395 170.585 45.725 170.785 ;
        RECT 45.895 170.365 46.065 170.995 ;
        RECT 48.150 170.975 48.490 171.605 ;
        RECT 48.660 170.975 48.910 171.775 ;
        RECT 49.100 171.125 49.430 171.605 ;
        RECT 49.600 171.315 49.825 171.775 ;
        RECT 49.995 171.125 50.325 171.605 ;
        RECT 46.250 170.535 46.600 170.785 ;
        RECT 39.410 169.225 42.920 170.315 ;
        RECT 43.090 169.395 43.430 170.365 ;
        RECT 43.600 169.225 43.770 170.365 ;
        RECT 43.960 170.195 46.395 170.365 ;
        RECT 44.040 169.225 44.290 170.025 ;
        RECT 44.935 169.395 45.265 170.195 ;
        RECT 45.565 169.225 45.895 170.025 ;
        RECT 46.065 169.395 46.395 170.195 ;
        RECT 47.690 169.225 47.980 170.390 ;
        RECT 48.150 170.365 48.325 170.975 ;
        RECT 49.100 170.955 50.325 171.125 ;
        RECT 50.955 170.995 51.455 171.605 ;
        RECT 51.830 171.005 53.500 171.775 ;
        RECT 53.730 171.295 54.010 171.775 ;
        RECT 54.180 171.125 54.440 171.515 ;
        RECT 54.615 171.295 54.870 171.775 ;
        RECT 55.040 171.125 55.335 171.515 ;
        RECT 55.515 171.295 55.790 171.775 ;
        RECT 55.960 171.275 56.260 171.605 ;
        RECT 48.495 170.615 49.190 170.785 ;
        RECT 49.020 170.365 49.190 170.615 ;
        RECT 49.365 170.585 49.785 170.785 ;
        RECT 49.955 170.585 50.285 170.785 ;
        RECT 50.455 170.585 50.785 170.785 ;
        RECT 50.955 170.365 51.125 170.995 ;
        RECT 51.310 170.535 51.660 170.785 ;
        RECT 48.150 169.395 48.490 170.365 ;
        RECT 48.660 169.225 48.830 170.365 ;
        RECT 49.020 170.195 51.455 170.365 ;
        RECT 49.100 169.225 49.350 170.025 ;
        RECT 49.995 169.395 50.325 170.195 ;
        RECT 50.625 169.225 50.955 170.025 ;
        RECT 51.125 169.395 51.455 170.195 ;
        RECT 51.830 170.315 52.580 170.835 ;
        RECT 52.750 170.485 53.500 171.005 ;
        RECT 53.685 170.955 55.335 171.125 ;
        RECT 53.685 170.445 54.090 170.955 ;
        RECT 54.260 170.615 55.400 170.785 ;
        RECT 51.830 169.225 53.500 170.315 ;
        RECT 53.685 170.275 54.440 170.445 ;
        RECT 53.725 169.225 54.010 170.095 ;
        RECT 54.180 170.025 54.440 170.275 ;
        RECT 55.230 170.365 55.400 170.615 ;
        RECT 55.570 170.535 55.920 171.105 ;
        RECT 56.090 170.365 56.260 171.275 ;
        RECT 57.440 171.225 57.610 171.605 ;
        RECT 57.825 171.395 58.155 171.775 ;
        RECT 57.440 171.055 58.155 171.225 ;
        RECT 57.350 170.505 57.705 170.875 ;
        RECT 57.985 170.865 58.155 171.055 ;
        RECT 58.325 171.030 58.580 171.605 ;
        RECT 57.985 170.535 58.240 170.865 ;
        RECT 55.230 170.195 56.260 170.365 ;
        RECT 57.985 170.325 58.155 170.535 ;
        RECT 54.180 169.855 55.300 170.025 ;
        RECT 54.180 169.395 54.440 169.855 ;
        RECT 54.615 169.225 54.870 169.685 ;
        RECT 55.040 169.395 55.300 169.855 ;
        RECT 55.470 169.225 55.780 170.025 ;
        RECT 55.950 169.395 56.260 170.195 ;
        RECT 57.440 170.155 58.155 170.325 ;
        RECT 58.410 170.300 58.580 171.030 ;
        RECT 58.755 170.935 59.015 171.775 ;
        RECT 59.460 171.380 59.790 171.775 ;
        RECT 59.960 171.205 60.160 171.560 ;
        RECT 60.330 171.375 60.660 171.775 ;
        RECT 60.830 171.205 61.030 171.550 ;
        RECT 59.190 171.035 61.030 171.205 ;
        RECT 61.200 171.035 61.530 171.775 ;
        RECT 61.765 171.205 61.935 171.455 ;
        RECT 61.765 171.035 62.240 171.205 ;
        RECT 57.440 169.395 57.610 170.155 ;
        RECT 57.825 169.225 58.155 169.985 ;
        RECT 58.325 169.395 58.580 170.300 ;
        RECT 58.755 169.225 59.015 170.375 ;
        RECT 59.190 169.410 59.450 171.035 ;
        RECT 59.630 170.065 59.850 170.865 ;
        RECT 60.090 170.245 60.390 170.865 ;
        RECT 60.560 170.245 60.890 170.865 ;
        RECT 61.060 170.245 61.380 170.865 ;
        RECT 61.550 170.245 61.900 170.865 ;
        RECT 62.070 170.065 62.240 171.035 ;
        RECT 62.410 171.025 63.620 171.775 ;
        RECT 59.630 169.855 62.240 170.065 ;
        RECT 62.410 170.315 62.930 170.855 ;
        RECT 63.100 170.485 63.620 171.025 ;
        RECT 63.790 171.275 64.050 171.605 ;
        RECT 64.360 171.395 64.690 171.775 ;
        RECT 64.870 171.435 66.350 171.605 ;
        RECT 63.790 170.575 63.960 171.275 ;
        RECT 64.870 171.105 65.270 171.435 ;
        RECT 64.310 170.915 64.520 171.095 ;
        RECT 64.310 170.745 64.930 170.915 ;
        RECT 65.100 170.625 65.270 171.105 ;
        RECT 65.460 170.935 66.010 171.265 ;
        RECT 63.790 170.405 64.920 170.575 ;
        RECT 65.100 170.455 65.670 170.625 ;
        RECT 61.200 169.225 61.530 169.675 ;
        RECT 62.410 169.225 63.620 170.315 ;
        RECT 63.790 169.725 63.960 170.405 ;
        RECT 64.750 170.285 64.920 170.405 ;
        RECT 64.130 169.905 64.480 170.235 ;
        RECT 64.750 170.115 65.330 170.285 ;
        RECT 65.500 169.945 65.670 170.455 ;
        RECT 64.930 169.775 65.670 169.945 ;
        RECT 65.840 169.945 66.010 170.935 ;
        RECT 66.180 170.535 66.350 171.435 ;
        RECT 66.600 170.865 66.785 171.445 ;
        RECT 67.055 170.865 67.250 171.440 ;
        RECT 67.460 171.395 67.790 171.775 ;
        RECT 66.600 170.535 66.830 170.865 ;
        RECT 67.055 170.535 67.310 170.865 ;
        RECT 66.600 170.225 66.785 170.535 ;
        RECT 67.055 170.225 67.250 170.535 ;
        RECT 67.620 169.945 67.790 170.865 ;
        RECT 65.840 169.775 67.790 169.945 ;
        RECT 63.790 169.395 64.050 169.725 ;
        RECT 64.360 169.225 64.690 169.605 ;
        RECT 64.930 169.395 65.120 169.775 ;
        RECT 65.370 169.225 65.700 169.605 ;
        RECT 65.910 169.395 66.080 169.775 ;
        RECT 66.275 169.225 66.605 169.605 ;
        RECT 66.865 169.395 67.035 169.775 ;
        RECT 67.460 169.225 67.790 169.605 ;
        RECT 67.960 169.395 68.220 171.605 ;
        RECT 68.695 171.205 68.865 171.455 ;
        RECT 68.390 171.035 68.865 171.205 ;
        RECT 69.100 171.035 69.430 171.775 ;
        RECT 69.600 171.205 69.800 171.550 ;
        RECT 69.970 171.375 70.300 171.775 ;
        RECT 70.470 171.205 70.670 171.560 ;
        RECT 70.840 171.380 71.170 171.775 ;
        RECT 72.160 171.225 72.330 171.605 ;
        RECT 72.510 171.395 72.840 171.775 ;
        RECT 69.600 171.035 71.440 171.205 ;
        RECT 72.160 171.055 72.825 171.225 ;
        RECT 73.020 171.100 73.280 171.605 ;
        RECT 68.390 170.065 68.560 171.035 ;
        RECT 68.730 170.245 69.080 170.865 ;
        RECT 69.250 170.245 69.570 170.865 ;
        RECT 69.740 170.245 70.070 170.865 ;
        RECT 70.240 170.245 70.540 170.865 ;
        RECT 70.780 170.065 71.000 170.865 ;
        RECT 68.390 169.855 71.000 170.065 ;
        RECT 69.100 169.225 69.430 169.675 ;
        RECT 71.180 169.410 71.440 171.035 ;
        RECT 72.090 170.505 72.420 170.875 ;
        RECT 72.655 170.800 72.825 171.055 ;
        RECT 72.655 170.470 72.940 170.800 ;
        RECT 72.655 170.325 72.825 170.470 ;
        RECT 72.160 170.155 72.825 170.325 ;
        RECT 73.110 170.300 73.280 171.100 ;
        RECT 73.450 171.050 73.740 171.775 ;
        RECT 74.000 171.225 74.170 171.515 ;
        RECT 74.340 171.395 74.670 171.775 ;
        RECT 74.000 171.055 74.665 171.225 ;
        RECT 72.160 169.395 72.330 170.155 ;
        RECT 72.510 169.225 72.840 169.985 ;
        RECT 73.010 169.395 73.280 170.300 ;
        RECT 73.450 169.225 73.740 170.390 ;
        RECT 73.915 170.235 74.265 170.885 ;
        RECT 74.435 170.065 74.665 171.055 ;
        RECT 74.000 169.895 74.665 170.065 ;
        RECT 74.000 169.395 74.170 169.895 ;
        RECT 74.340 169.225 74.670 169.725 ;
        RECT 74.840 169.395 75.065 171.515 ;
        RECT 75.280 171.395 75.610 171.775 ;
        RECT 75.780 171.225 75.950 171.555 ;
        RECT 76.250 171.395 77.265 171.595 ;
        RECT 75.255 171.035 75.950 171.225 ;
        RECT 75.255 170.065 75.425 171.035 ;
        RECT 75.595 170.235 76.005 170.855 ;
        RECT 76.175 170.285 76.395 171.155 ;
        RECT 76.575 170.845 76.925 171.215 ;
        RECT 77.095 170.665 77.265 171.395 ;
        RECT 77.435 171.335 77.845 171.775 ;
        RECT 78.135 171.135 78.385 171.565 ;
        RECT 78.585 171.315 78.905 171.775 ;
        RECT 79.465 171.385 80.315 171.555 ;
        RECT 77.435 170.795 77.845 171.125 ;
        RECT 78.135 170.795 78.555 171.135 ;
        RECT 76.845 170.625 77.265 170.665 ;
        RECT 76.845 170.455 78.195 170.625 ;
        RECT 75.255 169.895 75.950 170.065 ;
        RECT 76.175 169.905 76.675 170.285 ;
        RECT 75.280 169.225 75.610 169.725 ;
        RECT 75.780 169.395 75.950 169.895 ;
        RECT 76.845 169.610 77.015 170.455 ;
        RECT 77.945 170.295 78.195 170.455 ;
        RECT 77.185 170.025 77.435 170.285 ;
        RECT 78.365 170.025 78.555 170.795 ;
        RECT 77.185 169.775 78.555 170.025 ;
        RECT 78.725 170.965 79.975 171.135 ;
        RECT 78.725 170.205 78.895 170.965 ;
        RECT 79.645 170.845 79.975 170.965 ;
        RECT 79.065 170.385 79.245 170.795 ;
        RECT 80.145 170.625 80.315 171.385 ;
        RECT 80.515 171.295 81.175 171.775 ;
        RECT 81.355 171.180 81.675 171.510 ;
        RECT 80.505 170.855 81.165 171.125 ;
        RECT 80.505 170.795 80.835 170.855 ;
        RECT 80.985 170.625 81.315 170.685 ;
        RECT 79.415 170.455 81.315 170.625 ;
        RECT 78.725 169.895 79.245 170.205 ;
        RECT 79.415 169.945 79.585 170.455 ;
        RECT 81.485 170.285 81.675 171.180 ;
        RECT 79.755 170.115 81.675 170.285 ;
        RECT 81.355 170.095 81.675 170.115 ;
        RECT 81.875 170.865 82.125 171.515 ;
        RECT 82.305 171.315 82.590 171.775 ;
        RECT 82.770 171.065 83.025 171.595 ;
        RECT 81.875 170.535 82.675 170.865 ;
        RECT 79.415 169.775 80.625 169.945 ;
        RECT 76.185 169.440 77.015 169.610 ;
        RECT 77.255 169.225 77.635 169.605 ;
        RECT 77.815 169.485 77.985 169.775 ;
        RECT 79.415 169.695 79.585 169.775 ;
        RECT 78.155 169.225 78.485 169.605 ;
        RECT 78.955 169.445 79.585 169.695 ;
        RECT 79.765 169.225 80.185 169.605 ;
        RECT 80.385 169.485 80.625 169.775 ;
        RECT 80.855 169.225 81.185 169.915 ;
        RECT 81.355 169.485 81.525 170.095 ;
        RECT 81.875 169.945 82.125 170.535 ;
        RECT 82.845 170.205 83.025 171.065 ;
        RECT 83.845 170.965 84.090 171.570 ;
        RECT 84.310 171.240 84.820 171.775 ;
        RECT 81.795 169.435 82.125 169.945 ;
        RECT 82.305 169.225 82.590 170.025 ;
        RECT 82.770 169.735 83.025 170.205 ;
        RECT 83.570 170.795 84.800 170.965 ;
        RECT 83.570 169.985 83.910 170.795 ;
        RECT 84.080 170.230 84.830 170.420 ;
        RECT 82.770 169.565 83.110 169.735 ;
        RECT 83.570 169.575 84.085 169.985 ;
        RECT 82.770 169.535 83.025 169.565 ;
        RECT 84.320 169.225 84.490 169.985 ;
        RECT 84.660 169.565 84.830 170.230 ;
        RECT 85.000 170.245 85.190 171.605 ;
        RECT 85.360 170.755 85.635 171.605 ;
        RECT 85.825 171.240 86.355 171.605 ;
        RECT 86.780 171.375 87.110 171.775 ;
        RECT 86.180 171.205 86.355 171.240 ;
        RECT 85.360 170.585 85.640 170.755 ;
        RECT 85.360 170.445 85.635 170.585 ;
        RECT 85.840 170.245 86.010 171.045 ;
        RECT 85.000 170.075 86.010 170.245 ;
        RECT 86.180 171.035 87.110 171.205 ;
        RECT 87.280 171.035 87.535 171.605 ;
        RECT 86.180 169.905 86.350 171.035 ;
        RECT 86.940 170.865 87.110 171.035 ;
        RECT 85.225 169.735 86.350 169.905 ;
        RECT 86.520 170.535 86.715 170.865 ;
        RECT 86.940 170.535 87.195 170.865 ;
        RECT 86.520 169.565 86.690 170.535 ;
        RECT 87.365 170.365 87.535 171.035 ;
        RECT 87.825 171.145 88.110 171.605 ;
        RECT 88.280 171.315 88.550 171.775 ;
        RECT 87.825 170.975 88.780 171.145 ;
        RECT 84.660 169.395 86.690 169.565 ;
        RECT 86.860 169.225 87.030 170.365 ;
        RECT 87.200 169.395 87.535 170.365 ;
        RECT 87.710 170.245 88.400 170.805 ;
        RECT 88.570 170.075 88.780 170.975 ;
        RECT 87.825 169.855 88.780 170.075 ;
        RECT 88.950 170.805 89.350 171.605 ;
        RECT 89.540 171.145 89.820 171.605 ;
        RECT 90.340 171.315 90.665 171.775 ;
        RECT 89.540 170.975 90.665 171.145 ;
        RECT 90.835 171.035 91.220 171.605 ;
        RECT 90.215 170.865 90.665 170.975 ;
        RECT 88.950 170.245 90.045 170.805 ;
        RECT 90.215 170.535 90.770 170.865 ;
        RECT 87.825 169.395 88.110 169.855 ;
        RECT 88.280 169.225 88.550 169.685 ;
        RECT 88.950 169.395 89.350 170.245 ;
        RECT 90.215 170.075 90.665 170.535 ;
        RECT 90.940 170.365 91.220 171.035 ;
        RECT 91.665 170.965 91.910 171.570 ;
        RECT 92.130 171.240 92.640 171.775 ;
        RECT 89.540 169.855 90.665 170.075 ;
        RECT 89.540 169.395 89.820 169.855 ;
        RECT 90.340 169.225 90.665 169.685 ;
        RECT 90.835 169.395 91.220 170.365 ;
        RECT 91.390 170.795 92.620 170.965 ;
        RECT 91.390 169.985 91.730 170.795 ;
        RECT 91.900 170.230 92.650 170.420 ;
        RECT 91.390 169.575 91.905 169.985 ;
        RECT 92.140 169.225 92.310 169.985 ;
        RECT 92.480 169.565 92.650 170.230 ;
        RECT 92.820 170.245 93.010 171.605 ;
        RECT 93.180 171.095 93.455 171.605 ;
        RECT 93.645 171.240 94.175 171.605 ;
        RECT 94.600 171.375 94.930 171.775 ;
        RECT 94.000 171.205 94.175 171.240 ;
        RECT 93.180 170.925 93.460 171.095 ;
        RECT 93.180 170.445 93.455 170.925 ;
        RECT 93.660 170.245 93.830 171.045 ;
        RECT 92.820 170.075 93.830 170.245 ;
        RECT 94.000 171.035 94.930 171.205 ;
        RECT 95.100 171.035 95.355 171.605 ;
        RECT 94.000 169.905 94.170 171.035 ;
        RECT 94.760 170.865 94.930 171.035 ;
        RECT 93.045 169.735 94.170 169.905 ;
        RECT 94.340 170.535 94.535 170.865 ;
        RECT 94.760 170.535 95.015 170.865 ;
        RECT 94.340 169.565 94.510 170.535 ;
        RECT 95.185 170.365 95.355 171.035 ;
        RECT 92.480 169.395 94.510 169.565 ;
        RECT 94.680 169.225 94.850 170.365 ;
        RECT 95.020 169.395 95.355 170.365 ;
        RECT 95.530 171.100 95.790 171.605 ;
        RECT 95.970 171.395 96.300 171.775 ;
        RECT 96.480 171.225 96.650 171.605 ;
        RECT 95.530 170.300 95.700 171.100 ;
        RECT 95.985 171.055 96.650 171.225 ;
        RECT 96.910 171.100 97.170 171.605 ;
        RECT 97.350 171.395 97.680 171.775 ;
        RECT 97.860 171.225 98.030 171.605 ;
        RECT 95.985 170.800 96.155 171.055 ;
        RECT 95.870 170.470 96.155 170.800 ;
        RECT 96.390 170.505 96.720 170.875 ;
        RECT 95.985 170.325 96.155 170.470 ;
        RECT 95.530 169.395 95.800 170.300 ;
        RECT 95.985 170.155 96.650 170.325 ;
        RECT 95.970 169.225 96.300 169.985 ;
        RECT 96.480 169.395 96.650 170.155 ;
        RECT 96.910 170.300 97.080 171.100 ;
        RECT 97.365 171.055 98.030 171.225 ;
        RECT 97.365 170.800 97.535 171.055 ;
        RECT 99.210 171.050 99.500 171.775 ;
        RECT 100.865 170.965 101.110 171.570 ;
        RECT 101.330 171.240 101.840 171.775 ;
        RECT 97.250 170.470 97.535 170.800 ;
        RECT 97.770 170.505 98.100 170.875 ;
        RECT 100.590 170.795 101.820 170.965 ;
        RECT 97.365 170.325 97.535 170.470 ;
        RECT 96.910 169.395 97.180 170.300 ;
        RECT 97.365 170.155 98.030 170.325 ;
        RECT 97.350 169.225 97.680 169.985 ;
        RECT 97.860 169.395 98.030 170.155 ;
        RECT 99.210 169.225 99.500 170.390 ;
        RECT 100.590 169.985 100.930 170.795 ;
        RECT 101.100 170.230 101.850 170.420 ;
        RECT 100.590 169.575 101.105 169.985 ;
        RECT 101.340 169.225 101.510 169.985 ;
        RECT 101.680 169.565 101.850 170.230 ;
        RECT 102.020 170.245 102.210 171.605 ;
        RECT 102.380 170.755 102.655 171.605 ;
        RECT 102.845 171.240 103.375 171.605 ;
        RECT 103.800 171.375 104.130 171.775 ;
        RECT 103.200 171.205 103.375 171.240 ;
        RECT 102.380 170.585 102.660 170.755 ;
        RECT 102.380 170.445 102.655 170.585 ;
        RECT 102.860 170.245 103.030 171.045 ;
        RECT 102.020 170.075 103.030 170.245 ;
        RECT 103.200 171.035 104.130 171.205 ;
        RECT 104.300 171.035 104.555 171.605 ;
        RECT 103.200 169.905 103.370 171.035 ;
        RECT 103.960 170.865 104.130 171.035 ;
        RECT 102.245 169.735 103.370 169.905 ;
        RECT 103.540 170.535 103.735 170.865 ;
        RECT 103.960 170.535 104.215 170.865 ;
        RECT 103.540 169.565 103.710 170.535 ;
        RECT 104.385 170.365 104.555 171.035 ;
        RECT 101.680 169.395 103.710 169.565 ;
        RECT 103.880 169.225 104.050 170.365 ;
        RECT 104.220 169.395 104.555 170.365 ;
        RECT 104.735 171.035 104.990 171.605 ;
        RECT 105.160 171.375 105.490 171.775 ;
        RECT 105.915 171.240 106.445 171.605 ;
        RECT 105.915 171.205 106.090 171.240 ;
        RECT 105.160 171.035 106.090 171.205 ;
        RECT 106.635 171.095 106.910 171.605 ;
        RECT 104.735 170.365 104.905 171.035 ;
        RECT 105.160 170.865 105.330 171.035 ;
        RECT 105.075 170.535 105.330 170.865 ;
        RECT 105.555 170.535 105.750 170.865 ;
        RECT 104.735 169.395 105.070 170.365 ;
        RECT 105.240 169.225 105.410 170.365 ;
        RECT 105.580 169.565 105.750 170.535 ;
        RECT 105.920 169.905 106.090 171.035 ;
        RECT 106.260 170.245 106.430 171.045 ;
        RECT 106.630 170.925 106.910 171.095 ;
        RECT 106.635 170.445 106.910 170.925 ;
        RECT 107.080 170.245 107.270 171.605 ;
        RECT 107.450 171.240 107.960 171.775 ;
        RECT 108.180 170.965 108.425 171.570 ;
        RECT 109.330 171.005 111.000 171.775 ;
        RECT 111.170 171.025 112.380 171.775 ;
        RECT 107.470 170.795 108.700 170.965 ;
        RECT 106.260 170.075 107.270 170.245 ;
        RECT 107.440 170.230 108.190 170.420 ;
        RECT 105.920 169.735 107.045 169.905 ;
        RECT 107.440 169.565 107.610 170.230 ;
        RECT 108.360 169.985 108.700 170.795 ;
        RECT 105.580 169.395 107.610 169.565 ;
        RECT 107.780 169.225 107.950 169.985 ;
        RECT 108.185 169.575 108.700 169.985 ;
        RECT 109.330 170.315 110.080 170.835 ;
        RECT 110.250 170.485 111.000 171.005 ;
        RECT 111.170 170.315 111.690 170.855 ;
        RECT 111.860 170.485 112.380 171.025 ;
        RECT 109.330 169.225 111.000 170.315 ;
        RECT 111.170 169.225 112.380 170.315 ;
        RECT 18.165 169.055 112.465 169.225 ;
        RECT 18.250 167.965 19.460 169.055 ;
        RECT 18.250 167.255 18.770 167.795 ;
        RECT 18.940 167.425 19.460 167.965 ;
        RECT 20.090 167.965 21.760 169.055 ;
        RECT 20.090 167.445 20.840 167.965 ;
        RECT 21.970 167.915 22.200 169.055 ;
        RECT 22.370 167.905 22.700 168.885 ;
        RECT 22.870 167.915 23.080 169.055 ;
        RECT 23.310 167.980 23.580 168.885 ;
        RECT 23.750 168.295 24.080 169.055 ;
        RECT 24.260 168.125 24.430 168.885 ;
        RECT 21.010 167.275 21.760 167.795 ;
        RECT 21.950 167.495 22.280 167.745 ;
        RECT 18.250 166.505 19.460 167.255 ;
        RECT 20.090 166.505 21.760 167.275 ;
        RECT 21.970 166.505 22.200 167.325 ;
        RECT 22.450 167.305 22.700 167.905 ;
        RECT 22.370 166.675 22.700 167.305 ;
        RECT 22.870 166.505 23.080 167.325 ;
        RECT 23.310 167.180 23.480 167.980 ;
        RECT 23.765 167.955 24.430 168.125 ;
        RECT 23.765 167.810 23.935 167.955 ;
        RECT 23.650 167.480 23.935 167.810 ;
        RECT 24.695 167.915 25.030 168.885 ;
        RECT 25.200 167.915 25.370 169.055 ;
        RECT 25.540 168.715 27.570 168.885 ;
        RECT 23.765 167.225 23.935 167.480 ;
        RECT 24.170 167.405 24.500 167.775 ;
        RECT 24.695 167.245 24.865 167.915 ;
        RECT 25.540 167.745 25.710 168.715 ;
        RECT 25.035 167.415 25.290 167.745 ;
        RECT 25.515 167.415 25.710 167.745 ;
        RECT 25.880 168.375 27.005 168.545 ;
        RECT 25.120 167.245 25.290 167.415 ;
        RECT 25.880 167.245 26.050 168.375 ;
        RECT 23.310 166.675 23.570 167.180 ;
        RECT 23.765 167.055 24.430 167.225 ;
        RECT 23.750 166.505 24.080 166.885 ;
        RECT 24.260 166.675 24.430 167.055 ;
        RECT 24.695 166.675 24.950 167.245 ;
        RECT 25.120 167.075 26.050 167.245 ;
        RECT 26.220 168.035 27.230 168.205 ;
        RECT 26.220 167.235 26.390 168.035 ;
        RECT 25.875 167.040 26.050 167.075 ;
        RECT 25.120 166.505 25.450 166.905 ;
        RECT 25.875 166.675 26.405 167.040 ;
        RECT 26.595 167.015 26.870 167.835 ;
        RECT 26.590 166.845 26.870 167.015 ;
        RECT 26.595 166.675 26.870 166.845 ;
        RECT 27.040 166.675 27.230 168.035 ;
        RECT 27.400 168.050 27.570 168.715 ;
        RECT 27.740 168.295 27.910 169.055 ;
        RECT 28.145 168.295 28.660 168.705 ;
        RECT 27.400 167.860 28.150 168.050 ;
        RECT 28.320 167.485 28.660 168.295 ;
        RECT 28.920 168.125 29.090 168.885 ;
        RECT 29.270 168.295 29.600 169.055 ;
        RECT 28.920 167.955 29.585 168.125 ;
        RECT 29.770 167.980 30.040 168.885 ;
        RECT 29.415 167.810 29.585 167.955 ;
        RECT 27.430 167.315 28.660 167.485 ;
        RECT 28.850 167.405 29.180 167.775 ;
        RECT 29.415 167.480 29.700 167.810 ;
        RECT 27.410 166.505 27.920 167.040 ;
        RECT 28.140 166.710 28.385 167.315 ;
        RECT 29.415 167.225 29.585 167.480 ;
        RECT 28.920 167.055 29.585 167.225 ;
        RECT 29.870 167.180 30.040 167.980 ;
        RECT 31.335 168.085 31.665 168.885 ;
        RECT 31.835 168.255 32.165 169.055 ;
        RECT 32.465 168.085 32.795 168.885 ;
        RECT 33.440 168.255 33.690 169.055 ;
        RECT 31.335 167.915 33.770 168.085 ;
        RECT 33.960 167.915 34.130 169.055 ;
        RECT 34.300 167.915 34.640 168.885 ;
        RECT 31.130 167.495 31.480 167.745 ;
        RECT 31.665 167.285 31.835 167.915 ;
        RECT 32.005 167.495 32.335 167.695 ;
        RECT 32.505 167.495 32.835 167.695 ;
        RECT 33.005 167.495 33.425 167.695 ;
        RECT 33.600 167.665 33.770 167.915 ;
        RECT 33.600 167.495 34.295 167.665 ;
        RECT 34.465 167.355 34.640 167.915 ;
        RECT 34.810 167.890 35.100 169.055 ;
        RECT 35.270 167.915 35.610 168.885 ;
        RECT 35.780 167.915 35.950 169.055 ;
        RECT 36.220 168.255 36.470 169.055 ;
        RECT 37.115 168.085 37.445 168.885 ;
        RECT 37.745 168.255 38.075 169.055 ;
        RECT 38.245 168.085 38.575 168.885 ;
        RECT 36.140 167.915 38.575 168.085 ;
        RECT 38.990 167.915 39.220 169.055 ;
        RECT 28.920 166.675 29.090 167.055 ;
        RECT 29.270 166.505 29.600 166.885 ;
        RECT 29.780 166.675 30.040 167.180 ;
        RECT 31.335 166.675 31.835 167.285 ;
        RECT 32.465 167.155 33.690 167.325 ;
        RECT 34.410 167.305 34.640 167.355 ;
        RECT 32.465 166.675 32.795 167.155 ;
        RECT 32.965 166.505 33.190 166.965 ;
        RECT 33.360 166.675 33.690 167.155 ;
        RECT 33.880 166.505 34.130 167.305 ;
        RECT 34.300 166.675 34.640 167.305 ;
        RECT 35.270 167.305 35.445 167.915 ;
        RECT 36.140 167.665 36.310 167.915 ;
        RECT 35.615 167.495 36.310 167.665 ;
        RECT 36.485 167.495 36.905 167.695 ;
        RECT 37.075 167.495 37.405 167.695 ;
        RECT 37.575 167.495 37.905 167.695 ;
        RECT 34.810 166.505 35.100 167.230 ;
        RECT 35.270 166.675 35.610 167.305 ;
        RECT 35.780 166.505 36.030 167.305 ;
        RECT 36.220 167.155 37.445 167.325 ;
        RECT 36.220 166.675 36.550 167.155 ;
        RECT 36.720 166.505 36.945 166.965 ;
        RECT 37.115 166.675 37.445 167.155 ;
        RECT 38.075 167.285 38.245 167.915 ;
        RECT 39.390 167.905 39.720 168.885 ;
        RECT 39.890 167.915 40.100 169.055 ;
        RECT 40.535 168.085 40.865 168.885 ;
        RECT 41.035 168.255 41.365 169.055 ;
        RECT 41.665 168.085 41.995 168.885 ;
        RECT 42.640 168.255 42.890 169.055 ;
        RECT 40.535 167.915 42.970 168.085 ;
        RECT 43.160 167.915 43.330 169.055 ;
        RECT 43.500 167.915 43.840 168.885 ;
        RECT 38.430 167.495 38.780 167.745 ;
        RECT 38.970 167.495 39.300 167.745 ;
        RECT 38.075 166.675 38.575 167.285 ;
        RECT 38.990 166.505 39.220 167.325 ;
        RECT 39.470 167.305 39.720 167.905 ;
        RECT 40.330 167.495 40.680 167.745 ;
        RECT 39.390 166.675 39.720 167.305 ;
        RECT 39.890 166.505 40.100 167.325 ;
        RECT 40.865 167.285 41.035 167.915 ;
        RECT 41.205 167.495 41.535 167.695 ;
        RECT 41.705 167.495 42.035 167.695 ;
        RECT 42.205 167.495 42.625 167.695 ;
        RECT 42.800 167.665 42.970 167.915 ;
        RECT 42.800 167.495 43.495 167.665 ;
        RECT 40.535 166.675 41.035 167.285 ;
        RECT 41.665 167.155 42.890 167.325 ;
        RECT 43.665 167.305 43.840 167.915 ;
        RECT 41.665 166.675 41.995 167.155 ;
        RECT 42.165 166.505 42.390 166.965 ;
        RECT 42.560 166.675 42.890 167.155 ;
        RECT 43.080 166.505 43.330 167.305 ;
        RECT 43.500 166.675 43.840 167.305 ;
        RECT 44.010 167.915 44.395 168.885 ;
        RECT 44.565 168.595 44.890 169.055 ;
        RECT 45.410 168.425 45.690 168.885 ;
        RECT 44.565 168.205 45.690 168.425 ;
        RECT 44.010 167.245 44.290 167.915 ;
        RECT 44.565 167.745 45.015 168.205 ;
        RECT 45.880 168.035 46.280 168.885 ;
        RECT 46.680 168.595 46.950 169.055 ;
        RECT 47.120 168.425 47.405 168.885 ;
        RECT 44.460 167.415 45.015 167.745 ;
        RECT 45.185 167.475 46.280 168.035 ;
        RECT 44.565 167.305 45.015 167.415 ;
        RECT 44.010 166.675 44.395 167.245 ;
        RECT 44.565 167.135 45.690 167.305 ;
        RECT 44.565 166.505 44.890 166.965 ;
        RECT 45.410 166.675 45.690 167.135 ;
        RECT 45.880 166.675 46.280 167.475 ;
        RECT 46.450 168.205 47.405 168.425 ;
        RECT 46.450 167.305 46.660 168.205 ;
        RECT 47.895 168.085 48.225 168.885 ;
        RECT 48.395 168.255 48.725 169.055 ;
        RECT 49.025 168.085 49.355 168.885 ;
        RECT 50.000 168.255 50.250 169.055 ;
        RECT 46.830 167.475 47.520 168.035 ;
        RECT 47.895 167.915 50.330 168.085 ;
        RECT 50.520 167.915 50.690 169.055 ;
        RECT 50.860 167.915 51.200 168.885 ;
        RECT 47.690 167.495 48.040 167.745 ;
        RECT 46.450 167.135 47.405 167.305 ;
        RECT 48.225 167.285 48.395 167.915 ;
        RECT 48.565 167.495 48.895 167.695 ;
        RECT 49.065 167.495 49.395 167.695 ;
        RECT 49.565 167.495 49.985 167.695 ;
        RECT 50.160 167.665 50.330 167.915 ;
        RECT 50.160 167.495 50.855 167.665 ;
        RECT 46.680 166.505 46.950 166.965 ;
        RECT 47.120 166.675 47.405 167.135 ;
        RECT 47.895 166.675 48.395 167.285 ;
        RECT 49.025 167.155 50.250 167.325 ;
        RECT 51.025 167.305 51.200 167.915 ;
        RECT 52.290 167.965 55.800 169.055 ;
        RECT 52.290 167.445 53.980 167.965 ;
        RECT 55.975 167.905 56.235 169.055 ;
        RECT 56.410 167.980 56.665 168.885 ;
        RECT 56.835 168.295 57.165 169.055 ;
        RECT 57.380 168.125 57.550 168.885 ;
        RECT 49.025 166.675 49.355 167.155 ;
        RECT 49.525 166.505 49.750 166.965 ;
        RECT 49.920 166.675 50.250 167.155 ;
        RECT 50.440 166.505 50.690 167.305 ;
        RECT 50.860 166.675 51.200 167.305 ;
        RECT 54.150 167.275 55.800 167.795 ;
        RECT 52.290 166.505 55.800 167.275 ;
        RECT 55.975 166.505 56.235 167.345 ;
        RECT 56.410 167.250 56.580 167.980 ;
        RECT 56.835 167.955 57.550 168.125 ;
        RECT 57.820 167.995 58.150 169.055 ;
        RECT 56.835 167.745 57.005 167.955 ;
        RECT 56.750 167.415 57.005 167.745 ;
        RECT 56.410 166.675 56.665 167.250 ;
        RECT 56.835 167.225 57.005 167.415 ;
        RECT 57.285 167.405 57.640 167.775 ;
        RECT 58.330 167.745 58.500 168.715 ;
        RECT 58.670 168.465 59.000 168.865 ;
        RECT 59.170 168.695 59.500 169.055 ;
        RECT 59.700 168.465 60.400 168.885 ;
        RECT 58.670 168.235 60.400 168.465 ;
        RECT 58.670 168.015 59.000 168.235 ;
        RECT 59.195 167.745 59.520 168.035 ;
        RECT 57.810 167.415 58.120 167.745 ;
        RECT 58.330 167.415 58.705 167.745 ;
        RECT 59.025 167.415 59.520 167.745 ;
        RECT 59.695 167.495 60.025 168.035 ;
        RECT 60.195 167.265 60.400 168.235 ;
        RECT 60.570 167.890 60.860 169.055 ;
        RECT 62.660 168.605 62.990 169.055 ;
        RECT 61.950 168.215 64.560 168.425 ;
        RECT 56.835 167.055 57.550 167.225 ;
        RECT 56.835 166.505 57.165 166.885 ;
        RECT 57.380 166.675 57.550 167.055 ;
        RECT 57.820 167.035 59.180 167.245 ;
        RECT 57.820 166.675 58.150 167.035 ;
        RECT 58.320 166.505 58.650 166.865 ;
        RECT 58.850 166.675 59.180 167.035 ;
        RECT 59.690 166.675 60.400 167.265 ;
        RECT 61.950 167.245 62.120 168.215 ;
        RECT 62.290 167.415 62.640 168.035 ;
        RECT 62.810 167.415 63.130 168.035 ;
        RECT 63.300 167.415 63.630 168.035 ;
        RECT 63.800 167.415 64.100 168.035 ;
        RECT 64.340 167.415 64.560 168.215 ;
        RECT 64.740 167.245 65.000 168.870 ;
        RECT 65.180 167.995 65.510 169.055 ;
        RECT 65.690 167.745 65.860 168.715 ;
        RECT 66.030 168.465 66.360 168.865 ;
        RECT 66.530 168.695 66.860 169.055 ;
        RECT 67.060 168.465 67.760 168.885 ;
        RECT 66.030 168.235 67.760 168.465 ;
        RECT 66.030 168.015 66.360 168.235 ;
        RECT 66.555 167.745 66.880 168.035 ;
        RECT 65.170 167.415 65.480 167.745 ;
        RECT 65.690 167.415 66.065 167.745 ;
        RECT 66.385 167.415 66.880 167.745 ;
        RECT 67.055 167.495 67.385 168.035 ;
        RECT 67.555 167.265 67.760 168.235 ;
        RECT 67.970 167.915 68.200 169.055 ;
        RECT 68.370 167.905 68.700 168.885 ;
        RECT 68.870 167.915 69.080 169.055 ;
        RECT 70.340 168.255 70.510 169.055 ;
        RECT 70.680 168.035 71.010 168.885 ;
        RECT 71.180 168.255 71.350 169.055 ;
        RECT 71.520 168.035 71.850 168.885 ;
        RECT 72.020 168.255 72.190 169.055 ;
        RECT 72.360 168.035 72.690 168.885 ;
        RECT 72.860 168.255 73.030 169.055 ;
        RECT 73.200 168.035 73.530 168.885 ;
        RECT 73.700 168.255 73.870 169.055 ;
        RECT 74.040 168.035 74.370 168.885 ;
        RECT 74.540 168.255 74.710 169.055 ;
        RECT 74.880 168.035 75.210 168.885 ;
        RECT 75.380 168.255 75.550 169.055 ;
        RECT 75.720 168.035 76.050 168.885 ;
        RECT 76.220 168.255 76.390 169.055 ;
        RECT 76.560 168.035 76.890 168.885 ;
        RECT 77.060 168.255 77.230 169.055 ;
        RECT 77.400 168.035 77.730 168.885 ;
        RECT 77.900 168.255 78.070 169.055 ;
        RECT 78.240 168.035 78.570 168.885 ;
        RECT 78.740 168.255 78.910 169.055 ;
        RECT 79.080 168.035 79.410 168.885 ;
        RECT 79.580 168.205 79.750 169.055 ;
        RECT 79.920 168.035 80.250 168.885 ;
        RECT 80.420 168.205 80.590 169.055 ;
        RECT 80.760 168.035 81.090 168.885 ;
        RECT 67.950 167.495 68.280 167.745 ;
        RECT 60.570 166.505 60.860 167.230 ;
        RECT 61.950 167.075 62.425 167.245 ;
        RECT 62.255 166.825 62.425 167.075 ;
        RECT 62.660 166.505 62.990 167.245 ;
        RECT 63.160 167.075 65.000 167.245 ;
        RECT 63.160 166.730 63.360 167.075 ;
        RECT 63.530 166.505 63.860 166.905 ;
        RECT 64.030 166.720 64.230 167.075 ;
        RECT 65.180 167.035 66.540 167.245 ;
        RECT 64.400 166.505 64.730 166.900 ;
        RECT 65.180 166.675 65.510 167.035 ;
        RECT 65.680 166.505 66.010 166.865 ;
        RECT 66.210 166.675 66.540 167.035 ;
        RECT 67.050 166.675 67.760 167.265 ;
        RECT 67.970 166.505 68.200 167.325 ;
        RECT 68.450 167.305 68.700 167.905 ;
        RECT 70.230 167.865 76.890 168.035 ;
        RECT 77.060 167.865 79.410 168.035 ;
        RECT 79.580 167.865 81.090 168.035 ;
        RECT 81.270 168.295 81.785 168.705 ;
        RECT 82.020 168.295 82.190 169.055 ;
        RECT 82.360 168.715 84.390 168.885 ;
        RECT 70.230 167.325 70.505 167.865 ;
        RECT 77.060 167.695 77.235 167.865 ;
        RECT 79.580 167.695 79.750 167.865 ;
        RECT 70.675 167.495 77.235 167.695 ;
        RECT 77.440 167.495 79.750 167.695 ;
        RECT 79.920 167.495 81.095 167.695 ;
        RECT 77.060 167.325 77.235 167.495 ;
        RECT 79.580 167.325 79.750 167.495 ;
        RECT 81.270 167.485 81.610 168.295 ;
        RECT 82.360 168.050 82.530 168.715 ;
        RECT 82.925 168.375 84.050 168.545 ;
        RECT 81.780 167.860 82.530 168.050 ;
        RECT 82.700 168.035 83.710 168.205 ;
        RECT 68.370 166.675 68.700 167.305 ;
        RECT 68.870 166.505 69.080 167.325 ;
        RECT 70.230 167.155 76.890 167.325 ;
        RECT 77.060 167.155 79.410 167.325 ;
        RECT 79.580 167.155 81.090 167.325 ;
        RECT 81.270 167.315 82.500 167.485 ;
        RECT 70.340 166.505 70.510 166.985 ;
        RECT 70.680 166.680 71.010 167.155 ;
        RECT 71.180 166.505 71.350 166.985 ;
        RECT 71.520 166.680 71.850 167.155 ;
        RECT 72.020 166.505 72.190 166.985 ;
        RECT 72.360 166.680 72.690 167.155 ;
        RECT 72.860 166.505 73.030 166.985 ;
        RECT 73.200 166.680 73.530 167.155 ;
        RECT 73.700 166.505 73.870 166.985 ;
        RECT 74.040 166.680 74.370 167.155 ;
        RECT 74.540 166.505 74.710 166.985 ;
        RECT 74.880 166.680 75.210 167.155 ;
        RECT 74.960 166.675 75.130 166.680 ;
        RECT 75.380 166.505 75.550 166.985 ;
        RECT 75.720 166.680 76.050 167.155 ;
        RECT 75.800 166.675 75.970 166.680 ;
        RECT 76.220 166.505 76.390 166.985 ;
        RECT 76.560 166.680 76.890 167.155 ;
        RECT 76.640 166.675 76.890 166.680 ;
        RECT 77.060 166.505 77.230 166.985 ;
        RECT 77.400 166.680 77.730 167.155 ;
        RECT 77.900 166.505 78.070 166.985 ;
        RECT 78.240 166.680 78.570 167.155 ;
        RECT 78.740 166.505 78.910 166.985 ;
        RECT 79.080 166.680 79.410 167.155 ;
        RECT 79.580 166.505 79.750 166.985 ;
        RECT 79.920 166.680 80.250 167.155 ;
        RECT 80.420 166.505 80.590 166.985 ;
        RECT 80.760 166.680 81.090 167.155 ;
        RECT 81.545 166.710 81.790 167.315 ;
        RECT 82.010 166.505 82.520 167.040 ;
        RECT 82.700 166.675 82.890 168.035 ;
        RECT 83.060 167.015 83.335 167.835 ;
        RECT 83.540 167.235 83.710 168.035 ;
        RECT 83.880 167.245 84.050 168.375 ;
        RECT 84.220 167.745 84.390 168.715 ;
        RECT 84.560 167.915 84.730 169.055 ;
        RECT 84.900 167.915 85.235 168.885 ;
        RECT 84.220 167.415 84.415 167.745 ;
        RECT 84.640 167.415 84.895 167.745 ;
        RECT 84.640 167.245 84.810 167.415 ;
        RECT 85.065 167.245 85.235 167.915 ;
        RECT 86.330 167.890 86.620 169.055 ;
        RECT 86.995 168.085 87.325 168.885 ;
        RECT 87.495 168.255 87.825 169.055 ;
        RECT 88.125 168.085 88.455 168.885 ;
        RECT 89.100 168.255 89.350 169.055 ;
        RECT 86.995 167.915 89.430 168.085 ;
        RECT 89.620 167.915 89.790 169.055 ;
        RECT 89.960 167.915 90.300 168.885 ;
        RECT 90.675 168.085 91.005 168.885 ;
        RECT 91.175 168.255 91.505 169.055 ;
        RECT 91.805 168.085 92.135 168.885 ;
        RECT 92.780 168.255 93.030 169.055 ;
        RECT 90.675 167.915 93.110 168.085 ;
        RECT 93.300 167.915 93.470 169.055 ;
        RECT 93.640 167.915 93.980 168.885 ;
        RECT 94.355 168.085 94.685 168.885 ;
        RECT 94.855 168.255 95.185 169.055 ;
        RECT 95.485 168.085 95.815 168.885 ;
        RECT 96.460 168.255 96.710 169.055 ;
        RECT 94.355 167.915 96.790 168.085 ;
        RECT 96.980 167.915 97.150 169.055 ;
        RECT 97.320 167.915 97.660 168.885 ;
        RECT 86.790 167.495 87.140 167.745 ;
        RECT 87.325 167.285 87.495 167.915 ;
        RECT 87.665 167.495 87.995 167.695 ;
        RECT 88.165 167.495 88.495 167.695 ;
        RECT 88.665 167.495 89.085 167.695 ;
        RECT 89.260 167.665 89.430 167.915 ;
        RECT 89.260 167.495 89.955 167.665 ;
        RECT 83.880 167.075 84.810 167.245 ;
        RECT 83.880 167.040 84.055 167.075 ;
        RECT 83.060 166.845 83.340 167.015 ;
        RECT 83.060 166.675 83.335 166.845 ;
        RECT 83.525 166.675 84.055 167.040 ;
        RECT 84.480 166.505 84.810 166.905 ;
        RECT 84.980 166.675 85.235 167.245 ;
        RECT 86.330 166.505 86.620 167.230 ;
        RECT 86.995 166.675 87.495 167.285 ;
        RECT 88.125 167.155 89.350 167.325 ;
        RECT 90.125 167.305 90.300 167.915 ;
        RECT 90.470 167.495 90.820 167.745 ;
        RECT 88.125 166.675 88.455 167.155 ;
        RECT 88.625 166.505 88.850 166.965 ;
        RECT 89.020 166.675 89.350 167.155 ;
        RECT 89.540 166.505 89.790 167.305 ;
        RECT 89.960 166.675 90.300 167.305 ;
        RECT 91.005 167.285 91.175 167.915 ;
        RECT 91.345 167.495 91.675 167.695 ;
        RECT 91.845 167.495 92.175 167.695 ;
        RECT 92.345 167.495 92.765 167.695 ;
        RECT 92.940 167.665 93.110 167.915 ;
        RECT 92.940 167.495 93.635 167.665 ;
        RECT 90.675 166.675 91.175 167.285 ;
        RECT 91.805 167.155 93.030 167.325 ;
        RECT 93.805 167.305 93.980 167.915 ;
        RECT 94.150 167.495 94.500 167.745 ;
        RECT 91.805 166.675 92.135 167.155 ;
        RECT 92.305 166.505 92.530 166.965 ;
        RECT 92.700 166.675 93.030 167.155 ;
        RECT 93.220 166.505 93.470 167.305 ;
        RECT 93.640 166.675 93.980 167.305 ;
        RECT 94.685 167.285 94.855 167.915 ;
        RECT 95.025 167.495 95.355 167.695 ;
        RECT 95.525 167.495 95.855 167.695 ;
        RECT 96.025 167.495 96.445 167.695 ;
        RECT 96.620 167.665 96.790 167.915 ;
        RECT 96.620 167.495 97.315 167.665 ;
        RECT 94.355 166.675 94.855 167.285 ;
        RECT 95.485 167.155 96.710 167.325 ;
        RECT 97.485 167.305 97.660 167.915 ;
        RECT 98.290 167.965 100.880 169.055 ;
        RECT 101.050 168.295 101.565 168.705 ;
        RECT 101.800 168.295 101.970 169.055 ;
        RECT 102.140 168.715 104.170 168.885 ;
        RECT 98.290 167.445 99.500 167.965 ;
        RECT 95.485 166.675 95.815 167.155 ;
        RECT 95.985 166.505 96.210 166.965 ;
        RECT 96.380 166.675 96.710 167.155 ;
        RECT 96.900 166.505 97.150 167.305 ;
        RECT 97.320 166.675 97.660 167.305 ;
        RECT 99.670 167.275 100.880 167.795 ;
        RECT 101.050 167.485 101.390 168.295 ;
        RECT 102.140 168.050 102.310 168.715 ;
        RECT 102.705 168.375 103.830 168.545 ;
        RECT 101.560 167.860 102.310 168.050 ;
        RECT 102.480 168.035 103.490 168.205 ;
        RECT 101.050 167.315 102.280 167.485 ;
        RECT 98.290 166.505 100.880 167.275 ;
        RECT 101.325 166.710 101.570 167.315 ;
        RECT 101.790 166.505 102.300 167.040 ;
        RECT 102.480 166.675 102.670 168.035 ;
        RECT 102.840 167.015 103.115 167.835 ;
        RECT 103.320 167.235 103.490 168.035 ;
        RECT 103.660 167.245 103.830 168.375 ;
        RECT 104.000 167.745 104.170 168.715 ;
        RECT 104.340 167.915 104.510 169.055 ;
        RECT 104.680 167.915 105.015 168.885 ;
        RECT 105.740 168.125 105.910 168.885 ;
        RECT 106.090 168.295 106.420 169.055 ;
        RECT 105.740 167.955 106.405 168.125 ;
        RECT 106.590 167.980 106.860 168.885 ;
        RECT 104.000 167.415 104.195 167.745 ;
        RECT 104.420 167.415 104.675 167.745 ;
        RECT 104.420 167.245 104.590 167.415 ;
        RECT 104.845 167.245 105.015 167.915 ;
        RECT 106.235 167.810 106.405 167.955 ;
        RECT 105.670 167.405 106.000 167.775 ;
        RECT 106.235 167.480 106.520 167.810 ;
        RECT 103.660 167.075 104.590 167.245 ;
        RECT 103.660 167.040 103.835 167.075 ;
        RECT 102.840 166.845 103.120 167.015 ;
        RECT 102.840 166.675 103.115 166.845 ;
        RECT 103.305 166.675 103.835 167.040 ;
        RECT 104.260 166.505 104.590 166.905 ;
        RECT 104.760 166.675 105.015 167.245 ;
        RECT 106.235 167.225 106.405 167.480 ;
        RECT 105.740 167.055 106.405 167.225 ;
        RECT 106.690 167.180 106.860 167.980 ;
        RECT 107.490 167.965 111.000 169.055 ;
        RECT 111.170 167.965 112.380 169.055 ;
        RECT 107.490 167.445 109.180 167.965 ;
        RECT 109.350 167.275 111.000 167.795 ;
        RECT 111.170 167.425 111.690 167.965 ;
        RECT 105.740 166.675 105.910 167.055 ;
        RECT 106.090 166.505 106.420 166.885 ;
        RECT 106.600 166.675 106.860 167.180 ;
        RECT 107.490 166.505 111.000 167.275 ;
        RECT 111.860 167.255 112.380 167.795 ;
        RECT 111.170 166.505 112.380 167.255 ;
        RECT 18.165 166.335 112.465 166.505 ;
        RECT 18.250 165.585 19.460 166.335 ;
        RECT 18.250 165.045 18.770 165.585 ;
        RECT 20.090 165.565 21.760 166.335 ;
        RECT 21.930 165.610 22.220 166.335 ;
        RECT 22.395 165.625 22.650 166.155 ;
        RECT 22.820 165.875 23.125 166.335 ;
        RECT 23.370 165.955 24.440 166.125 ;
        RECT 18.940 164.875 19.460 165.415 ;
        RECT 18.250 163.785 19.460 164.875 ;
        RECT 20.090 164.875 20.840 165.395 ;
        RECT 21.010 165.045 21.760 165.565 ;
        RECT 22.395 164.975 22.605 165.625 ;
        RECT 23.370 165.600 23.690 165.955 ;
        RECT 23.365 165.425 23.690 165.600 ;
        RECT 22.775 165.125 23.690 165.425 ;
        RECT 23.860 165.385 24.100 165.785 ;
        RECT 24.270 165.725 24.440 165.955 ;
        RECT 24.610 165.895 24.800 166.335 ;
        RECT 24.970 165.885 25.920 166.165 ;
        RECT 26.140 165.975 26.490 166.145 ;
        RECT 24.270 165.555 24.800 165.725 ;
        RECT 22.775 165.095 23.515 165.125 ;
        RECT 20.090 163.785 21.760 164.875 ;
        RECT 21.930 163.785 22.220 164.950 ;
        RECT 22.395 164.095 22.650 164.975 ;
        RECT 22.820 163.785 23.125 164.925 ;
        RECT 23.345 164.505 23.515 165.095 ;
        RECT 23.860 165.015 24.400 165.385 ;
        RECT 24.580 165.275 24.800 165.555 ;
        RECT 24.970 165.105 25.140 165.885 ;
        RECT 24.735 164.935 25.140 165.105 ;
        RECT 25.310 165.095 25.660 165.715 ;
        RECT 24.735 164.845 24.905 164.935 ;
        RECT 25.830 164.925 26.040 165.715 ;
        RECT 23.685 164.675 24.905 164.845 ;
        RECT 25.365 164.765 26.040 164.925 ;
        RECT 23.345 164.335 24.145 164.505 ;
        RECT 23.465 163.785 23.795 164.165 ;
        RECT 23.975 164.045 24.145 164.335 ;
        RECT 24.735 164.295 24.905 164.675 ;
        RECT 25.075 164.755 26.040 164.765 ;
        RECT 26.230 165.585 26.490 165.975 ;
        RECT 26.700 165.875 27.030 166.335 ;
        RECT 27.905 165.945 28.760 166.115 ;
        RECT 28.965 165.945 29.460 166.115 ;
        RECT 29.630 165.975 29.960 166.335 ;
        RECT 26.230 164.895 26.400 165.585 ;
        RECT 26.570 165.235 26.740 165.415 ;
        RECT 26.910 165.405 27.700 165.655 ;
        RECT 27.905 165.235 28.075 165.945 ;
        RECT 28.245 165.435 28.600 165.655 ;
        RECT 26.570 165.065 28.260 165.235 ;
        RECT 25.075 164.465 25.535 164.755 ;
        RECT 26.230 164.725 27.730 164.895 ;
        RECT 26.230 164.585 26.400 164.725 ;
        RECT 25.840 164.415 26.400 164.585 ;
        RECT 24.315 163.785 24.565 164.245 ;
        RECT 24.735 163.955 25.605 164.295 ;
        RECT 25.840 163.955 26.010 164.415 ;
        RECT 26.845 164.385 27.920 164.555 ;
        RECT 26.180 163.785 26.550 164.245 ;
        RECT 26.845 164.045 27.015 164.385 ;
        RECT 27.185 163.785 27.515 164.215 ;
        RECT 27.750 164.045 27.920 164.385 ;
        RECT 28.090 164.285 28.260 165.065 ;
        RECT 28.430 164.845 28.600 165.435 ;
        RECT 28.770 165.035 29.120 165.655 ;
        RECT 28.430 164.455 28.895 164.845 ;
        RECT 29.290 164.585 29.460 165.945 ;
        RECT 29.630 164.755 30.090 165.805 ;
        RECT 29.065 164.415 29.460 164.585 ;
        RECT 29.065 164.285 29.235 164.415 ;
        RECT 28.090 163.955 28.770 164.285 ;
        RECT 28.985 163.955 29.235 164.285 ;
        RECT 29.405 163.785 29.655 164.245 ;
        RECT 29.825 163.970 30.150 164.755 ;
        RECT 30.320 163.955 30.490 166.075 ;
        RECT 30.660 165.955 30.990 166.335 ;
        RECT 31.160 165.785 31.415 166.075 ;
        RECT 30.665 165.615 31.415 165.785 ;
        RECT 30.665 164.625 30.895 165.615 ;
        RECT 31.590 165.585 32.800 166.335 ;
        RECT 31.065 164.795 31.415 165.445 ;
        RECT 31.590 164.875 32.110 165.415 ;
        RECT 32.280 165.045 32.800 165.585 ;
        RECT 33.245 165.525 33.490 166.130 ;
        RECT 33.710 165.800 34.220 166.335 ;
        RECT 32.970 165.355 34.200 165.525 ;
        RECT 30.665 164.455 31.415 164.625 ;
        RECT 30.660 163.785 30.990 164.285 ;
        RECT 31.160 163.955 31.415 164.455 ;
        RECT 31.590 163.785 32.800 164.875 ;
        RECT 32.970 164.545 33.310 165.355 ;
        RECT 33.480 164.790 34.230 164.980 ;
        RECT 32.970 164.135 33.485 164.545 ;
        RECT 33.720 163.785 33.890 164.545 ;
        RECT 34.060 164.125 34.230 164.790 ;
        RECT 34.400 164.805 34.590 166.165 ;
        RECT 34.760 165.655 35.035 166.165 ;
        RECT 35.225 165.800 35.755 166.165 ;
        RECT 36.180 165.935 36.510 166.335 ;
        RECT 35.580 165.765 35.755 165.800 ;
        RECT 34.760 165.485 35.040 165.655 ;
        RECT 34.760 165.005 35.035 165.485 ;
        RECT 35.240 164.805 35.410 165.605 ;
        RECT 34.400 164.635 35.410 164.805 ;
        RECT 35.580 165.595 36.510 165.765 ;
        RECT 36.680 165.595 36.935 166.165 ;
        RECT 35.580 164.465 35.750 165.595 ;
        RECT 36.340 165.425 36.510 165.595 ;
        RECT 34.625 164.295 35.750 164.465 ;
        RECT 35.920 165.095 36.115 165.425 ;
        RECT 36.340 165.095 36.595 165.425 ;
        RECT 35.920 164.125 36.090 165.095 ;
        RECT 36.765 164.925 36.935 165.595 ;
        RECT 34.060 163.955 36.090 164.125 ;
        RECT 36.260 163.785 36.430 164.925 ;
        RECT 36.600 163.955 36.935 164.925 ;
        RECT 37.485 165.625 37.740 166.155 ;
        RECT 37.920 165.875 38.205 166.335 ;
        RECT 37.485 164.765 37.665 165.625 ;
        RECT 38.385 165.425 38.635 166.075 ;
        RECT 37.835 165.095 38.635 165.425 ;
        RECT 37.485 164.635 37.740 164.765 ;
        RECT 37.400 164.465 37.740 164.635 ;
        RECT 37.485 164.095 37.740 164.465 ;
        RECT 37.920 163.785 38.205 164.585 ;
        RECT 38.385 164.505 38.635 165.095 ;
        RECT 38.835 165.740 39.155 166.070 ;
        RECT 39.335 165.855 39.995 166.335 ;
        RECT 40.195 165.945 41.045 166.115 ;
        RECT 38.835 164.845 39.025 165.740 ;
        RECT 39.345 165.415 40.005 165.685 ;
        RECT 39.675 165.355 40.005 165.415 ;
        RECT 39.195 165.185 39.525 165.245 ;
        RECT 40.195 165.185 40.365 165.945 ;
        RECT 41.605 165.875 41.925 166.335 ;
        RECT 42.125 165.695 42.375 166.125 ;
        RECT 42.665 165.895 43.075 166.335 ;
        RECT 43.245 165.955 44.260 166.155 ;
        RECT 40.535 165.525 41.785 165.695 ;
        RECT 40.535 165.405 40.865 165.525 ;
        RECT 39.195 165.015 41.095 165.185 ;
        RECT 38.835 164.675 40.755 164.845 ;
        RECT 38.835 164.655 39.155 164.675 ;
        RECT 38.385 163.995 38.715 164.505 ;
        RECT 38.985 164.045 39.155 164.655 ;
        RECT 40.925 164.505 41.095 165.015 ;
        RECT 41.265 164.945 41.445 165.355 ;
        RECT 41.615 164.765 41.785 165.525 ;
        RECT 39.325 163.785 39.655 164.475 ;
        RECT 39.885 164.335 41.095 164.505 ;
        RECT 41.265 164.455 41.785 164.765 ;
        RECT 41.955 165.355 42.375 165.695 ;
        RECT 42.665 165.355 43.075 165.685 ;
        RECT 41.955 164.585 42.145 165.355 ;
        RECT 43.245 165.225 43.415 165.955 ;
        RECT 44.560 165.785 44.730 166.115 ;
        RECT 44.900 165.955 45.230 166.335 ;
        RECT 43.585 165.405 43.935 165.775 ;
        RECT 43.245 165.185 43.665 165.225 ;
        RECT 42.315 165.015 43.665 165.185 ;
        RECT 42.315 164.855 42.565 165.015 ;
        RECT 43.075 164.585 43.325 164.845 ;
        RECT 41.955 164.335 43.325 164.585 ;
        RECT 39.885 164.045 40.125 164.335 ;
        RECT 40.925 164.255 41.095 164.335 ;
        RECT 40.325 163.785 40.745 164.165 ;
        RECT 40.925 164.005 41.555 164.255 ;
        RECT 42.025 163.785 42.355 164.165 ;
        RECT 42.525 164.045 42.695 164.335 ;
        RECT 43.495 164.170 43.665 165.015 ;
        RECT 44.115 164.845 44.335 165.715 ;
        RECT 44.560 165.595 45.255 165.785 ;
        RECT 43.835 164.465 44.335 164.845 ;
        RECT 44.505 164.795 44.915 165.415 ;
        RECT 45.085 164.625 45.255 165.595 ;
        RECT 44.560 164.455 45.255 164.625 ;
        RECT 42.875 163.785 43.255 164.165 ;
        RECT 43.495 164.000 44.325 164.170 ;
        RECT 44.560 163.955 44.730 164.455 ;
        RECT 44.900 163.785 45.230 164.285 ;
        RECT 45.445 163.955 45.670 166.075 ;
        RECT 45.840 165.955 46.170 166.335 ;
        RECT 46.340 165.785 46.510 166.075 ;
        RECT 45.845 165.615 46.510 165.785 ;
        RECT 45.845 164.625 46.075 165.615 ;
        RECT 47.690 165.610 47.980 166.335 ;
        RECT 48.150 165.660 48.410 166.165 ;
        RECT 48.590 165.955 48.920 166.335 ;
        RECT 49.100 165.785 49.270 166.165 ;
        RECT 46.245 164.795 46.595 165.445 ;
        RECT 45.845 164.455 46.510 164.625 ;
        RECT 45.840 163.785 46.170 164.285 ;
        RECT 46.340 163.955 46.510 164.455 ;
        RECT 47.690 163.785 47.980 164.950 ;
        RECT 48.150 164.860 48.320 165.660 ;
        RECT 48.605 165.615 49.270 165.785 ;
        RECT 48.605 165.360 48.775 165.615 ;
        RECT 49.570 165.515 49.800 166.335 ;
        RECT 49.970 165.535 50.300 166.165 ;
        RECT 48.490 165.030 48.775 165.360 ;
        RECT 49.010 165.065 49.340 165.435 ;
        RECT 49.550 165.095 49.880 165.345 ;
        RECT 48.605 164.885 48.775 165.030 ;
        RECT 50.050 164.935 50.300 165.535 ;
        RECT 50.470 165.515 50.680 166.335 ;
        RECT 51.185 165.525 51.430 166.130 ;
        RECT 51.650 165.800 52.160 166.335 ;
        RECT 48.150 163.955 48.420 164.860 ;
        RECT 48.605 164.715 49.270 164.885 ;
        RECT 48.590 163.785 48.920 164.545 ;
        RECT 49.100 163.955 49.270 164.715 ;
        RECT 49.570 163.785 49.800 164.925 ;
        RECT 49.970 163.955 50.300 164.935 ;
        RECT 50.910 165.355 52.140 165.525 ;
        RECT 50.470 163.785 50.680 164.925 ;
        RECT 50.910 164.545 51.250 165.355 ;
        RECT 51.420 164.790 52.170 164.980 ;
        RECT 50.910 164.135 51.425 164.545 ;
        RECT 51.660 163.785 51.830 164.545 ;
        RECT 52.000 164.125 52.170 164.790 ;
        RECT 52.340 164.805 52.530 166.165 ;
        RECT 52.700 165.995 52.975 166.165 ;
        RECT 52.700 165.825 52.980 165.995 ;
        RECT 52.700 165.005 52.975 165.825 ;
        RECT 53.165 165.800 53.695 166.165 ;
        RECT 54.120 165.935 54.450 166.335 ;
        RECT 53.520 165.765 53.695 165.800 ;
        RECT 53.180 164.805 53.350 165.605 ;
        RECT 52.340 164.635 53.350 164.805 ;
        RECT 53.520 165.595 54.450 165.765 ;
        RECT 54.620 165.595 54.875 166.165 ;
        RECT 56.060 165.785 56.230 166.165 ;
        RECT 56.410 165.955 56.740 166.335 ;
        RECT 56.060 165.615 56.725 165.785 ;
        RECT 56.920 165.660 57.180 166.165 ;
        RECT 53.520 164.465 53.690 165.595 ;
        RECT 54.280 165.425 54.450 165.595 ;
        RECT 52.565 164.295 53.690 164.465 ;
        RECT 53.860 165.095 54.055 165.425 ;
        RECT 54.280 165.095 54.535 165.425 ;
        RECT 53.860 164.125 54.030 165.095 ;
        RECT 54.705 164.925 54.875 165.595 ;
        RECT 55.990 165.065 56.320 165.435 ;
        RECT 56.555 165.360 56.725 165.615 ;
        RECT 52.000 163.955 54.030 164.125 ;
        RECT 54.200 163.785 54.370 164.925 ;
        RECT 54.540 163.955 54.875 164.925 ;
        RECT 56.555 165.030 56.840 165.360 ;
        RECT 56.555 164.885 56.725 165.030 ;
        RECT 56.060 164.715 56.725 164.885 ;
        RECT 57.010 164.860 57.180 165.660 ;
        RECT 57.440 165.785 57.610 166.165 ;
        RECT 57.825 165.955 58.155 166.335 ;
        RECT 57.440 165.615 58.155 165.785 ;
        RECT 57.350 165.065 57.705 165.435 ;
        RECT 57.985 165.425 58.155 165.615 ;
        RECT 58.325 165.590 58.580 166.165 ;
        RECT 57.985 165.095 58.240 165.425 ;
        RECT 57.985 164.885 58.155 165.095 ;
        RECT 56.060 163.955 56.230 164.715 ;
        RECT 56.410 163.785 56.740 164.545 ;
        RECT 56.910 163.955 57.180 164.860 ;
        RECT 57.440 164.715 58.155 164.885 ;
        RECT 58.410 164.860 58.580 165.590 ;
        RECT 58.755 165.495 59.015 166.335 ;
        RECT 59.280 165.785 59.450 166.165 ;
        RECT 59.665 165.955 59.995 166.335 ;
        RECT 59.280 165.615 59.995 165.785 ;
        RECT 59.190 165.065 59.545 165.435 ;
        RECT 59.825 165.425 59.995 165.615 ;
        RECT 60.165 165.590 60.420 166.165 ;
        RECT 59.825 165.095 60.080 165.425 ;
        RECT 57.440 163.955 57.610 164.715 ;
        RECT 57.825 163.785 58.155 164.545 ;
        RECT 58.325 163.955 58.580 164.860 ;
        RECT 58.755 163.785 59.015 164.935 ;
        RECT 59.825 164.885 59.995 165.095 ;
        RECT 59.280 164.715 59.995 164.885 ;
        RECT 60.250 164.860 60.420 165.590 ;
        RECT 60.595 165.495 60.855 166.335 ;
        RECT 61.090 165.855 61.370 166.335 ;
        RECT 61.540 165.685 61.800 166.075 ;
        RECT 61.975 165.855 62.230 166.335 ;
        RECT 62.400 165.685 62.695 166.075 ;
        RECT 62.875 165.855 63.150 166.335 ;
        RECT 63.320 165.835 63.620 166.165 ;
        RECT 61.045 165.515 62.695 165.685 ;
        RECT 61.045 165.005 61.450 165.515 ;
        RECT 61.620 165.175 62.760 165.345 ;
        RECT 59.280 163.955 59.450 164.715 ;
        RECT 59.665 163.785 59.995 164.545 ;
        RECT 60.165 163.955 60.420 164.860 ;
        RECT 60.595 163.785 60.855 164.935 ;
        RECT 61.045 164.835 61.800 165.005 ;
        RECT 61.085 163.785 61.370 164.655 ;
        RECT 61.540 164.585 61.800 164.835 ;
        RECT 62.590 164.925 62.760 165.175 ;
        RECT 62.930 165.095 63.280 165.665 ;
        RECT 63.450 164.925 63.620 165.835 ;
        RECT 62.590 164.755 63.620 164.925 ;
        RECT 61.540 164.415 62.660 164.585 ;
        RECT 61.540 163.955 61.800 164.415 ;
        RECT 61.975 163.785 62.230 164.245 ;
        RECT 62.400 163.955 62.660 164.415 ;
        RECT 62.830 163.785 63.140 164.585 ;
        RECT 63.310 163.955 63.620 164.755 ;
        RECT 63.790 165.660 64.050 166.165 ;
        RECT 64.230 165.955 64.560 166.335 ;
        RECT 64.740 165.785 64.910 166.165 ;
        RECT 63.790 164.860 63.960 165.660 ;
        RECT 64.245 165.615 64.910 165.785 ;
        RECT 64.245 165.360 64.415 165.615 ;
        RECT 65.835 165.555 66.335 166.165 ;
        RECT 64.130 165.030 64.415 165.360 ;
        RECT 64.650 165.065 64.980 165.435 ;
        RECT 65.630 165.095 65.980 165.345 ;
        RECT 64.245 164.885 64.415 165.030 ;
        RECT 66.165 164.925 66.335 165.555 ;
        RECT 66.965 165.685 67.295 166.165 ;
        RECT 67.465 165.875 67.690 166.335 ;
        RECT 67.860 165.685 68.190 166.165 ;
        RECT 66.965 165.515 68.190 165.685 ;
        RECT 68.380 165.535 68.630 166.335 ;
        RECT 68.800 165.535 69.140 166.165 ;
        RECT 66.505 165.145 66.835 165.345 ;
        RECT 67.005 165.145 67.335 165.345 ;
        RECT 67.505 165.145 67.925 165.345 ;
        RECT 68.100 165.175 68.795 165.345 ;
        RECT 68.100 164.925 68.270 165.175 ;
        RECT 68.965 164.925 69.140 165.535 ;
        RECT 69.585 165.525 69.830 166.130 ;
        RECT 70.050 165.800 70.560 166.335 ;
        RECT 63.790 163.955 64.060 164.860 ;
        RECT 64.245 164.715 64.910 164.885 ;
        RECT 64.230 163.785 64.560 164.545 ;
        RECT 64.740 163.955 64.910 164.715 ;
        RECT 65.835 164.755 68.270 164.925 ;
        RECT 65.835 163.955 66.165 164.755 ;
        RECT 66.335 163.785 66.665 164.585 ;
        RECT 66.965 163.955 67.295 164.755 ;
        RECT 67.940 163.785 68.190 164.585 ;
        RECT 68.460 163.785 68.630 164.925 ;
        RECT 68.800 163.955 69.140 164.925 ;
        RECT 69.310 165.355 70.540 165.525 ;
        RECT 69.310 164.545 69.650 165.355 ;
        RECT 69.820 164.790 70.570 164.980 ;
        RECT 69.310 164.135 69.825 164.545 ;
        RECT 70.060 163.785 70.230 164.545 ;
        RECT 70.400 164.125 70.570 164.790 ;
        RECT 70.740 164.805 70.930 166.165 ;
        RECT 71.100 165.655 71.375 166.165 ;
        RECT 71.565 165.800 72.095 166.165 ;
        RECT 72.520 165.935 72.850 166.335 ;
        RECT 71.920 165.765 72.095 165.800 ;
        RECT 71.100 165.485 71.380 165.655 ;
        RECT 71.100 165.005 71.375 165.485 ;
        RECT 71.580 164.805 71.750 165.605 ;
        RECT 70.740 164.635 71.750 164.805 ;
        RECT 71.920 165.595 72.850 165.765 ;
        RECT 73.020 165.595 73.275 166.165 ;
        RECT 73.450 165.610 73.740 166.335 ;
        RECT 73.910 165.825 74.215 166.335 ;
        RECT 71.920 164.465 72.090 165.595 ;
        RECT 72.680 165.425 72.850 165.595 ;
        RECT 70.965 164.295 72.090 164.465 ;
        RECT 72.260 165.095 72.455 165.425 ;
        RECT 72.680 165.095 72.935 165.425 ;
        RECT 72.260 164.125 72.430 165.095 ;
        RECT 73.105 164.925 73.275 165.595 ;
        RECT 73.910 165.095 74.225 165.655 ;
        RECT 74.395 165.345 74.645 166.155 ;
        RECT 74.815 165.810 75.075 166.335 ;
        RECT 75.255 165.345 75.505 166.155 ;
        RECT 75.675 165.775 75.935 166.335 ;
        RECT 76.105 165.685 76.365 166.140 ;
        RECT 76.535 165.855 76.795 166.335 ;
        RECT 76.965 165.685 77.225 166.140 ;
        RECT 77.395 165.855 77.655 166.335 ;
        RECT 77.825 165.685 78.085 166.140 ;
        RECT 78.255 165.855 78.500 166.335 ;
        RECT 78.670 165.685 78.945 166.140 ;
        RECT 79.115 165.855 79.360 166.335 ;
        RECT 79.530 165.685 79.790 166.140 ;
        RECT 79.970 165.855 80.220 166.335 ;
        RECT 80.390 165.685 80.650 166.140 ;
        RECT 80.830 165.855 81.080 166.335 ;
        RECT 81.250 165.685 81.510 166.140 ;
        RECT 81.690 165.855 81.950 166.335 ;
        RECT 82.120 165.685 82.380 166.140 ;
        RECT 82.550 165.855 82.850 166.335 ;
        RECT 76.105 165.515 82.850 165.685 ;
        RECT 74.395 165.095 81.515 165.345 ;
        RECT 70.400 163.955 72.430 164.125 ;
        RECT 72.600 163.785 72.770 164.925 ;
        RECT 72.940 163.955 73.275 164.925 ;
        RECT 73.450 163.785 73.740 164.950 ;
        RECT 73.920 163.785 74.215 164.595 ;
        RECT 74.395 163.955 74.640 165.095 ;
        RECT 74.815 163.785 75.075 164.595 ;
        RECT 75.255 163.960 75.505 165.095 ;
        RECT 81.685 164.975 82.850 165.515 ;
        RECT 83.945 165.625 84.200 166.155 ;
        RECT 84.380 165.875 84.665 166.335 ;
        RECT 81.685 164.925 82.880 164.975 ;
        RECT 76.105 164.805 82.880 164.925 ;
        RECT 76.105 164.700 82.850 164.805 ;
        RECT 83.945 164.765 84.125 165.625 ;
        RECT 84.845 165.425 85.095 166.075 ;
        RECT 84.295 165.095 85.095 165.425 ;
        RECT 76.105 164.685 81.510 164.700 ;
        RECT 75.675 163.790 75.935 164.585 ;
        RECT 76.105 163.960 76.365 164.685 ;
        RECT 76.535 163.790 76.795 164.515 ;
        RECT 76.965 163.960 77.225 164.685 ;
        RECT 77.395 163.790 77.655 164.515 ;
        RECT 77.825 163.960 78.085 164.685 ;
        RECT 78.255 163.790 78.515 164.515 ;
        RECT 78.685 163.960 78.945 164.685 ;
        RECT 79.115 163.790 79.360 164.515 ;
        RECT 79.530 163.960 79.790 164.685 ;
        RECT 79.975 163.790 80.220 164.515 ;
        RECT 80.390 163.960 80.650 164.685 ;
        RECT 80.835 163.790 81.080 164.515 ;
        RECT 81.250 163.960 81.510 164.685 ;
        RECT 81.695 163.790 81.950 164.515 ;
        RECT 82.120 163.960 82.410 164.700 ;
        RECT 75.675 163.785 81.950 163.790 ;
        RECT 82.580 163.785 82.850 164.530 ;
        RECT 83.945 164.295 84.200 164.765 ;
        RECT 83.860 164.125 84.200 164.295 ;
        RECT 83.945 164.095 84.200 164.125 ;
        RECT 84.380 163.785 84.665 164.585 ;
        RECT 84.845 164.505 85.095 165.095 ;
        RECT 85.295 165.740 85.615 166.070 ;
        RECT 85.795 165.855 86.455 166.335 ;
        RECT 86.655 165.945 87.505 166.115 ;
        RECT 85.295 164.845 85.485 165.740 ;
        RECT 85.805 165.415 86.465 165.685 ;
        RECT 86.135 165.355 86.465 165.415 ;
        RECT 85.655 165.185 85.985 165.245 ;
        RECT 86.655 165.185 86.825 165.945 ;
        RECT 88.065 165.875 88.385 166.335 ;
        RECT 88.585 165.695 88.835 166.125 ;
        RECT 89.125 165.895 89.535 166.335 ;
        RECT 89.705 165.955 90.720 166.155 ;
        RECT 86.995 165.525 88.245 165.695 ;
        RECT 86.995 165.405 87.325 165.525 ;
        RECT 85.655 165.015 87.555 165.185 ;
        RECT 85.295 164.675 87.215 164.845 ;
        RECT 85.295 164.655 85.615 164.675 ;
        RECT 84.845 163.995 85.175 164.505 ;
        RECT 85.445 164.045 85.615 164.655 ;
        RECT 87.385 164.505 87.555 165.015 ;
        RECT 87.725 164.945 87.905 165.355 ;
        RECT 88.075 164.765 88.245 165.525 ;
        RECT 85.785 163.785 86.115 164.475 ;
        RECT 86.345 164.335 87.555 164.505 ;
        RECT 87.725 164.455 88.245 164.765 ;
        RECT 88.415 165.355 88.835 165.695 ;
        RECT 89.125 165.355 89.535 165.685 ;
        RECT 88.415 164.585 88.605 165.355 ;
        RECT 89.705 165.225 89.875 165.955 ;
        RECT 91.020 165.785 91.190 166.115 ;
        RECT 91.360 165.955 91.690 166.335 ;
        RECT 90.045 165.405 90.395 165.775 ;
        RECT 89.705 165.185 90.125 165.225 ;
        RECT 88.775 165.015 90.125 165.185 ;
        RECT 88.775 164.855 89.025 165.015 ;
        RECT 89.535 164.585 89.785 164.845 ;
        RECT 88.415 164.335 89.785 164.585 ;
        RECT 86.345 164.045 86.585 164.335 ;
        RECT 87.385 164.255 87.555 164.335 ;
        RECT 86.785 163.785 87.205 164.165 ;
        RECT 87.385 164.005 88.015 164.255 ;
        RECT 88.485 163.785 88.815 164.165 ;
        RECT 88.985 164.045 89.155 164.335 ;
        RECT 89.955 164.170 90.125 165.015 ;
        RECT 90.575 164.845 90.795 165.715 ;
        RECT 91.020 165.595 91.715 165.785 ;
        RECT 90.295 164.465 90.795 164.845 ;
        RECT 90.965 164.795 91.375 165.415 ;
        RECT 91.545 164.625 91.715 165.595 ;
        RECT 91.020 164.455 91.715 164.625 ;
        RECT 89.335 163.785 89.715 164.165 ;
        RECT 89.955 164.000 90.785 164.170 ;
        RECT 91.020 163.955 91.190 164.455 ;
        RECT 91.360 163.785 91.690 164.285 ;
        RECT 91.905 163.955 92.130 166.075 ;
        RECT 92.300 165.955 92.630 166.335 ;
        RECT 92.800 165.785 92.970 166.075 ;
        RECT 92.305 165.615 92.970 165.785 ;
        RECT 92.305 164.625 92.535 165.615 ;
        RECT 93.230 165.585 94.440 166.335 ;
        RECT 92.705 164.795 93.055 165.445 ;
        RECT 93.230 164.875 93.750 165.415 ;
        RECT 93.920 165.045 94.440 165.585 ;
        RECT 94.610 165.535 94.950 166.165 ;
        RECT 95.120 165.535 95.370 166.335 ;
        RECT 95.560 165.685 95.890 166.165 ;
        RECT 96.060 165.875 96.285 166.335 ;
        RECT 96.455 165.685 96.785 166.165 ;
        RECT 94.610 164.925 94.785 165.535 ;
        RECT 95.560 165.515 96.785 165.685 ;
        RECT 97.415 165.555 97.915 166.165 ;
        RECT 99.210 165.610 99.500 166.335 ;
        RECT 100.135 165.625 100.390 166.155 ;
        RECT 100.560 165.875 100.865 166.335 ;
        RECT 101.110 165.955 102.180 166.125 ;
        RECT 94.955 165.175 95.650 165.345 ;
        RECT 95.480 164.925 95.650 165.175 ;
        RECT 95.825 165.145 96.245 165.345 ;
        RECT 96.415 165.145 96.745 165.345 ;
        RECT 96.915 165.145 97.245 165.345 ;
        RECT 97.415 164.925 97.585 165.555 ;
        RECT 97.770 165.095 98.120 165.345 ;
        RECT 100.135 164.975 100.345 165.625 ;
        RECT 101.110 165.600 101.430 165.955 ;
        RECT 101.105 165.425 101.430 165.600 ;
        RECT 100.515 165.125 101.430 165.425 ;
        RECT 101.600 165.385 101.840 165.785 ;
        RECT 102.010 165.725 102.180 165.955 ;
        RECT 102.350 165.895 102.540 166.335 ;
        RECT 102.710 165.885 103.660 166.165 ;
        RECT 103.880 165.975 104.230 166.145 ;
        RECT 102.010 165.555 102.540 165.725 ;
        RECT 100.515 165.095 101.255 165.125 ;
        RECT 92.305 164.455 92.970 164.625 ;
        RECT 92.300 163.785 92.630 164.285 ;
        RECT 92.800 163.955 92.970 164.455 ;
        RECT 93.230 163.785 94.440 164.875 ;
        RECT 94.610 163.955 94.950 164.925 ;
        RECT 95.120 163.785 95.290 164.925 ;
        RECT 95.480 164.755 97.915 164.925 ;
        RECT 95.560 163.785 95.810 164.585 ;
        RECT 96.455 163.955 96.785 164.755 ;
        RECT 97.085 163.785 97.415 164.585 ;
        RECT 97.585 163.955 97.915 164.755 ;
        RECT 99.210 163.785 99.500 164.950 ;
        RECT 100.135 164.095 100.390 164.975 ;
        RECT 100.560 163.785 100.865 164.925 ;
        RECT 101.085 164.505 101.255 165.095 ;
        RECT 101.600 165.015 102.140 165.385 ;
        RECT 102.320 165.275 102.540 165.555 ;
        RECT 102.710 165.105 102.880 165.885 ;
        RECT 102.475 164.935 102.880 165.105 ;
        RECT 103.050 165.095 103.400 165.715 ;
        RECT 102.475 164.845 102.645 164.935 ;
        RECT 103.570 164.925 103.780 165.715 ;
        RECT 101.425 164.675 102.645 164.845 ;
        RECT 103.105 164.765 103.780 164.925 ;
        RECT 101.085 164.335 101.885 164.505 ;
        RECT 101.205 163.785 101.535 164.165 ;
        RECT 101.715 164.045 101.885 164.335 ;
        RECT 102.475 164.295 102.645 164.675 ;
        RECT 102.815 164.755 103.780 164.765 ;
        RECT 103.970 165.585 104.230 165.975 ;
        RECT 104.440 165.875 104.770 166.335 ;
        RECT 105.645 165.945 106.500 166.115 ;
        RECT 106.705 165.945 107.200 166.115 ;
        RECT 107.370 165.975 107.700 166.335 ;
        RECT 103.970 164.895 104.140 165.585 ;
        RECT 104.310 165.235 104.480 165.415 ;
        RECT 104.650 165.405 105.440 165.655 ;
        RECT 105.645 165.235 105.815 165.945 ;
        RECT 105.985 165.435 106.340 165.655 ;
        RECT 104.310 165.065 106.000 165.235 ;
        RECT 102.815 164.465 103.275 164.755 ;
        RECT 103.970 164.725 105.470 164.895 ;
        RECT 103.970 164.585 104.140 164.725 ;
        RECT 103.580 164.415 104.140 164.585 ;
        RECT 102.055 163.785 102.305 164.245 ;
        RECT 102.475 163.955 103.345 164.295 ;
        RECT 103.580 163.955 103.750 164.415 ;
        RECT 104.585 164.385 105.660 164.555 ;
        RECT 103.920 163.785 104.290 164.245 ;
        RECT 104.585 164.045 104.755 164.385 ;
        RECT 104.925 163.785 105.255 164.215 ;
        RECT 105.490 164.045 105.660 164.385 ;
        RECT 105.830 164.285 106.000 165.065 ;
        RECT 106.170 164.845 106.340 165.435 ;
        RECT 106.510 165.035 106.860 165.655 ;
        RECT 106.170 164.455 106.635 164.845 ;
        RECT 107.030 164.585 107.200 165.945 ;
        RECT 107.370 164.755 107.830 165.805 ;
        RECT 106.805 164.415 107.200 164.585 ;
        RECT 106.805 164.285 106.975 164.415 ;
        RECT 105.830 163.955 106.510 164.285 ;
        RECT 106.725 163.955 106.975 164.285 ;
        RECT 107.145 163.785 107.395 164.245 ;
        RECT 107.565 163.970 107.890 164.755 ;
        RECT 108.060 163.955 108.230 166.075 ;
        RECT 108.400 165.955 108.730 166.335 ;
        RECT 108.900 165.785 109.155 166.075 ;
        RECT 108.405 165.615 109.155 165.785 ;
        RECT 108.405 164.625 108.635 165.615 ;
        RECT 109.330 165.565 111.000 166.335 ;
        RECT 111.170 165.585 112.380 166.335 ;
        RECT 108.805 164.795 109.155 165.445 ;
        RECT 109.330 164.875 110.080 165.395 ;
        RECT 110.250 165.045 111.000 165.565 ;
        RECT 111.170 164.875 111.690 165.415 ;
        RECT 111.860 165.045 112.380 165.585 ;
        RECT 108.405 164.455 109.155 164.625 ;
        RECT 108.400 163.785 108.730 164.285 ;
        RECT 108.900 163.955 109.155 164.455 ;
        RECT 109.330 163.785 111.000 164.875 ;
        RECT 111.170 163.785 112.380 164.875 ;
        RECT 18.165 163.615 112.465 163.785 ;
        RECT 18.250 162.525 19.460 163.615 ;
        RECT 18.250 161.815 18.770 162.355 ;
        RECT 18.940 161.985 19.460 162.525 ;
        RECT 19.690 162.475 19.900 163.615 ;
        RECT 20.070 162.465 20.400 163.445 ;
        RECT 20.570 162.475 20.800 163.615 ;
        RECT 21.100 162.685 21.270 163.445 ;
        RECT 21.450 162.855 21.780 163.615 ;
        RECT 21.100 162.515 21.765 162.685 ;
        RECT 21.950 162.540 22.220 163.445 ;
        RECT 18.250 161.065 19.460 161.815 ;
        RECT 19.690 161.065 19.900 161.885 ;
        RECT 20.070 161.865 20.320 162.465 ;
        RECT 21.595 162.370 21.765 162.515 ;
        RECT 20.490 162.055 20.820 162.305 ;
        RECT 21.030 161.965 21.360 162.335 ;
        RECT 21.595 162.040 21.880 162.370 ;
        RECT 20.070 161.235 20.400 161.865 ;
        RECT 20.570 161.065 20.800 161.885 ;
        RECT 21.595 161.785 21.765 162.040 ;
        RECT 21.100 161.615 21.765 161.785 ;
        RECT 22.050 161.740 22.220 162.540 ;
        RECT 21.100 161.235 21.270 161.615 ;
        RECT 21.450 161.065 21.780 161.445 ;
        RECT 21.960 161.235 22.220 161.740 ;
        RECT 22.395 162.425 22.650 163.305 ;
        RECT 22.820 162.475 23.125 163.615 ;
        RECT 23.465 163.235 23.795 163.615 ;
        RECT 23.975 163.065 24.145 163.355 ;
        RECT 24.315 163.155 24.565 163.615 ;
        RECT 23.345 162.895 24.145 163.065 ;
        RECT 24.735 163.105 25.605 163.445 ;
        RECT 22.395 161.775 22.605 162.425 ;
        RECT 23.345 162.305 23.515 162.895 ;
        RECT 24.735 162.725 24.905 163.105 ;
        RECT 25.840 162.985 26.010 163.445 ;
        RECT 26.180 163.155 26.550 163.615 ;
        RECT 26.845 163.015 27.015 163.355 ;
        RECT 27.185 163.185 27.515 163.615 ;
        RECT 27.750 163.015 27.920 163.355 ;
        RECT 23.685 162.555 24.905 162.725 ;
        RECT 25.075 162.645 25.535 162.935 ;
        RECT 25.840 162.815 26.400 162.985 ;
        RECT 26.845 162.845 27.920 163.015 ;
        RECT 28.090 163.115 28.770 163.445 ;
        RECT 28.985 163.115 29.235 163.445 ;
        RECT 29.405 163.155 29.655 163.615 ;
        RECT 26.230 162.675 26.400 162.815 ;
        RECT 25.075 162.635 26.040 162.645 ;
        RECT 24.735 162.465 24.905 162.555 ;
        RECT 25.365 162.475 26.040 162.635 ;
        RECT 22.775 162.275 23.515 162.305 ;
        RECT 22.775 161.975 23.690 162.275 ;
        RECT 23.365 161.800 23.690 161.975 ;
        RECT 22.395 161.245 22.650 161.775 ;
        RECT 22.820 161.065 23.125 161.525 ;
        RECT 23.370 161.445 23.690 161.800 ;
        RECT 23.860 162.015 24.400 162.385 ;
        RECT 24.735 162.295 25.140 162.465 ;
        RECT 23.860 161.615 24.100 162.015 ;
        RECT 24.580 161.845 24.800 162.125 ;
        RECT 24.270 161.675 24.800 161.845 ;
        RECT 24.270 161.445 24.440 161.675 ;
        RECT 24.970 161.515 25.140 162.295 ;
        RECT 25.310 161.685 25.660 162.305 ;
        RECT 25.830 161.685 26.040 162.475 ;
        RECT 26.230 162.505 27.730 162.675 ;
        RECT 26.230 161.815 26.400 162.505 ;
        RECT 28.090 162.335 28.260 163.115 ;
        RECT 29.065 162.985 29.235 163.115 ;
        RECT 26.570 162.165 28.260 162.335 ;
        RECT 28.430 162.555 28.895 162.945 ;
        RECT 29.065 162.815 29.460 162.985 ;
        RECT 26.570 161.985 26.740 162.165 ;
        RECT 23.370 161.275 24.440 161.445 ;
        RECT 24.610 161.065 24.800 161.505 ;
        RECT 24.970 161.235 25.920 161.515 ;
        RECT 26.230 161.425 26.490 161.815 ;
        RECT 26.910 161.745 27.700 161.995 ;
        RECT 26.140 161.255 26.490 161.425 ;
        RECT 26.700 161.065 27.030 161.525 ;
        RECT 27.905 161.455 28.075 162.165 ;
        RECT 28.430 161.965 28.600 162.555 ;
        RECT 28.245 161.745 28.600 161.965 ;
        RECT 28.770 161.745 29.120 162.365 ;
        RECT 29.290 161.455 29.460 162.815 ;
        RECT 29.825 162.645 30.150 163.430 ;
        RECT 29.630 161.595 30.090 162.645 ;
        RECT 27.905 161.285 28.760 161.455 ;
        RECT 28.965 161.285 29.460 161.455 ;
        RECT 29.630 161.065 29.960 161.425 ;
        RECT 30.320 161.325 30.490 163.445 ;
        RECT 30.660 163.115 30.990 163.615 ;
        RECT 31.160 162.945 31.415 163.445 ;
        RECT 30.665 162.775 31.415 162.945 ;
        RECT 30.665 161.785 30.895 162.775 ;
        RECT 31.065 161.955 31.415 162.605 ;
        RECT 32.050 162.525 34.640 163.615 ;
        RECT 32.050 162.005 33.260 162.525 ;
        RECT 34.810 162.450 35.100 163.615 ;
        RECT 35.270 162.525 36.940 163.615 ;
        RECT 37.200 162.870 37.470 163.615 ;
        RECT 38.100 163.610 44.375 163.615 ;
        RECT 37.640 162.700 37.930 163.440 ;
        RECT 38.100 162.885 38.355 163.610 ;
        RECT 38.540 162.715 38.800 163.440 ;
        RECT 38.970 162.885 39.215 163.610 ;
        RECT 39.400 162.715 39.660 163.440 ;
        RECT 39.830 162.885 40.075 163.610 ;
        RECT 40.260 162.715 40.520 163.440 ;
        RECT 40.690 162.885 40.935 163.610 ;
        RECT 41.105 162.715 41.365 163.440 ;
        RECT 41.535 162.885 41.795 163.610 ;
        RECT 41.965 162.715 42.225 163.440 ;
        RECT 42.395 162.885 42.655 163.610 ;
        RECT 42.825 162.715 43.085 163.440 ;
        RECT 43.255 162.885 43.515 163.610 ;
        RECT 43.685 162.715 43.945 163.440 ;
        RECT 44.115 162.815 44.375 163.610 ;
        RECT 38.540 162.700 43.945 162.715 ;
        RECT 33.430 161.835 34.640 162.355 ;
        RECT 35.270 162.005 36.020 162.525 ;
        RECT 37.200 162.475 43.945 162.700 ;
        RECT 36.190 161.835 36.940 162.355 ;
        RECT 30.665 161.615 31.415 161.785 ;
        RECT 30.660 161.065 30.990 161.445 ;
        RECT 31.160 161.325 31.415 161.615 ;
        RECT 32.050 161.065 34.640 161.835 ;
        RECT 34.810 161.065 35.100 161.790 ;
        RECT 35.270 161.065 36.940 161.835 ;
        RECT 37.200 161.885 38.365 162.475 ;
        RECT 44.545 162.305 44.795 163.440 ;
        RECT 44.975 162.805 45.235 163.615 ;
        RECT 45.410 162.305 45.655 163.445 ;
        RECT 45.835 162.805 46.130 163.615 ;
        RECT 46.410 163.155 46.580 163.615 ;
        RECT 46.750 162.665 47.080 163.445 ;
        RECT 47.250 162.815 47.420 163.615 ;
        RECT 46.310 162.645 47.080 162.665 ;
        RECT 47.590 162.645 47.920 163.445 ;
        RECT 48.090 162.815 48.260 163.615 ;
        RECT 48.430 162.645 48.760 163.445 ;
        RECT 46.310 162.475 48.760 162.645 ;
        RECT 49.020 162.475 49.315 163.615 ;
        RECT 38.535 162.055 45.655 162.305 ;
        RECT 37.200 161.715 43.945 161.885 ;
        RECT 37.200 161.065 37.500 161.545 ;
        RECT 37.670 161.260 37.930 161.715 ;
        RECT 38.100 161.065 38.360 161.545 ;
        RECT 38.540 161.260 38.800 161.715 ;
        RECT 38.970 161.065 39.220 161.545 ;
        RECT 39.400 161.260 39.660 161.715 ;
        RECT 39.830 161.065 40.080 161.545 ;
        RECT 40.260 161.260 40.520 161.715 ;
        RECT 40.690 161.065 40.935 161.545 ;
        RECT 41.105 161.260 41.380 161.715 ;
        RECT 41.550 161.065 41.795 161.545 ;
        RECT 41.965 161.260 42.225 161.715 ;
        RECT 42.395 161.065 42.655 161.545 ;
        RECT 42.825 161.260 43.085 161.715 ;
        RECT 43.255 161.065 43.515 161.545 ;
        RECT 43.685 161.260 43.945 161.715 ;
        RECT 44.115 161.065 44.375 161.625 ;
        RECT 44.545 161.245 44.795 162.055 ;
        RECT 44.975 161.065 45.235 161.590 ;
        RECT 45.405 161.245 45.655 162.055 ;
        RECT 45.825 161.745 46.140 162.305 ;
        RECT 46.310 161.885 46.660 162.475 ;
        RECT 49.535 162.425 49.790 163.305 ;
        RECT 49.960 162.475 50.265 163.615 ;
        RECT 50.605 163.235 50.935 163.615 ;
        RECT 51.115 163.065 51.285 163.355 ;
        RECT 51.455 163.155 51.705 163.615 ;
        RECT 50.485 162.895 51.285 163.065 ;
        RECT 51.875 163.105 52.745 163.445 ;
        RECT 46.830 162.055 49.340 162.305 ;
        RECT 46.310 161.705 48.680 161.885 ;
        RECT 45.835 161.065 46.140 161.575 ;
        RECT 46.410 161.065 46.660 161.530 ;
        RECT 46.830 161.235 47.000 161.705 ;
        RECT 47.250 161.065 47.420 161.525 ;
        RECT 47.670 161.235 47.840 161.705 ;
        RECT 48.090 161.065 48.260 161.525 ;
        RECT 48.510 161.235 48.680 161.705 ;
        RECT 49.535 161.775 49.745 162.425 ;
        RECT 50.485 162.305 50.655 162.895 ;
        RECT 51.875 162.725 52.045 163.105 ;
        RECT 52.980 162.985 53.150 163.445 ;
        RECT 53.320 163.155 53.690 163.615 ;
        RECT 53.985 163.015 54.155 163.355 ;
        RECT 54.325 163.185 54.655 163.615 ;
        RECT 54.890 163.015 55.060 163.355 ;
        RECT 50.825 162.555 52.045 162.725 ;
        RECT 52.215 162.645 52.675 162.935 ;
        RECT 52.980 162.815 53.540 162.985 ;
        RECT 53.985 162.845 55.060 163.015 ;
        RECT 55.230 163.115 55.910 163.445 ;
        RECT 56.125 163.115 56.375 163.445 ;
        RECT 56.545 163.155 56.795 163.615 ;
        RECT 53.370 162.675 53.540 162.815 ;
        RECT 52.215 162.635 53.180 162.645 ;
        RECT 51.875 162.465 52.045 162.555 ;
        RECT 52.505 162.475 53.180 162.635 ;
        RECT 49.915 162.275 50.655 162.305 ;
        RECT 49.915 161.975 50.830 162.275 ;
        RECT 50.505 161.800 50.830 161.975 ;
        RECT 49.050 161.065 49.315 161.525 ;
        RECT 49.535 161.245 49.790 161.775 ;
        RECT 49.960 161.065 50.265 161.525 ;
        RECT 50.510 161.445 50.830 161.800 ;
        RECT 51.000 162.015 51.540 162.385 ;
        RECT 51.875 162.295 52.280 162.465 ;
        RECT 51.000 161.615 51.240 162.015 ;
        RECT 51.720 161.845 51.940 162.125 ;
        RECT 51.410 161.675 51.940 161.845 ;
        RECT 51.410 161.445 51.580 161.675 ;
        RECT 52.110 161.515 52.280 162.295 ;
        RECT 52.450 161.685 52.800 162.305 ;
        RECT 52.970 161.685 53.180 162.475 ;
        RECT 53.370 162.505 54.870 162.675 ;
        RECT 53.370 161.815 53.540 162.505 ;
        RECT 55.230 162.335 55.400 163.115 ;
        RECT 56.205 162.985 56.375 163.115 ;
        RECT 53.710 162.165 55.400 162.335 ;
        RECT 55.570 162.555 56.035 162.945 ;
        RECT 56.205 162.815 56.600 162.985 ;
        RECT 53.710 161.985 53.880 162.165 ;
        RECT 50.510 161.275 51.580 161.445 ;
        RECT 51.750 161.065 51.940 161.505 ;
        RECT 52.110 161.235 53.060 161.515 ;
        RECT 53.370 161.425 53.630 161.815 ;
        RECT 54.050 161.745 54.840 161.995 ;
        RECT 53.280 161.255 53.630 161.425 ;
        RECT 53.840 161.065 54.170 161.525 ;
        RECT 55.045 161.455 55.215 162.165 ;
        RECT 55.570 161.965 55.740 162.555 ;
        RECT 55.385 161.745 55.740 161.965 ;
        RECT 55.910 161.745 56.260 162.365 ;
        RECT 56.430 161.455 56.600 162.815 ;
        RECT 56.965 162.645 57.290 163.430 ;
        RECT 56.770 161.595 57.230 162.645 ;
        RECT 55.045 161.285 55.900 161.455 ;
        RECT 56.105 161.285 56.600 161.455 ;
        RECT 56.770 161.065 57.100 161.425 ;
        RECT 57.460 161.325 57.630 163.445 ;
        RECT 57.800 163.115 58.130 163.615 ;
        RECT 58.300 162.945 58.555 163.445 ;
        RECT 57.805 162.775 58.555 162.945 ;
        RECT 57.805 161.785 58.035 162.775 ;
        RECT 58.205 161.955 58.555 162.605 ;
        RECT 58.730 162.525 60.400 163.615 ;
        RECT 58.730 162.005 59.480 162.525 ;
        RECT 60.570 162.450 60.860 163.615 ;
        RECT 61.490 162.525 63.160 163.615 ;
        RECT 59.650 161.835 60.400 162.355 ;
        RECT 61.490 162.005 62.240 162.525 ;
        RECT 63.335 162.465 63.595 163.615 ;
        RECT 63.770 162.540 64.025 163.445 ;
        RECT 64.195 162.855 64.525 163.615 ;
        RECT 64.740 162.685 64.910 163.445 ;
        RECT 62.410 161.835 63.160 162.355 ;
        RECT 57.805 161.615 58.555 161.785 ;
        RECT 57.800 161.065 58.130 161.445 ;
        RECT 58.300 161.325 58.555 161.615 ;
        RECT 58.730 161.065 60.400 161.835 ;
        RECT 60.570 161.065 60.860 161.790 ;
        RECT 61.490 161.065 63.160 161.835 ;
        RECT 63.335 161.065 63.595 161.905 ;
        RECT 63.770 161.810 63.940 162.540 ;
        RECT 64.195 162.515 64.910 162.685 ;
        RECT 65.170 162.525 67.760 163.615 ;
        RECT 67.930 162.540 68.200 163.445 ;
        RECT 68.370 162.855 68.700 163.615 ;
        RECT 68.880 162.685 69.050 163.445 ;
        RECT 64.195 162.305 64.365 162.515 ;
        RECT 64.110 161.975 64.365 162.305 ;
        RECT 63.770 161.235 64.025 161.810 ;
        RECT 64.195 161.785 64.365 161.975 ;
        RECT 64.645 161.965 65.000 162.335 ;
        RECT 65.170 162.005 66.380 162.525 ;
        RECT 66.550 161.835 67.760 162.355 ;
        RECT 64.195 161.615 64.910 161.785 ;
        RECT 64.195 161.065 64.525 161.445 ;
        RECT 64.740 161.235 64.910 161.615 ;
        RECT 65.170 161.065 67.760 161.835 ;
        RECT 67.930 161.740 68.100 162.540 ;
        RECT 68.385 162.515 69.050 162.685 ;
        RECT 69.310 162.525 70.520 163.615 ;
        RECT 68.385 162.370 68.555 162.515 ;
        RECT 68.270 162.040 68.555 162.370 ;
        RECT 68.385 161.785 68.555 162.040 ;
        RECT 68.790 161.965 69.120 162.335 ;
        RECT 69.310 161.985 69.830 162.525 ;
        RECT 70.690 162.475 71.030 163.445 ;
        RECT 71.200 162.475 71.370 163.615 ;
        RECT 71.640 162.815 71.890 163.615 ;
        RECT 72.535 162.645 72.865 163.445 ;
        RECT 73.165 162.815 73.495 163.615 ;
        RECT 73.665 162.645 73.995 163.445 ;
        RECT 71.560 162.475 73.995 162.645 ;
        RECT 74.375 162.475 74.710 163.445 ;
        RECT 74.880 162.475 75.050 163.615 ;
        RECT 75.220 163.275 77.250 163.445 ;
        RECT 70.690 162.425 70.920 162.475 ;
        RECT 70.000 161.815 70.520 162.355 ;
        RECT 67.930 161.235 68.190 161.740 ;
        RECT 68.385 161.615 69.050 161.785 ;
        RECT 68.370 161.065 68.700 161.445 ;
        RECT 68.880 161.235 69.050 161.615 ;
        RECT 69.310 161.065 70.520 161.815 ;
        RECT 70.690 161.865 70.865 162.425 ;
        RECT 71.560 162.225 71.730 162.475 ;
        RECT 71.035 162.055 71.730 162.225 ;
        RECT 71.905 162.055 72.325 162.255 ;
        RECT 72.495 162.055 72.825 162.255 ;
        RECT 72.995 162.055 73.325 162.255 ;
        RECT 70.690 161.235 71.030 161.865 ;
        RECT 71.200 161.065 71.450 161.865 ;
        RECT 71.640 161.715 72.865 161.885 ;
        RECT 71.640 161.235 71.970 161.715 ;
        RECT 72.140 161.065 72.365 161.525 ;
        RECT 72.535 161.235 72.865 161.715 ;
        RECT 73.495 161.845 73.665 162.475 ;
        RECT 73.850 162.055 74.200 162.305 ;
        RECT 73.495 161.235 73.995 161.845 ;
        RECT 74.375 161.805 74.545 162.475 ;
        RECT 75.220 162.305 75.390 163.275 ;
        RECT 74.715 161.975 74.970 162.305 ;
        RECT 75.195 161.975 75.390 162.305 ;
        RECT 75.560 162.935 76.685 163.105 ;
        RECT 74.800 161.805 74.970 161.975 ;
        RECT 75.560 161.805 75.730 162.935 ;
        RECT 74.375 161.235 74.630 161.805 ;
        RECT 74.800 161.635 75.730 161.805 ;
        RECT 75.900 162.595 76.910 162.765 ;
        RECT 75.900 161.795 76.070 162.595 ;
        RECT 76.275 161.915 76.550 162.395 ;
        RECT 76.270 161.745 76.550 161.915 ;
        RECT 75.555 161.600 75.730 161.635 ;
        RECT 74.800 161.065 75.130 161.465 ;
        RECT 75.555 161.235 76.085 161.600 ;
        RECT 76.275 161.235 76.550 161.745 ;
        RECT 76.720 161.235 76.910 162.595 ;
        RECT 77.080 162.610 77.250 163.275 ;
        RECT 77.420 162.855 77.590 163.615 ;
        RECT 77.825 162.855 78.340 163.265 ;
        RECT 77.080 162.420 77.830 162.610 ;
        RECT 78.000 162.045 78.340 162.855 ;
        RECT 77.110 161.875 78.340 162.045 ;
        RECT 78.510 162.855 79.025 163.265 ;
        RECT 79.260 162.855 79.430 163.615 ;
        RECT 79.600 163.275 81.630 163.445 ;
        RECT 78.510 162.045 78.850 162.855 ;
        RECT 79.600 162.610 79.770 163.275 ;
        RECT 80.165 162.935 81.290 163.105 ;
        RECT 79.020 162.420 79.770 162.610 ;
        RECT 79.940 162.595 80.950 162.765 ;
        RECT 78.510 161.875 79.740 162.045 ;
        RECT 77.090 161.065 77.600 161.600 ;
        RECT 77.820 161.270 78.065 161.875 ;
        RECT 78.785 161.270 79.030 161.875 ;
        RECT 79.250 161.065 79.760 161.600 ;
        RECT 79.940 161.235 80.130 162.595 ;
        RECT 80.300 161.575 80.575 162.395 ;
        RECT 80.780 161.795 80.950 162.595 ;
        RECT 81.120 161.805 81.290 162.935 ;
        RECT 81.460 162.305 81.630 163.275 ;
        RECT 81.800 162.475 81.970 163.615 ;
        RECT 82.140 162.475 82.475 163.445 ;
        RECT 83.610 162.475 83.840 163.615 ;
        RECT 81.460 161.975 81.655 162.305 ;
        RECT 81.880 161.975 82.135 162.305 ;
        RECT 81.880 161.805 82.050 161.975 ;
        RECT 82.305 161.805 82.475 162.475 ;
        RECT 84.010 162.465 84.340 163.445 ;
        RECT 84.510 162.475 84.720 163.615 ;
        RECT 84.950 162.540 85.220 163.445 ;
        RECT 85.390 162.855 85.720 163.615 ;
        RECT 85.900 162.685 86.070 163.445 ;
        RECT 83.590 162.055 83.920 162.305 ;
        RECT 81.120 161.635 82.050 161.805 ;
        RECT 81.120 161.600 81.295 161.635 ;
        RECT 80.300 161.405 80.580 161.575 ;
        RECT 80.300 161.235 80.575 161.405 ;
        RECT 80.765 161.235 81.295 161.600 ;
        RECT 81.720 161.065 82.050 161.465 ;
        RECT 82.220 161.235 82.475 161.805 ;
        RECT 83.610 161.065 83.840 161.885 ;
        RECT 84.090 161.865 84.340 162.465 ;
        RECT 84.010 161.235 84.340 161.865 ;
        RECT 84.510 161.065 84.720 161.885 ;
        RECT 84.950 161.740 85.120 162.540 ;
        RECT 85.405 162.515 86.070 162.685 ;
        RECT 85.405 162.370 85.575 162.515 ;
        RECT 86.330 162.450 86.620 163.615 ;
        RECT 87.710 162.855 88.225 163.265 ;
        RECT 88.460 162.855 88.630 163.615 ;
        RECT 88.800 163.275 90.830 163.445 ;
        RECT 85.290 162.040 85.575 162.370 ;
        RECT 85.405 161.785 85.575 162.040 ;
        RECT 85.810 161.965 86.140 162.335 ;
        RECT 87.710 162.045 88.050 162.855 ;
        RECT 88.800 162.610 88.970 163.275 ;
        RECT 89.365 162.935 90.490 163.105 ;
        RECT 88.220 162.420 88.970 162.610 ;
        RECT 89.140 162.595 90.150 162.765 ;
        RECT 87.710 161.875 88.940 162.045 ;
        RECT 84.950 161.235 85.210 161.740 ;
        RECT 85.405 161.615 86.070 161.785 ;
        RECT 85.390 161.065 85.720 161.445 ;
        RECT 85.900 161.235 86.070 161.615 ;
        RECT 86.330 161.065 86.620 161.790 ;
        RECT 87.985 161.270 88.230 161.875 ;
        RECT 88.450 161.065 88.960 161.600 ;
        RECT 89.140 161.235 89.330 162.595 ;
        RECT 89.500 161.575 89.775 162.395 ;
        RECT 89.980 161.795 90.150 162.595 ;
        RECT 90.320 161.805 90.490 162.935 ;
        RECT 90.660 162.305 90.830 163.275 ;
        RECT 91.000 162.475 91.170 163.615 ;
        RECT 91.340 162.475 91.675 163.445 ;
        RECT 90.660 161.975 90.855 162.305 ;
        RECT 91.080 161.975 91.335 162.305 ;
        RECT 91.080 161.805 91.250 161.975 ;
        RECT 91.505 161.805 91.675 162.475 ;
        RECT 90.320 161.635 91.250 161.805 ;
        RECT 90.320 161.600 90.495 161.635 ;
        RECT 89.500 161.405 89.780 161.575 ;
        RECT 89.500 161.235 89.775 161.405 ;
        RECT 89.965 161.235 90.495 161.600 ;
        RECT 90.920 161.065 91.250 161.465 ;
        RECT 91.420 161.235 91.675 161.805 ;
        RECT 91.850 162.540 92.120 163.445 ;
        RECT 92.290 162.855 92.620 163.615 ;
        RECT 92.800 162.685 92.970 163.445 ;
        RECT 91.850 161.740 92.020 162.540 ;
        RECT 92.305 162.515 92.970 162.685 ;
        RECT 93.230 162.525 94.440 163.615 ;
        RECT 92.305 162.370 92.475 162.515 ;
        RECT 92.190 162.040 92.475 162.370 ;
        RECT 92.305 161.785 92.475 162.040 ;
        RECT 92.710 161.965 93.040 162.335 ;
        RECT 93.230 161.985 93.750 162.525 ;
        RECT 94.610 162.475 94.950 163.445 ;
        RECT 95.120 162.475 95.290 163.615 ;
        RECT 95.560 162.815 95.810 163.615 ;
        RECT 96.455 162.645 96.785 163.445 ;
        RECT 97.085 162.815 97.415 163.615 ;
        RECT 97.585 162.645 97.915 163.445 ;
        RECT 95.480 162.475 97.915 162.645 ;
        RECT 98.750 162.525 100.420 163.615 ;
        RECT 100.590 162.855 101.105 163.265 ;
        RECT 101.340 162.855 101.510 163.615 ;
        RECT 101.680 163.275 103.710 163.445 ;
        RECT 94.610 162.425 94.840 162.475 ;
        RECT 93.920 161.815 94.440 162.355 ;
        RECT 91.850 161.235 92.110 161.740 ;
        RECT 92.305 161.615 92.970 161.785 ;
        RECT 92.290 161.065 92.620 161.445 ;
        RECT 92.800 161.235 92.970 161.615 ;
        RECT 93.230 161.065 94.440 161.815 ;
        RECT 94.610 161.865 94.785 162.425 ;
        RECT 95.480 162.225 95.650 162.475 ;
        RECT 94.955 162.055 95.650 162.225 ;
        RECT 95.825 162.055 96.245 162.255 ;
        RECT 96.415 162.055 96.745 162.255 ;
        RECT 96.915 162.055 97.245 162.255 ;
        RECT 94.610 161.235 94.950 161.865 ;
        RECT 95.120 161.065 95.370 161.865 ;
        RECT 95.560 161.715 96.785 161.885 ;
        RECT 95.560 161.235 95.890 161.715 ;
        RECT 96.060 161.065 96.285 161.525 ;
        RECT 96.455 161.235 96.785 161.715 ;
        RECT 97.415 161.845 97.585 162.475 ;
        RECT 97.770 162.055 98.120 162.305 ;
        RECT 98.750 162.005 99.500 162.525 ;
        RECT 97.415 161.235 97.915 161.845 ;
        RECT 99.670 161.835 100.420 162.355 ;
        RECT 100.590 162.045 100.930 162.855 ;
        RECT 101.680 162.610 101.850 163.275 ;
        RECT 102.245 162.935 103.370 163.105 ;
        RECT 101.100 162.420 101.850 162.610 ;
        RECT 102.020 162.595 103.030 162.765 ;
        RECT 100.590 161.875 101.820 162.045 ;
        RECT 98.750 161.065 100.420 161.835 ;
        RECT 100.865 161.270 101.110 161.875 ;
        RECT 101.330 161.065 101.840 161.600 ;
        RECT 102.020 161.235 102.210 162.595 ;
        RECT 102.380 162.255 102.655 162.395 ;
        RECT 102.380 162.085 102.660 162.255 ;
        RECT 102.380 161.235 102.655 162.085 ;
        RECT 102.860 161.795 103.030 162.595 ;
        RECT 103.200 161.805 103.370 162.935 ;
        RECT 103.540 162.305 103.710 163.275 ;
        RECT 103.880 162.475 104.050 163.615 ;
        RECT 104.220 162.475 104.555 163.445 ;
        RECT 104.770 162.475 105.000 163.615 ;
        RECT 103.540 161.975 103.735 162.305 ;
        RECT 103.960 161.975 104.215 162.305 ;
        RECT 103.960 161.805 104.130 161.975 ;
        RECT 104.385 161.805 104.555 162.475 ;
        RECT 105.170 162.465 105.500 163.445 ;
        RECT 105.670 162.475 105.880 163.615 ;
        RECT 107.035 163.190 107.370 163.615 ;
        RECT 107.540 163.010 107.725 163.415 ;
        RECT 107.060 162.835 107.725 163.010 ;
        RECT 107.930 162.835 108.260 163.615 ;
        RECT 104.750 162.055 105.080 162.305 ;
        RECT 103.200 161.635 104.130 161.805 ;
        RECT 103.200 161.600 103.375 161.635 ;
        RECT 102.845 161.235 103.375 161.600 ;
        RECT 103.800 161.065 104.130 161.465 ;
        RECT 104.300 161.235 104.555 161.805 ;
        RECT 104.770 161.065 105.000 161.885 ;
        RECT 105.250 161.865 105.500 162.465 ;
        RECT 105.170 161.235 105.500 161.865 ;
        RECT 105.670 161.065 105.880 161.885 ;
        RECT 107.060 161.805 107.400 162.835 ;
        RECT 108.430 162.645 108.700 163.415 ;
        RECT 107.570 162.475 108.700 162.645 ;
        RECT 108.960 162.685 109.130 163.445 ;
        RECT 109.310 162.855 109.640 163.615 ;
        RECT 108.960 162.515 109.625 162.685 ;
        RECT 109.810 162.540 110.080 163.445 ;
        RECT 107.570 161.975 107.820 162.475 ;
        RECT 107.060 161.635 107.745 161.805 ;
        RECT 108.000 161.725 108.360 162.305 ;
        RECT 107.035 161.065 107.370 161.465 ;
        RECT 107.540 161.235 107.745 161.635 ;
        RECT 108.530 161.565 108.700 162.475 ;
        RECT 109.455 162.370 109.625 162.515 ;
        RECT 108.890 161.965 109.220 162.335 ;
        RECT 109.455 162.040 109.740 162.370 ;
        RECT 109.455 161.785 109.625 162.040 ;
        RECT 107.955 161.065 108.230 161.545 ;
        RECT 108.440 161.235 108.700 161.565 ;
        RECT 108.960 161.615 109.625 161.785 ;
        RECT 109.910 161.740 110.080 162.540 ;
        RECT 111.170 162.525 112.380 163.615 ;
        RECT 111.170 161.985 111.690 162.525 ;
        RECT 111.860 161.815 112.380 162.355 ;
        RECT 108.960 161.235 109.130 161.615 ;
        RECT 109.310 161.065 109.640 161.445 ;
        RECT 109.820 161.235 110.080 161.740 ;
        RECT 111.170 161.065 112.380 161.815 ;
        RECT 18.165 160.895 112.465 161.065 ;
        RECT 18.250 160.145 19.460 160.895 ;
        RECT 18.250 159.605 18.770 160.145 ;
        RECT 20.090 160.125 21.760 160.895 ;
        RECT 21.930 160.170 22.220 160.895 ;
        RECT 18.940 159.435 19.460 159.975 ;
        RECT 18.250 158.345 19.460 159.435 ;
        RECT 20.090 159.435 20.840 159.955 ;
        RECT 21.010 159.605 21.760 160.125 ;
        RECT 22.390 160.095 22.730 160.725 ;
        RECT 22.900 160.095 23.150 160.895 ;
        RECT 23.340 160.245 23.670 160.725 ;
        RECT 23.840 160.435 24.065 160.895 ;
        RECT 24.235 160.245 24.565 160.725 ;
        RECT 20.090 158.345 21.760 159.435 ;
        RECT 21.930 158.345 22.220 159.510 ;
        RECT 22.390 159.485 22.565 160.095 ;
        RECT 23.340 160.075 24.565 160.245 ;
        RECT 25.195 160.115 25.695 160.725 ;
        RECT 22.735 159.735 23.430 159.905 ;
        RECT 23.260 159.485 23.430 159.735 ;
        RECT 23.605 159.705 24.025 159.905 ;
        RECT 24.195 159.705 24.525 159.905 ;
        RECT 24.695 159.705 25.025 159.905 ;
        RECT 25.195 159.485 25.365 160.115 ;
        RECT 26.345 160.085 26.590 160.690 ;
        RECT 26.810 160.360 27.320 160.895 ;
        RECT 26.070 159.915 27.300 160.085 ;
        RECT 25.550 159.655 25.900 159.905 ;
        RECT 22.390 158.515 22.730 159.485 ;
        RECT 22.900 158.345 23.070 159.485 ;
        RECT 23.260 159.315 25.695 159.485 ;
        RECT 23.340 158.345 23.590 159.145 ;
        RECT 24.235 158.515 24.565 159.315 ;
        RECT 24.865 158.345 25.195 159.145 ;
        RECT 25.365 158.515 25.695 159.315 ;
        RECT 26.070 159.105 26.410 159.915 ;
        RECT 26.580 159.350 27.330 159.540 ;
        RECT 26.070 158.695 26.585 159.105 ;
        RECT 26.820 158.345 26.990 159.105 ;
        RECT 27.160 158.685 27.330 159.350 ;
        RECT 27.500 159.365 27.690 160.725 ;
        RECT 27.860 159.875 28.135 160.725 ;
        RECT 28.325 160.360 28.855 160.725 ;
        RECT 29.280 160.495 29.610 160.895 ;
        RECT 28.680 160.325 28.855 160.360 ;
        RECT 27.860 159.705 28.140 159.875 ;
        RECT 27.860 159.565 28.135 159.705 ;
        RECT 28.340 159.365 28.510 160.165 ;
        RECT 27.500 159.195 28.510 159.365 ;
        RECT 28.680 160.155 29.610 160.325 ;
        RECT 29.780 160.155 30.035 160.725 ;
        RECT 30.320 160.415 30.490 160.895 ;
        RECT 30.660 160.245 30.990 160.720 ;
        RECT 31.160 160.415 31.330 160.895 ;
        RECT 31.500 160.245 31.830 160.720 ;
        RECT 32.000 160.415 32.170 160.895 ;
        RECT 32.340 160.245 32.670 160.720 ;
        RECT 32.840 160.415 33.010 160.895 ;
        RECT 33.180 160.245 33.510 160.720 ;
        RECT 33.680 160.415 33.850 160.895 ;
        RECT 34.020 160.245 34.350 160.720 ;
        RECT 34.520 160.415 34.690 160.895 ;
        RECT 34.940 160.720 35.110 160.725 ;
        RECT 34.860 160.245 35.190 160.720 ;
        RECT 35.360 160.415 35.530 160.895 ;
        RECT 35.780 160.720 35.950 160.725 ;
        RECT 35.700 160.245 36.030 160.720 ;
        RECT 36.200 160.415 36.370 160.895 ;
        RECT 36.620 160.720 36.870 160.725 ;
        RECT 36.540 160.245 36.870 160.720 ;
        RECT 37.040 160.415 37.210 160.895 ;
        RECT 37.380 160.245 37.710 160.720 ;
        RECT 37.880 160.415 38.050 160.895 ;
        RECT 38.220 160.245 38.550 160.720 ;
        RECT 38.720 160.415 38.890 160.895 ;
        RECT 39.060 160.245 39.390 160.720 ;
        RECT 39.560 160.415 39.730 160.895 ;
        RECT 39.900 160.245 40.230 160.720 ;
        RECT 40.400 160.415 40.570 160.895 ;
        RECT 40.740 160.245 41.070 160.720 ;
        RECT 28.680 159.025 28.850 160.155 ;
        RECT 29.440 159.985 29.610 160.155 ;
        RECT 27.725 158.855 28.850 159.025 ;
        RECT 29.020 159.655 29.215 159.985 ;
        RECT 29.440 159.655 29.695 159.985 ;
        RECT 29.020 158.685 29.190 159.655 ;
        RECT 29.865 159.485 30.035 160.155 ;
        RECT 27.160 158.515 29.190 158.685 ;
        RECT 29.360 158.345 29.530 159.485 ;
        RECT 29.700 158.515 30.035 159.485 ;
        RECT 30.210 160.075 36.870 160.245 ;
        RECT 37.040 160.075 39.390 160.245 ;
        RECT 39.560 160.075 41.070 160.245 ;
        RECT 41.710 160.125 43.380 160.895 ;
        RECT 30.210 159.535 30.485 160.075 ;
        RECT 37.040 159.905 37.215 160.075 ;
        RECT 39.560 159.905 39.730 160.075 ;
        RECT 30.655 159.705 37.215 159.905 ;
        RECT 37.420 159.705 39.730 159.905 ;
        RECT 39.900 159.705 41.075 159.905 ;
        RECT 37.040 159.535 37.215 159.705 ;
        RECT 39.560 159.535 39.730 159.705 ;
        RECT 30.210 159.365 36.870 159.535 ;
        RECT 37.040 159.365 39.390 159.535 ;
        RECT 39.560 159.365 41.070 159.535 ;
        RECT 30.320 158.345 30.490 159.145 ;
        RECT 30.660 158.515 30.990 159.365 ;
        RECT 31.160 158.345 31.330 159.145 ;
        RECT 31.500 158.515 31.830 159.365 ;
        RECT 32.000 158.345 32.170 159.145 ;
        RECT 32.340 158.515 32.670 159.365 ;
        RECT 32.840 158.345 33.010 159.145 ;
        RECT 33.180 158.515 33.510 159.365 ;
        RECT 33.680 158.345 33.850 159.145 ;
        RECT 34.020 158.515 34.350 159.365 ;
        RECT 34.520 158.345 34.690 159.145 ;
        RECT 34.860 158.515 35.190 159.365 ;
        RECT 35.360 158.345 35.530 159.145 ;
        RECT 35.700 158.515 36.030 159.365 ;
        RECT 36.200 158.345 36.370 159.145 ;
        RECT 36.540 158.515 36.870 159.365 ;
        RECT 37.040 158.345 37.210 159.145 ;
        RECT 37.380 158.515 37.710 159.365 ;
        RECT 37.880 158.345 38.050 159.145 ;
        RECT 38.220 158.515 38.550 159.365 ;
        RECT 38.720 158.345 38.890 159.145 ;
        RECT 39.060 158.515 39.390 159.365 ;
        RECT 39.560 158.345 39.730 159.195 ;
        RECT 39.900 158.515 40.230 159.365 ;
        RECT 40.400 158.345 40.570 159.195 ;
        RECT 40.740 158.515 41.070 159.365 ;
        RECT 41.710 159.435 42.460 159.955 ;
        RECT 42.630 159.605 43.380 160.125 ;
        RECT 43.825 160.085 44.070 160.690 ;
        RECT 44.290 160.360 44.800 160.895 ;
        RECT 43.550 159.915 44.780 160.085 ;
        RECT 41.710 158.345 43.380 159.435 ;
        RECT 43.550 159.105 43.890 159.915 ;
        RECT 44.060 159.350 44.810 159.540 ;
        RECT 43.550 158.695 44.065 159.105 ;
        RECT 44.300 158.345 44.470 159.105 ;
        RECT 44.640 158.685 44.810 159.350 ;
        RECT 44.980 159.365 45.170 160.725 ;
        RECT 45.340 160.555 45.615 160.725 ;
        RECT 45.340 160.385 45.620 160.555 ;
        RECT 45.340 159.565 45.615 160.385 ;
        RECT 45.805 160.360 46.335 160.725 ;
        RECT 46.760 160.495 47.090 160.895 ;
        RECT 46.160 160.325 46.335 160.360 ;
        RECT 45.820 159.365 45.990 160.165 ;
        RECT 44.980 159.195 45.990 159.365 ;
        RECT 46.160 160.155 47.090 160.325 ;
        RECT 47.260 160.155 47.515 160.725 ;
        RECT 47.690 160.170 47.980 160.895 ;
        RECT 46.160 159.025 46.330 160.155 ;
        RECT 46.920 159.985 47.090 160.155 ;
        RECT 45.205 158.855 46.330 159.025 ;
        RECT 46.500 159.655 46.695 159.985 ;
        RECT 46.920 159.655 47.175 159.985 ;
        RECT 46.500 158.685 46.670 159.655 ;
        RECT 47.345 159.485 47.515 160.155 ;
        RECT 48.150 160.095 48.490 160.725 ;
        RECT 48.660 160.095 48.910 160.895 ;
        RECT 49.100 160.245 49.430 160.725 ;
        RECT 49.600 160.435 49.825 160.895 ;
        RECT 49.995 160.245 50.325 160.725 ;
        RECT 44.640 158.515 46.670 158.685 ;
        RECT 46.840 158.345 47.010 159.485 ;
        RECT 47.180 158.515 47.515 159.485 ;
        RECT 47.690 158.345 47.980 159.510 ;
        RECT 48.150 159.485 48.325 160.095 ;
        RECT 49.100 160.075 50.325 160.245 ;
        RECT 50.955 160.115 51.455 160.725 ;
        RECT 48.495 159.735 49.190 159.905 ;
        RECT 49.020 159.485 49.190 159.735 ;
        RECT 49.365 159.705 49.785 159.905 ;
        RECT 49.955 159.705 50.285 159.905 ;
        RECT 50.455 159.705 50.785 159.905 ;
        RECT 50.955 159.485 51.125 160.115 ;
        RECT 51.830 160.095 52.170 160.725 ;
        RECT 52.340 160.095 52.590 160.895 ;
        RECT 52.780 160.245 53.110 160.725 ;
        RECT 53.280 160.435 53.505 160.895 ;
        RECT 53.675 160.245 54.005 160.725 ;
        RECT 51.310 159.655 51.660 159.905 ;
        RECT 51.830 159.485 52.005 160.095 ;
        RECT 52.780 160.075 54.005 160.245 ;
        RECT 54.635 160.115 55.135 160.725 ;
        RECT 52.175 159.735 52.870 159.905 ;
        RECT 52.700 159.485 52.870 159.735 ;
        RECT 53.045 159.705 53.465 159.905 ;
        RECT 53.635 159.705 53.965 159.905 ;
        RECT 54.135 159.705 54.465 159.905 ;
        RECT 54.635 159.485 54.805 160.115 ;
        RECT 55.660 160.095 55.990 160.895 ;
        RECT 56.160 160.245 56.330 160.725 ;
        RECT 56.500 160.415 56.830 160.895 ;
        RECT 57.000 160.245 57.170 160.725 ;
        RECT 57.420 160.415 57.660 160.895 ;
        RECT 57.840 160.245 58.010 160.725 ;
        RECT 56.160 160.075 57.170 160.245 ;
        RECT 57.375 160.075 58.010 160.245 ;
        RECT 58.270 160.220 58.530 160.725 ;
        RECT 58.710 160.515 59.040 160.895 ;
        RECT 59.220 160.345 59.390 160.725 ;
        RECT 56.160 160.045 56.660 160.075 ;
        RECT 54.990 159.655 55.340 159.905 ;
        RECT 56.160 159.535 56.655 160.045 ;
        RECT 57.375 159.905 57.545 160.075 ;
        RECT 57.045 159.735 57.545 159.905 ;
        RECT 48.150 158.515 48.490 159.485 ;
        RECT 48.660 158.345 48.830 159.485 ;
        RECT 49.020 159.315 51.455 159.485 ;
        RECT 49.100 158.345 49.350 159.145 ;
        RECT 49.995 158.515 50.325 159.315 ;
        RECT 50.625 158.345 50.955 159.145 ;
        RECT 51.125 158.515 51.455 159.315 ;
        RECT 51.830 158.515 52.170 159.485 ;
        RECT 52.340 158.345 52.510 159.485 ;
        RECT 52.700 159.315 55.135 159.485 ;
        RECT 52.780 158.345 53.030 159.145 ;
        RECT 53.675 158.515 54.005 159.315 ;
        RECT 54.305 158.345 54.635 159.145 ;
        RECT 54.805 158.515 55.135 159.315 ;
        RECT 55.660 158.345 55.990 159.495 ;
        RECT 56.160 159.365 57.170 159.535 ;
        RECT 56.160 158.515 56.330 159.365 ;
        RECT 56.500 158.345 56.830 159.145 ;
        RECT 57.000 158.515 57.170 159.365 ;
        RECT 57.375 159.495 57.545 159.735 ;
        RECT 57.715 159.665 58.095 159.905 ;
        RECT 57.375 159.325 58.090 159.495 ;
        RECT 57.350 158.345 57.590 159.145 ;
        RECT 57.760 158.515 58.090 159.325 ;
        RECT 58.270 159.420 58.440 160.220 ;
        RECT 58.725 160.175 59.390 160.345 ;
        RECT 58.725 159.920 58.895 160.175 ;
        RECT 59.655 160.055 59.915 160.895 ;
        RECT 60.090 160.150 60.345 160.725 ;
        RECT 60.515 160.515 60.845 160.895 ;
        RECT 61.060 160.345 61.230 160.725 ;
        RECT 60.515 160.175 61.230 160.345 ;
        RECT 58.610 159.590 58.895 159.920 ;
        RECT 59.130 159.625 59.460 159.995 ;
        RECT 58.725 159.445 58.895 159.590 ;
        RECT 58.270 158.515 58.540 159.420 ;
        RECT 58.725 159.275 59.390 159.445 ;
        RECT 58.710 158.345 59.040 159.105 ;
        RECT 59.220 158.515 59.390 159.275 ;
        RECT 59.655 158.345 59.915 159.495 ;
        RECT 60.090 159.420 60.260 160.150 ;
        RECT 60.515 159.985 60.685 160.175 ;
        RECT 61.495 160.055 61.755 160.895 ;
        RECT 61.930 160.150 62.185 160.725 ;
        RECT 62.355 160.515 62.685 160.895 ;
        RECT 62.900 160.345 63.070 160.725 ;
        RECT 62.355 160.175 63.070 160.345 ;
        RECT 60.430 159.655 60.685 159.985 ;
        RECT 60.515 159.445 60.685 159.655 ;
        RECT 60.965 159.625 61.320 159.995 ;
        RECT 60.090 158.515 60.345 159.420 ;
        RECT 60.515 159.275 61.230 159.445 ;
        RECT 60.515 158.345 60.845 159.105 ;
        RECT 61.060 158.515 61.230 159.275 ;
        RECT 61.495 158.345 61.755 159.495 ;
        RECT 61.930 159.420 62.100 160.150 ;
        RECT 62.355 159.985 62.525 160.175 ;
        RECT 63.335 160.055 63.595 160.895 ;
        RECT 63.770 160.150 64.025 160.725 ;
        RECT 64.195 160.515 64.525 160.895 ;
        RECT 64.740 160.345 64.910 160.725 ;
        RECT 64.195 160.175 64.910 160.345 ;
        RECT 62.270 159.655 62.525 159.985 ;
        RECT 62.355 159.445 62.525 159.655 ;
        RECT 62.805 159.625 63.160 159.995 ;
        RECT 61.930 158.515 62.185 159.420 ;
        RECT 62.355 159.275 63.070 159.445 ;
        RECT 62.355 158.345 62.685 159.105 ;
        RECT 62.900 158.515 63.070 159.275 ;
        RECT 63.335 158.345 63.595 159.495 ;
        RECT 63.770 159.420 63.940 160.150 ;
        RECT 64.195 159.985 64.365 160.175 ;
        RECT 65.175 160.055 65.435 160.895 ;
        RECT 65.610 160.150 65.865 160.725 ;
        RECT 66.035 160.515 66.365 160.895 ;
        RECT 66.580 160.345 66.750 160.725 ;
        RECT 66.035 160.175 66.750 160.345 ;
        RECT 64.110 159.655 64.365 159.985 ;
        RECT 64.195 159.445 64.365 159.655 ;
        RECT 64.645 159.625 65.000 159.995 ;
        RECT 63.770 158.515 64.025 159.420 ;
        RECT 64.195 159.275 64.910 159.445 ;
        RECT 64.195 158.345 64.525 159.105 ;
        RECT 64.740 158.515 64.910 159.275 ;
        RECT 65.175 158.345 65.435 159.495 ;
        RECT 65.610 159.420 65.780 160.150 ;
        RECT 66.035 159.985 66.205 160.175 ;
        RECT 67.010 160.125 69.600 160.895 ;
        RECT 65.950 159.655 66.205 159.985 ;
        RECT 66.035 159.445 66.205 159.655 ;
        RECT 66.485 159.625 66.840 159.995 ;
        RECT 65.610 158.515 65.865 159.420 ;
        RECT 66.035 159.275 66.750 159.445 ;
        RECT 66.035 158.345 66.365 159.105 ;
        RECT 66.580 158.515 66.750 159.275 ;
        RECT 67.010 159.435 68.220 159.955 ;
        RECT 68.390 159.605 69.600 160.125 ;
        RECT 69.770 160.095 70.110 160.725 ;
        RECT 70.280 160.095 70.530 160.895 ;
        RECT 70.720 160.245 71.050 160.725 ;
        RECT 71.220 160.435 71.445 160.895 ;
        RECT 71.615 160.245 71.945 160.725 ;
        RECT 69.770 159.485 69.945 160.095 ;
        RECT 70.720 160.075 71.945 160.245 ;
        RECT 72.575 160.115 73.075 160.725 ;
        RECT 73.450 160.170 73.740 160.895 ;
        RECT 70.115 159.735 70.810 159.905 ;
        RECT 70.640 159.485 70.810 159.735 ;
        RECT 70.985 159.705 71.405 159.905 ;
        RECT 71.575 159.705 71.905 159.905 ;
        RECT 72.075 159.705 72.405 159.905 ;
        RECT 72.575 159.485 72.745 160.115 ;
        RECT 73.970 160.075 74.180 160.895 ;
        RECT 74.350 160.095 74.680 160.725 ;
        RECT 72.930 159.655 73.280 159.905 ;
        RECT 67.010 158.345 69.600 159.435 ;
        RECT 69.770 158.515 70.110 159.485 ;
        RECT 70.280 158.345 70.450 159.485 ;
        RECT 70.640 159.315 73.075 159.485 ;
        RECT 70.720 158.345 70.970 159.145 ;
        RECT 71.615 158.515 71.945 159.315 ;
        RECT 72.245 158.345 72.575 159.145 ;
        RECT 72.745 158.515 73.075 159.315 ;
        RECT 73.450 158.345 73.740 159.510 ;
        RECT 74.350 159.495 74.600 160.095 ;
        RECT 74.850 160.075 75.080 160.895 ;
        RECT 75.380 160.345 75.550 160.725 ;
        RECT 75.730 160.515 76.060 160.895 ;
        RECT 75.380 160.175 76.045 160.345 ;
        RECT 76.240 160.220 76.500 160.725 ;
        RECT 74.770 159.655 75.100 159.905 ;
        RECT 75.310 159.625 75.640 159.995 ;
        RECT 75.875 159.920 76.045 160.175 ;
        RECT 75.875 159.590 76.160 159.920 ;
        RECT 73.970 158.345 74.180 159.485 ;
        RECT 74.350 158.515 74.680 159.495 ;
        RECT 74.850 158.345 75.080 159.485 ;
        RECT 75.875 159.445 76.045 159.590 ;
        RECT 75.380 159.275 76.045 159.445 ;
        RECT 76.330 159.420 76.500 160.220 ;
        RECT 77.045 160.185 77.300 160.715 ;
        RECT 77.480 160.435 77.765 160.895 ;
        RECT 77.045 159.875 77.225 160.185 ;
        RECT 77.945 159.985 78.195 160.635 ;
        RECT 76.960 159.705 77.225 159.875 ;
        RECT 75.380 158.515 75.550 159.275 ;
        RECT 75.730 158.345 76.060 159.105 ;
        RECT 76.230 158.515 76.500 159.420 ;
        RECT 77.045 159.325 77.225 159.705 ;
        RECT 77.395 159.655 78.195 159.985 ;
        RECT 77.045 158.655 77.300 159.325 ;
        RECT 77.480 158.345 77.765 159.145 ;
        RECT 77.945 159.065 78.195 159.655 ;
        RECT 78.395 160.300 78.715 160.630 ;
        RECT 78.895 160.415 79.555 160.895 ;
        RECT 79.755 160.505 80.605 160.675 ;
        RECT 78.395 159.405 78.585 160.300 ;
        RECT 78.905 159.975 79.565 160.245 ;
        RECT 79.235 159.915 79.565 159.975 ;
        RECT 78.755 159.745 79.085 159.805 ;
        RECT 79.755 159.745 79.925 160.505 ;
        RECT 81.165 160.435 81.485 160.895 ;
        RECT 81.685 160.255 81.935 160.685 ;
        RECT 82.225 160.455 82.635 160.895 ;
        RECT 82.805 160.515 83.820 160.715 ;
        RECT 80.095 160.085 81.345 160.255 ;
        RECT 80.095 159.965 80.425 160.085 ;
        RECT 78.755 159.575 80.655 159.745 ;
        RECT 78.395 159.235 80.315 159.405 ;
        RECT 78.395 159.215 78.715 159.235 ;
        RECT 77.945 158.555 78.275 159.065 ;
        RECT 78.545 158.605 78.715 159.215 ;
        RECT 80.485 159.065 80.655 159.575 ;
        RECT 80.825 159.505 81.005 159.915 ;
        RECT 81.175 159.325 81.345 160.085 ;
        RECT 78.885 158.345 79.215 159.035 ;
        RECT 79.445 158.895 80.655 159.065 ;
        RECT 80.825 159.015 81.345 159.325 ;
        RECT 81.515 159.915 81.935 160.255 ;
        RECT 82.225 159.915 82.635 160.245 ;
        RECT 81.515 159.145 81.705 159.915 ;
        RECT 82.805 159.785 82.975 160.515 ;
        RECT 84.120 160.345 84.290 160.675 ;
        RECT 84.460 160.515 84.790 160.895 ;
        RECT 83.145 159.965 83.495 160.335 ;
        RECT 82.805 159.745 83.225 159.785 ;
        RECT 81.875 159.575 83.225 159.745 ;
        RECT 81.875 159.415 82.125 159.575 ;
        RECT 82.635 159.145 82.885 159.405 ;
        RECT 81.515 158.895 82.885 159.145 ;
        RECT 79.445 158.605 79.685 158.895 ;
        RECT 80.485 158.815 80.655 158.895 ;
        RECT 79.885 158.345 80.305 158.725 ;
        RECT 80.485 158.565 81.115 158.815 ;
        RECT 81.585 158.345 81.915 158.725 ;
        RECT 82.085 158.605 82.255 158.895 ;
        RECT 83.055 158.730 83.225 159.575 ;
        RECT 83.675 159.405 83.895 160.275 ;
        RECT 84.120 160.155 84.815 160.345 ;
        RECT 83.395 159.025 83.895 159.405 ;
        RECT 84.065 159.355 84.475 159.975 ;
        RECT 84.645 159.185 84.815 160.155 ;
        RECT 84.120 159.015 84.815 159.185 ;
        RECT 82.435 158.345 82.815 158.725 ;
        RECT 83.055 158.560 83.885 158.730 ;
        RECT 84.120 158.515 84.290 159.015 ;
        RECT 84.460 158.345 84.790 158.845 ;
        RECT 85.005 158.515 85.230 160.635 ;
        RECT 85.400 160.515 85.730 160.895 ;
        RECT 85.900 160.345 86.070 160.635 ;
        RECT 86.420 160.415 86.720 160.895 ;
        RECT 85.405 160.175 86.070 160.345 ;
        RECT 86.890 160.245 87.150 160.700 ;
        RECT 87.320 160.415 87.580 160.895 ;
        RECT 87.760 160.245 88.020 160.700 ;
        RECT 88.190 160.415 88.440 160.895 ;
        RECT 88.620 160.245 88.880 160.700 ;
        RECT 89.050 160.415 89.300 160.895 ;
        RECT 89.480 160.245 89.740 160.700 ;
        RECT 89.910 160.415 90.155 160.895 ;
        RECT 90.325 160.245 90.600 160.700 ;
        RECT 90.770 160.415 91.015 160.895 ;
        RECT 91.185 160.245 91.445 160.700 ;
        RECT 91.615 160.415 91.875 160.895 ;
        RECT 92.045 160.245 92.305 160.700 ;
        RECT 92.475 160.415 92.735 160.895 ;
        RECT 92.905 160.245 93.165 160.700 ;
        RECT 93.335 160.335 93.595 160.895 ;
        RECT 85.405 159.185 85.635 160.175 ;
        RECT 86.420 160.075 93.165 160.245 ;
        RECT 85.805 159.355 86.155 160.005 ;
        RECT 86.420 159.485 87.585 160.075 ;
        RECT 93.765 159.905 94.015 160.715 ;
        RECT 94.195 160.370 94.455 160.895 ;
        RECT 94.625 159.905 94.875 160.715 ;
        RECT 95.055 160.385 95.360 160.895 ;
        RECT 87.755 159.655 94.875 159.905 ;
        RECT 95.045 159.655 95.360 160.215 ;
        RECT 95.530 160.095 95.870 160.725 ;
        RECT 96.040 160.095 96.290 160.895 ;
        RECT 96.480 160.245 96.810 160.725 ;
        RECT 96.980 160.435 97.205 160.895 ;
        RECT 97.375 160.245 97.705 160.725 ;
        RECT 86.420 159.260 93.165 159.485 ;
        RECT 85.405 159.015 86.070 159.185 ;
        RECT 85.400 158.345 85.730 158.845 ;
        RECT 85.900 158.515 86.070 159.015 ;
        RECT 86.420 158.345 86.690 159.090 ;
        RECT 86.860 158.520 87.150 159.260 ;
        RECT 87.760 159.245 93.165 159.260 ;
        RECT 87.320 158.350 87.575 159.075 ;
        RECT 87.760 158.520 88.020 159.245 ;
        RECT 88.190 158.350 88.435 159.075 ;
        RECT 88.620 158.520 88.880 159.245 ;
        RECT 89.050 158.350 89.295 159.075 ;
        RECT 89.480 158.520 89.740 159.245 ;
        RECT 89.910 158.350 90.155 159.075 ;
        RECT 90.325 158.520 90.585 159.245 ;
        RECT 90.755 158.350 91.015 159.075 ;
        RECT 91.185 158.520 91.445 159.245 ;
        RECT 91.615 158.350 91.875 159.075 ;
        RECT 92.045 158.520 92.305 159.245 ;
        RECT 92.475 158.350 92.735 159.075 ;
        RECT 92.905 158.520 93.165 159.245 ;
        RECT 93.335 158.350 93.595 159.145 ;
        RECT 93.765 158.520 94.015 159.655 ;
        RECT 87.320 158.345 93.595 158.350 ;
        RECT 94.195 158.345 94.455 159.155 ;
        RECT 94.630 158.515 94.875 159.655 ;
        RECT 95.530 159.485 95.705 160.095 ;
        RECT 96.480 160.075 97.705 160.245 ;
        RECT 98.335 160.115 98.835 160.725 ;
        RECT 99.210 160.170 99.500 160.895 ;
        RECT 99.670 160.125 101.340 160.895 ;
        RECT 101.885 160.555 102.140 160.715 ;
        RECT 101.800 160.385 102.140 160.555 ;
        RECT 102.320 160.435 102.605 160.895 ;
        RECT 95.875 159.735 96.570 159.905 ;
        RECT 96.400 159.485 96.570 159.735 ;
        RECT 96.745 159.705 97.165 159.905 ;
        RECT 97.335 159.705 97.665 159.905 ;
        RECT 97.835 159.705 98.165 159.905 ;
        RECT 98.335 159.485 98.505 160.115 ;
        RECT 98.690 159.655 99.040 159.905 ;
        RECT 95.055 158.345 95.350 159.155 ;
        RECT 95.530 158.515 95.870 159.485 ;
        RECT 96.040 158.345 96.210 159.485 ;
        RECT 96.400 159.315 98.835 159.485 ;
        RECT 96.480 158.345 96.730 159.145 ;
        RECT 97.375 158.515 97.705 159.315 ;
        RECT 98.005 158.345 98.335 159.145 ;
        RECT 98.505 158.515 98.835 159.315 ;
        RECT 99.210 158.345 99.500 159.510 ;
        RECT 99.670 159.435 100.420 159.955 ;
        RECT 100.590 159.605 101.340 160.125 ;
        RECT 101.885 160.185 102.140 160.385 ;
        RECT 99.670 158.345 101.340 159.435 ;
        RECT 101.885 159.325 102.065 160.185 ;
        RECT 102.785 159.985 103.035 160.635 ;
        RECT 102.235 159.655 103.035 159.985 ;
        RECT 101.885 158.655 102.140 159.325 ;
        RECT 102.320 158.345 102.605 159.145 ;
        RECT 102.785 159.065 103.035 159.655 ;
        RECT 103.235 160.300 103.555 160.630 ;
        RECT 103.735 160.415 104.395 160.895 ;
        RECT 104.595 160.505 105.445 160.675 ;
        RECT 103.235 159.405 103.425 160.300 ;
        RECT 103.745 159.975 104.405 160.245 ;
        RECT 104.075 159.915 104.405 159.975 ;
        RECT 103.595 159.745 103.925 159.805 ;
        RECT 104.595 159.745 104.765 160.505 ;
        RECT 106.005 160.435 106.325 160.895 ;
        RECT 106.525 160.255 106.775 160.685 ;
        RECT 107.065 160.455 107.475 160.895 ;
        RECT 107.645 160.515 108.660 160.715 ;
        RECT 104.935 160.085 106.185 160.255 ;
        RECT 104.935 159.965 105.265 160.085 ;
        RECT 103.595 159.575 105.495 159.745 ;
        RECT 103.235 159.235 105.155 159.405 ;
        RECT 103.235 159.215 103.555 159.235 ;
        RECT 102.785 158.555 103.115 159.065 ;
        RECT 103.385 158.605 103.555 159.215 ;
        RECT 105.325 159.065 105.495 159.575 ;
        RECT 105.665 159.505 105.845 159.915 ;
        RECT 106.015 159.325 106.185 160.085 ;
        RECT 103.725 158.345 104.055 159.035 ;
        RECT 104.285 158.895 105.495 159.065 ;
        RECT 105.665 159.015 106.185 159.325 ;
        RECT 106.355 159.915 106.775 160.255 ;
        RECT 107.065 159.915 107.475 160.245 ;
        RECT 106.355 159.145 106.545 159.915 ;
        RECT 107.645 159.785 107.815 160.515 ;
        RECT 108.960 160.345 109.130 160.675 ;
        RECT 109.300 160.515 109.630 160.895 ;
        RECT 107.985 159.965 108.335 160.335 ;
        RECT 107.645 159.745 108.065 159.785 ;
        RECT 106.715 159.575 108.065 159.745 ;
        RECT 106.715 159.415 106.965 159.575 ;
        RECT 107.475 159.145 107.725 159.405 ;
        RECT 106.355 158.895 107.725 159.145 ;
        RECT 104.285 158.605 104.525 158.895 ;
        RECT 105.325 158.815 105.495 158.895 ;
        RECT 104.725 158.345 105.145 158.725 ;
        RECT 105.325 158.565 105.955 158.815 ;
        RECT 106.425 158.345 106.755 158.725 ;
        RECT 106.925 158.605 107.095 158.895 ;
        RECT 107.895 158.730 108.065 159.575 ;
        RECT 108.515 159.405 108.735 160.275 ;
        RECT 108.960 160.155 109.655 160.345 ;
        RECT 108.235 159.025 108.735 159.405 ;
        RECT 108.905 159.355 109.315 159.975 ;
        RECT 109.485 159.185 109.655 160.155 ;
        RECT 108.960 159.015 109.655 159.185 ;
        RECT 107.275 158.345 107.655 158.725 ;
        RECT 107.895 158.560 108.725 158.730 ;
        RECT 108.960 158.515 109.130 159.015 ;
        RECT 109.300 158.345 109.630 158.845 ;
        RECT 109.845 158.515 110.070 160.635 ;
        RECT 110.240 160.515 110.570 160.895 ;
        RECT 110.740 160.345 110.910 160.635 ;
        RECT 110.245 160.175 110.910 160.345 ;
        RECT 110.245 159.185 110.475 160.175 ;
        RECT 111.170 160.145 112.380 160.895 ;
        RECT 110.645 159.355 110.995 160.005 ;
        RECT 111.170 159.435 111.690 159.975 ;
        RECT 111.860 159.605 112.380 160.145 ;
        RECT 110.245 159.015 110.910 159.185 ;
        RECT 110.240 158.345 110.570 158.845 ;
        RECT 110.740 158.515 110.910 159.015 ;
        RECT 111.170 158.345 112.380 159.435 ;
        RECT 18.165 158.175 112.465 158.345 ;
        RECT 18.250 157.085 19.460 158.175 ;
        RECT 18.250 156.375 18.770 156.915 ;
        RECT 18.940 156.545 19.460 157.085 ;
        RECT 20.150 157.035 20.360 158.175 ;
        RECT 20.530 157.025 20.860 158.005 ;
        RECT 21.030 157.035 21.260 158.175 ;
        RECT 21.475 157.035 21.810 158.005 ;
        RECT 21.980 157.035 22.150 158.175 ;
        RECT 22.320 157.835 24.350 158.005 ;
        RECT 18.250 155.625 19.460 156.375 ;
        RECT 20.150 155.625 20.360 156.445 ;
        RECT 20.530 156.425 20.780 157.025 ;
        RECT 20.950 156.615 21.280 156.865 ;
        RECT 20.530 155.795 20.860 156.425 ;
        RECT 21.030 155.625 21.260 156.445 ;
        RECT 21.475 156.365 21.645 157.035 ;
        RECT 22.320 156.865 22.490 157.835 ;
        RECT 21.815 156.535 22.070 156.865 ;
        RECT 22.295 156.535 22.490 156.865 ;
        RECT 22.660 157.495 23.785 157.665 ;
        RECT 21.900 156.365 22.070 156.535 ;
        RECT 22.660 156.365 22.830 157.495 ;
        RECT 21.475 155.795 21.730 156.365 ;
        RECT 21.900 156.195 22.830 156.365 ;
        RECT 23.000 157.155 24.010 157.325 ;
        RECT 23.000 156.355 23.170 157.155 ;
        RECT 22.655 156.160 22.830 156.195 ;
        RECT 21.900 155.625 22.230 156.025 ;
        RECT 22.655 155.795 23.185 156.160 ;
        RECT 23.375 156.135 23.650 156.955 ;
        RECT 23.370 155.965 23.650 156.135 ;
        RECT 23.375 155.795 23.650 155.965 ;
        RECT 23.820 155.795 24.010 157.155 ;
        RECT 24.180 157.170 24.350 157.835 ;
        RECT 24.520 157.415 24.690 158.175 ;
        RECT 24.925 157.415 25.440 157.825 ;
        RECT 24.180 156.980 24.930 157.170 ;
        RECT 25.100 156.605 25.440 157.415 ;
        RECT 24.210 156.435 25.440 156.605 ;
        RECT 25.615 156.985 25.870 157.865 ;
        RECT 26.040 157.035 26.345 158.175 ;
        RECT 26.685 157.795 27.015 158.175 ;
        RECT 27.195 157.625 27.365 157.915 ;
        RECT 27.535 157.715 27.785 158.175 ;
        RECT 26.565 157.455 27.365 157.625 ;
        RECT 27.955 157.665 28.825 158.005 ;
        RECT 24.190 155.625 24.700 156.160 ;
        RECT 24.920 155.830 25.165 156.435 ;
        RECT 25.615 156.335 25.825 156.985 ;
        RECT 26.565 156.865 26.735 157.455 ;
        RECT 27.955 157.285 28.125 157.665 ;
        RECT 29.060 157.545 29.230 158.005 ;
        RECT 29.400 157.715 29.770 158.175 ;
        RECT 30.065 157.575 30.235 157.915 ;
        RECT 30.405 157.745 30.735 158.175 ;
        RECT 30.970 157.575 31.140 157.915 ;
        RECT 26.905 157.115 28.125 157.285 ;
        RECT 28.295 157.205 28.755 157.495 ;
        RECT 29.060 157.375 29.620 157.545 ;
        RECT 30.065 157.405 31.140 157.575 ;
        RECT 31.310 157.675 31.990 158.005 ;
        RECT 32.205 157.675 32.455 158.005 ;
        RECT 32.625 157.715 32.875 158.175 ;
        RECT 29.450 157.235 29.620 157.375 ;
        RECT 28.295 157.195 29.260 157.205 ;
        RECT 27.955 157.025 28.125 157.115 ;
        RECT 28.585 157.035 29.260 157.195 ;
        RECT 25.995 156.835 26.735 156.865 ;
        RECT 25.995 156.535 26.910 156.835 ;
        RECT 26.585 156.360 26.910 156.535 ;
        RECT 25.615 155.805 25.870 156.335 ;
        RECT 26.040 155.625 26.345 156.085 ;
        RECT 26.590 156.005 26.910 156.360 ;
        RECT 27.080 156.575 27.620 156.945 ;
        RECT 27.955 156.855 28.360 157.025 ;
        RECT 27.080 156.175 27.320 156.575 ;
        RECT 27.800 156.405 28.020 156.685 ;
        RECT 27.490 156.235 28.020 156.405 ;
        RECT 27.490 156.005 27.660 156.235 ;
        RECT 28.190 156.075 28.360 156.855 ;
        RECT 28.530 156.245 28.880 156.865 ;
        RECT 29.050 156.245 29.260 157.035 ;
        RECT 29.450 157.065 30.950 157.235 ;
        RECT 29.450 156.375 29.620 157.065 ;
        RECT 31.310 156.895 31.480 157.675 ;
        RECT 32.285 157.545 32.455 157.675 ;
        RECT 29.790 156.725 31.480 156.895 ;
        RECT 31.650 157.115 32.115 157.505 ;
        RECT 32.285 157.375 32.680 157.545 ;
        RECT 29.790 156.545 29.960 156.725 ;
        RECT 26.590 155.835 27.660 156.005 ;
        RECT 27.830 155.625 28.020 156.065 ;
        RECT 28.190 155.795 29.140 156.075 ;
        RECT 29.450 155.985 29.710 156.375 ;
        RECT 30.130 156.305 30.920 156.555 ;
        RECT 29.360 155.815 29.710 155.985 ;
        RECT 29.920 155.625 30.250 156.085 ;
        RECT 31.125 156.015 31.295 156.725 ;
        RECT 31.650 156.525 31.820 157.115 ;
        RECT 31.465 156.305 31.820 156.525 ;
        RECT 31.990 156.305 32.340 156.925 ;
        RECT 32.510 156.015 32.680 157.375 ;
        RECT 33.045 157.205 33.370 157.990 ;
        RECT 32.850 156.155 33.310 157.205 ;
        RECT 31.125 155.845 31.980 156.015 ;
        RECT 32.185 155.845 32.680 156.015 ;
        RECT 32.850 155.625 33.180 155.985 ;
        RECT 33.540 155.885 33.710 158.005 ;
        RECT 33.880 157.675 34.210 158.175 ;
        RECT 34.380 157.505 34.635 158.005 ;
        RECT 33.885 157.335 34.635 157.505 ;
        RECT 33.885 156.345 34.115 157.335 ;
        RECT 34.285 156.515 34.635 157.165 ;
        RECT 34.810 157.010 35.100 158.175 ;
        RECT 35.275 156.985 35.530 157.865 ;
        RECT 35.700 157.035 36.005 158.175 ;
        RECT 36.345 157.795 36.675 158.175 ;
        RECT 36.855 157.625 37.025 157.915 ;
        RECT 37.195 157.715 37.445 158.175 ;
        RECT 36.225 157.455 37.025 157.625 ;
        RECT 37.615 157.665 38.485 158.005 ;
        RECT 33.885 156.175 34.635 156.345 ;
        RECT 33.880 155.625 34.210 156.005 ;
        RECT 34.380 155.885 34.635 156.175 ;
        RECT 34.810 155.625 35.100 156.350 ;
        RECT 35.275 156.335 35.485 156.985 ;
        RECT 36.225 156.865 36.395 157.455 ;
        RECT 37.615 157.285 37.785 157.665 ;
        RECT 38.720 157.545 38.890 158.005 ;
        RECT 39.060 157.715 39.430 158.175 ;
        RECT 39.725 157.575 39.895 157.915 ;
        RECT 40.065 157.745 40.395 158.175 ;
        RECT 40.630 157.575 40.800 157.915 ;
        RECT 36.565 157.115 37.785 157.285 ;
        RECT 37.955 157.205 38.415 157.495 ;
        RECT 38.720 157.375 39.280 157.545 ;
        RECT 39.725 157.405 40.800 157.575 ;
        RECT 40.970 157.675 41.650 158.005 ;
        RECT 41.865 157.675 42.115 158.005 ;
        RECT 42.285 157.715 42.535 158.175 ;
        RECT 39.110 157.235 39.280 157.375 ;
        RECT 37.955 157.195 38.920 157.205 ;
        RECT 37.615 157.025 37.785 157.115 ;
        RECT 38.245 157.035 38.920 157.195 ;
        RECT 35.655 156.835 36.395 156.865 ;
        RECT 35.655 156.535 36.570 156.835 ;
        RECT 36.245 156.360 36.570 156.535 ;
        RECT 35.275 155.805 35.530 156.335 ;
        RECT 35.700 155.625 36.005 156.085 ;
        RECT 36.250 156.005 36.570 156.360 ;
        RECT 36.740 156.575 37.280 156.945 ;
        RECT 37.615 156.855 38.020 157.025 ;
        RECT 36.740 156.175 36.980 156.575 ;
        RECT 37.460 156.405 37.680 156.685 ;
        RECT 37.150 156.235 37.680 156.405 ;
        RECT 37.150 156.005 37.320 156.235 ;
        RECT 37.850 156.075 38.020 156.855 ;
        RECT 38.190 156.245 38.540 156.865 ;
        RECT 38.710 156.245 38.920 157.035 ;
        RECT 39.110 157.065 40.610 157.235 ;
        RECT 39.110 156.375 39.280 157.065 ;
        RECT 40.970 156.895 41.140 157.675 ;
        RECT 41.945 157.545 42.115 157.675 ;
        RECT 39.450 156.725 41.140 156.895 ;
        RECT 41.310 157.115 41.775 157.505 ;
        RECT 41.945 157.375 42.340 157.545 ;
        RECT 39.450 156.545 39.620 156.725 ;
        RECT 36.250 155.835 37.320 156.005 ;
        RECT 37.490 155.625 37.680 156.065 ;
        RECT 37.850 155.795 38.800 156.075 ;
        RECT 39.110 155.985 39.370 156.375 ;
        RECT 39.790 156.305 40.580 156.555 ;
        RECT 39.020 155.815 39.370 155.985 ;
        RECT 39.580 155.625 39.910 156.085 ;
        RECT 40.785 156.015 40.955 156.725 ;
        RECT 41.310 156.525 41.480 157.115 ;
        RECT 41.125 156.305 41.480 156.525 ;
        RECT 41.650 156.305 42.000 156.925 ;
        RECT 42.170 156.015 42.340 157.375 ;
        RECT 42.705 157.205 43.030 157.990 ;
        RECT 42.510 156.155 42.970 157.205 ;
        RECT 40.785 155.845 41.640 156.015 ;
        RECT 41.845 155.845 42.340 156.015 ;
        RECT 42.510 155.625 42.840 155.985 ;
        RECT 43.200 155.885 43.370 158.005 ;
        RECT 43.540 157.675 43.870 158.175 ;
        RECT 44.040 157.505 44.295 158.005 ;
        RECT 43.545 157.335 44.295 157.505 ;
        RECT 43.545 156.345 43.775 157.335 ;
        RECT 43.945 156.515 44.295 157.165 ;
        RECT 45.390 157.035 45.730 158.005 ;
        RECT 45.900 157.035 46.070 158.175 ;
        RECT 46.340 157.375 46.590 158.175 ;
        RECT 47.235 157.205 47.565 158.005 ;
        RECT 47.865 157.375 48.195 158.175 ;
        RECT 48.365 157.205 48.695 158.005 ;
        RECT 46.260 157.035 48.695 157.205 ;
        RECT 49.275 157.205 49.605 158.005 ;
        RECT 49.775 157.375 50.105 158.175 ;
        RECT 50.405 157.205 50.735 158.005 ;
        RECT 51.380 157.375 51.630 158.175 ;
        RECT 49.275 157.035 51.710 157.205 ;
        RECT 51.900 157.035 52.070 158.175 ;
        RECT 52.240 157.035 52.580 158.005 ;
        RECT 45.390 156.425 45.565 157.035 ;
        RECT 46.260 156.785 46.430 157.035 ;
        RECT 45.735 156.615 46.430 156.785 ;
        RECT 46.605 156.615 47.025 156.815 ;
        RECT 47.195 156.615 47.525 156.815 ;
        RECT 47.695 156.615 48.025 156.815 ;
        RECT 43.545 156.175 44.295 156.345 ;
        RECT 43.540 155.625 43.870 156.005 ;
        RECT 44.040 155.885 44.295 156.175 ;
        RECT 45.390 155.795 45.730 156.425 ;
        RECT 45.900 155.625 46.150 156.425 ;
        RECT 46.340 156.275 47.565 156.445 ;
        RECT 46.340 155.795 46.670 156.275 ;
        RECT 46.840 155.625 47.065 156.085 ;
        RECT 47.235 155.795 47.565 156.275 ;
        RECT 48.195 156.405 48.365 157.035 ;
        RECT 48.550 156.615 48.900 156.865 ;
        RECT 49.070 156.615 49.420 156.865 ;
        RECT 49.605 156.405 49.775 157.035 ;
        RECT 49.945 156.615 50.275 156.815 ;
        RECT 50.445 156.615 50.775 156.815 ;
        RECT 50.945 156.615 51.365 156.815 ;
        RECT 51.540 156.785 51.710 157.035 ;
        RECT 51.540 156.615 52.235 156.785 ;
        RECT 48.195 155.795 48.695 156.405 ;
        RECT 49.275 155.795 49.775 156.405 ;
        RECT 50.405 156.275 51.630 156.445 ;
        RECT 52.405 156.425 52.580 157.035 ;
        RECT 52.900 157.025 53.230 158.175 ;
        RECT 53.400 157.155 53.570 158.005 ;
        RECT 53.740 157.375 54.070 158.175 ;
        RECT 54.240 157.155 54.410 158.005 ;
        RECT 54.590 157.375 54.830 158.175 ;
        RECT 55.000 157.195 55.330 158.005 ;
        RECT 53.400 156.985 54.410 157.155 ;
        RECT 54.615 157.025 55.330 157.195 ;
        RECT 55.510 157.085 57.180 158.175 ;
        RECT 53.400 156.445 53.895 156.985 ;
        RECT 54.615 156.785 54.785 157.025 ;
        RECT 54.285 156.615 54.785 156.785 ;
        RECT 54.955 156.615 55.335 156.855 ;
        RECT 54.615 156.445 54.785 156.615 ;
        RECT 55.510 156.565 56.260 157.085 ;
        RECT 57.390 157.035 57.620 158.175 ;
        RECT 57.790 157.025 58.120 158.005 ;
        RECT 58.290 157.035 58.500 158.175 ;
        RECT 58.735 157.025 58.995 158.175 ;
        RECT 59.170 157.100 59.425 158.005 ;
        RECT 59.595 157.415 59.925 158.175 ;
        RECT 60.140 157.245 60.310 158.005 ;
        RECT 50.405 155.795 50.735 156.275 ;
        RECT 50.905 155.625 51.130 156.085 ;
        RECT 51.300 155.795 51.630 156.275 ;
        RECT 51.820 155.625 52.070 156.425 ;
        RECT 52.240 155.795 52.580 156.425 ;
        RECT 52.900 155.625 53.230 156.425 ;
        RECT 53.400 156.275 54.410 156.445 ;
        RECT 54.615 156.275 55.250 156.445 ;
        RECT 56.430 156.395 57.180 156.915 ;
        RECT 57.370 156.615 57.700 156.865 ;
        RECT 53.400 155.795 53.570 156.275 ;
        RECT 53.740 155.625 54.070 156.105 ;
        RECT 54.240 155.795 54.410 156.275 ;
        RECT 54.660 155.625 54.900 156.105 ;
        RECT 55.080 155.795 55.250 156.275 ;
        RECT 55.510 155.625 57.180 156.395 ;
        RECT 57.390 155.625 57.620 156.445 ;
        RECT 57.870 156.425 58.120 157.025 ;
        RECT 57.790 155.795 58.120 156.425 ;
        RECT 58.290 155.625 58.500 156.445 ;
        RECT 58.735 155.625 58.995 156.465 ;
        RECT 59.170 156.370 59.340 157.100 ;
        RECT 59.595 157.075 60.310 157.245 ;
        RECT 59.595 156.865 59.765 157.075 ;
        RECT 60.570 157.010 60.860 158.175 ;
        RECT 61.085 157.305 61.370 158.175 ;
        RECT 61.540 157.545 61.800 158.005 ;
        RECT 61.975 157.715 62.230 158.175 ;
        RECT 62.400 157.545 62.660 158.005 ;
        RECT 61.540 157.375 62.660 157.545 ;
        RECT 62.830 157.375 63.140 158.175 ;
        RECT 61.540 157.125 61.800 157.375 ;
        RECT 63.310 157.205 63.620 158.005 ;
        RECT 61.045 156.955 61.800 157.125 ;
        RECT 62.590 157.035 63.620 157.205 ;
        RECT 59.510 156.535 59.765 156.865 ;
        RECT 59.170 155.795 59.425 156.370 ;
        RECT 59.595 156.345 59.765 156.535 ;
        RECT 60.045 156.525 60.400 156.895 ;
        RECT 61.045 156.445 61.450 156.955 ;
        RECT 62.590 156.785 62.760 157.035 ;
        RECT 61.620 156.615 62.760 156.785 ;
        RECT 59.595 156.175 60.310 156.345 ;
        RECT 59.595 155.625 59.925 156.005 ;
        RECT 60.140 155.795 60.310 156.175 ;
        RECT 60.570 155.625 60.860 156.350 ;
        RECT 61.045 156.275 62.695 156.445 ;
        RECT 62.930 156.295 63.280 156.865 ;
        RECT 61.090 155.625 61.370 156.105 ;
        RECT 61.540 155.885 61.800 156.275 ;
        RECT 61.975 155.625 62.230 156.105 ;
        RECT 62.400 155.885 62.695 156.275 ;
        RECT 63.450 156.125 63.620 157.035 ;
        RECT 63.790 157.085 65.000 158.175 ;
        RECT 65.180 157.195 65.510 158.005 ;
        RECT 65.680 157.375 65.920 158.175 ;
        RECT 63.790 156.545 64.310 157.085 ;
        RECT 65.180 157.025 65.895 157.195 ;
        RECT 64.480 156.375 65.000 156.915 ;
        RECT 65.175 156.615 65.555 156.855 ;
        RECT 65.725 156.785 65.895 157.025 ;
        RECT 66.100 157.155 66.270 158.005 ;
        RECT 66.440 157.375 66.770 158.175 ;
        RECT 66.940 157.155 67.110 158.005 ;
        RECT 66.100 156.985 67.110 157.155 ;
        RECT 67.280 157.025 67.610 158.175 ;
        RECT 68.020 157.245 68.190 158.005 ;
        RECT 68.405 157.415 68.735 158.175 ;
        RECT 68.020 157.075 68.735 157.245 ;
        RECT 68.905 157.100 69.160 158.005 ;
        RECT 65.725 156.615 66.225 156.785 ;
        RECT 65.725 156.445 65.895 156.615 ;
        RECT 66.615 156.445 67.110 156.985 ;
        RECT 67.930 156.525 68.285 156.895 ;
        RECT 68.565 156.865 68.735 157.075 ;
        RECT 68.565 156.535 68.820 156.865 ;
        RECT 62.875 155.625 63.150 156.105 ;
        RECT 63.320 155.795 63.620 156.125 ;
        RECT 63.790 155.625 65.000 156.375 ;
        RECT 65.260 156.275 65.895 156.445 ;
        RECT 66.100 156.275 67.110 156.445 ;
        RECT 65.260 155.795 65.430 156.275 ;
        RECT 65.610 155.625 65.850 156.105 ;
        RECT 66.100 155.795 66.270 156.275 ;
        RECT 66.440 155.625 66.770 156.105 ;
        RECT 66.940 155.795 67.110 156.275 ;
        RECT 67.280 155.625 67.610 156.425 ;
        RECT 68.565 156.345 68.735 156.535 ;
        RECT 68.990 156.370 69.160 157.100 ;
        RECT 69.335 157.025 69.595 158.175 ;
        RECT 69.770 157.035 70.110 158.005 ;
        RECT 70.280 157.035 70.450 158.175 ;
        RECT 70.720 157.375 70.970 158.175 ;
        RECT 71.615 157.205 71.945 158.005 ;
        RECT 72.245 157.375 72.575 158.175 ;
        RECT 72.745 157.205 73.075 158.005 ;
        RECT 73.825 157.835 74.080 157.865 ;
        RECT 73.740 157.665 74.080 157.835 ;
        RECT 70.640 157.035 73.075 157.205 ;
        RECT 73.825 157.195 74.080 157.665 ;
        RECT 74.260 157.375 74.545 158.175 ;
        RECT 74.725 157.455 75.055 157.965 ;
        RECT 68.020 156.175 68.735 156.345 ;
        RECT 68.020 155.795 68.190 156.175 ;
        RECT 68.405 155.625 68.735 156.005 ;
        RECT 68.905 155.795 69.160 156.370 ;
        RECT 69.335 155.625 69.595 156.465 ;
        RECT 69.770 156.425 69.945 157.035 ;
        RECT 70.640 156.785 70.810 157.035 ;
        RECT 70.115 156.615 70.810 156.785 ;
        RECT 70.985 156.615 71.405 156.815 ;
        RECT 71.575 156.615 71.905 156.815 ;
        RECT 72.075 156.615 72.405 156.815 ;
        RECT 69.770 155.795 70.110 156.425 ;
        RECT 70.280 155.625 70.530 156.425 ;
        RECT 70.720 156.275 71.945 156.445 ;
        RECT 70.720 155.795 71.050 156.275 ;
        RECT 71.220 155.625 71.445 156.085 ;
        RECT 71.615 155.795 71.945 156.275 ;
        RECT 72.575 156.405 72.745 157.035 ;
        RECT 72.930 156.615 73.280 156.865 ;
        RECT 72.575 155.795 73.075 156.405 ;
        RECT 73.825 156.335 74.005 157.195 ;
        RECT 74.725 156.865 74.975 157.455 ;
        RECT 75.325 157.305 75.495 157.915 ;
        RECT 75.665 157.485 75.995 158.175 ;
        RECT 76.225 157.625 76.465 157.915 ;
        RECT 76.665 157.795 77.085 158.175 ;
        RECT 77.265 157.705 77.895 157.955 ;
        RECT 78.365 157.795 78.695 158.175 ;
        RECT 77.265 157.625 77.435 157.705 ;
        RECT 78.865 157.625 79.035 157.915 ;
        RECT 79.215 157.795 79.595 158.175 ;
        RECT 79.835 157.790 80.665 157.960 ;
        RECT 76.225 157.455 77.435 157.625 ;
        RECT 74.175 156.535 74.975 156.865 ;
        RECT 73.825 155.805 74.080 156.335 ;
        RECT 74.260 155.625 74.545 156.085 ;
        RECT 74.725 155.885 74.975 156.535 ;
        RECT 75.175 157.285 75.495 157.305 ;
        RECT 75.175 157.115 77.095 157.285 ;
        RECT 75.175 156.220 75.365 157.115 ;
        RECT 77.265 156.945 77.435 157.455 ;
        RECT 77.605 157.195 78.125 157.505 ;
        RECT 75.535 156.775 77.435 156.945 ;
        RECT 75.535 156.715 75.865 156.775 ;
        RECT 76.015 156.545 76.345 156.605 ;
        RECT 75.685 156.275 76.345 156.545 ;
        RECT 75.175 155.890 75.495 156.220 ;
        RECT 75.675 155.625 76.335 156.105 ;
        RECT 76.535 156.015 76.705 156.775 ;
        RECT 77.605 156.605 77.785 157.015 ;
        RECT 76.875 156.435 77.205 156.555 ;
        RECT 77.955 156.435 78.125 157.195 ;
        RECT 76.875 156.265 78.125 156.435 ;
        RECT 78.295 157.375 79.665 157.625 ;
        RECT 78.295 156.605 78.485 157.375 ;
        RECT 79.415 157.115 79.665 157.375 ;
        RECT 78.655 156.945 78.905 157.105 ;
        RECT 79.835 156.945 80.005 157.790 ;
        RECT 80.900 157.505 81.070 158.005 ;
        RECT 81.240 157.675 81.570 158.175 ;
        RECT 80.175 157.115 80.675 157.495 ;
        RECT 80.900 157.335 81.595 157.505 ;
        RECT 78.655 156.775 80.005 156.945 ;
        RECT 79.585 156.735 80.005 156.775 ;
        RECT 78.295 156.265 78.715 156.605 ;
        RECT 79.005 156.275 79.415 156.605 ;
        RECT 76.535 155.845 77.385 156.015 ;
        RECT 77.945 155.625 78.265 156.085 ;
        RECT 78.465 155.835 78.715 156.265 ;
        RECT 79.005 155.625 79.415 156.065 ;
        RECT 79.585 156.005 79.755 156.735 ;
        RECT 79.925 156.185 80.275 156.555 ;
        RECT 80.455 156.245 80.675 157.115 ;
        RECT 80.845 156.545 81.255 157.165 ;
        RECT 81.425 156.365 81.595 157.335 ;
        RECT 80.900 156.175 81.595 156.365 ;
        RECT 79.585 155.805 80.600 156.005 ;
        RECT 80.900 155.845 81.070 156.175 ;
        RECT 81.240 155.625 81.570 156.005 ;
        RECT 81.785 155.885 82.010 158.005 ;
        RECT 82.180 157.675 82.510 158.175 ;
        RECT 82.680 157.505 82.850 158.005 ;
        RECT 82.185 157.335 82.850 157.505 ;
        RECT 82.185 156.345 82.415 157.335 ;
        RECT 82.585 156.515 82.935 157.165 ;
        RECT 83.570 157.085 86.160 158.175 ;
        RECT 83.570 156.565 84.780 157.085 ;
        RECT 86.330 157.010 86.620 158.175 ;
        RECT 87.310 157.340 87.565 158.175 ;
        RECT 87.735 157.170 87.995 157.975 ;
        RECT 88.165 157.340 88.425 158.175 ;
        RECT 88.595 157.170 88.850 157.975 ;
        RECT 87.250 157.000 88.850 157.170 ;
        RECT 89.090 157.035 89.430 158.005 ;
        RECT 89.600 157.035 89.770 158.175 ;
        RECT 90.040 157.375 90.290 158.175 ;
        RECT 90.935 157.205 91.265 158.005 ;
        RECT 91.565 157.375 91.895 158.175 ;
        RECT 92.065 157.205 92.395 158.005 ;
        RECT 89.960 157.035 92.395 157.205 ;
        RECT 93.435 157.205 93.765 158.005 ;
        RECT 93.935 157.375 94.265 158.175 ;
        RECT 94.565 157.205 94.895 158.005 ;
        RECT 95.540 157.375 95.790 158.175 ;
        RECT 93.435 157.035 95.870 157.205 ;
        RECT 96.060 157.035 96.230 158.175 ;
        RECT 96.400 157.035 96.740 158.005 ;
        RECT 84.950 156.395 86.160 156.915 ;
        RECT 82.185 156.175 82.850 156.345 ;
        RECT 82.180 155.625 82.510 156.005 ;
        RECT 82.680 155.885 82.850 156.175 ;
        RECT 83.570 155.625 86.160 156.395 ;
        RECT 87.250 156.435 87.530 157.000 ;
        RECT 87.700 156.605 88.920 156.830 ;
        RECT 86.330 155.625 86.620 156.350 ;
        RECT 87.250 156.265 87.980 156.435 ;
        RECT 87.255 155.625 87.585 156.095 ;
        RECT 87.755 155.820 87.980 156.265 ;
        RECT 89.090 156.425 89.265 157.035 ;
        RECT 89.960 156.785 90.130 157.035 ;
        RECT 89.435 156.615 90.130 156.785 ;
        RECT 90.305 156.615 90.725 156.815 ;
        RECT 90.895 156.615 91.225 156.815 ;
        RECT 91.395 156.615 91.725 156.815 ;
        RECT 88.150 155.625 88.445 156.150 ;
        RECT 89.090 155.795 89.430 156.425 ;
        RECT 89.600 155.625 89.850 156.425 ;
        RECT 90.040 156.275 91.265 156.445 ;
        RECT 90.040 155.795 90.370 156.275 ;
        RECT 90.540 155.625 90.765 156.085 ;
        RECT 90.935 155.795 91.265 156.275 ;
        RECT 91.895 156.405 92.065 157.035 ;
        RECT 92.250 156.615 92.600 156.865 ;
        RECT 93.230 156.615 93.580 156.865 ;
        RECT 93.765 156.405 93.935 157.035 ;
        RECT 94.105 156.615 94.435 156.815 ;
        RECT 94.605 156.615 94.935 156.815 ;
        RECT 95.105 156.615 95.525 156.815 ;
        RECT 95.700 156.785 95.870 157.035 ;
        RECT 95.700 156.615 96.395 156.785 ;
        RECT 91.895 155.795 92.395 156.405 ;
        RECT 93.435 155.795 93.935 156.405 ;
        RECT 94.565 156.275 95.790 156.445 ;
        RECT 96.565 156.425 96.740 157.035 ;
        RECT 94.565 155.795 94.895 156.275 ;
        RECT 95.065 155.625 95.290 156.085 ;
        RECT 95.460 155.795 95.790 156.275 ;
        RECT 95.980 155.625 96.230 156.425 ;
        RECT 96.400 155.795 96.740 156.425 ;
        RECT 96.910 157.035 97.250 158.005 ;
        RECT 97.420 157.035 97.590 158.175 ;
        RECT 97.860 157.375 98.110 158.175 ;
        RECT 98.755 157.205 99.085 158.005 ;
        RECT 99.385 157.375 99.715 158.175 ;
        RECT 99.885 157.205 100.215 158.005 ;
        RECT 97.780 157.035 100.215 157.205 ;
        RECT 101.050 157.085 102.720 158.175 ;
        RECT 96.910 156.475 97.085 157.035 ;
        RECT 97.780 156.785 97.950 157.035 ;
        RECT 97.255 156.615 97.950 156.785 ;
        RECT 98.125 156.615 98.545 156.815 ;
        RECT 98.715 156.615 99.045 156.815 ;
        RECT 99.215 156.615 99.545 156.815 ;
        RECT 96.910 156.425 97.140 156.475 ;
        RECT 96.910 155.795 97.250 156.425 ;
        RECT 97.420 155.625 97.670 156.425 ;
        RECT 97.860 156.275 99.085 156.445 ;
        RECT 97.860 155.795 98.190 156.275 ;
        RECT 98.360 155.625 98.585 156.085 ;
        RECT 98.755 155.795 99.085 156.275 ;
        RECT 99.715 156.405 99.885 157.035 ;
        RECT 100.070 156.615 100.420 156.865 ;
        RECT 101.050 156.565 101.800 157.085 ;
        RECT 103.040 157.025 103.370 158.175 ;
        RECT 103.540 157.155 103.710 158.005 ;
        RECT 103.880 157.375 104.210 158.175 ;
        RECT 104.380 157.155 104.550 158.005 ;
        RECT 104.730 157.375 104.970 158.175 ;
        RECT 105.140 157.195 105.470 158.005 ;
        RECT 105.655 157.740 111.000 158.175 ;
        RECT 103.540 156.985 104.550 157.155 ;
        RECT 104.755 157.025 105.470 157.195 ;
        RECT 99.715 155.795 100.215 156.405 ;
        RECT 101.970 156.395 102.720 156.915 ;
        RECT 103.540 156.445 104.035 156.985 ;
        RECT 104.755 156.785 104.925 157.025 ;
        RECT 104.425 156.615 104.925 156.785 ;
        RECT 105.095 156.615 105.475 156.855 ;
        RECT 104.755 156.445 104.925 156.615 ;
        RECT 107.245 156.490 107.595 157.740 ;
        RECT 111.170 157.085 112.380 158.175 ;
        RECT 101.050 155.625 102.720 156.395 ;
        RECT 103.040 155.625 103.370 156.425 ;
        RECT 103.540 156.275 104.550 156.445 ;
        RECT 104.755 156.275 105.390 156.445 ;
        RECT 103.540 155.795 103.710 156.275 ;
        RECT 103.880 155.625 104.210 156.105 ;
        RECT 104.380 155.795 104.550 156.275 ;
        RECT 104.800 155.625 105.040 156.105 ;
        RECT 105.220 155.795 105.390 156.275 ;
        RECT 109.075 156.170 109.415 157.000 ;
        RECT 111.170 156.545 111.690 157.085 ;
        RECT 111.860 156.375 112.380 156.915 ;
        RECT 105.655 155.625 111.000 156.170 ;
        RECT 111.170 155.625 112.380 156.375 ;
        RECT 18.165 155.455 112.465 155.625 ;
        RECT 18.250 154.705 19.460 155.455 ;
        RECT 18.250 154.165 18.770 154.705 ;
        RECT 20.610 154.635 20.820 155.455 ;
        RECT 20.990 154.655 21.320 155.285 ;
        RECT 18.940 153.995 19.460 154.535 ;
        RECT 20.990 154.055 21.240 154.655 ;
        RECT 21.490 154.635 21.720 155.455 ;
        RECT 21.930 154.730 22.220 155.455 ;
        RECT 22.890 154.635 23.120 155.455 ;
        RECT 23.290 154.655 23.620 155.285 ;
        RECT 21.410 154.215 21.740 154.465 ;
        RECT 22.870 154.215 23.200 154.465 ;
        RECT 18.250 152.905 19.460 153.995 ;
        RECT 20.610 152.905 20.820 154.045 ;
        RECT 20.990 153.075 21.320 154.055 ;
        RECT 21.490 152.905 21.720 154.045 ;
        RECT 21.930 152.905 22.220 154.070 ;
        RECT 23.370 154.055 23.620 154.655 ;
        RECT 23.790 154.635 24.000 155.455 ;
        RECT 24.345 154.825 24.630 155.285 ;
        RECT 24.800 154.995 25.070 155.455 ;
        RECT 24.345 154.655 25.300 154.825 ;
        RECT 22.890 152.905 23.120 154.045 ;
        RECT 23.290 153.075 23.620 154.055 ;
        RECT 23.790 152.905 24.000 154.045 ;
        RECT 24.230 153.925 24.920 154.485 ;
        RECT 25.090 153.755 25.300 154.655 ;
        RECT 24.345 153.535 25.300 153.755 ;
        RECT 25.470 154.485 25.870 155.285 ;
        RECT 26.060 154.825 26.340 155.285 ;
        RECT 26.860 154.995 27.185 155.455 ;
        RECT 26.060 154.655 27.185 154.825 ;
        RECT 27.355 154.715 27.740 155.285 ;
        RECT 26.735 154.545 27.185 154.655 ;
        RECT 25.470 153.925 26.565 154.485 ;
        RECT 26.735 154.215 27.290 154.545 ;
        RECT 24.345 153.075 24.630 153.535 ;
        RECT 24.800 152.905 25.070 153.365 ;
        RECT 25.470 153.075 25.870 153.925 ;
        RECT 26.735 153.755 27.185 154.215 ;
        RECT 27.460 154.045 27.740 154.715 ;
        RECT 28.185 154.645 28.430 155.250 ;
        RECT 28.650 154.920 29.160 155.455 ;
        RECT 26.060 153.535 27.185 153.755 ;
        RECT 26.060 153.075 26.340 153.535 ;
        RECT 26.860 152.905 27.185 153.365 ;
        RECT 27.355 153.075 27.740 154.045 ;
        RECT 27.910 154.475 29.140 154.645 ;
        RECT 27.910 153.665 28.250 154.475 ;
        RECT 28.420 153.910 29.170 154.100 ;
        RECT 27.910 153.255 28.425 153.665 ;
        RECT 28.660 152.905 28.830 153.665 ;
        RECT 29.000 153.245 29.170 153.910 ;
        RECT 29.340 153.925 29.530 155.285 ;
        RECT 29.700 154.775 29.975 155.285 ;
        RECT 30.165 154.920 30.695 155.285 ;
        RECT 31.120 155.055 31.450 155.455 ;
        RECT 30.520 154.885 30.695 154.920 ;
        RECT 29.700 154.605 29.980 154.775 ;
        RECT 29.700 154.125 29.975 154.605 ;
        RECT 30.180 153.925 30.350 154.725 ;
        RECT 29.340 153.755 30.350 153.925 ;
        RECT 30.520 154.715 31.450 154.885 ;
        RECT 31.620 154.715 31.875 155.285 ;
        RECT 32.140 154.975 32.440 155.455 ;
        RECT 32.610 154.805 32.870 155.260 ;
        RECT 33.040 154.975 33.300 155.455 ;
        RECT 33.480 154.805 33.740 155.260 ;
        RECT 33.910 154.975 34.160 155.455 ;
        RECT 34.340 154.805 34.600 155.260 ;
        RECT 34.770 154.975 35.020 155.455 ;
        RECT 35.200 154.805 35.460 155.260 ;
        RECT 35.630 154.975 35.875 155.455 ;
        RECT 36.045 154.805 36.320 155.260 ;
        RECT 36.490 154.975 36.735 155.455 ;
        RECT 36.905 154.805 37.165 155.260 ;
        RECT 37.335 154.975 37.595 155.455 ;
        RECT 37.765 154.805 38.025 155.260 ;
        RECT 38.195 154.975 38.455 155.455 ;
        RECT 38.625 154.805 38.885 155.260 ;
        RECT 39.055 154.895 39.315 155.455 ;
        RECT 30.520 153.585 30.690 154.715 ;
        RECT 31.280 154.545 31.450 154.715 ;
        RECT 29.565 153.415 30.690 153.585 ;
        RECT 30.860 154.215 31.055 154.545 ;
        RECT 31.280 154.215 31.535 154.545 ;
        RECT 30.860 153.245 31.030 154.215 ;
        RECT 31.705 154.045 31.875 154.715 ;
        RECT 29.000 153.075 31.030 153.245 ;
        RECT 31.200 152.905 31.370 154.045 ;
        RECT 31.540 153.075 31.875 154.045 ;
        RECT 32.140 154.635 38.885 154.805 ;
        RECT 32.140 154.045 33.305 154.635 ;
        RECT 39.485 154.465 39.735 155.275 ;
        RECT 39.915 154.930 40.175 155.455 ;
        RECT 40.345 154.465 40.595 155.275 ;
        RECT 40.775 154.945 41.080 155.455 ;
        RECT 41.340 154.905 41.510 155.285 ;
        RECT 41.690 155.075 42.020 155.455 ;
        RECT 33.475 154.215 40.595 154.465 ;
        RECT 40.765 154.215 41.080 154.775 ;
        RECT 41.340 154.735 42.005 154.905 ;
        RECT 42.200 154.780 42.460 155.285 ;
        RECT 32.140 153.820 38.885 154.045 ;
        RECT 32.140 152.905 32.410 153.650 ;
        RECT 32.580 153.080 32.870 153.820 ;
        RECT 33.480 153.805 38.885 153.820 ;
        RECT 33.040 152.910 33.295 153.635 ;
        RECT 33.480 153.080 33.740 153.805 ;
        RECT 33.910 152.910 34.155 153.635 ;
        RECT 34.340 153.080 34.600 153.805 ;
        RECT 34.770 152.910 35.015 153.635 ;
        RECT 35.200 153.080 35.460 153.805 ;
        RECT 35.630 152.910 35.875 153.635 ;
        RECT 36.045 153.080 36.305 153.805 ;
        RECT 36.475 152.910 36.735 153.635 ;
        RECT 36.905 153.080 37.165 153.805 ;
        RECT 37.335 152.910 37.595 153.635 ;
        RECT 37.765 153.080 38.025 153.805 ;
        RECT 38.195 152.910 38.455 153.635 ;
        RECT 38.625 153.080 38.885 153.805 ;
        RECT 39.055 152.910 39.315 153.705 ;
        RECT 39.485 153.080 39.735 154.215 ;
        RECT 33.040 152.905 39.315 152.910 ;
        RECT 39.915 152.905 40.175 153.715 ;
        RECT 40.350 153.075 40.595 154.215 ;
        RECT 41.270 154.185 41.600 154.555 ;
        RECT 41.835 154.480 42.005 154.735 ;
        RECT 41.835 154.150 42.120 154.480 ;
        RECT 41.835 154.005 42.005 154.150 ;
        RECT 41.340 153.835 42.005 154.005 ;
        RECT 42.290 153.980 42.460 154.780 ;
        RECT 42.630 154.705 43.840 155.455 ;
        RECT 40.775 152.905 41.070 153.715 ;
        RECT 41.340 153.075 41.510 153.835 ;
        RECT 41.690 152.905 42.020 153.665 ;
        RECT 42.190 153.075 42.460 153.980 ;
        RECT 42.630 153.995 43.150 154.535 ;
        RECT 43.320 154.165 43.840 154.705 ;
        RECT 44.215 154.675 44.715 155.285 ;
        RECT 44.010 154.215 44.360 154.465 ;
        RECT 44.545 154.045 44.715 154.675 ;
        RECT 45.345 154.805 45.675 155.285 ;
        RECT 45.845 154.995 46.070 155.455 ;
        RECT 46.240 154.805 46.570 155.285 ;
        RECT 45.345 154.635 46.570 154.805 ;
        RECT 46.760 154.655 47.010 155.455 ;
        RECT 47.180 154.655 47.520 155.285 ;
        RECT 47.690 154.730 47.980 155.455 ;
        RECT 48.150 154.685 49.820 155.455 ;
        RECT 49.995 154.910 55.340 155.455 ;
        RECT 44.885 154.265 45.215 154.465 ;
        RECT 45.385 154.265 45.715 154.465 ;
        RECT 45.885 154.265 46.305 154.465 ;
        RECT 46.480 154.295 47.175 154.465 ;
        RECT 46.480 154.045 46.650 154.295 ;
        RECT 47.345 154.045 47.520 154.655 ;
        RECT 42.630 152.905 43.840 153.995 ;
        RECT 44.215 153.875 46.650 154.045 ;
        RECT 44.215 153.075 44.545 153.875 ;
        RECT 44.715 152.905 45.045 153.705 ;
        RECT 45.345 153.075 45.675 153.875 ;
        RECT 46.320 152.905 46.570 153.705 ;
        RECT 46.840 152.905 47.010 154.045 ;
        RECT 47.180 153.075 47.520 154.045 ;
        RECT 47.690 152.905 47.980 154.070 ;
        RECT 48.150 153.995 48.900 154.515 ;
        RECT 49.070 154.165 49.820 154.685 ;
        RECT 48.150 152.905 49.820 153.995 ;
        RECT 51.585 153.340 51.935 154.590 ;
        RECT 53.415 154.080 53.755 154.910 ;
        RECT 55.885 154.745 56.140 155.275 ;
        RECT 56.320 154.995 56.605 155.455 ;
        RECT 55.885 153.885 56.065 154.745 ;
        RECT 56.785 154.545 57.035 155.195 ;
        RECT 56.235 154.215 57.035 154.545 ;
        RECT 55.885 153.415 56.140 153.885 ;
        RECT 49.995 152.905 55.340 153.340 ;
        RECT 55.800 153.245 56.140 153.415 ;
        RECT 55.885 153.215 56.140 153.245 ;
        RECT 56.320 152.905 56.605 153.705 ;
        RECT 56.785 153.625 57.035 154.215 ;
        RECT 57.235 154.860 57.555 155.190 ;
        RECT 57.735 154.975 58.395 155.455 ;
        RECT 58.595 155.065 59.445 155.235 ;
        RECT 57.235 153.965 57.425 154.860 ;
        RECT 57.745 154.535 58.405 154.805 ;
        RECT 58.075 154.475 58.405 154.535 ;
        RECT 57.595 154.305 57.925 154.365 ;
        RECT 58.595 154.305 58.765 155.065 ;
        RECT 60.005 154.995 60.325 155.455 ;
        RECT 60.525 154.815 60.775 155.245 ;
        RECT 61.065 155.015 61.475 155.455 ;
        RECT 61.645 155.075 62.660 155.275 ;
        RECT 58.935 154.645 60.185 154.815 ;
        RECT 58.935 154.525 59.265 154.645 ;
        RECT 57.595 154.135 59.495 154.305 ;
        RECT 57.235 153.795 59.155 153.965 ;
        RECT 57.235 153.775 57.555 153.795 ;
        RECT 56.785 153.115 57.115 153.625 ;
        RECT 57.385 153.165 57.555 153.775 ;
        RECT 59.325 153.625 59.495 154.135 ;
        RECT 59.665 154.065 59.845 154.475 ;
        RECT 60.015 153.885 60.185 154.645 ;
        RECT 57.725 152.905 58.055 153.595 ;
        RECT 58.285 153.455 59.495 153.625 ;
        RECT 59.665 153.575 60.185 153.885 ;
        RECT 60.355 154.475 60.775 154.815 ;
        RECT 61.065 154.475 61.475 154.805 ;
        RECT 60.355 153.705 60.545 154.475 ;
        RECT 61.645 154.345 61.815 155.075 ;
        RECT 62.960 154.905 63.130 155.235 ;
        RECT 63.300 155.075 63.630 155.455 ;
        RECT 61.985 154.525 62.335 154.895 ;
        RECT 61.645 154.305 62.065 154.345 ;
        RECT 60.715 154.135 62.065 154.305 ;
        RECT 60.715 153.975 60.965 154.135 ;
        RECT 61.475 153.705 61.725 153.965 ;
        RECT 60.355 153.455 61.725 153.705 ;
        RECT 58.285 153.165 58.525 153.455 ;
        RECT 59.325 153.375 59.495 153.455 ;
        RECT 58.725 152.905 59.145 153.285 ;
        RECT 59.325 153.125 59.955 153.375 ;
        RECT 60.425 152.905 60.755 153.285 ;
        RECT 60.925 153.165 61.095 153.455 ;
        RECT 61.895 153.290 62.065 154.135 ;
        RECT 62.515 153.965 62.735 154.835 ;
        RECT 62.960 154.715 63.655 154.905 ;
        RECT 62.235 153.585 62.735 153.965 ;
        RECT 62.905 153.915 63.315 154.535 ;
        RECT 63.485 153.745 63.655 154.715 ;
        RECT 62.960 153.575 63.655 153.745 ;
        RECT 61.275 152.905 61.655 153.285 ;
        RECT 61.895 153.120 62.725 153.290 ;
        RECT 62.960 153.075 63.130 153.575 ;
        RECT 63.300 152.905 63.630 153.405 ;
        RECT 63.845 153.075 64.070 155.195 ;
        RECT 64.240 155.075 64.570 155.455 ;
        RECT 64.740 154.905 64.910 155.195 ;
        RECT 64.245 154.735 64.910 154.905 ;
        RECT 66.100 154.925 66.430 155.285 ;
        RECT 66.600 155.095 66.930 155.455 ;
        RECT 67.130 154.925 67.460 155.285 ;
        RECT 64.245 153.745 64.475 154.735 ;
        RECT 66.100 154.715 67.460 154.925 ;
        RECT 67.970 154.695 68.680 155.285 ;
        RECT 68.940 154.905 69.110 155.285 ;
        RECT 69.325 155.075 69.655 155.455 ;
        RECT 68.940 154.735 69.655 154.905 ;
        RECT 64.645 153.915 64.995 154.565 ;
        RECT 66.090 154.215 66.400 154.545 ;
        RECT 66.610 154.215 66.985 154.545 ;
        RECT 67.305 154.215 67.800 154.545 ;
        RECT 64.245 153.575 64.910 153.745 ;
        RECT 64.240 152.905 64.570 153.405 ;
        RECT 64.740 153.075 64.910 153.575 ;
        RECT 66.100 152.905 66.430 153.965 ;
        RECT 66.610 153.290 66.780 154.215 ;
        RECT 66.950 153.725 67.280 153.945 ;
        RECT 67.475 153.925 67.800 154.215 ;
        RECT 67.975 153.925 68.305 154.465 ;
        RECT 68.475 153.725 68.680 154.695 ;
        RECT 68.850 154.185 69.205 154.555 ;
        RECT 69.485 154.545 69.655 154.735 ;
        RECT 69.825 154.710 70.080 155.285 ;
        RECT 69.485 154.215 69.740 154.545 ;
        RECT 69.485 154.005 69.655 154.215 ;
        RECT 66.950 153.495 68.680 153.725 ;
        RECT 66.950 153.095 67.280 153.495 ;
        RECT 67.450 152.905 67.780 153.265 ;
        RECT 67.980 153.075 68.680 153.495 ;
        RECT 68.940 153.835 69.655 154.005 ;
        RECT 69.910 153.980 70.080 154.710 ;
        RECT 70.255 154.615 70.515 155.455 ;
        RECT 70.690 154.685 73.280 155.455 ;
        RECT 73.450 154.730 73.740 155.455 ;
        RECT 74.370 154.955 74.670 155.285 ;
        RECT 74.840 154.975 75.115 155.455 ;
        RECT 68.940 153.075 69.110 153.835 ;
        RECT 69.325 152.905 69.655 153.665 ;
        RECT 69.825 153.075 70.080 153.980 ;
        RECT 70.255 152.905 70.515 154.055 ;
        RECT 70.690 153.995 71.900 154.515 ;
        RECT 72.070 154.165 73.280 154.685 ;
        RECT 70.690 152.905 73.280 153.995 ;
        RECT 73.450 152.905 73.740 154.070 ;
        RECT 74.370 154.045 74.540 154.955 ;
        RECT 75.295 154.805 75.590 155.195 ;
        RECT 75.760 154.975 76.015 155.455 ;
        RECT 76.190 154.805 76.450 155.195 ;
        RECT 76.620 154.975 76.900 155.455 ;
        RECT 74.710 154.215 75.060 154.785 ;
        RECT 75.295 154.635 76.945 154.805 ;
        RECT 78.110 154.635 78.320 155.455 ;
        RECT 78.490 154.655 78.820 155.285 ;
        RECT 75.230 154.295 76.370 154.465 ;
        RECT 75.230 154.045 75.400 154.295 ;
        RECT 76.540 154.125 76.945 154.635 ;
        RECT 74.370 153.875 75.400 154.045 ;
        RECT 76.190 153.955 76.945 154.125 ;
        RECT 78.490 154.055 78.740 154.655 ;
        RECT 78.990 154.635 79.220 155.455 ;
        RECT 79.890 154.685 82.480 155.455 ;
        RECT 82.655 154.910 88.000 155.455 ;
        RECT 78.910 154.215 79.240 154.465 ;
        RECT 74.370 153.075 74.680 153.875 ;
        RECT 76.190 153.705 76.450 153.955 ;
        RECT 74.850 152.905 75.160 153.705 ;
        RECT 75.330 153.535 76.450 153.705 ;
        RECT 75.330 153.075 75.590 153.535 ;
        RECT 75.760 152.905 76.015 153.365 ;
        RECT 76.190 153.075 76.450 153.535 ;
        RECT 76.620 152.905 76.905 153.775 ;
        RECT 78.110 152.905 78.320 154.045 ;
        RECT 78.490 153.075 78.820 154.055 ;
        RECT 78.990 152.905 79.220 154.045 ;
        RECT 79.890 153.995 81.100 154.515 ;
        RECT 81.270 154.165 82.480 154.685 ;
        RECT 79.890 152.905 82.480 153.995 ;
        RECT 84.245 153.340 84.595 154.590 ;
        RECT 86.075 154.080 86.415 154.910 ;
        RECT 88.170 154.655 88.510 155.285 ;
        RECT 88.680 154.655 88.930 155.455 ;
        RECT 89.120 154.805 89.450 155.285 ;
        RECT 89.620 154.995 89.845 155.455 ;
        RECT 90.015 154.805 90.345 155.285 ;
        RECT 88.170 154.045 88.345 154.655 ;
        RECT 89.120 154.635 90.345 154.805 ;
        RECT 90.975 154.675 91.475 155.285 ;
        RECT 88.515 154.295 89.210 154.465 ;
        RECT 89.040 154.045 89.210 154.295 ;
        RECT 89.385 154.265 89.805 154.465 ;
        RECT 89.975 154.265 90.305 154.465 ;
        RECT 90.475 154.265 90.805 154.465 ;
        RECT 90.975 154.045 91.145 154.675 ;
        RECT 92.310 154.655 92.650 155.285 ;
        RECT 92.820 154.655 93.070 155.455 ;
        RECT 93.260 154.805 93.590 155.285 ;
        RECT 93.760 154.995 93.985 155.455 ;
        RECT 94.155 154.805 94.485 155.285 ;
        RECT 91.330 154.215 91.680 154.465 ;
        RECT 92.310 154.045 92.485 154.655 ;
        RECT 93.260 154.635 94.485 154.805 ;
        RECT 95.115 154.675 95.615 155.285 ;
        RECT 96.450 154.685 99.040 155.455 ;
        RECT 99.210 154.730 99.500 155.455 ;
        RECT 99.670 154.685 102.260 155.455 ;
        RECT 92.655 154.295 93.350 154.465 ;
        RECT 93.180 154.045 93.350 154.295 ;
        RECT 93.525 154.265 93.945 154.465 ;
        RECT 94.115 154.265 94.445 154.465 ;
        RECT 94.615 154.265 94.945 154.465 ;
        RECT 95.115 154.045 95.285 154.675 ;
        RECT 95.470 154.215 95.820 154.465 ;
        RECT 82.655 152.905 88.000 153.340 ;
        RECT 88.170 153.075 88.510 154.045 ;
        RECT 88.680 152.905 88.850 154.045 ;
        RECT 89.040 153.875 91.475 154.045 ;
        RECT 89.120 152.905 89.370 153.705 ;
        RECT 90.015 153.075 90.345 153.875 ;
        RECT 90.645 152.905 90.975 153.705 ;
        RECT 91.145 153.075 91.475 153.875 ;
        RECT 92.310 153.075 92.650 154.045 ;
        RECT 92.820 152.905 92.990 154.045 ;
        RECT 93.180 153.875 95.615 154.045 ;
        RECT 93.260 152.905 93.510 153.705 ;
        RECT 94.155 153.075 94.485 153.875 ;
        RECT 94.785 152.905 95.115 153.705 ;
        RECT 95.285 153.075 95.615 153.875 ;
        RECT 96.450 153.995 97.660 154.515 ;
        RECT 97.830 154.165 99.040 154.685 ;
        RECT 96.450 152.905 99.040 153.995 ;
        RECT 99.210 152.905 99.500 154.070 ;
        RECT 99.670 153.995 100.880 154.515 ;
        RECT 101.050 154.165 102.260 154.685 ;
        RECT 102.520 154.805 102.690 155.285 ;
        RECT 102.870 154.975 103.110 155.455 ;
        RECT 103.360 154.805 103.530 155.285 ;
        RECT 103.700 154.975 104.030 155.455 ;
        RECT 104.200 154.805 104.370 155.285 ;
        RECT 102.520 154.635 103.155 154.805 ;
        RECT 103.360 154.635 104.370 154.805 ;
        RECT 104.540 154.655 104.870 155.455 ;
        RECT 105.740 154.905 105.910 155.285 ;
        RECT 106.090 155.075 106.420 155.455 ;
        RECT 105.740 154.735 106.405 154.905 ;
        RECT 106.600 154.780 106.860 155.285 ;
        RECT 102.985 154.465 103.155 154.635 ;
        RECT 103.870 154.605 104.370 154.635 ;
        RECT 102.435 154.225 102.815 154.465 ;
        RECT 102.985 154.295 103.485 154.465 ;
        RECT 102.985 154.055 103.155 154.295 ;
        RECT 103.875 154.095 104.370 154.605 ;
        RECT 105.670 154.185 106.000 154.555 ;
        RECT 106.235 154.480 106.405 154.735 ;
        RECT 99.670 152.905 102.260 153.995 ;
        RECT 102.440 153.885 103.155 154.055 ;
        RECT 103.360 153.925 104.370 154.095 ;
        RECT 106.235 154.150 106.520 154.480 ;
        RECT 102.440 153.075 102.770 153.885 ;
        RECT 102.940 152.905 103.180 153.705 ;
        RECT 103.360 153.075 103.530 153.925 ;
        RECT 103.700 152.905 104.030 153.705 ;
        RECT 104.200 153.075 104.370 153.925 ;
        RECT 104.540 152.905 104.870 154.055 ;
        RECT 106.235 154.005 106.405 154.150 ;
        RECT 105.740 153.835 106.405 154.005 ;
        RECT 106.690 153.980 106.860 154.780 ;
        RECT 107.490 154.685 111.000 155.455 ;
        RECT 111.170 154.705 112.380 155.455 ;
        RECT 105.740 153.075 105.910 153.835 ;
        RECT 106.090 152.905 106.420 153.665 ;
        RECT 106.590 153.075 106.860 153.980 ;
        RECT 107.490 153.995 109.180 154.515 ;
        RECT 109.350 154.165 111.000 154.685 ;
        RECT 111.170 153.995 111.690 154.535 ;
        RECT 111.860 154.165 112.380 154.705 ;
        RECT 107.490 152.905 111.000 153.995 ;
        RECT 111.170 152.905 112.380 153.995 ;
        RECT 18.165 152.735 112.465 152.905 ;
        RECT 18.250 151.645 19.460 152.735 ;
        RECT 18.250 150.935 18.770 151.475 ;
        RECT 18.940 151.105 19.460 151.645 ;
        RECT 20.095 151.545 20.350 152.425 ;
        RECT 20.520 151.595 20.825 152.735 ;
        RECT 21.165 152.355 21.495 152.735 ;
        RECT 21.675 152.185 21.845 152.475 ;
        RECT 22.015 152.275 22.265 152.735 ;
        RECT 21.045 152.015 21.845 152.185 ;
        RECT 22.435 152.225 23.305 152.565 ;
        RECT 18.250 150.185 19.460 150.935 ;
        RECT 20.095 150.895 20.305 151.545 ;
        RECT 21.045 151.425 21.215 152.015 ;
        RECT 22.435 151.845 22.605 152.225 ;
        RECT 23.540 152.105 23.710 152.565 ;
        RECT 23.880 152.275 24.250 152.735 ;
        RECT 24.545 152.135 24.715 152.475 ;
        RECT 24.885 152.305 25.215 152.735 ;
        RECT 25.450 152.135 25.620 152.475 ;
        RECT 21.385 151.675 22.605 151.845 ;
        RECT 22.775 151.765 23.235 152.055 ;
        RECT 23.540 151.935 24.100 152.105 ;
        RECT 24.545 151.965 25.620 152.135 ;
        RECT 25.790 152.235 26.470 152.565 ;
        RECT 26.685 152.235 26.935 152.565 ;
        RECT 27.105 152.275 27.355 152.735 ;
        RECT 23.930 151.795 24.100 151.935 ;
        RECT 22.775 151.755 23.740 151.765 ;
        RECT 22.435 151.585 22.605 151.675 ;
        RECT 23.065 151.595 23.740 151.755 ;
        RECT 20.475 151.395 21.215 151.425 ;
        RECT 20.475 151.095 21.390 151.395 ;
        RECT 21.065 150.920 21.390 151.095 ;
        RECT 20.095 150.365 20.350 150.895 ;
        RECT 20.520 150.185 20.825 150.645 ;
        RECT 21.070 150.565 21.390 150.920 ;
        RECT 21.560 151.135 22.100 151.505 ;
        RECT 22.435 151.415 22.840 151.585 ;
        RECT 21.560 150.735 21.800 151.135 ;
        RECT 22.280 150.965 22.500 151.245 ;
        RECT 21.970 150.795 22.500 150.965 ;
        RECT 21.970 150.565 22.140 150.795 ;
        RECT 22.670 150.635 22.840 151.415 ;
        RECT 23.010 150.805 23.360 151.425 ;
        RECT 23.530 150.805 23.740 151.595 ;
        RECT 23.930 151.625 25.430 151.795 ;
        RECT 23.930 150.935 24.100 151.625 ;
        RECT 25.790 151.455 25.960 152.235 ;
        RECT 26.765 152.105 26.935 152.235 ;
        RECT 24.270 151.285 25.960 151.455 ;
        RECT 26.130 151.675 26.595 152.065 ;
        RECT 26.765 151.935 27.160 152.105 ;
        RECT 24.270 151.105 24.440 151.285 ;
        RECT 21.070 150.395 22.140 150.565 ;
        RECT 22.310 150.185 22.500 150.625 ;
        RECT 22.670 150.355 23.620 150.635 ;
        RECT 23.930 150.545 24.190 150.935 ;
        RECT 24.610 150.865 25.400 151.115 ;
        RECT 23.840 150.375 24.190 150.545 ;
        RECT 24.400 150.185 24.730 150.645 ;
        RECT 25.605 150.575 25.775 151.285 ;
        RECT 26.130 151.085 26.300 151.675 ;
        RECT 25.945 150.865 26.300 151.085 ;
        RECT 26.470 150.865 26.820 151.485 ;
        RECT 26.990 150.575 27.160 151.935 ;
        RECT 27.525 151.765 27.850 152.550 ;
        RECT 27.330 150.715 27.790 151.765 ;
        RECT 25.605 150.405 26.460 150.575 ;
        RECT 26.665 150.405 27.160 150.575 ;
        RECT 27.330 150.185 27.660 150.545 ;
        RECT 28.020 150.445 28.190 152.565 ;
        RECT 28.360 152.235 28.690 152.735 ;
        RECT 28.860 152.065 29.115 152.565 ;
        RECT 28.365 151.895 29.115 152.065 ;
        RECT 28.365 150.905 28.595 151.895 ;
        RECT 28.765 151.075 29.115 151.725 ;
        RECT 29.290 151.660 29.560 152.565 ;
        RECT 29.730 151.975 30.060 152.735 ;
        RECT 30.240 151.805 30.410 152.565 ;
        RECT 28.365 150.735 29.115 150.905 ;
        RECT 28.360 150.185 28.690 150.565 ;
        RECT 28.860 150.445 29.115 150.735 ;
        RECT 29.290 150.860 29.460 151.660 ;
        RECT 29.745 151.635 30.410 151.805 ;
        RECT 30.760 151.805 30.930 152.565 ;
        RECT 31.110 151.975 31.440 152.735 ;
        RECT 30.760 151.635 31.425 151.805 ;
        RECT 31.610 151.660 31.880 152.565 ;
        RECT 29.745 151.490 29.915 151.635 ;
        RECT 29.630 151.160 29.915 151.490 ;
        RECT 31.255 151.490 31.425 151.635 ;
        RECT 29.745 150.905 29.915 151.160 ;
        RECT 30.150 151.085 30.480 151.455 ;
        RECT 30.690 151.085 31.020 151.455 ;
        RECT 31.255 151.160 31.540 151.490 ;
        RECT 31.255 150.905 31.425 151.160 ;
        RECT 29.290 150.355 29.550 150.860 ;
        RECT 29.745 150.735 30.410 150.905 ;
        RECT 29.730 150.185 30.060 150.565 ;
        RECT 30.240 150.355 30.410 150.735 ;
        RECT 30.760 150.735 31.425 150.905 ;
        RECT 31.710 150.860 31.880 151.660 ;
        RECT 30.760 150.355 30.930 150.735 ;
        RECT 31.110 150.185 31.440 150.565 ;
        RECT 31.620 150.355 31.880 150.860 ;
        RECT 32.050 151.595 32.320 152.565 ;
        RECT 32.530 151.935 32.810 152.735 ;
        RECT 32.980 152.225 34.635 152.515 ;
        RECT 33.045 151.885 34.635 152.055 ;
        RECT 33.045 151.765 33.215 151.885 ;
        RECT 32.490 151.595 33.215 151.765 ;
        RECT 32.050 150.860 32.220 151.595 ;
        RECT 32.490 151.425 32.660 151.595 ;
        RECT 33.405 151.545 34.120 151.715 ;
        RECT 34.315 151.595 34.635 151.885 ;
        RECT 34.810 151.570 35.100 152.735 ;
        RECT 35.270 151.595 35.610 152.565 ;
        RECT 35.780 151.595 35.950 152.735 ;
        RECT 36.220 151.935 36.470 152.735 ;
        RECT 37.115 151.765 37.445 152.565 ;
        RECT 37.745 151.935 38.075 152.735 ;
        RECT 38.245 151.765 38.575 152.565 ;
        RECT 36.140 151.595 38.575 151.765 ;
        RECT 39.410 151.645 42.920 152.735 ;
        RECT 35.270 151.545 35.500 151.595 ;
        RECT 32.390 151.095 32.660 151.425 ;
        RECT 32.830 151.095 33.235 151.425 ;
        RECT 33.405 151.095 34.115 151.545 ;
        RECT 32.490 150.925 32.660 151.095 ;
        RECT 32.050 150.515 32.320 150.860 ;
        RECT 32.490 150.755 34.100 150.925 ;
        RECT 34.285 150.855 34.635 151.425 ;
        RECT 35.270 150.985 35.445 151.545 ;
        RECT 36.140 151.345 36.310 151.595 ;
        RECT 35.615 151.175 36.310 151.345 ;
        RECT 36.485 151.175 36.905 151.375 ;
        RECT 37.075 151.175 37.405 151.375 ;
        RECT 37.575 151.175 37.905 151.375 ;
        RECT 32.510 150.185 32.890 150.585 ;
        RECT 33.060 150.405 33.230 150.755 ;
        RECT 33.400 150.185 33.730 150.585 ;
        RECT 33.930 150.405 34.100 150.755 ;
        RECT 34.300 150.185 34.630 150.685 ;
        RECT 34.810 150.185 35.100 150.910 ;
        RECT 35.270 150.355 35.610 150.985 ;
        RECT 35.780 150.185 36.030 150.985 ;
        RECT 36.220 150.835 37.445 151.005 ;
        RECT 36.220 150.355 36.550 150.835 ;
        RECT 36.720 150.185 36.945 150.645 ;
        RECT 37.115 150.355 37.445 150.835 ;
        RECT 38.075 150.965 38.245 151.595 ;
        RECT 38.430 151.175 38.780 151.425 ;
        RECT 39.410 151.125 41.100 151.645 ;
        RECT 43.090 151.595 43.360 152.565 ;
        RECT 43.570 151.935 43.850 152.735 ;
        RECT 44.020 152.225 45.675 152.515 ;
        RECT 44.085 151.885 45.675 152.055 ;
        RECT 44.085 151.765 44.255 151.885 ;
        RECT 43.530 151.595 44.255 151.765 ;
        RECT 38.075 150.355 38.575 150.965 ;
        RECT 41.270 150.955 42.920 151.475 ;
        RECT 39.410 150.185 42.920 150.955 ;
        RECT 43.090 150.860 43.260 151.595 ;
        RECT 43.530 151.425 43.700 151.595 ;
        RECT 44.445 151.545 45.160 151.715 ;
        RECT 45.355 151.595 45.675 151.885 ;
        RECT 45.850 151.595 46.120 152.565 ;
        RECT 46.330 151.935 46.610 152.735 ;
        RECT 46.780 152.225 48.435 152.515 ;
        RECT 46.845 151.885 48.435 152.055 ;
        RECT 46.845 151.765 47.015 151.885 ;
        RECT 46.290 151.595 47.015 151.765 ;
        RECT 43.430 151.095 43.700 151.425 ;
        RECT 43.870 151.095 44.275 151.425 ;
        RECT 44.445 151.095 45.155 151.545 ;
        RECT 43.530 150.925 43.700 151.095 ;
        RECT 43.090 150.515 43.360 150.860 ;
        RECT 43.530 150.755 45.140 150.925 ;
        RECT 45.325 150.855 45.675 151.425 ;
        RECT 45.850 150.860 46.020 151.595 ;
        RECT 46.290 151.425 46.460 151.595 ;
        RECT 47.205 151.545 47.920 151.715 ;
        RECT 48.115 151.595 48.435 151.885 ;
        RECT 48.610 151.595 48.950 152.565 ;
        RECT 49.120 151.595 49.290 152.735 ;
        RECT 49.560 151.935 49.810 152.735 ;
        RECT 50.455 151.765 50.785 152.565 ;
        RECT 51.085 151.935 51.415 152.735 ;
        RECT 51.585 151.765 51.915 152.565 ;
        RECT 49.480 151.595 51.915 151.765 ;
        RECT 52.290 151.975 52.805 152.385 ;
        RECT 53.040 151.975 53.210 152.735 ;
        RECT 53.380 152.395 55.410 152.565 ;
        RECT 48.610 151.545 48.840 151.595 ;
        RECT 46.190 151.095 46.460 151.425 ;
        RECT 46.630 151.095 47.035 151.425 ;
        RECT 47.205 151.095 47.915 151.545 ;
        RECT 46.290 150.925 46.460 151.095 ;
        RECT 43.550 150.185 43.930 150.585 ;
        RECT 44.100 150.405 44.270 150.755 ;
        RECT 44.440 150.185 44.770 150.585 ;
        RECT 44.970 150.405 45.140 150.755 ;
        RECT 45.340 150.185 45.670 150.685 ;
        RECT 45.850 150.515 46.120 150.860 ;
        RECT 46.290 150.755 47.900 150.925 ;
        RECT 48.085 150.855 48.435 151.425 ;
        RECT 48.610 150.985 48.785 151.545 ;
        RECT 49.480 151.345 49.650 151.595 ;
        RECT 48.955 151.175 49.650 151.345 ;
        RECT 49.825 151.175 50.245 151.375 ;
        RECT 50.415 151.175 50.745 151.375 ;
        RECT 50.915 151.175 51.245 151.375 ;
        RECT 46.310 150.185 46.690 150.585 ;
        RECT 46.860 150.405 47.030 150.755 ;
        RECT 47.200 150.185 47.530 150.585 ;
        RECT 47.730 150.405 47.900 150.755 ;
        RECT 48.100 150.185 48.430 150.685 ;
        RECT 48.610 150.355 48.950 150.985 ;
        RECT 49.120 150.185 49.370 150.985 ;
        RECT 49.560 150.835 50.785 151.005 ;
        RECT 49.560 150.355 49.890 150.835 ;
        RECT 50.060 150.185 50.285 150.645 ;
        RECT 50.455 150.355 50.785 150.835 ;
        RECT 51.415 150.965 51.585 151.595 ;
        RECT 51.770 151.175 52.120 151.425 ;
        RECT 52.290 151.165 52.630 151.975 ;
        RECT 53.380 151.730 53.550 152.395 ;
        RECT 53.945 152.055 55.070 152.225 ;
        RECT 52.800 151.540 53.550 151.730 ;
        RECT 53.720 151.715 54.730 151.885 ;
        RECT 52.290 150.995 53.520 151.165 ;
        RECT 51.415 150.355 51.915 150.965 ;
        RECT 52.565 150.390 52.810 150.995 ;
        RECT 53.030 150.185 53.540 150.720 ;
        RECT 53.720 150.355 53.910 151.715 ;
        RECT 54.080 150.695 54.355 151.515 ;
        RECT 54.560 150.915 54.730 151.715 ;
        RECT 54.900 150.925 55.070 152.055 ;
        RECT 55.240 151.425 55.410 152.395 ;
        RECT 55.580 151.595 55.750 152.735 ;
        RECT 55.920 151.595 56.255 152.565 ;
        RECT 57.005 152.105 57.290 152.565 ;
        RECT 57.460 152.275 57.730 152.735 ;
        RECT 57.005 151.885 57.960 152.105 ;
        RECT 55.240 151.095 55.435 151.425 ;
        RECT 55.660 151.095 55.915 151.425 ;
        RECT 55.660 150.925 55.830 151.095 ;
        RECT 56.085 150.925 56.255 151.595 ;
        RECT 56.890 151.155 57.580 151.715 ;
        RECT 57.750 150.985 57.960 151.885 ;
        RECT 54.900 150.755 55.830 150.925 ;
        RECT 54.900 150.720 55.075 150.755 ;
        RECT 54.080 150.525 54.360 150.695 ;
        RECT 54.080 150.355 54.355 150.525 ;
        RECT 54.545 150.355 55.075 150.720 ;
        RECT 55.500 150.185 55.830 150.585 ;
        RECT 56.000 150.355 56.255 150.925 ;
        RECT 57.005 150.815 57.960 150.985 ;
        RECT 58.130 151.715 58.530 152.565 ;
        RECT 58.720 152.105 59.000 152.565 ;
        RECT 59.520 152.275 59.845 152.735 ;
        RECT 58.720 151.885 59.845 152.105 ;
        RECT 58.130 151.155 59.225 151.715 ;
        RECT 59.395 151.425 59.845 151.885 ;
        RECT 60.015 151.595 60.400 152.565 ;
        RECT 57.005 150.355 57.290 150.815 ;
        RECT 57.460 150.185 57.730 150.645 ;
        RECT 58.130 150.355 58.530 151.155 ;
        RECT 59.395 151.095 59.950 151.425 ;
        RECT 59.395 150.985 59.845 151.095 ;
        RECT 58.720 150.815 59.845 150.985 ;
        RECT 60.120 150.925 60.400 151.595 ;
        RECT 60.570 151.570 60.860 152.735 ;
        RECT 62.040 151.805 62.210 152.565 ;
        RECT 62.425 151.975 62.755 152.735 ;
        RECT 62.040 151.635 62.755 151.805 ;
        RECT 62.925 151.660 63.180 152.565 ;
        RECT 61.950 151.085 62.305 151.455 ;
        RECT 62.585 151.425 62.755 151.635 ;
        RECT 62.585 151.095 62.840 151.425 ;
        RECT 58.720 150.355 59.000 150.815 ;
        RECT 59.520 150.185 59.845 150.645 ;
        RECT 60.015 150.355 60.400 150.925 ;
        RECT 60.570 150.185 60.860 150.910 ;
        RECT 62.585 150.905 62.755 151.095 ;
        RECT 63.010 150.930 63.180 151.660 ;
        RECT 63.355 151.585 63.615 152.735 ;
        RECT 63.845 151.865 64.130 152.735 ;
        RECT 64.300 152.105 64.560 152.565 ;
        RECT 64.735 152.275 64.990 152.735 ;
        RECT 65.160 152.105 65.420 152.565 ;
        RECT 64.300 151.935 65.420 152.105 ;
        RECT 65.590 151.935 65.900 152.735 ;
        RECT 64.300 151.685 64.560 151.935 ;
        RECT 66.070 151.765 66.380 152.565 ;
        RECT 63.805 151.515 64.560 151.685 ;
        RECT 65.350 151.595 66.380 151.765 ;
        RECT 66.640 151.805 66.810 152.565 ;
        RECT 67.025 151.975 67.355 152.735 ;
        RECT 66.640 151.635 67.355 151.805 ;
        RECT 67.525 151.660 67.780 152.565 ;
        RECT 62.040 150.735 62.755 150.905 ;
        RECT 62.040 150.355 62.210 150.735 ;
        RECT 62.425 150.185 62.755 150.565 ;
        RECT 62.925 150.355 63.180 150.930 ;
        RECT 63.355 150.185 63.615 151.025 ;
        RECT 63.805 151.005 64.210 151.515 ;
        RECT 65.350 151.345 65.520 151.595 ;
        RECT 64.380 151.175 65.520 151.345 ;
        RECT 63.805 150.835 65.455 151.005 ;
        RECT 65.690 150.855 66.040 151.425 ;
        RECT 63.850 150.185 64.130 150.665 ;
        RECT 64.300 150.445 64.560 150.835 ;
        RECT 64.735 150.185 64.990 150.665 ;
        RECT 65.160 150.445 65.455 150.835 ;
        RECT 66.210 150.685 66.380 151.595 ;
        RECT 66.550 151.085 66.905 151.455 ;
        RECT 67.185 151.425 67.355 151.635 ;
        RECT 67.185 151.095 67.440 151.425 ;
        RECT 67.185 150.905 67.355 151.095 ;
        RECT 67.610 150.930 67.780 151.660 ;
        RECT 67.955 151.585 68.215 152.735 ;
        RECT 68.480 151.805 68.650 152.565 ;
        RECT 68.865 151.975 69.195 152.735 ;
        RECT 68.480 151.635 69.195 151.805 ;
        RECT 69.365 151.660 69.620 152.565 ;
        RECT 68.390 151.085 68.745 151.455 ;
        RECT 69.025 151.425 69.195 151.635 ;
        RECT 69.025 151.095 69.280 151.425 ;
        RECT 65.635 150.185 65.910 150.665 ;
        RECT 66.080 150.355 66.380 150.685 ;
        RECT 66.640 150.735 67.355 150.905 ;
        RECT 66.640 150.355 66.810 150.735 ;
        RECT 67.025 150.185 67.355 150.565 ;
        RECT 67.525 150.355 67.780 150.930 ;
        RECT 67.955 150.185 68.215 151.025 ;
        RECT 69.025 150.905 69.195 151.095 ;
        RECT 69.450 150.930 69.620 151.660 ;
        RECT 69.795 151.585 70.055 152.735 ;
        RECT 70.690 151.645 72.360 152.735 ;
        RECT 70.690 151.125 71.440 151.645 ;
        RECT 72.530 151.595 72.870 152.565 ;
        RECT 73.040 151.595 73.210 152.735 ;
        RECT 73.480 151.935 73.730 152.735 ;
        RECT 74.375 151.765 74.705 152.565 ;
        RECT 75.005 151.935 75.335 152.735 ;
        RECT 75.505 151.765 75.835 152.565 ;
        RECT 73.400 151.595 75.835 151.765 ;
        RECT 76.210 151.595 76.550 152.565 ;
        RECT 76.720 151.595 76.890 152.735 ;
        RECT 77.160 151.935 77.410 152.735 ;
        RECT 78.055 151.765 78.385 152.565 ;
        RECT 78.685 151.935 79.015 152.735 ;
        RECT 79.185 151.765 79.515 152.565 ;
        RECT 77.080 151.595 79.515 151.765 ;
        RECT 80.850 151.595 81.080 152.735 ;
        RECT 68.480 150.735 69.195 150.905 ;
        RECT 68.480 150.355 68.650 150.735 ;
        RECT 68.865 150.185 69.195 150.565 ;
        RECT 69.365 150.355 69.620 150.930 ;
        RECT 69.795 150.185 70.055 151.025 ;
        RECT 71.610 150.955 72.360 151.475 ;
        RECT 70.690 150.185 72.360 150.955 ;
        RECT 72.530 150.985 72.705 151.595 ;
        RECT 73.400 151.345 73.570 151.595 ;
        RECT 72.875 151.175 73.570 151.345 ;
        RECT 73.745 151.175 74.165 151.375 ;
        RECT 74.335 151.175 74.665 151.375 ;
        RECT 74.835 151.175 75.165 151.375 ;
        RECT 72.530 150.355 72.870 150.985 ;
        RECT 73.040 150.185 73.290 150.985 ;
        RECT 73.480 150.835 74.705 151.005 ;
        RECT 73.480 150.355 73.810 150.835 ;
        RECT 73.980 150.185 74.205 150.645 ;
        RECT 74.375 150.355 74.705 150.835 ;
        RECT 75.335 150.965 75.505 151.595 ;
        RECT 75.690 151.175 76.040 151.425 ;
        RECT 76.210 150.985 76.385 151.595 ;
        RECT 77.080 151.345 77.250 151.595 ;
        RECT 76.555 151.175 77.250 151.345 ;
        RECT 77.425 151.175 77.845 151.375 ;
        RECT 78.015 151.175 78.345 151.375 ;
        RECT 78.515 151.175 78.845 151.375 ;
        RECT 75.335 150.355 75.835 150.965 ;
        RECT 76.210 150.355 76.550 150.985 ;
        RECT 76.720 150.185 76.970 150.985 ;
        RECT 77.160 150.835 78.385 151.005 ;
        RECT 77.160 150.355 77.490 150.835 ;
        RECT 77.660 150.185 77.885 150.645 ;
        RECT 78.055 150.355 78.385 150.835 ;
        RECT 79.015 150.965 79.185 151.595 ;
        RECT 81.250 151.585 81.580 152.565 ;
        RECT 81.750 151.595 81.960 152.735 ;
        RECT 82.190 151.975 82.705 152.385 ;
        RECT 82.940 151.975 83.110 152.735 ;
        RECT 83.280 152.395 85.310 152.565 ;
        RECT 79.370 151.175 79.720 151.425 ;
        RECT 80.830 151.175 81.160 151.425 ;
        RECT 79.015 150.355 79.515 150.965 ;
        RECT 80.850 150.185 81.080 151.005 ;
        RECT 81.330 150.985 81.580 151.585 ;
        RECT 82.190 151.165 82.530 151.975 ;
        RECT 83.280 151.730 83.450 152.395 ;
        RECT 83.845 152.055 84.970 152.225 ;
        RECT 82.700 151.540 83.450 151.730 ;
        RECT 83.620 151.715 84.630 151.885 ;
        RECT 81.250 150.355 81.580 150.985 ;
        RECT 81.750 150.185 81.960 151.005 ;
        RECT 82.190 150.995 83.420 151.165 ;
        RECT 82.465 150.390 82.710 150.995 ;
        RECT 82.930 150.185 83.440 150.720 ;
        RECT 83.620 150.355 83.810 151.715 ;
        RECT 83.980 151.035 84.255 151.515 ;
        RECT 83.980 150.865 84.260 151.035 ;
        RECT 84.460 150.915 84.630 151.715 ;
        RECT 84.800 150.925 84.970 152.055 ;
        RECT 85.140 151.425 85.310 152.395 ;
        RECT 85.480 151.595 85.650 152.735 ;
        RECT 85.820 151.595 86.155 152.565 ;
        RECT 85.140 151.095 85.335 151.425 ;
        RECT 85.560 151.095 85.815 151.425 ;
        RECT 85.560 150.925 85.730 151.095 ;
        RECT 85.985 150.925 86.155 151.595 ;
        RECT 86.330 151.570 86.620 152.735 ;
        RECT 87.800 151.805 87.970 152.565 ;
        RECT 88.150 151.975 88.480 152.735 ;
        RECT 87.800 151.635 88.465 151.805 ;
        RECT 88.650 151.660 88.920 152.565 ;
        RECT 88.295 151.490 88.465 151.635 ;
        RECT 87.730 151.085 88.060 151.455 ;
        RECT 88.295 151.160 88.580 151.490 ;
        RECT 83.980 150.355 84.255 150.865 ;
        RECT 84.800 150.755 85.730 150.925 ;
        RECT 84.800 150.720 84.975 150.755 ;
        RECT 84.445 150.355 84.975 150.720 ;
        RECT 85.400 150.185 85.730 150.585 ;
        RECT 85.900 150.355 86.155 150.925 ;
        RECT 86.330 150.185 86.620 150.910 ;
        RECT 88.295 150.905 88.465 151.160 ;
        RECT 87.800 150.735 88.465 150.905 ;
        RECT 88.750 150.860 88.920 151.660 ;
        RECT 89.090 151.645 91.680 152.735 ;
        RECT 92.055 151.765 92.385 152.565 ;
        RECT 92.555 151.935 92.885 152.735 ;
        RECT 93.185 151.765 93.515 152.565 ;
        RECT 94.160 151.935 94.410 152.735 ;
        RECT 89.090 151.125 90.300 151.645 ;
        RECT 92.055 151.595 94.490 151.765 ;
        RECT 94.680 151.595 94.850 152.735 ;
        RECT 95.020 151.595 95.360 152.565 ;
        RECT 90.470 150.955 91.680 151.475 ;
        RECT 91.850 151.175 92.200 151.425 ;
        RECT 92.385 150.965 92.555 151.595 ;
        RECT 92.725 151.175 93.055 151.375 ;
        RECT 93.225 151.175 93.555 151.375 ;
        RECT 93.725 151.175 94.145 151.375 ;
        RECT 94.320 151.345 94.490 151.595 ;
        RECT 94.320 151.175 95.015 151.345 ;
        RECT 87.800 150.355 87.970 150.735 ;
        RECT 88.150 150.185 88.480 150.565 ;
        RECT 88.660 150.355 88.920 150.860 ;
        RECT 89.090 150.185 91.680 150.955 ;
        RECT 92.055 150.355 92.555 150.965 ;
        RECT 93.185 150.835 94.410 151.005 ;
        RECT 95.185 150.985 95.360 151.595 ;
        RECT 93.185 150.355 93.515 150.835 ;
        RECT 93.685 150.185 93.910 150.645 ;
        RECT 94.080 150.355 94.410 150.835 ;
        RECT 94.600 150.185 94.850 150.985 ;
        RECT 95.020 150.355 95.360 150.985 ;
        RECT 95.530 151.595 95.870 152.565 ;
        RECT 96.040 151.595 96.210 152.735 ;
        RECT 96.480 151.935 96.730 152.735 ;
        RECT 97.375 151.765 97.705 152.565 ;
        RECT 98.005 151.935 98.335 152.735 ;
        RECT 98.505 151.765 98.835 152.565 ;
        RECT 96.400 151.595 98.835 151.765 ;
        RECT 99.710 151.595 99.940 152.735 ;
        RECT 95.530 150.985 95.705 151.595 ;
        RECT 96.400 151.345 96.570 151.595 ;
        RECT 95.875 151.175 96.570 151.345 ;
        RECT 96.745 151.175 97.165 151.375 ;
        RECT 97.335 151.175 97.665 151.375 ;
        RECT 97.835 151.175 98.165 151.375 ;
        RECT 95.530 150.355 95.870 150.985 ;
        RECT 96.040 150.185 96.290 150.985 ;
        RECT 96.480 150.835 97.705 151.005 ;
        RECT 96.480 150.355 96.810 150.835 ;
        RECT 96.980 150.185 97.205 150.645 ;
        RECT 97.375 150.355 97.705 150.835 ;
        RECT 98.335 150.965 98.505 151.595 ;
        RECT 100.110 151.585 100.440 152.565 ;
        RECT 100.610 151.595 100.820 152.735 ;
        RECT 98.690 151.175 99.040 151.425 ;
        RECT 99.690 151.175 100.020 151.425 ;
        RECT 98.335 150.355 98.835 150.965 ;
        RECT 99.710 150.185 99.940 151.005 ;
        RECT 100.190 150.985 100.440 151.585 ;
        RECT 101.055 151.545 101.310 152.425 ;
        RECT 101.480 151.595 101.785 152.735 ;
        RECT 102.125 152.355 102.455 152.735 ;
        RECT 102.635 152.185 102.805 152.475 ;
        RECT 102.975 152.275 103.225 152.735 ;
        RECT 102.005 152.015 102.805 152.185 ;
        RECT 103.395 152.225 104.265 152.565 ;
        RECT 100.110 150.355 100.440 150.985 ;
        RECT 100.610 150.185 100.820 151.005 ;
        RECT 101.055 150.895 101.265 151.545 ;
        RECT 102.005 151.425 102.175 152.015 ;
        RECT 103.395 151.845 103.565 152.225 ;
        RECT 104.500 152.105 104.670 152.565 ;
        RECT 104.840 152.275 105.210 152.735 ;
        RECT 105.505 152.135 105.675 152.475 ;
        RECT 105.845 152.305 106.175 152.735 ;
        RECT 106.410 152.135 106.580 152.475 ;
        RECT 102.345 151.675 103.565 151.845 ;
        RECT 103.735 151.765 104.195 152.055 ;
        RECT 104.500 151.935 105.060 152.105 ;
        RECT 105.505 151.965 106.580 152.135 ;
        RECT 106.750 152.235 107.430 152.565 ;
        RECT 107.645 152.235 107.895 152.565 ;
        RECT 108.065 152.275 108.315 152.735 ;
        RECT 104.890 151.795 105.060 151.935 ;
        RECT 103.735 151.755 104.700 151.765 ;
        RECT 103.395 151.585 103.565 151.675 ;
        RECT 104.025 151.595 104.700 151.755 ;
        RECT 101.435 151.395 102.175 151.425 ;
        RECT 101.435 151.095 102.350 151.395 ;
        RECT 102.025 150.920 102.350 151.095 ;
        RECT 101.055 150.365 101.310 150.895 ;
        RECT 101.480 150.185 101.785 150.645 ;
        RECT 102.030 150.565 102.350 150.920 ;
        RECT 102.520 151.135 103.060 151.505 ;
        RECT 103.395 151.415 103.800 151.585 ;
        RECT 102.520 150.735 102.760 151.135 ;
        RECT 103.240 150.965 103.460 151.245 ;
        RECT 102.930 150.795 103.460 150.965 ;
        RECT 102.930 150.565 103.100 150.795 ;
        RECT 103.630 150.635 103.800 151.415 ;
        RECT 103.970 150.805 104.320 151.425 ;
        RECT 104.490 150.805 104.700 151.595 ;
        RECT 104.890 151.625 106.390 151.795 ;
        RECT 104.890 150.935 105.060 151.625 ;
        RECT 106.750 151.455 106.920 152.235 ;
        RECT 107.725 152.105 107.895 152.235 ;
        RECT 105.230 151.285 106.920 151.455 ;
        RECT 107.090 151.675 107.555 152.065 ;
        RECT 107.725 151.935 108.120 152.105 ;
        RECT 105.230 151.105 105.400 151.285 ;
        RECT 102.030 150.395 103.100 150.565 ;
        RECT 103.270 150.185 103.460 150.625 ;
        RECT 103.630 150.355 104.580 150.635 ;
        RECT 104.890 150.545 105.150 150.935 ;
        RECT 105.570 150.865 106.360 151.115 ;
        RECT 104.800 150.375 105.150 150.545 ;
        RECT 105.360 150.185 105.690 150.645 ;
        RECT 106.565 150.575 106.735 151.285 ;
        RECT 107.090 151.085 107.260 151.675 ;
        RECT 106.905 150.865 107.260 151.085 ;
        RECT 107.430 150.865 107.780 151.485 ;
        RECT 107.950 150.575 108.120 151.935 ;
        RECT 108.485 151.765 108.810 152.550 ;
        RECT 108.290 150.715 108.750 151.765 ;
        RECT 106.565 150.405 107.420 150.575 ;
        RECT 107.625 150.405 108.120 150.575 ;
        RECT 108.290 150.185 108.620 150.545 ;
        RECT 108.980 150.445 109.150 152.565 ;
        RECT 109.320 152.235 109.650 152.735 ;
        RECT 109.820 152.065 110.075 152.565 ;
        RECT 109.325 151.895 110.075 152.065 ;
        RECT 109.325 150.905 109.555 151.895 ;
        RECT 109.725 151.075 110.075 151.725 ;
        RECT 111.170 151.645 112.380 152.735 ;
        RECT 111.170 151.105 111.690 151.645 ;
        RECT 111.860 150.935 112.380 151.475 ;
        RECT 109.325 150.735 110.075 150.905 ;
        RECT 109.320 150.185 109.650 150.565 ;
        RECT 109.820 150.445 110.075 150.735 ;
        RECT 111.170 150.185 112.380 150.935 ;
        RECT 18.165 150.015 112.465 150.185 ;
        RECT 18.250 149.265 19.460 150.015 ;
        RECT 18.250 148.725 18.770 149.265 ;
        RECT 20.090 149.245 21.760 150.015 ;
        RECT 21.930 149.290 22.220 150.015 ;
        RECT 22.390 149.265 23.600 150.015 ;
        RECT 18.940 148.555 19.460 149.095 ;
        RECT 18.250 147.465 19.460 148.555 ;
        RECT 20.090 148.555 20.840 149.075 ;
        RECT 21.010 148.725 21.760 149.245 ;
        RECT 20.090 147.465 21.760 148.555 ;
        RECT 21.930 147.465 22.220 148.630 ;
        RECT 22.390 148.555 22.910 149.095 ;
        RECT 23.080 148.725 23.600 149.265 ;
        RECT 24.045 149.205 24.290 149.810 ;
        RECT 24.510 149.480 25.020 150.015 ;
        RECT 23.770 149.035 25.000 149.205 ;
        RECT 22.390 147.465 23.600 148.555 ;
        RECT 23.770 148.225 24.110 149.035 ;
        RECT 24.280 148.470 25.030 148.660 ;
        RECT 23.770 147.815 24.285 148.225 ;
        RECT 24.520 147.465 24.690 148.225 ;
        RECT 24.860 147.805 25.030 148.470 ;
        RECT 25.200 148.485 25.390 149.845 ;
        RECT 25.560 148.995 25.835 149.845 ;
        RECT 26.025 149.480 26.555 149.845 ;
        RECT 26.980 149.615 27.310 150.015 ;
        RECT 26.380 149.445 26.555 149.480 ;
        RECT 25.560 148.825 25.840 148.995 ;
        RECT 25.560 148.685 25.835 148.825 ;
        RECT 26.040 148.485 26.210 149.285 ;
        RECT 25.200 148.315 26.210 148.485 ;
        RECT 26.380 149.275 27.310 149.445 ;
        RECT 27.480 149.275 27.735 149.845 ;
        RECT 26.380 148.145 26.550 149.275 ;
        RECT 27.140 149.105 27.310 149.275 ;
        RECT 25.425 147.975 26.550 148.145 ;
        RECT 26.720 148.775 26.915 149.105 ;
        RECT 27.140 148.775 27.395 149.105 ;
        RECT 26.720 147.805 26.890 148.775 ;
        RECT 27.565 148.605 27.735 149.275 ;
        RECT 28.370 149.245 30.040 150.015 ;
        RECT 24.860 147.635 26.890 147.805 ;
        RECT 27.060 147.465 27.230 148.605 ;
        RECT 27.400 147.635 27.735 148.605 ;
        RECT 28.370 148.555 29.120 149.075 ;
        RECT 29.290 148.725 30.040 149.245 ;
        RECT 30.270 149.195 30.480 150.015 ;
        RECT 30.650 149.215 30.980 149.845 ;
        RECT 30.650 148.615 30.900 149.215 ;
        RECT 31.150 149.195 31.380 150.015 ;
        RECT 31.590 149.215 31.930 149.845 ;
        RECT 32.100 149.215 32.350 150.015 ;
        RECT 32.540 149.365 32.870 149.845 ;
        RECT 33.040 149.555 33.265 150.015 ;
        RECT 33.435 149.365 33.765 149.845 ;
        RECT 31.070 148.775 31.400 149.025 ;
        RECT 28.370 147.465 30.040 148.555 ;
        RECT 30.270 147.465 30.480 148.605 ;
        RECT 30.650 147.635 30.980 148.615 ;
        RECT 31.590 148.605 31.765 149.215 ;
        RECT 32.540 149.195 33.765 149.365 ;
        RECT 34.395 149.235 34.895 149.845 ;
        RECT 31.935 148.855 32.630 149.025 ;
        RECT 32.460 148.605 32.630 148.855 ;
        RECT 32.805 148.825 33.225 149.025 ;
        RECT 33.395 148.825 33.725 149.025 ;
        RECT 33.895 148.825 34.225 149.025 ;
        RECT 34.395 148.605 34.565 149.235 ;
        RECT 36.190 149.215 36.530 149.845 ;
        RECT 36.700 149.215 36.950 150.015 ;
        RECT 37.140 149.365 37.470 149.845 ;
        RECT 37.640 149.555 37.865 150.015 ;
        RECT 38.035 149.365 38.365 149.845 ;
        RECT 34.750 148.775 35.100 149.025 ;
        RECT 36.190 148.605 36.365 149.215 ;
        RECT 37.140 149.195 38.365 149.365 ;
        RECT 38.995 149.235 39.495 149.845 ;
        RECT 39.985 149.385 40.270 149.845 ;
        RECT 40.440 149.555 40.710 150.015 ;
        RECT 36.535 148.855 37.230 149.025 ;
        RECT 37.060 148.605 37.230 148.855 ;
        RECT 37.405 148.825 37.825 149.025 ;
        RECT 37.995 148.825 38.325 149.025 ;
        RECT 38.495 148.825 38.825 149.025 ;
        RECT 38.995 148.605 39.165 149.235 ;
        RECT 39.985 149.215 40.940 149.385 ;
        RECT 39.350 148.775 39.700 149.025 ;
        RECT 31.150 147.465 31.380 148.605 ;
        RECT 31.590 147.635 31.930 148.605 ;
        RECT 32.100 147.465 32.270 148.605 ;
        RECT 32.460 148.435 34.895 148.605 ;
        RECT 32.540 147.465 32.790 148.265 ;
        RECT 33.435 147.635 33.765 148.435 ;
        RECT 34.065 147.465 34.395 148.265 ;
        RECT 34.565 147.635 34.895 148.435 ;
        RECT 36.190 147.635 36.530 148.605 ;
        RECT 36.700 147.465 36.870 148.605 ;
        RECT 37.060 148.435 39.495 148.605 ;
        RECT 39.870 148.485 40.560 149.045 ;
        RECT 37.140 147.465 37.390 148.265 ;
        RECT 38.035 147.635 38.365 148.435 ;
        RECT 38.665 147.465 38.995 148.265 ;
        RECT 39.165 147.635 39.495 148.435 ;
        RECT 40.730 148.315 40.940 149.215 ;
        RECT 39.985 148.095 40.940 148.315 ;
        RECT 41.110 149.045 41.510 149.845 ;
        RECT 41.700 149.385 41.980 149.845 ;
        RECT 42.500 149.555 42.825 150.015 ;
        RECT 41.700 149.215 42.825 149.385 ;
        RECT 42.995 149.275 43.380 149.845 ;
        RECT 42.375 149.105 42.825 149.215 ;
        RECT 41.110 148.485 42.205 149.045 ;
        RECT 42.375 148.775 42.930 149.105 ;
        RECT 39.985 147.635 40.270 148.095 ;
        RECT 40.440 147.465 40.710 147.925 ;
        RECT 41.110 147.635 41.510 148.485 ;
        RECT 42.375 148.315 42.825 148.775 ;
        RECT 43.100 148.605 43.380 149.275 ;
        RECT 43.825 149.205 44.070 149.810 ;
        RECT 44.290 149.480 44.800 150.015 ;
        RECT 41.700 148.095 42.825 148.315 ;
        RECT 41.700 147.635 41.980 148.095 ;
        RECT 42.500 147.465 42.825 147.925 ;
        RECT 42.995 147.635 43.380 148.605 ;
        RECT 43.550 149.035 44.780 149.205 ;
        RECT 43.550 148.225 43.890 149.035 ;
        RECT 44.060 148.470 44.810 148.660 ;
        RECT 43.550 147.815 44.065 148.225 ;
        RECT 44.300 147.465 44.470 148.225 ;
        RECT 44.640 147.805 44.810 148.470 ;
        RECT 44.980 148.485 45.170 149.845 ;
        RECT 45.340 148.995 45.615 149.845 ;
        RECT 45.805 149.480 46.335 149.845 ;
        RECT 46.760 149.615 47.090 150.015 ;
        RECT 46.160 149.445 46.335 149.480 ;
        RECT 45.340 148.825 45.620 148.995 ;
        RECT 45.340 148.685 45.615 148.825 ;
        RECT 45.820 148.485 45.990 149.285 ;
        RECT 44.980 148.315 45.990 148.485 ;
        RECT 46.160 149.275 47.090 149.445 ;
        RECT 47.260 149.275 47.515 149.845 ;
        RECT 47.690 149.290 47.980 150.015 ;
        RECT 48.615 149.305 48.870 149.835 ;
        RECT 49.040 149.555 49.345 150.015 ;
        RECT 49.590 149.635 50.660 149.805 ;
        RECT 46.160 148.145 46.330 149.275 ;
        RECT 46.920 149.105 47.090 149.275 ;
        RECT 45.205 147.975 46.330 148.145 ;
        RECT 46.500 148.775 46.695 149.105 ;
        RECT 46.920 148.775 47.175 149.105 ;
        RECT 46.500 147.805 46.670 148.775 ;
        RECT 47.345 148.605 47.515 149.275 ;
        RECT 48.615 148.655 48.825 149.305 ;
        RECT 49.590 149.280 49.910 149.635 ;
        RECT 49.585 149.105 49.910 149.280 ;
        RECT 48.995 148.805 49.910 149.105 ;
        RECT 50.080 149.065 50.320 149.465 ;
        RECT 50.490 149.405 50.660 149.635 ;
        RECT 50.830 149.575 51.020 150.015 ;
        RECT 51.190 149.565 52.140 149.845 ;
        RECT 52.360 149.655 52.710 149.825 ;
        RECT 50.490 149.235 51.020 149.405 ;
        RECT 48.995 148.775 49.735 148.805 ;
        RECT 44.640 147.635 46.670 147.805 ;
        RECT 46.840 147.465 47.010 148.605 ;
        RECT 47.180 147.635 47.515 148.605 ;
        RECT 47.690 147.465 47.980 148.630 ;
        RECT 48.615 147.775 48.870 148.655 ;
        RECT 49.040 147.465 49.345 148.605 ;
        RECT 49.565 148.185 49.735 148.775 ;
        RECT 50.080 148.695 50.620 149.065 ;
        RECT 50.800 148.955 51.020 149.235 ;
        RECT 51.190 148.785 51.360 149.565 ;
        RECT 50.955 148.615 51.360 148.785 ;
        RECT 51.530 148.775 51.880 149.395 ;
        RECT 50.955 148.525 51.125 148.615 ;
        RECT 52.050 148.605 52.260 149.395 ;
        RECT 49.905 148.355 51.125 148.525 ;
        RECT 51.585 148.445 52.260 148.605 ;
        RECT 49.565 148.015 50.365 148.185 ;
        RECT 49.685 147.465 50.015 147.845 ;
        RECT 50.195 147.725 50.365 148.015 ;
        RECT 50.955 147.975 51.125 148.355 ;
        RECT 51.295 148.435 52.260 148.445 ;
        RECT 52.450 149.265 52.710 149.655 ;
        RECT 52.920 149.555 53.250 150.015 ;
        RECT 54.125 149.625 54.980 149.795 ;
        RECT 55.185 149.625 55.680 149.795 ;
        RECT 55.850 149.655 56.180 150.015 ;
        RECT 52.450 148.575 52.620 149.265 ;
        RECT 52.790 148.915 52.960 149.095 ;
        RECT 53.130 149.085 53.920 149.335 ;
        RECT 54.125 148.915 54.295 149.625 ;
        RECT 54.465 149.115 54.820 149.335 ;
        RECT 52.790 148.745 54.480 148.915 ;
        RECT 51.295 148.145 51.755 148.435 ;
        RECT 52.450 148.405 53.950 148.575 ;
        RECT 52.450 148.265 52.620 148.405 ;
        RECT 52.060 148.095 52.620 148.265 ;
        RECT 50.535 147.465 50.785 147.925 ;
        RECT 50.955 147.635 51.825 147.975 ;
        RECT 52.060 147.635 52.230 148.095 ;
        RECT 53.065 148.065 54.140 148.235 ;
        RECT 52.400 147.465 52.770 147.925 ;
        RECT 53.065 147.725 53.235 148.065 ;
        RECT 53.405 147.465 53.735 147.895 ;
        RECT 53.970 147.725 54.140 148.065 ;
        RECT 54.310 147.965 54.480 148.745 ;
        RECT 54.650 148.525 54.820 149.115 ;
        RECT 54.990 148.715 55.340 149.335 ;
        RECT 54.650 148.135 55.115 148.525 ;
        RECT 55.510 148.265 55.680 149.625 ;
        RECT 55.850 148.435 56.310 149.485 ;
        RECT 55.285 148.095 55.680 148.265 ;
        RECT 55.285 147.965 55.455 148.095 ;
        RECT 54.310 147.635 54.990 147.965 ;
        RECT 55.205 147.635 55.455 147.965 ;
        RECT 55.625 147.465 55.875 147.925 ;
        RECT 56.045 147.650 56.370 148.435 ;
        RECT 56.540 147.635 56.710 149.755 ;
        RECT 56.880 149.635 57.210 150.015 ;
        RECT 57.380 149.465 57.635 149.755 ;
        RECT 56.885 149.295 57.635 149.465 ;
        RECT 57.810 149.340 58.070 149.845 ;
        RECT 58.250 149.635 58.580 150.015 ;
        RECT 58.760 149.465 58.930 149.845 ;
        RECT 56.885 148.305 57.115 149.295 ;
        RECT 57.285 148.475 57.635 149.125 ;
        RECT 57.810 148.540 57.980 149.340 ;
        RECT 58.265 149.295 58.930 149.465 ;
        RECT 58.265 149.040 58.435 149.295 ;
        RECT 59.190 149.215 59.530 149.845 ;
        RECT 59.700 149.215 59.950 150.015 ;
        RECT 60.140 149.365 60.470 149.845 ;
        RECT 60.640 149.555 60.865 150.015 ;
        RECT 61.035 149.365 61.365 149.845 ;
        RECT 59.190 149.165 59.420 149.215 ;
        RECT 60.140 149.195 61.365 149.365 ;
        RECT 61.995 149.235 62.495 149.845 ;
        RECT 62.870 149.515 63.130 149.845 ;
        RECT 63.300 149.655 63.630 150.015 ;
        RECT 63.885 149.635 65.185 149.845 ;
        RECT 62.870 149.505 63.100 149.515 ;
        RECT 58.150 148.710 58.435 149.040 ;
        RECT 58.670 148.745 59.000 149.115 ;
        RECT 58.265 148.565 58.435 148.710 ;
        RECT 59.190 148.605 59.365 149.165 ;
        RECT 59.535 148.855 60.230 149.025 ;
        RECT 60.060 148.605 60.230 148.855 ;
        RECT 60.405 148.825 60.825 149.025 ;
        RECT 60.995 148.825 61.325 149.025 ;
        RECT 61.495 148.825 61.825 149.025 ;
        RECT 61.995 148.605 62.165 149.235 ;
        RECT 62.350 148.775 62.700 149.025 ;
        RECT 56.885 148.135 57.635 148.305 ;
        RECT 56.880 147.465 57.210 147.965 ;
        RECT 57.380 147.635 57.635 148.135 ;
        RECT 57.810 147.635 58.080 148.540 ;
        RECT 58.265 148.395 58.930 148.565 ;
        RECT 58.250 147.465 58.580 148.225 ;
        RECT 58.760 147.635 58.930 148.395 ;
        RECT 59.190 147.635 59.530 148.605 ;
        RECT 59.700 147.465 59.870 148.605 ;
        RECT 60.060 148.435 62.495 148.605 ;
        RECT 60.140 147.465 60.390 148.265 ;
        RECT 61.035 147.635 61.365 148.435 ;
        RECT 61.665 147.465 61.995 148.265 ;
        RECT 62.165 147.635 62.495 148.435 ;
        RECT 62.870 148.315 63.040 149.505 ;
        RECT 63.885 149.485 64.055 149.635 ;
        RECT 63.300 149.360 64.055 149.485 ;
        RECT 63.210 149.315 64.055 149.360 ;
        RECT 63.210 149.195 63.480 149.315 ;
        RECT 63.210 148.620 63.380 149.195 ;
        RECT 63.610 148.755 64.020 149.060 ;
        RECT 64.310 149.025 64.520 149.425 ;
        RECT 64.190 148.815 64.520 149.025 ;
        RECT 64.765 149.025 64.985 149.425 ;
        RECT 65.460 149.250 65.915 150.015 ;
        RECT 66.180 149.465 66.350 149.845 ;
        RECT 66.565 149.635 66.895 150.015 ;
        RECT 66.180 149.295 66.895 149.465 ;
        RECT 64.765 148.815 65.240 149.025 ;
        RECT 65.430 148.825 65.920 149.025 ;
        RECT 66.090 148.745 66.445 149.115 ;
        RECT 66.725 149.105 66.895 149.295 ;
        RECT 67.065 149.270 67.320 149.845 ;
        RECT 66.725 148.775 66.980 149.105 ;
        RECT 63.210 148.585 63.410 148.620 ;
        RECT 64.740 148.585 65.915 148.645 ;
        RECT 63.210 148.475 65.915 148.585 ;
        RECT 66.725 148.565 66.895 148.775 ;
        RECT 63.270 148.415 65.070 148.475 ;
        RECT 64.740 148.385 65.070 148.415 ;
        RECT 62.870 147.635 63.130 148.315 ;
        RECT 63.300 147.465 63.550 148.245 ;
        RECT 63.800 148.215 64.635 148.225 ;
        RECT 65.225 148.215 65.410 148.305 ;
        RECT 63.800 148.015 65.410 148.215 ;
        RECT 63.800 147.635 64.050 148.015 ;
        RECT 65.180 147.975 65.410 148.015 ;
        RECT 65.660 147.855 65.915 148.475 ;
        RECT 64.220 147.465 64.575 147.845 ;
        RECT 65.580 147.635 65.915 147.855 ;
        RECT 66.180 148.395 66.895 148.565 ;
        RECT 67.150 148.540 67.320 149.270 ;
        RECT 67.495 149.175 67.755 150.015 ;
        RECT 68.020 149.465 68.190 149.845 ;
        RECT 68.405 149.635 68.735 150.015 ;
        RECT 68.020 149.295 68.735 149.465 ;
        RECT 67.930 148.745 68.285 149.115 ;
        RECT 68.565 149.105 68.735 149.295 ;
        RECT 68.905 149.270 69.160 149.845 ;
        RECT 68.565 148.775 68.820 149.105 ;
        RECT 66.180 147.635 66.350 148.395 ;
        RECT 66.565 147.465 66.895 148.225 ;
        RECT 67.065 147.635 67.320 148.540 ;
        RECT 67.495 147.465 67.755 148.615 ;
        RECT 68.565 148.565 68.735 148.775 ;
        RECT 68.020 148.395 68.735 148.565 ;
        RECT 68.990 148.540 69.160 149.270 ;
        RECT 69.335 149.175 69.595 150.015 ;
        RECT 69.975 149.235 70.475 149.845 ;
        RECT 69.770 148.775 70.120 149.025 ;
        RECT 68.020 147.635 68.190 148.395 ;
        RECT 68.405 147.465 68.735 148.225 ;
        RECT 68.905 147.635 69.160 148.540 ;
        RECT 69.335 147.465 69.595 148.615 ;
        RECT 70.305 148.605 70.475 149.235 ;
        RECT 71.105 149.365 71.435 149.845 ;
        RECT 71.605 149.555 71.830 150.015 ;
        RECT 72.000 149.365 72.330 149.845 ;
        RECT 71.105 149.195 72.330 149.365 ;
        RECT 72.520 149.215 72.770 150.015 ;
        RECT 72.940 149.215 73.280 149.845 ;
        RECT 73.450 149.290 73.740 150.015 ;
        RECT 70.645 148.825 70.975 149.025 ;
        RECT 71.145 148.825 71.475 149.025 ;
        RECT 71.645 148.825 72.065 149.025 ;
        RECT 72.240 148.855 72.935 149.025 ;
        RECT 72.240 148.605 72.410 148.855 ;
        RECT 73.105 148.655 73.280 149.215 ;
        RECT 73.050 148.605 73.280 148.655 ;
        RECT 73.910 149.215 74.250 149.845 ;
        RECT 74.420 149.215 74.670 150.015 ;
        RECT 74.860 149.365 75.190 149.845 ;
        RECT 75.360 149.555 75.585 150.015 ;
        RECT 75.755 149.365 76.085 149.845 ;
        RECT 69.975 148.435 72.410 148.605 ;
        RECT 69.975 147.635 70.305 148.435 ;
        RECT 70.475 147.465 70.805 148.265 ;
        RECT 71.105 147.635 71.435 148.435 ;
        RECT 72.080 147.465 72.330 148.265 ;
        RECT 72.600 147.465 72.770 148.605 ;
        RECT 72.940 147.635 73.280 148.605 ;
        RECT 73.450 147.465 73.740 148.630 ;
        RECT 73.910 148.605 74.085 149.215 ;
        RECT 74.860 149.195 76.085 149.365 ;
        RECT 76.715 149.235 77.215 149.845 ;
        RECT 78.510 149.245 82.020 150.015 ;
        RECT 74.255 148.855 74.950 149.025 ;
        RECT 74.780 148.605 74.950 148.855 ;
        RECT 75.125 148.825 75.545 149.025 ;
        RECT 75.715 148.825 76.045 149.025 ;
        RECT 76.215 148.825 76.545 149.025 ;
        RECT 76.715 148.605 76.885 149.235 ;
        RECT 77.070 148.775 77.420 149.025 ;
        RECT 73.910 147.635 74.250 148.605 ;
        RECT 74.420 147.465 74.590 148.605 ;
        RECT 74.780 148.435 77.215 148.605 ;
        RECT 74.860 147.465 75.110 148.265 ;
        RECT 75.755 147.635 76.085 148.435 ;
        RECT 76.385 147.465 76.715 148.265 ;
        RECT 76.885 147.635 77.215 148.435 ;
        RECT 78.510 148.555 80.200 149.075 ;
        RECT 80.370 148.725 82.020 149.245 ;
        RECT 82.195 149.305 82.450 149.835 ;
        RECT 82.620 149.555 82.925 150.015 ;
        RECT 83.170 149.635 84.240 149.805 ;
        RECT 82.195 148.655 82.405 149.305 ;
        RECT 83.170 149.280 83.490 149.635 ;
        RECT 83.165 149.105 83.490 149.280 ;
        RECT 82.575 148.805 83.490 149.105 ;
        RECT 83.660 149.065 83.900 149.465 ;
        RECT 84.070 149.405 84.240 149.635 ;
        RECT 84.410 149.575 84.600 150.015 ;
        RECT 84.770 149.565 85.720 149.845 ;
        RECT 85.940 149.655 86.290 149.825 ;
        RECT 84.070 149.235 84.600 149.405 ;
        RECT 82.575 148.775 83.315 148.805 ;
        RECT 78.510 147.465 82.020 148.555 ;
        RECT 82.195 147.775 82.450 148.655 ;
        RECT 82.620 147.465 82.925 148.605 ;
        RECT 83.145 148.185 83.315 148.775 ;
        RECT 83.660 148.695 84.200 149.065 ;
        RECT 84.380 148.955 84.600 149.235 ;
        RECT 84.770 148.785 84.940 149.565 ;
        RECT 84.535 148.615 84.940 148.785 ;
        RECT 85.110 148.775 85.460 149.395 ;
        RECT 84.535 148.525 84.705 148.615 ;
        RECT 85.630 148.605 85.840 149.395 ;
        RECT 83.485 148.355 84.705 148.525 ;
        RECT 85.165 148.445 85.840 148.605 ;
        RECT 83.145 148.015 83.945 148.185 ;
        RECT 83.265 147.465 83.595 147.845 ;
        RECT 83.775 147.725 83.945 148.015 ;
        RECT 84.535 147.975 84.705 148.355 ;
        RECT 84.875 148.435 85.840 148.445 ;
        RECT 86.030 149.265 86.290 149.655 ;
        RECT 86.500 149.555 86.830 150.015 ;
        RECT 87.705 149.625 88.560 149.795 ;
        RECT 88.765 149.625 89.260 149.795 ;
        RECT 89.430 149.655 89.760 150.015 ;
        RECT 86.030 148.575 86.200 149.265 ;
        RECT 86.370 148.915 86.540 149.095 ;
        RECT 86.710 149.085 87.500 149.335 ;
        RECT 87.705 148.915 87.875 149.625 ;
        RECT 88.045 149.115 88.400 149.335 ;
        RECT 86.370 148.745 88.060 148.915 ;
        RECT 84.875 148.145 85.335 148.435 ;
        RECT 86.030 148.405 87.530 148.575 ;
        RECT 86.030 148.265 86.200 148.405 ;
        RECT 85.640 148.095 86.200 148.265 ;
        RECT 84.115 147.465 84.365 147.925 ;
        RECT 84.535 147.635 85.405 147.975 ;
        RECT 85.640 147.635 85.810 148.095 ;
        RECT 86.645 148.065 87.720 148.235 ;
        RECT 85.980 147.465 86.350 147.925 ;
        RECT 86.645 147.725 86.815 148.065 ;
        RECT 86.985 147.465 87.315 147.895 ;
        RECT 87.550 147.725 87.720 148.065 ;
        RECT 87.890 147.965 88.060 148.745 ;
        RECT 88.230 148.525 88.400 149.115 ;
        RECT 88.570 148.715 88.920 149.335 ;
        RECT 88.230 148.135 88.695 148.525 ;
        RECT 89.090 148.265 89.260 149.625 ;
        RECT 89.430 148.435 89.890 149.485 ;
        RECT 88.865 148.095 89.260 148.265 ;
        RECT 88.865 147.965 89.035 148.095 ;
        RECT 87.890 147.635 88.570 147.965 ;
        RECT 88.785 147.635 89.035 147.965 ;
        RECT 89.205 147.465 89.455 147.925 ;
        RECT 89.625 147.650 89.950 148.435 ;
        RECT 90.120 147.635 90.290 149.755 ;
        RECT 90.460 149.635 90.790 150.015 ;
        RECT 90.960 149.465 91.215 149.755 ;
        RECT 90.465 149.295 91.215 149.465 ;
        RECT 90.465 148.305 90.695 149.295 ;
        RECT 91.595 149.235 92.095 149.845 ;
        RECT 90.865 148.475 91.215 149.125 ;
        RECT 91.390 148.775 91.740 149.025 ;
        RECT 91.925 148.605 92.095 149.235 ;
        RECT 92.725 149.365 93.055 149.845 ;
        RECT 93.225 149.555 93.450 150.015 ;
        RECT 93.620 149.365 93.950 149.845 ;
        RECT 92.725 149.195 93.950 149.365 ;
        RECT 94.140 149.215 94.390 150.015 ;
        RECT 94.560 149.215 94.900 149.845 ;
        RECT 92.265 148.825 92.595 149.025 ;
        RECT 92.765 148.825 93.095 149.025 ;
        RECT 93.265 148.825 93.685 149.025 ;
        RECT 93.860 148.855 94.555 149.025 ;
        RECT 93.860 148.605 94.030 148.855 ;
        RECT 94.725 148.605 94.900 149.215 ;
        RECT 95.345 149.205 95.590 149.810 ;
        RECT 95.810 149.480 96.320 150.015 ;
        RECT 91.595 148.435 94.030 148.605 ;
        RECT 90.465 148.135 91.215 148.305 ;
        RECT 90.460 147.465 90.790 147.965 ;
        RECT 90.960 147.635 91.215 148.135 ;
        RECT 91.595 147.635 91.925 148.435 ;
        RECT 92.095 147.465 92.425 148.265 ;
        RECT 92.725 147.635 93.055 148.435 ;
        RECT 93.700 147.465 93.950 148.265 ;
        RECT 94.220 147.465 94.390 148.605 ;
        RECT 94.560 147.635 94.900 148.605 ;
        RECT 95.070 149.035 96.300 149.205 ;
        RECT 95.070 148.225 95.410 149.035 ;
        RECT 95.580 148.470 96.330 148.660 ;
        RECT 95.070 147.815 95.585 148.225 ;
        RECT 95.820 147.465 95.990 148.225 ;
        RECT 96.160 147.805 96.330 148.470 ;
        RECT 96.500 148.485 96.690 149.845 ;
        RECT 96.860 149.675 97.135 149.845 ;
        RECT 96.860 149.505 97.140 149.675 ;
        RECT 96.860 148.685 97.135 149.505 ;
        RECT 97.325 149.480 97.855 149.845 ;
        RECT 98.280 149.615 98.610 150.015 ;
        RECT 97.680 149.445 97.855 149.480 ;
        RECT 97.340 148.485 97.510 149.285 ;
        RECT 96.500 148.315 97.510 148.485 ;
        RECT 97.680 149.275 98.610 149.445 ;
        RECT 98.780 149.275 99.035 149.845 ;
        RECT 99.210 149.290 99.500 150.015 ;
        RECT 97.680 148.145 97.850 149.275 ;
        RECT 98.440 149.105 98.610 149.275 ;
        RECT 96.725 147.975 97.850 148.145 ;
        RECT 98.020 148.775 98.215 149.105 ;
        RECT 98.440 148.775 98.695 149.105 ;
        RECT 98.020 147.805 98.190 148.775 ;
        RECT 98.865 148.605 99.035 149.275 ;
        RECT 99.670 149.245 101.340 150.015 ;
        RECT 96.160 147.635 98.190 147.805 ;
        RECT 98.360 147.465 98.530 148.605 ;
        RECT 98.700 147.635 99.035 148.605 ;
        RECT 99.210 147.465 99.500 148.630 ;
        RECT 99.670 148.555 100.420 149.075 ;
        RECT 100.590 148.725 101.340 149.245 ;
        RECT 101.885 149.305 102.140 149.835 ;
        RECT 102.320 149.555 102.605 150.015 ;
        RECT 99.670 147.465 101.340 148.555 ;
        RECT 101.885 148.445 102.065 149.305 ;
        RECT 102.785 149.105 103.035 149.755 ;
        RECT 102.235 148.775 103.035 149.105 ;
        RECT 101.885 147.975 102.140 148.445 ;
        RECT 101.800 147.805 102.140 147.975 ;
        RECT 101.885 147.775 102.140 147.805 ;
        RECT 102.320 147.465 102.605 148.265 ;
        RECT 102.785 148.185 103.035 148.775 ;
        RECT 103.235 149.420 103.555 149.750 ;
        RECT 103.735 149.535 104.395 150.015 ;
        RECT 104.595 149.625 105.445 149.795 ;
        RECT 103.235 148.525 103.425 149.420 ;
        RECT 103.745 149.095 104.405 149.365 ;
        RECT 104.075 149.035 104.405 149.095 ;
        RECT 103.595 148.865 103.925 148.925 ;
        RECT 104.595 148.865 104.765 149.625 ;
        RECT 106.005 149.555 106.325 150.015 ;
        RECT 106.525 149.375 106.775 149.805 ;
        RECT 107.065 149.575 107.475 150.015 ;
        RECT 107.645 149.635 108.660 149.835 ;
        RECT 104.935 149.205 106.185 149.375 ;
        RECT 104.935 149.085 105.265 149.205 ;
        RECT 103.595 148.695 105.495 148.865 ;
        RECT 103.235 148.355 105.155 148.525 ;
        RECT 103.235 148.335 103.555 148.355 ;
        RECT 102.785 147.675 103.115 148.185 ;
        RECT 103.385 147.725 103.555 148.335 ;
        RECT 105.325 148.185 105.495 148.695 ;
        RECT 105.665 148.625 105.845 149.035 ;
        RECT 106.015 148.445 106.185 149.205 ;
        RECT 103.725 147.465 104.055 148.155 ;
        RECT 104.285 148.015 105.495 148.185 ;
        RECT 105.665 148.135 106.185 148.445 ;
        RECT 106.355 149.035 106.775 149.375 ;
        RECT 107.065 149.035 107.475 149.365 ;
        RECT 106.355 148.265 106.545 149.035 ;
        RECT 107.645 148.905 107.815 149.635 ;
        RECT 108.960 149.465 109.130 149.795 ;
        RECT 109.300 149.635 109.630 150.015 ;
        RECT 107.985 149.085 108.335 149.455 ;
        RECT 107.645 148.865 108.065 148.905 ;
        RECT 106.715 148.695 108.065 148.865 ;
        RECT 106.715 148.535 106.965 148.695 ;
        RECT 107.475 148.265 107.725 148.525 ;
        RECT 106.355 148.015 107.725 148.265 ;
        RECT 104.285 147.725 104.525 148.015 ;
        RECT 105.325 147.935 105.495 148.015 ;
        RECT 104.725 147.465 105.145 147.845 ;
        RECT 105.325 147.685 105.955 147.935 ;
        RECT 106.425 147.465 106.755 147.845 ;
        RECT 106.925 147.725 107.095 148.015 ;
        RECT 107.895 147.850 108.065 148.695 ;
        RECT 108.515 148.525 108.735 149.395 ;
        RECT 108.960 149.275 109.655 149.465 ;
        RECT 108.235 148.145 108.735 148.525 ;
        RECT 108.905 148.475 109.315 149.095 ;
        RECT 109.485 148.305 109.655 149.275 ;
        RECT 108.960 148.135 109.655 148.305 ;
        RECT 107.275 147.465 107.655 147.845 ;
        RECT 107.895 147.680 108.725 147.850 ;
        RECT 108.960 147.635 109.130 148.135 ;
        RECT 109.300 147.465 109.630 147.965 ;
        RECT 109.845 147.635 110.070 149.755 ;
        RECT 110.240 149.635 110.570 150.015 ;
        RECT 110.740 149.465 110.910 149.755 ;
        RECT 110.245 149.295 110.910 149.465 ;
        RECT 110.245 148.305 110.475 149.295 ;
        RECT 111.170 149.265 112.380 150.015 ;
        RECT 110.645 148.475 110.995 149.125 ;
        RECT 111.170 148.555 111.690 149.095 ;
        RECT 111.860 148.725 112.380 149.265 ;
        RECT 110.245 148.135 110.910 148.305 ;
        RECT 110.240 147.465 110.570 147.965 ;
        RECT 110.740 147.635 110.910 148.135 ;
        RECT 111.170 147.465 112.380 148.555 ;
        RECT 18.165 147.295 112.465 147.465 ;
        RECT 18.250 146.205 19.460 147.295 ;
        RECT 18.250 145.495 18.770 146.035 ;
        RECT 18.940 145.665 19.460 146.205 ;
        RECT 19.635 146.105 19.890 146.985 ;
        RECT 20.060 146.155 20.365 147.295 ;
        RECT 20.705 146.915 21.035 147.295 ;
        RECT 21.215 146.745 21.385 147.035 ;
        RECT 21.555 146.835 21.805 147.295 ;
        RECT 20.585 146.575 21.385 146.745 ;
        RECT 21.975 146.785 22.845 147.125 ;
        RECT 18.250 144.745 19.460 145.495 ;
        RECT 19.635 145.455 19.845 146.105 ;
        RECT 20.585 145.985 20.755 146.575 ;
        RECT 21.975 146.405 22.145 146.785 ;
        RECT 23.080 146.665 23.250 147.125 ;
        RECT 23.420 146.835 23.790 147.295 ;
        RECT 24.085 146.695 24.255 147.035 ;
        RECT 24.425 146.865 24.755 147.295 ;
        RECT 24.990 146.695 25.160 147.035 ;
        RECT 20.925 146.235 22.145 146.405 ;
        RECT 22.315 146.325 22.775 146.615 ;
        RECT 23.080 146.495 23.640 146.665 ;
        RECT 24.085 146.525 25.160 146.695 ;
        RECT 25.330 146.795 26.010 147.125 ;
        RECT 26.225 146.795 26.475 147.125 ;
        RECT 26.645 146.835 26.895 147.295 ;
        RECT 23.470 146.355 23.640 146.495 ;
        RECT 22.315 146.315 23.280 146.325 ;
        RECT 21.975 146.145 22.145 146.235 ;
        RECT 22.605 146.155 23.280 146.315 ;
        RECT 20.015 145.955 20.755 145.985 ;
        RECT 20.015 145.655 20.930 145.955 ;
        RECT 20.605 145.480 20.930 145.655 ;
        RECT 19.635 144.925 19.890 145.455 ;
        RECT 20.060 144.745 20.365 145.205 ;
        RECT 20.610 145.125 20.930 145.480 ;
        RECT 21.100 145.695 21.640 146.065 ;
        RECT 21.975 145.975 22.380 146.145 ;
        RECT 21.100 145.295 21.340 145.695 ;
        RECT 21.820 145.525 22.040 145.805 ;
        RECT 21.510 145.355 22.040 145.525 ;
        RECT 21.510 145.125 21.680 145.355 ;
        RECT 22.210 145.195 22.380 145.975 ;
        RECT 22.550 145.365 22.900 145.985 ;
        RECT 23.070 145.365 23.280 146.155 ;
        RECT 23.470 146.185 24.970 146.355 ;
        RECT 23.470 145.495 23.640 146.185 ;
        RECT 25.330 146.015 25.500 146.795 ;
        RECT 26.305 146.665 26.475 146.795 ;
        RECT 23.810 145.845 25.500 146.015 ;
        RECT 25.670 146.235 26.135 146.625 ;
        RECT 26.305 146.495 26.700 146.665 ;
        RECT 23.810 145.665 23.980 145.845 ;
        RECT 20.610 144.955 21.680 145.125 ;
        RECT 21.850 144.745 22.040 145.185 ;
        RECT 22.210 144.915 23.160 145.195 ;
        RECT 23.470 145.105 23.730 145.495 ;
        RECT 24.150 145.425 24.940 145.675 ;
        RECT 23.380 144.935 23.730 145.105 ;
        RECT 23.940 144.745 24.270 145.205 ;
        RECT 25.145 145.135 25.315 145.845 ;
        RECT 25.670 145.645 25.840 146.235 ;
        RECT 25.485 145.425 25.840 145.645 ;
        RECT 26.010 145.425 26.360 146.045 ;
        RECT 26.530 145.135 26.700 146.495 ;
        RECT 27.065 146.325 27.390 147.110 ;
        RECT 26.870 145.275 27.330 146.325 ;
        RECT 25.145 144.965 26.000 145.135 ;
        RECT 26.205 144.965 26.700 145.135 ;
        RECT 26.870 144.745 27.200 145.105 ;
        RECT 27.560 145.005 27.730 147.125 ;
        RECT 27.900 146.795 28.230 147.295 ;
        RECT 28.400 146.625 28.655 147.125 ;
        RECT 27.905 146.455 28.655 146.625 ;
        RECT 27.905 145.465 28.135 146.455 ;
        RECT 28.920 146.365 29.090 147.125 ;
        RECT 29.270 146.535 29.600 147.295 ;
        RECT 28.305 145.635 28.655 146.285 ;
        RECT 28.920 146.195 29.585 146.365 ;
        RECT 29.770 146.220 30.040 147.125 ;
        RECT 29.415 146.050 29.585 146.195 ;
        RECT 28.850 145.645 29.180 146.015 ;
        RECT 29.415 145.720 29.700 146.050 ;
        RECT 29.415 145.465 29.585 145.720 ;
        RECT 27.905 145.295 28.655 145.465 ;
        RECT 27.900 144.745 28.230 145.125 ;
        RECT 28.400 145.005 28.655 145.295 ;
        RECT 28.920 145.295 29.585 145.465 ;
        RECT 29.870 145.420 30.040 146.220 ;
        RECT 31.335 146.325 31.665 147.125 ;
        RECT 31.835 146.495 32.165 147.295 ;
        RECT 32.465 146.325 32.795 147.125 ;
        RECT 33.440 146.495 33.690 147.295 ;
        RECT 31.335 146.155 33.770 146.325 ;
        RECT 33.960 146.155 34.130 147.295 ;
        RECT 34.300 146.155 34.640 147.125 ;
        RECT 31.130 145.735 31.480 145.985 ;
        RECT 31.665 145.525 31.835 146.155 ;
        RECT 32.005 145.735 32.335 145.935 ;
        RECT 32.505 145.735 32.835 145.935 ;
        RECT 33.005 145.735 33.425 145.935 ;
        RECT 33.600 145.905 33.770 146.155 ;
        RECT 33.600 145.735 34.295 145.905 ;
        RECT 34.465 145.595 34.640 146.155 ;
        RECT 34.810 146.130 35.100 147.295 ;
        RECT 35.270 146.155 35.610 147.125 ;
        RECT 35.780 146.155 35.950 147.295 ;
        RECT 36.220 146.495 36.470 147.295 ;
        RECT 37.115 146.325 37.445 147.125 ;
        RECT 37.745 146.495 38.075 147.295 ;
        RECT 38.245 146.325 38.575 147.125 ;
        RECT 36.140 146.155 38.575 146.325 ;
        RECT 39.785 146.315 40.040 146.985 ;
        RECT 40.220 146.495 40.505 147.295 ;
        RECT 40.685 146.575 41.015 147.085 ;
        RECT 39.785 146.275 39.965 146.315 ;
        RECT 28.920 144.915 29.090 145.295 ;
        RECT 29.270 144.745 29.600 145.125 ;
        RECT 29.780 144.915 30.040 145.420 ;
        RECT 31.335 144.915 31.835 145.525 ;
        RECT 32.465 145.395 33.690 145.565 ;
        RECT 34.410 145.545 34.640 145.595 ;
        RECT 32.465 144.915 32.795 145.395 ;
        RECT 32.965 144.745 33.190 145.205 ;
        RECT 33.360 144.915 33.690 145.395 ;
        RECT 33.880 144.745 34.130 145.545 ;
        RECT 34.300 144.915 34.640 145.545 ;
        RECT 35.270 145.545 35.445 146.155 ;
        RECT 36.140 145.905 36.310 146.155 ;
        RECT 35.615 145.735 36.310 145.905 ;
        RECT 36.485 145.735 36.905 145.935 ;
        RECT 37.075 145.735 37.405 145.935 ;
        RECT 37.575 145.735 37.905 145.935 ;
        RECT 34.810 144.745 35.100 145.470 ;
        RECT 35.270 144.915 35.610 145.545 ;
        RECT 35.780 144.745 36.030 145.545 ;
        RECT 36.220 145.395 37.445 145.565 ;
        RECT 36.220 144.915 36.550 145.395 ;
        RECT 36.720 144.745 36.945 145.205 ;
        RECT 37.115 144.915 37.445 145.395 ;
        RECT 38.075 145.525 38.245 146.155 ;
        RECT 39.700 146.105 39.965 146.275 ;
        RECT 38.430 145.735 38.780 145.985 ;
        RECT 38.075 144.915 38.575 145.525 ;
        RECT 39.785 145.455 39.965 146.105 ;
        RECT 40.685 145.985 40.935 146.575 ;
        RECT 41.285 146.425 41.455 147.035 ;
        RECT 41.625 146.605 41.955 147.295 ;
        RECT 42.185 146.745 42.425 147.035 ;
        RECT 42.625 146.915 43.045 147.295 ;
        RECT 43.225 146.825 43.855 147.075 ;
        RECT 44.325 146.915 44.655 147.295 ;
        RECT 43.225 146.745 43.395 146.825 ;
        RECT 44.825 146.745 44.995 147.035 ;
        RECT 45.175 146.915 45.555 147.295 ;
        RECT 45.795 146.910 46.625 147.080 ;
        RECT 42.185 146.575 43.395 146.745 ;
        RECT 40.135 145.655 40.935 145.985 ;
        RECT 39.785 144.925 40.040 145.455 ;
        RECT 40.220 144.745 40.505 145.205 ;
        RECT 40.685 145.005 40.935 145.655 ;
        RECT 41.135 146.405 41.455 146.425 ;
        RECT 41.135 146.235 43.055 146.405 ;
        RECT 41.135 145.340 41.325 146.235 ;
        RECT 43.225 146.065 43.395 146.575 ;
        RECT 43.565 146.315 44.085 146.625 ;
        RECT 41.495 145.895 43.395 146.065 ;
        RECT 41.495 145.835 41.825 145.895 ;
        RECT 41.975 145.665 42.305 145.725 ;
        RECT 41.645 145.395 42.305 145.665 ;
        RECT 41.135 145.010 41.455 145.340 ;
        RECT 41.635 144.745 42.295 145.225 ;
        RECT 42.495 145.135 42.665 145.895 ;
        RECT 43.565 145.725 43.745 146.135 ;
        RECT 42.835 145.555 43.165 145.675 ;
        RECT 43.915 145.555 44.085 146.315 ;
        RECT 42.835 145.385 44.085 145.555 ;
        RECT 44.255 146.495 45.625 146.745 ;
        RECT 44.255 145.725 44.445 146.495 ;
        RECT 45.375 146.235 45.625 146.495 ;
        RECT 44.615 146.065 44.865 146.225 ;
        RECT 45.795 146.065 45.965 146.910 ;
        RECT 46.860 146.625 47.030 147.125 ;
        RECT 47.200 146.795 47.530 147.295 ;
        RECT 46.135 146.235 46.635 146.615 ;
        RECT 46.860 146.455 47.555 146.625 ;
        RECT 44.615 145.895 45.965 146.065 ;
        RECT 45.545 145.855 45.965 145.895 ;
        RECT 44.255 145.385 44.675 145.725 ;
        RECT 44.965 145.395 45.375 145.725 ;
        RECT 42.495 144.965 43.345 145.135 ;
        RECT 43.905 144.745 44.225 145.205 ;
        RECT 44.425 144.955 44.675 145.385 ;
        RECT 44.965 144.745 45.375 145.185 ;
        RECT 45.545 145.125 45.715 145.855 ;
        RECT 45.885 145.305 46.235 145.675 ;
        RECT 46.415 145.365 46.635 146.235 ;
        RECT 46.805 145.665 47.215 146.285 ;
        RECT 47.385 145.485 47.555 146.455 ;
        RECT 46.860 145.295 47.555 145.485 ;
        RECT 45.545 144.925 46.560 145.125 ;
        RECT 46.860 144.965 47.030 145.295 ;
        RECT 47.200 144.745 47.530 145.125 ;
        RECT 47.745 145.005 47.970 147.125 ;
        RECT 48.140 146.795 48.470 147.295 ;
        RECT 48.640 146.625 48.810 147.125 ;
        RECT 48.145 146.455 48.810 146.625 ;
        RECT 48.145 145.465 48.375 146.455 ;
        RECT 48.545 145.635 48.895 146.285 ;
        RECT 49.070 146.220 49.340 147.125 ;
        RECT 49.510 146.535 49.840 147.295 ;
        RECT 50.020 146.365 50.190 147.125 ;
        RECT 48.145 145.295 48.810 145.465 ;
        RECT 48.140 144.745 48.470 145.125 ;
        RECT 48.640 145.005 48.810 145.295 ;
        RECT 49.070 145.420 49.240 146.220 ;
        RECT 49.525 146.195 50.190 146.365 ;
        RECT 49.525 146.050 49.695 146.195 ;
        RECT 50.950 146.155 51.180 147.295 ;
        RECT 51.350 146.145 51.680 147.125 ;
        RECT 51.850 146.155 52.060 147.295 ;
        RECT 52.750 146.155 53.090 147.125 ;
        RECT 53.260 146.155 53.430 147.295 ;
        RECT 53.700 146.495 53.950 147.295 ;
        RECT 54.595 146.325 54.925 147.125 ;
        RECT 55.225 146.495 55.555 147.295 ;
        RECT 55.725 146.325 56.055 147.125 ;
        RECT 53.620 146.155 56.055 146.325 ;
        RECT 56.430 146.535 56.945 146.945 ;
        RECT 57.180 146.535 57.350 147.295 ;
        RECT 57.520 146.955 59.550 147.125 ;
        RECT 49.410 145.720 49.695 146.050 ;
        RECT 49.525 145.465 49.695 145.720 ;
        RECT 49.930 145.645 50.260 146.015 ;
        RECT 50.930 145.735 51.260 145.985 ;
        RECT 49.070 144.915 49.330 145.420 ;
        RECT 49.525 145.295 50.190 145.465 ;
        RECT 49.510 144.745 49.840 145.125 ;
        RECT 50.020 144.915 50.190 145.295 ;
        RECT 50.950 144.745 51.180 145.565 ;
        RECT 51.430 145.545 51.680 146.145 ;
        RECT 51.350 144.915 51.680 145.545 ;
        RECT 51.850 144.745 52.060 145.565 ;
        RECT 52.750 145.545 52.925 146.155 ;
        RECT 53.620 145.905 53.790 146.155 ;
        RECT 53.095 145.735 53.790 145.905 ;
        RECT 53.965 145.735 54.385 145.935 ;
        RECT 54.555 145.735 54.885 145.935 ;
        RECT 55.055 145.735 55.385 145.935 ;
        RECT 52.750 144.915 53.090 145.545 ;
        RECT 53.260 144.745 53.510 145.545 ;
        RECT 53.700 145.395 54.925 145.565 ;
        RECT 53.700 144.915 54.030 145.395 ;
        RECT 54.200 144.745 54.425 145.205 ;
        RECT 54.595 144.915 54.925 145.395 ;
        RECT 55.555 145.525 55.725 146.155 ;
        RECT 55.910 145.735 56.260 145.985 ;
        RECT 56.430 145.725 56.770 146.535 ;
        RECT 57.520 146.290 57.690 146.955 ;
        RECT 58.085 146.615 59.210 146.785 ;
        RECT 56.940 146.100 57.690 146.290 ;
        RECT 57.860 146.275 58.870 146.445 ;
        RECT 56.430 145.555 57.660 145.725 ;
        RECT 55.555 144.915 56.055 145.525 ;
        RECT 56.705 144.950 56.950 145.555 ;
        RECT 57.170 144.745 57.680 145.280 ;
        RECT 57.860 144.915 58.050 146.275 ;
        RECT 58.220 145.255 58.495 146.075 ;
        RECT 58.700 145.475 58.870 146.275 ;
        RECT 59.040 145.485 59.210 146.615 ;
        RECT 59.380 145.985 59.550 146.955 ;
        RECT 59.720 146.155 59.890 147.295 ;
        RECT 60.060 146.155 60.395 147.125 ;
        RECT 59.380 145.655 59.575 145.985 ;
        RECT 59.800 145.655 60.055 145.985 ;
        RECT 59.800 145.485 59.970 145.655 ;
        RECT 60.225 145.485 60.395 146.155 ;
        RECT 60.570 146.130 60.860 147.295 ;
        RECT 61.490 146.205 63.160 147.295 ;
        RECT 63.420 146.365 63.590 147.125 ;
        RECT 63.805 146.535 64.135 147.295 ;
        RECT 61.490 145.685 62.240 146.205 ;
        RECT 63.420 146.195 64.135 146.365 ;
        RECT 64.305 146.220 64.560 147.125 ;
        RECT 62.410 145.515 63.160 146.035 ;
        RECT 63.330 145.645 63.685 146.015 ;
        RECT 63.965 145.985 64.135 146.195 ;
        RECT 63.965 145.655 64.220 145.985 ;
        RECT 59.040 145.315 59.970 145.485 ;
        RECT 59.040 145.280 59.215 145.315 ;
        RECT 58.220 145.085 58.500 145.255 ;
        RECT 58.220 144.915 58.495 145.085 ;
        RECT 58.685 144.915 59.215 145.280 ;
        RECT 59.640 144.745 59.970 145.145 ;
        RECT 60.140 144.915 60.395 145.485 ;
        RECT 60.570 144.745 60.860 145.470 ;
        RECT 61.490 144.745 63.160 145.515 ;
        RECT 63.965 145.465 64.135 145.655 ;
        RECT 64.390 145.490 64.560 146.220 ;
        RECT 64.735 146.145 64.995 147.295 ;
        RECT 65.230 146.155 65.440 147.295 ;
        RECT 65.610 146.145 65.940 147.125 ;
        RECT 66.110 146.155 66.340 147.295 ;
        RECT 66.640 146.365 66.810 147.125 ;
        RECT 66.990 146.535 67.320 147.295 ;
        RECT 66.640 146.195 67.305 146.365 ;
        RECT 67.490 146.220 67.760 147.125 ;
        RECT 63.420 145.295 64.135 145.465 ;
        RECT 63.420 144.915 63.590 145.295 ;
        RECT 63.805 144.745 64.135 145.125 ;
        RECT 64.305 144.915 64.560 145.490 ;
        RECT 64.735 144.745 64.995 145.585 ;
        RECT 65.230 144.745 65.440 145.565 ;
        RECT 65.610 145.545 65.860 146.145 ;
        RECT 67.135 146.050 67.305 146.195 ;
        RECT 66.030 145.735 66.360 145.985 ;
        RECT 66.570 145.645 66.900 146.015 ;
        RECT 67.135 145.720 67.420 146.050 ;
        RECT 65.610 144.915 65.940 145.545 ;
        RECT 66.110 144.745 66.340 145.565 ;
        RECT 67.135 145.465 67.305 145.720 ;
        RECT 66.640 145.295 67.305 145.465 ;
        RECT 67.590 145.420 67.760 146.220 ;
        RECT 68.390 146.205 70.060 147.295 ;
        RECT 68.390 145.685 69.140 146.205 ;
        RECT 70.230 146.155 70.500 147.125 ;
        RECT 70.710 146.495 70.990 147.295 ;
        RECT 71.160 146.785 72.815 147.075 ;
        RECT 71.225 146.445 72.815 146.615 ;
        RECT 71.225 146.325 71.395 146.445 ;
        RECT 70.670 146.155 71.395 146.325 ;
        RECT 69.310 145.515 70.060 146.035 ;
        RECT 66.640 144.915 66.810 145.295 ;
        RECT 66.990 144.745 67.320 145.125 ;
        RECT 67.500 144.915 67.760 145.420 ;
        RECT 68.390 144.745 70.060 145.515 ;
        RECT 70.230 145.420 70.400 146.155 ;
        RECT 70.670 145.985 70.840 146.155 ;
        RECT 71.585 146.105 72.300 146.275 ;
        RECT 72.495 146.155 72.815 146.445 ;
        RECT 72.990 146.155 73.330 147.125 ;
        RECT 73.500 146.155 73.670 147.295 ;
        RECT 73.940 146.495 74.190 147.295 ;
        RECT 74.835 146.325 75.165 147.125 ;
        RECT 75.465 146.495 75.795 147.295 ;
        RECT 75.965 146.325 76.295 147.125 ;
        RECT 77.045 146.955 77.300 146.985 ;
        RECT 76.960 146.785 77.300 146.955 ;
        RECT 73.860 146.155 76.295 146.325 ;
        RECT 77.045 146.315 77.300 146.785 ;
        RECT 77.480 146.495 77.765 147.295 ;
        RECT 77.945 146.575 78.275 147.085 ;
        RECT 70.570 145.655 70.840 145.985 ;
        RECT 71.010 145.655 71.415 145.985 ;
        RECT 71.585 145.655 72.295 146.105 ;
        RECT 70.670 145.485 70.840 145.655 ;
        RECT 70.230 145.075 70.500 145.420 ;
        RECT 70.670 145.315 72.280 145.485 ;
        RECT 72.465 145.415 72.815 145.985 ;
        RECT 72.990 145.595 73.165 146.155 ;
        RECT 73.860 145.905 74.030 146.155 ;
        RECT 73.335 145.735 74.030 145.905 ;
        RECT 74.205 145.735 74.625 145.935 ;
        RECT 74.795 145.735 75.125 145.935 ;
        RECT 75.295 145.735 75.625 145.935 ;
        RECT 72.990 145.545 73.220 145.595 ;
        RECT 70.690 144.745 71.070 145.145 ;
        RECT 71.240 144.965 71.410 145.315 ;
        RECT 71.580 144.745 71.910 145.145 ;
        RECT 72.110 144.965 72.280 145.315 ;
        RECT 72.480 144.745 72.810 145.245 ;
        RECT 72.990 144.915 73.330 145.545 ;
        RECT 73.500 144.745 73.750 145.545 ;
        RECT 73.940 145.395 75.165 145.565 ;
        RECT 73.940 144.915 74.270 145.395 ;
        RECT 74.440 144.745 74.665 145.205 ;
        RECT 74.835 144.915 75.165 145.395 ;
        RECT 75.795 145.525 75.965 146.155 ;
        RECT 76.150 145.735 76.500 145.985 ;
        RECT 75.795 144.915 76.295 145.525 ;
        RECT 77.045 145.455 77.225 146.315 ;
        RECT 77.945 145.985 78.195 146.575 ;
        RECT 78.545 146.425 78.715 147.035 ;
        RECT 78.885 146.605 79.215 147.295 ;
        RECT 79.445 146.745 79.685 147.035 ;
        RECT 79.885 146.915 80.305 147.295 ;
        RECT 80.485 146.825 81.115 147.075 ;
        RECT 81.585 146.915 81.915 147.295 ;
        RECT 80.485 146.745 80.655 146.825 ;
        RECT 82.085 146.745 82.255 147.035 ;
        RECT 82.435 146.915 82.815 147.295 ;
        RECT 83.055 146.910 83.885 147.080 ;
        RECT 79.445 146.575 80.655 146.745 ;
        RECT 77.395 145.655 78.195 145.985 ;
        RECT 77.045 144.925 77.300 145.455 ;
        RECT 77.480 144.745 77.765 145.205 ;
        RECT 77.945 145.005 78.195 145.655 ;
        RECT 78.395 146.405 78.715 146.425 ;
        RECT 78.395 146.235 80.315 146.405 ;
        RECT 78.395 145.340 78.585 146.235 ;
        RECT 80.485 146.065 80.655 146.575 ;
        RECT 80.825 146.315 81.345 146.625 ;
        RECT 78.755 145.895 80.655 146.065 ;
        RECT 78.755 145.835 79.085 145.895 ;
        RECT 79.235 145.665 79.565 145.725 ;
        RECT 78.905 145.395 79.565 145.665 ;
        RECT 78.395 145.010 78.715 145.340 ;
        RECT 78.895 144.745 79.555 145.225 ;
        RECT 79.755 145.135 79.925 145.895 ;
        RECT 80.825 145.725 81.005 146.135 ;
        RECT 80.095 145.555 80.425 145.675 ;
        RECT 81.175 145.555 81.345 146.315 ;
        RECT 80.095 145.385 81.345 145.555 ;
        RECT 81.515 146.495 82.885 146.745 ;
        RECT 81.515 145.725 81.705 146.495 ;
        RECT 82.635 146.235 82.885 146.495 ;
        RECT 81.875 146.065 82.125 146.225 ;
        RECT 83.055 146.065 83.225 146.910 ;
        RECT 84.120 146.625 84.290 147.125 ;
        RECT 84.460 146.795 84.790 147.295 ;
        RECT 83.395 146.235 83.895 146.615 ;
        RECT 84.120 146.455 84.815 146.625 ;
        RECT 81.875 145.895 83.225 146.065 ;
        RECT 82.805 145.855 83.225 145.895 ;
        RECT 81.515 145.385 81.935 145.725 ;
        RECT 82.225 145.395 82.635 145.725 ;
        RECT 79.755 144.965 80.605 145.135 ;
        RECT 81.165 144.745 81.485 145.205 ;
        RECT 81.685 144.955 81.935 145.385 ;
        RECT 82.225 144.745 82.635 145.185 ;
        RECT 82.805 145.125 82.975 145.855 ;
        RECT 83.145 145.305 83.495 145.675 ;
        RECT 83.675 145.365 83.895 146.235 ;
        RECT 84.065 145.665 84.475 146.285 ;
        RECT 84.645 145.485 84.815 146.455 ;
        RECT 84.120 145.295 84.815 145.485 ;
        RECT 82.805 144.925 83.820 145.125 ;
        RECT 84.120 144.965 84.290 145.295 ;
        RECT 84.460 144.745 84.790 145.125 ;
        RECT 85.005 145.005 85.230 147.125 ;
        RECT 85.400 146.795 85.730 147.295 ;
        RECT 85.900 146.625 86.070 147.125 ;
        RECT 85.405 146.455 86.070 146.625 ;
        RECT 85.405 145.465 85.635 146.455 ;
        RECT 85.805 145.635 86.155 146.285 ;
        RECT 86.330 146.130 86.620 147.295 ;
        RECT 86.850 146.155 87.060 147.295 ;
        RECT 87.230 146.145 87.560 147.125 ;
        RECT 87.730 146.155 87.960 147.295 ;
        RECT 88.170 146.205 91.680 147.295 ;
        RECT 85.405 145.295 86.070 145.465 ;
        RECT 85.400 144.745 85.730 145.125 ;
        RECT 85.900 145.005 86.070 145.295 ;
        RECT 86.330 144.745 86.620 145.470 ;
        RECT 86.850 144.745 87.060 145.565 ;
        RECT 87.230 145.545 87.480 146.145 ;
        RECT 87.650 145.735 87.980 145.985 ;
        RECT 88.170 145.685 89.860 146.205 ;
        RECT 91.850 146.155 92.120 147.125 ;
        RECT 92.330 146.495 92.610 147.295 ;
        RECT 92.780 146.785 94.435 147.075 ;
        RECT 94.615 146.785 96.270 147.075 ;
        RECT 92.845 146.445 94.435 146.615 ;
        RECT 92.845 146.325 93.015 146.445 ;
        RECT 92.290 146.155 93.015 146.325 ;
        RECT 87.230 144.915 87.560 145.545 ;
        RECT 87.730 144.745 87.960 145.565 ;
        RECT 90.030 145.515 91.680 146.035 ;
        RECT 88.170 144.745 91.680 145.515 ;
        RECT 91.850 145.420 92.020 146.155 ;
        RECT 92.290 145.985 92.460 146.155 ;
        RECT 92.190 145.655 92.460 145.985 ;
        RECT 92.630 145.655 93.035 145.985 ;
        RECT 93.205 145.655 93.915 146.275 ;
        RECT 94.115 146.155 94.435 146.445 ;
        RECT 94.615 146.445 96.205 146.615 ;
        RECT 96.440 146.495 96.720 147.295 ;
        RECT 94.615 146.155 94.935 146.445 ;
        RECT 96.035 146.325 96.205 146.445 ;
        RECT 95.130 146.105 95.845 146.275 ;
        RECT 96.035 146.155 96.760 146.325 ;
        RECT 96.930 146.155 97.200 147.125 ;
        RECT 92.290 145.485 92.460 145.655 ;
        RECT 91.850 145.075 92.120 145.420 ;
        RECT 92.290 145.315 93.900 145.485 ;
        RECT 94.085 145.415 94.435 145.985 ;
        RECT 94.615 145.415 94.965 145.985 ;
        RECT 95.135 145.655 95.845 146.105 ;
        RECT 96.590 145.985 96.760 146.155 ;
        RECT 96.015 145.655 96.420 145.985 ;
        RECT 96.590 145.655 96.860 145.985 ;
        RECT 96.590 145.485 96.760 145.655 ;
        RECT 92.310 144.745 92.690 145.145 ;
        RECT 92.860 144.965 93.030 145.315 ;
        RECT 93.200 144.745 93.530 145.145 ;
        RECT 93.730 144.965 93.900 145.315 ;
        RECT 95.150 145.315 96.760 145.485 ;
        RECT 97.030 145.420 97.200 146.155 ;
        RECT 97.830 146.205 100.420 147.295 ;
        RECT 100.590 146.535 101.105 146.945 ;
        RECT 101.340 146.535 101.510 147.295 ;
        RECT 101.680 146.955 103.710 147.125 ;
        RECT 97.830 145.685 99.040 146.205 ;
        RECT 99.210 145.515 100.420 146.035 ;
        RECT 100.590 145.725 100.930 146.535 ;
        RECT 101.680 146.290 101.850 146.955 ;
        RECT 102.245 146.615 103.370 146.785 ;
        RECT 101.100 146.100 101.850 146.290 ;
        RECT 102.020 146.275 103.030 146.445 ;
        RECT 100.590 145.555 101.820 145.725 ;
        RECT 94.100 144.745 94.430 145.245 ;
        RECT 94.620 144.745 94.950 145.245 ;
        RECT 95.150 144.965 95.320 145.315 ;
        RECT 95.520 144.745 95.850 145.145 ;
        RECT 96.020 144.965 96.190 145.315 ;
        RECT 96.360 144.745 96.740 145.145 ;
        RECT 96.930 145.075 97.200 145.420 ;
        RECT 97.830 144.745 100.420 145.515 ;
        RECT 100.865 144.950 101.110 145.555 ;
        RECT 101.330 144.745 101.840 145.280 ;
        RECT 102.020 144.915 102.210 146.275 ;
        RECT 102.380 145.935 102.655 146.075 ;
        RECT 102.380 145.765 102.660 145.935 ;
        RECT 102.380 144.915 102.655 145.765 ;
        RECT 102.860 145.475 103.030 146.275 ;
        RECT 103.200 145.485 103.370 146.615 ;
        RECT 103.540 145.985 103.710 146.955 ;
        RECT 103.880 146.155 104.050 147.295 ;
        RECT 104.220 146.155 104.555 147.125 ;
        RECT 104.770 146.155 105.000 147.295 ;
        RECT 103.540 145.655 103.735 145.985 ;
        RECT 103.960 145.655 104.215 145.985 ;
        RECT 103.960 145.485 104.130 145.655 ;
        RECT 104.385 145.485 104.555 146.155 ;
        RECT 105.170 146.145 105.500 147.125 ;
        RECT 105.670 146.155 105.880 147.295 ;
        RECT 106.660 146.365 106.830 147.125 ;
        RECT 107.010 146.535 107.340 147.295 ;
        RECT 106.660 146.195 107.325 146.365 ;
        RECT 107.510 146.220 107.780 147.125 ;
        RECT 104.750 145.735 105.080 145.985 ;
        RECT 103.200 145.315 104.130 145.485 ;
        RECT 103.200 145.280 103.375 145.315 ;
        RECT 102.845 144.915 103.375 145.280 ;
        RECT 103.800 144.745 104.130 145.145 ;
        RECT 104.300 144.915 104.555 145.485 ;
        RECT 104.770 144.745 105.000 145.565 ;
        RECT 105.250 145.545 105.500 146.145 ;
        RECT 107.155 146.050 107.325 146.195 ;
        RECT 106.590 145.645 106.920 146.015 ;
        RECT 107.155 145.720 107.440 146.050 ;
        RECT 105.170 144.915 105.500 145.545 ;
        RECT 105.670 144.745 105.880 145.565 ;
        RECT 107.155 145.465 107.325 145.720 ;
        RECT 106.660 145.295 107.325 145.465 ;
        RECT 107.610 145.420 107.780 146.220 ;
        RECT 108.410 146.205 111.000 147.295 ;
        RECT 111.170 146.205 112.380 147.295 ;
        RECT 108.410 145.685 109.620 146.205 ;
        RECT 109.790 145.515 111.000 146.035 ;
        RECT 111.170 145.665 111.690 146.205 ;
        RECT 106.660 144.915 106.830 145.295 ;
        RECT 107.010 144.745 107.340 145.125 ;
        RECT 107.520 144.915 107.780 145.420 ;
        RECT 108.410 144.745 111.000 145.515 ;
        RECT 111.860 145.495 112.380 146.035 ;
        RECT 111.170 144.745 112.380 145.495 ;
        RECT 18.165 144.575 112.465 144.745 ;
        RECT 18.250 143.825 19.460 144.575 ;
        RECT 20.640 144.025 20.810 144.405 ;
        RECT 20.990 144.195 21.320 144.575 ;
        RECT 20.640 143.855 21.305 144.025 ;
        RECT 21.500 143.900 21.760 144.405 ;
        RECT 18.250 143.285 18.770 143.825 ;
        RECT 18.940 143.115 19.460 143.655 ;
        RECT 20.570 143.305 20.900 143.675 ;
        RECT 21.135 143.600 21.305 143.855 ;
        RECT 21.135 143.270 21.420 143.600 ;
        RECT 21.135 143.125 21.305 143.270 ;
        RECT 18.250 142.025 19.460 143.115 ;
        RECT 20.640 142.955 21.305 143.125 ;
        RECT 21.590 143.100 21.760 143.900 ;
        RECT 21.930 143.850 22.220 144.575 ;
        RECT 22.395 143.865 22.650 144.395 ;
        RECT 22.820 144.115 23.125 144.575 ;
        RECT 23.370 144.195 24.440 144.365 ;
        RECT 22.395 143.215 22.605 143.865 ;
        RECT 23.370 143.840 23.690 144.195 ;
        RECT 23.365 143.665 23.690 143.840 ;
        RECT 22.775 143.365 23.690 143.665 ;
        RECT 23.860 143.625 24.100 144.025 ;
        RECT 24.270 143.965 24.440 144.195 ;
        RECT 24.610 144.135 24.800 144.575 ;
        RECT 24.970 144.125 25.920 144.405 ;
        RECT 26.140 144.215 26.490 144.385 ;
        RECT 24.270 143.795 24.800 143.965 ;
        RECT 22.775 143.335 23.515 143.365 ;
        RECT 20.640 142.195 20.810 142.955 ;
        RECT 20.990 142.025 21.320 142.785 ;
        RECT 21.490 142.195 21.760 143.100 ;
        RECT 21.930 142.025 22.220 143.190 ;
        RECT 22.395 142.335 22.650 143.215 ;
        RECT 22.820 142.025 23.125 143.165 ;
        RECT 23.345 142.745 23.515 143.335 ;
        RECT 23.860 143.255 24.400 143.625 ;
        RECT 24.580 143.515 24.800 143.795 ;
        RECT 24.970 143.345 25.140 144.125 ;
        RECT 24.735 143.175 25.140 143.345 ;
        RECT 25.310 143.335 25.660 143.955 ;
        RECT 24.735 143.085 24.905 143.175 ;
        RECT 25.830 143.165 26.040 143.955 ;
        RECT 23.685 142.915 24.905 143.085 ;
        RECT 25.365 143.005 26.040 143.165 ;
        RECT 23.345 142.575 24.145 142.745 ;
        RECT 23.465 142.025 23.795 142.405 ;
        RECT 23.975 142.285 24.145 142.575 ;
        RECT 24.735 142.535 24.905 142.915 ;
        RECT 25.075 142.995 26.040 143.005 ;
        RECT 26.230 143.825 26.490 144.215 ;
        RECT 26.700 144.115 27.030 144.575 ;
        RECT 27.905 144.185 28.760 144.355 ;
        RECT 28.965 144.185 29.460 144.355 ;
        RECT 29.630 144.215 29.960 144.575 ;
        RECT 26.230 143.135 26.400 143.825 ;
        RECT 26.570 143.475 26.740 143.655 ;
        RECT 26.910 143.645 27.700 143.895 ;
        RECT 27.905 143.475 28.075 144.185 ;
        RECT 28.245 143.675 28.600 143.895 ;
        RECT 26.570 143.305 28.260 143.475 ;
        RECT 25.075 142.705 25.535 142.995 ;
        RECT 26.230 142.965 27.730 143.135 ;
        RECT 26.230 142.825 26.400 142.965 ;
        RECT 25.840 142.655 26.400 142.825 ;
        RECT 24.315 142.025 24.565 142.485 ;
        RECT 24.735 142.195 25.605 142.535 ;
        RECT 25.840 142.195 26.010 142.655 ;
        RECT 26.845 142.625 27.920 142.795 ;
        RECT 26.180 142.025 26.550 142.485 ;
        RECT 26.845 142.285 27.015 142.625 ;
        RECT 27.185 142.025 27.515 142.455 ;
        RECT 27.750 142.285 27.920 142.625 ;
        RECT 28.090 142.525 28.260 143.305 ;
        RECT 28.430 143.085 28.600 143.675 ;
        RECT 28.770 143.275 29.120 143.895 ;
        RECT 28.430 142.695 28.895 143.085 ;
        RECT 29.290 142.825 29.460 144.185 ;
        RECT 29.630 142.995 30.090 144.045 ;
        RECT 29.065 142.655 29.460 142.825 ;
        RECT 29.065 142.525 29.235 142.655 ;
        RECT 28.090 142.195 28.770 142.525 ;
        RECT 28.985 142.195 29.235 142.525 ;
        RECT 29.405 142.025 29.655 142.485 ;
        RECT 29.825 142.210 30.150 142.995 ;
        RECT 30.320 142.195 30.490 144.315 ;
        RECT 30.660 144.195 30.990 144.575 ;
        RECT 31.160 144.025 31.415 144.315 ;
        RECT 30.665 143.855 31.415 144.025 ;
        RECT 30.665 142.865 30.895 143.855 ;
        RECT 32.715 143.795 33.215 144.405 ;
        RECT 31.065 143.035 31.415 143.685 ;
        RECT 32.510 143.335 32.860 143.585 ;
        RECT 33.045 143.165 33.215 143.795 ;
        RECT 33.845 143.925 34.175 144.405 ;
        RECT 34.345 144.115 34.570 144.575 ;
        RECT 34.740 143.925 35.070 144.405 ;
        RECT 33.845 143.755 35.070 143.925 ;
        RECT 35.260 143.775 35.510 144.575 ;
        RECT 35.680 143.775 36.020 144.405 ;
        RECT 36.190 143.825 37.400 144.575 ;
        RECT 33.385 143.385 33.715 143.585 ;
        RECT 33.885 143.385 34.215 143.585 ;
        RECT 34.385 143.385 34.805 143.585 ;
        RECT 34.980 143.415 35.675 143.585 ;
        RECT 34.980 143.165 35.150 143.415 ;
        RECT 35.845 143.165 36.020 143.775 ;
        RECT 32.715 142.995 35.150 143.165 ;
        RECT 30.665 142.695 31.415 142.865 ;
        RECT 30.660 142.025 30.990 142.525 ;
        RECT 31.160 142.195 31.415 142.695 ;
        RECT 32.715 142.195 33.045 142.995 ;
        RECT 33.215 142.025 33.545 142.825 ;
        RECT 33.845 142.195 34.175 142.995 ;
        RECT 34.820 142.025 35.070 142.825 ;
        RECT 35.340 142.025 35.510 143.165 ;
        RECT 35.680 142.195 36.020 143.165 ;
        RECT 36.190 143.115 36.710 143.655 ;
        RECT 36.880 143.285 37.400 143.825 ;
        RECT 37.570 143.775 37.910 144.405 ;
        RECT 38.080 143.775 38.330 144.575 ;
        RECT 38.520 143.925 38.850 144.405 ;
        RECT 39.020 144.115 39.245 144.575 ;
        RECT 39.415 143.925 39.745 144.405 ;
        RECT 37.570 143.165 37.745 143.775 ;
        RECT 38.520 143.755 39.745 143.925 ;
        RECT 40.375 143.795 40.875 144.405 ;
        RECT 41.710 143.805 43.380 144.575 ;
        RECT 37.915 143.415 38.610 143.585 ;
        RECT 38.440 143.165 38.610 143.415 ;
        RECT 38.785 143.385 39.205 143.585 ;
        RECT 39.375 143.385 39.705 143.585 ;
        RECT 39.875 143.385 40.205 143.585 ;
        RECT 40.375 143.165 40.545 143.795 ;
        RECT 40.730 143.335 41.080 143.585 ;
        RECT 36.190 142.025 37.400 143.115 ;
        RECT 37.570 142.195 37.910 143.165 ;
        RECT 38.080 142.025 38.250 143.165 ;
        RECT 38.440 142.995 40.875 143.165 ;
        RECT 38.520 142.025 38.770 142.825 ;
        RECT 39.415 142.195 39.745 142.995 ;
        RECT 40.045 142.025 40.375 142.825 ;
        RECT 40.545 142.195 40.875 142.995 ;
        RECT 41.710 143.115 42.460 143.635 ;
        RECT 42.630 143.285 43.380 143.805 ;
        RECT 43.555 143.835 43.810 144.405 ;
        RECT 43.980 144.175 44.310 144.575 ;
        RECT 44.735 144.040 45.265 144.405 ;
        RECT 45.455 144.235 45.730 144.405 ;
        RECT 45.450 144.065 45.730 144.235 ;
        RECT 44.735 144.005 44.910 144.040 ;
        RECT 43.980 143.835 44.910 144.005 ;
        RECT 43.555 143.165 43.725 143.835 ;
        RECT 43.980 143.665 44.150 143.835 ;
        RECT 43.895 143.335 44.150 143.665 ;
        RECT 44.375 143.335 44.570 143.665 ;
        RECT 41.710 142.025 43.380 143.115 ;
        RECT 43.555 142.195 43.890 143.165 ;
        RECT 44.060 142.025 44.230 143.165 ;
        RECT 44.400 142.365 44.570 143.335 ;
        RECT 44.740 142.705 44.910 143.835 ;
        RECT 45.080 143.045 45.250 143.845 ;
        RECT 45.455 143.245 45.730 144.065 ;
        RECT 45.900 143.045 46.090 144.405 ;
        RECT 46.270 144.040 46.780 144.575 ;
        RECT 47.000 143.765 47.245 144.370 ;
        RECT 47.690 143.850 47.980 144.575 ;
        RECT 48.610 143.805 52.120 144.575 ;
        RECT 52.380 144.095 52.680 144.575 ;
        RECT 52.850 143.925 53.110 144.380 ;
        RECT 53.280 144.095 53.540 144.575 ;
        RECT 53.720 143.925 53.980 144.380 ;
        RECT 54.150 144.095 54.400 144.575 ;
        RECT 54.580 143.925 54.840 144.380 ;
        RECT 55.010 144.095 55.260 144.575 ;
        RECT 55.440 143.925 55.700 144.380 ;
        RECT 55.870 144.095 56.115 144.575 ;
        RECT 56.285 143.925 56.560 144.380 ;
        RECT 56.730 144.095 56.975 144.575 ;
        RECT 57.145 143.925 57.405 144.380 ;
        RECT 57.575 144.095 57.835 144.575 ;
        RECT 58.005 143.925 58.265 144.380 ;
        RECT 58.435 144.095 58.695 144.575 ;
        RECT 58.865 143.925 59.125 144.380 ;
        RECT 59.295 144.015 59.555 144.575 ;
        RECT 46.290 143.595 47.520 143.765 ;
        RECT 45.080 142.875 46.090 143.045 ;
        RECT 46.260 143.030 47.010 143.220 ;
        RECT 44.740 142.535 45.865 142.705 ;
        RECT 46.260 142.365 46.430 143.030 ;
        RECT 47.180 142.785 47.520 143.595 ;
        RECT 44.400 142.195 46.430 142.365 ;
        RECT 46.600 142.025 46.770 142.785 ;
        RECT 47.005 142.375 47.520 142.785 ;
        RECT 47.690 142.025 47.980 143.190 ;
        RECT 48.610 143.115 50.300 143.635 ;
        RECT 50.470 143.285 52.120 143.805 ;
        RECT 52.380 143.755 59.125 143.925 ;
        RECT 52.380 143.165 53.545 143.755 ;
        RECT 59.725 143.585 59.975 144.395 ;
        RECT 60.155 144.050 60.415 144.575 ;
        RECT 60.585 143.585 60.835 144.395 ;
        RECT 61.015 144.065 61.320 144.575 ;
        RECT 61.865 144.235 62.120 144.395 ;
        RECT 61.780 144.065 62.120 144.235 ;
        RECT 62.300 144.115 62.585 144.575 ;
        RECT 53.715 143.335 60.835 143.585 ;
        RECT 61.005 143.335 61.320 143.895 ;
        RECT 61.865 143.865 62.120 144.065 ;
        RECT 48.610 142.025 52.120 143.115 ;
        RECT 52.380 142.940 59.125 143.165 ;
        RECT 52.380 142.025 52.650 142.770 ;
        RECT 52.820 142.200 53.110 142.940 ;
        RECT 53.720 142.925 59.125 142.940 ;
        RECT 53.280 142.030 53.535 142.755 ;
        RECT 53.720 142.200 53.980 142.925 ;
        RECT 54.150 142.030 54.395 142.755 ;
        RECT 54.580 142.200 54.840 142.925 ;
        RECT 55.010 142.030 55.255 142.755 ;
        RECT 55.440 142.200 55.700 142.925 ;
        RECT 55.870 142.030 56.115 142.755 ;
        RECT 56.285 142.200 56.545 142.925 ;
        RECT 56.715 142.030 56.975 142.755 ;
        RECT 57.145 142.200 57.405 142.925 ;
        RECT 57.575 142.030 57.835 142.755 ;
        RECT 58.005 142.200 58.265 142.925 ;
        RECT 58.435 142.030 58.695 142.755 ;
        RECT 58.865 142.200 59.125 142.925 ;
        RECT 59.295 142.030 59.555 142.825 ;
        RECT 59.725 142.200 59.975 143.335 ;
        RECT 53.280 142.025 59.555 142.030 ;
        RECT 60.155 142.025 60.415 142.835 ;
        RECT 60.590 142.195 60.835 143.335 ;
        RECT 61.865 143.005 62.045 143.865 ;
        RECT 62.765 143.665 63.015 144.315 ;
        RECT 62.215 143.335 63.015 143.665 ;
        RECT 61.015 142.025 61.310 142.835 ;
        RECT 61.865 142.335 62.120 143.005 ;
        RECT 62.300 142.025 62.585 142.825 ;
        RECT 62.765 142.745 63.015 143.335 ;
        RECT 63.215 143.980 63.535 144.310 ;
        RECT 63.715 144.095 64.375 144.575 ;
        RECT 64.575 144.185 65.425 144.355 ;
        RECT 63.215 143.085 63.405 143.980 ;
        RECT 63.725 143.655 64.385 143.925 ;
        RECT 64.055 143.595 64.385 143.655 ;
        RECT 63.575 143.425 63.905 143.485 ;
        RECT 64.575 143.425 64.745 144.185 ;
        RECT 65.985 144.115 66.305 144.575 ;
        RECT 66.505 143.935 66.755 144.365 ;
        RECT 67.045 144.135 67.455 144.575 ;
        RECT 67.625 144.195 68.640 144.395 ;
        RECT 64.915 143.765 66.165 143.935 ;
        RECT 64.915 143.645 65.245 143.765 ;
        RECT 63.575 143.255 65.475 143.425 ;
        RECT 63.215 142.915 65.135 143.085 ;
        RECT 63.215 142.895 63.535 142.915 ;
        RECT 62.765 142.235 63.095 142.745 ;
        RECT 63.365 142.285 63.535 142.895 ;
        RECT 65.305 142.745 65.475 143.255 ;
        RECT 65.645 143.185 65.825 143.595 ;
        RECT 65.995 143.005 66.165 143.765 ;
        RECT 63.705 142.025 64.035 142.715 ;
        RECT 64.265 142.575 65.475 142.745 ;
        RECT 65.645 142.695 66.165 143.005 ;
        RECT 66.335 143.595 66.755 143.935 ;
        RECT 67.045 143.595 67.455 143.925 ;
        RECT 66.335 142.825 66.525 143.595 ;
        RECT 67.625 143.465 67.795 144.195 ;
        RECT 68.940 144.025 69.110 144.355 ;
        RECT 69.280 144.195 69.610 144.575 ;
        RECT 67.965 143.645 68.315 144.015 ;
        RECT 67.625 143.425 68.045 143.465 ;
        RECT 66.695 143.255 68.045 143.425 ;
        RECT 66.695 143.095 66.945 143.255 ;
        RECT 67.455 142.825 67.705 143.085 ;
        RECT 66.335 142.575 67.705 142.825 ;
        RECT 64.265 142.285 64.505 142.575 ;
        RECT 65.305 142.495 65.475 142.575 ;
        RECT 64.705 142.025 65.125 142.405 ;
        RECT 65.305 142.245 65.935 142.495 ;
        RECT 66.405 142.025 66.735 142.405 ;
        RECT 66.905 142.285 67.075 142.575 ;
        RECT 67.875 142.410 68.045 143.255 ;
        RECT 68.495 143.085 68.715 143.955 ;
        RECT 68.940 143.835 69.635 144.025 ;
        RECT 68.215 142.705 68.715 143.085 ;
        RECT 68.885 143.035 69.295 143.655 ;
        RECT 69.465 142.865 69.635 143.835 ;
        RECT 68.940 142.695 69.635 142.865 ;
        RECT 67.255 142.025 67.635 142.405 ;
        RECT 67.875 142.240 68.705 142.410 ;
        RECT 68.940 142.195 69.110 142.695 ;
        RECT 69.280 142.025 69.610 142.525 ;
        RECT 69.825 142.195 70.050 144.315 ;
        RECT 70.220 144.195 70.550 144.575 ;
        RECT 70.720 144.025 70.890 144.315 ;
        RECT 70.225 143.855 70.890 144.025 ;
        RECT 70.225 142.865 70.455 143.855 ;
        RECT 71.610 143.805 73.280 144.575 ;
        RECT 73.450 143.850 73.740 144.575 ;
        RECT 73.915 144.030 79.260 144.575 ;
        RECT 70.625 143.035 70.975 143.685 ;
        RECT 71.610 143.115 72.360 143.635 ;
        RECT 72.530 143.285 73.280 143.805 ;
        RECT 70.225 142.695 70.890 142.865 ;
        RECT 70.220 142.025 70.550 142.525 ;
        RECT 70.720 142.195 70.890 142.695 ;
        RECT 71.610 142.025 73.280 143.115 ;
        RECT 73.450 142.025 73.740 143.190 ;
        RECT 75.505 142.460 75.855 143.710 ;
        RECT 77.335 143.200 77.675 144.030 ;
        RECT 79.705 143.765 79.950 144.370 ;
        RECT 80.170 144.040 80.680 144.575 ;
        RECT 79.430 143.595 80.660 143.765 ;
        RECT 79.430 142.785 79.770 143.595 ;
        RECT 79.940 143.030 80.690 143.220 ;
        RECT 73.915 142.025 79.260 142.460 ;
        RECT 79.430 142.375 79.945 142.785 ;
        RECT 80.180 142.025 80.350 142.785 ;
        RECT 80.520 142.365 80.690 143.030 ;
        RECT 80.860 143.045 81.050 144.405 ;
        RECT 81.220 143.555 81.495 144.405 ;
        RECT 81.685 144.040 82.215 144.405 ;
        RECT 82.640 144.175 82.970 144.575 ;
        RECT 82.040 144.005 82.215 144.040 ;
        RECT 81.220 143.385 81.500 143.555 ;
        RECT 81.220 143.245 81.495 143.385 ;
        RECT 81.700 143.045 81.870 143.845 ;
        RECT 80.860 142.875 81.870 143.045 ;
        RECT 82.040 143.835 82.970 144.005 ;
        RECT 83.140 143.835 83.395 144.405 ;
        RECT 82.040 142.705 82.210 143.835 ;
        RECT 82.800 143.665 82.970 143.835 ;
        RECT 81.085 142.535 82.210 142.705 ;
        RECT 82.380 143.335 82.575 143.665 ;
        RECT 82.800 143.335 83.055 143.665 ;
        RECT 82.380 142.365 82.550 143.335 ;
        RECT 83.225 143.165 83.395 143.835 ;
        RECT 80.520 142.195 82.550 142.365 ;
        RECT 82.720 142.025 82.890 143.165 ;
        RECT 83.060 142.195 83.395 143.165 ;
        RECT 84.490 143.900 84.750 144.405 ;
        RECT 84.930 144.195 85.260 144.575 ;
        RECT 85.440 144.025 85.610 144.405 ;
        RECT 84.490 143.100 84.660 143.900 ;
        RECT 84.945 143.855 85.610 144.025 ;
        RECT 84.945 143.600 85.115 143.855 ;
        RECT 85.870 143.825 87.080 144.575 ;
        RECT 87.255 144.030 92.600 144.575 ;
        RECT 84.830 143.270 85.115 143.600 ;
        RECT 85.350 143.305 85.680 143.675 ;
        RECT 84.945 143.125 85.115 143.270 ;
        RECT 84.490 142.195 84.760 143.100 ;
        RECT 84.945 142.955 85.610 143.125 ;
        RECT 84.930 142.025 85.260 142.785 ;
        RECT 85.440 142.195 85.610 142.955 ;
        RECT 85.870 143.115 86.390 143.655 ;
        RECT 86.560 143.285 87.080 143.825 ;
        RECT 85.870 142.025 87.080 143.115 ;
        RECT 88.845 142.460 89.195 143.710 ;
        RECT 90.675 143.200 91.015 144.030 ;
        RECT 92.770 143.900 93.040 144.245 ;
        RECT 93.230 144.175 93.610 144.575 ;
        RECT 93.780 144.005 93.950 144.355 ;
        RECT 94.120 144.175 94.450 144.575 ;
        RECT 94.650 144.005 94.820 144.355 ;
        RECT 95.020 144.075 95.350 144.575 ;
        RECT 92.770 143.165 92.940 143.900 ;
        RECT 93.210 143.835 94.820 144.005 ;
        RECT 93.210 143.665 93.380 143.835 ;
        RECT 93.110 143.335 93.380 143.665 ;
        RECT 93.550 143.335 93.955 143.665 ;
        RECT 93.210 143.165 93.380 143.335 ;
        RECT 94.125 143.215 94.835 143.665 ;
        RECT 95.005 143.335 95.355 143.905 ;
        RECT 95.530 143.775 95.870 144.405 ;
        RECT 96.040 143.775 96.290 144.575 ;
        RECT 96.480 143.925 96.810 144.405 ;
        RECT 96.980 144.115 97.205 144.575 ;
        RECT 97.375 143.925 97.705 144.405 ;
        RECT 95.530 143.725 95.760 143.775 ;
        RECT 96.480 143.755 97.705 143.925 ;
        RECT 98.335 143.795 98.835 144.405 ;
        RECT 99.210 143.850 99.500 144.575 ;
        RECT 99.675 144.030 105.020 144.575 ;
        RECT 87.255 142.025 92.600 142.460 ;
        RECT 92.770 142.195 93.040 143.165 ;
        RECT 93.210 142.995 93.935 143.165 ;
        RECT 94.125 143.045 94.840 143.215 ;
        RECT 95.530 143.165 95.705 143.725 ;
        RECT 95.875 143.415 96.570 143.585 ;
        RECT 96.400 143.165 96.570 143.415 ;
        RECT 96.745 143.385 97.165 143.585 ;
        RECT 97.335 143.385 97.665 143.585 ;
        RECT 97.835 143.385 98.165 143.585 ;
        RECT 98.335 143.165 98.505 143.795 ;
        RECT 98.690 143.335 99.040 143.585 ;
        RECT 93.765 142.875 93.935 142.995 ;
        RECT 95.035 142.875 95.355 143.165 ;
        RECT 93.250 142.025 93.530 142.825 ;
        RECT 93.765 142.705 95.355 142.875 ;
        RECT 93.700 142.245 95.355 142.535 ;
        RECT 95.530 142.195 95.870 143.165 ;
        RECT 96.040 142.025 96.210 143.165 ;
        RECT 96.400 142.995 98.835 143.165 ;
        RECT 96.480 142.025 96.730 142.825 ;
        RECT 97.375 142.195 97.705 142.995 ;
        RECT 98.005 142.025 98.335 142.825 ;
        RECT 98.505 142.195 98.835 142.995 ;
        RECT 99.210 142.025 99.500 143.190 ;
        RECT 101.265 142.460 101.615 143.710 ;
        RECT 103.095 143.200 103.435 144.030 ;
        RECT 105.230 143.755 105.460 144.575 ;
        RECT 105.630 143.775 105.960 144.405 ;
        RECT 105.210 143.335 105.540 143.585 ;
        RECT 105.710 143.175 105.960 143.775 ;
        RECT 106.130 143.755 106.340 144.575 ;
        RECT 106.660 144.025 106.830 144.405 ;
        RECT 107.010 144.195 107.340 144.575 ;
        RECT 106.660 143.855 107.325 144.025 ;
        RECT 107.520 143.900 107.780 144.405 ;
        RECT 106.590 143.305 106.920 143.675 ;
        RECT 107.155 143.600 107.325 143.855 ;
        RECT 99.675 142.025 105.020 142.460 ;
        RECT 105.230 142.025 105.460 143.165 ;
        RECT 105.630 142.195 105.960 143.175 ;
        RECT 107.155 143.270 107.440 143.600 ;
        RECT 106.130 142.025 106.340 143.165 ;
        RECT 107.155 143.125 107.325 143.270 ;
        RECT 106.660 142.955 107.325 143.125 ;
        RECT 107.610 143.100 107.780 143.900 ;
        RECT 108.410 143.805 111.000 144.575 ;
        RECT 111.170 143.825 112.380 144.575 ;
        RECT 106.660 142.195 106.830 142.955 ;
        RECT 107.010 142.025 107.340 142.785 ;
        RECT 107.510 142.195 107.780 143.100 ;
        RECT 108.410 143.115 109.620 143.635 ;
        RECT 109.790 143.285 111.000 143.805 ;
        RECT 111.170 143.115 111.690 143.655 ;
        RECT 111.860 143.285 112.380 143.825 ;
        RECT 108.410 142.025 111.000 143.115 ;
        RECT 111.170 142.025 112.380 143.115 ;
        RECT 18.165 141.855 112.465 142.025 ;
        RECT 18.250 140.765 19.460 141.855 ;
        RECT 18.250 140.055 18.770 140.595 ;
        RECT 18.940 140.225 19.460 140.765 ;
        RECT 20.150 140.715 20.360 141.855 ;
        RECT 20.530 140.705 20.860 141.685 ;
        RECT 21.030 140.715 21.260 141.855 ;
        RECT 21.510 140.715 21.740 141.855 ;
        RECT 21.910 140.705 22.240 141.685 ;
        RECT 22.410 140.715 22.620 141.855 ;
        RECT 22.855 140.715 23.190 141.685 ;
        RECT 23.360 140.715 23.530 141.855 ;
        RECT 23.700 141.515 25.730 141.685 ;
        RECT 18.250 139.305 19.460 140.055 ;
        RECT 20.150 139.305 20.360 140.125 ;
        RECT 20.530 140.105 20.780 140.705 ;
        RECT 20.950 140.295 21.280 140.545 ;
        RECT 21.490 140.295 21.820 140.545 ;
        RECT 20.530 139.475 20.860 140.105 ;
        RECT 21.030 139.305 21.260 140.125 ;
        RECT 21.510 139.305 21.740 140.125 ;
        RECT 21.990 140.105 22.240 140.705 ;
        RECT 21.910 139.475 22.240 140.105 ;
        RECT 22.410 139.305 22.620 140.125 ;
        RECT 22.855 140.045 23.025 140.715 ;
        RECT 23.700 140.545 23.870 141.515 ;
        RECT 23.195 140.215 23.450 140.545 ;
        RECT 23.675 140.215 23.870 140.545 ;
        RECT 24.040 141.175 25.165 141.345 ;
        RECT 23.280 140.045 23.450 140.215 ;
        RECT 24.040 140.045 24.210 141.175 ;
        RECT 22.855 139.475 23.110 140.045 ;
        RECT 23.280 139.875 24.210 140.045 ;
        RECT 24.380 140.835 25.390 141.005 ;
        RECT 24.380 140.035 24.550 140.835 ;
        RECT 24.755 140.495 25.030 140.635 ;
        RECT 24.750 140.325 25.030 140.495 ;
        RECT 24.035 139.840 24.210 139.875 ;
        RECT 23.280 139.305 23.610 139.705 ;
        RECT 24.035 139.475 24.565 139.840 ;
        RECT 24.755 139.475 25.030 140.325 ;
        RECT 25.200 139.475 25.390 140.835 ;
        RECT 25.560 140.850 25.730 141.515 ;
        RECT 25.900 141.095 26.070 141.855 ;
        RECT 26.305 141.095 26.820 141.505 ;
        RECT 25.560 140.660 26.310 140.850 ;
        RECT 26.480 140.285 26.820 141.095 ;
        RECT 25.590 140.115 26.820 140.285 ;
        RECT 26.990 141.095 27.505 141.505 ;
        RECT 27.740 141.095 27.910 141.855 ;
        RECT 28.080 141.515 30.110 141.685 ;
        RECT 26.990 140.285 27.330 141.095 ;
        RECT 28.080 140.850 28.250 141.515 ;
        RECT 28.645 141.175 29.770 141.345 ;
        RECT 27.500 140.660 28.250 140.850 ;
        RECT 28.420 140.835 29.430 141.005 ;
        RECT 26.990 140.115 28.220 140.285 ;
        RECT 25.570 139.305 26.080 139.840 ;
        RECT 26.300 139.510 26.545 140.115 ;
        RECT 27.265 139.510 27.510 140.115 ;
        RECT 27.730 139.305 28.240 139.840 ;
        RECT 28.420 139.475 28.610 140.835 ;
        RECT 28.780 140.155 29.055 140.635 ;
        RECT 28.780 139.985 29.060 140.155 ;
        RECT 29.260 140.035 29.430 140.835 ;
        RECT 29.600 140.045 29.770 141.175 ;
        RECT 29.940 140.545 30.110 141.515 ;
        RECT 30.280 140.715 30.450 141.855 ;
        RECT 30.620 140.715 30.955 141.685 ;
        RECT 29.940 140.215 30.135 140.545 ;
        RECT 30.360 140.215 30.615 140.545 ;
        RECT 30.360 140.045 30.530 140.215 ;
        RECT 30.785 140.045 30.955 140.715 ;
        RECT 28.780 139.475 29.055 139.985 ;
        RECT 29.600 139.875 30.530 140.045 ;
        RECT 29.600 139.840 29.775 139.875 ;
        RECT 29.245 139.475 29.775 139.840 ;
        RECT 30.200 139.305 30.530 139.705 ;
        RECT 30.700 139.475 30.955 140.045 ;
        RECT 32.050 140.715 32.320 141.685 ;
        RECT 32.530 141.055 32.810 141.855 ;
        RECT 32.980 141.345 34.635 141.635 ;
        RECT 33.045 141.005 34.635 141.175 ;
        RECT 33.045 140.885 33.215 141.005 ;
        RECT 32.490 140.715 33.215 140.885 ;
        RECT 32.050 139.980 32.220 140.715 ;
        RECT 32.490 140.545 32.660 140.715 ;
        RECT 33.405 140.665 34.120 140.835 ;
        RECT 34.315 140.715 34.635 141.005 ;
        RECT 34.810 140.690 35.100 141.855 ;
        RECT 36.190 140.765 39.700 141.855 ;
        RECT 32.390 140.215 32.660 140.545 ;
        RECT 32.830 140.215 33.235 140.545 ;
        RECT 33.405 140.215 34.115 140.665 ;
        RECT 32.490 140.045 32.660 140.215 ;
        RECT 32.050 139.635 32.320 139.980 ;
        RECT 32.490 139.875 34.100 140.045 ;
        RECT 34.285 139.975 34.635 140.545 ;
        RECT 36.190 140.245 37.880 140.765 ;
        RECT 39.910 140.715 40.140 141.855 ;
        RECT 40.310 140.705 40.640 141.685 ;
        RECT 40.810 140.715 41.020 141.855 ;
        RECT 41.625 140.875 41.880 141.545 ;
        RECT 42.060 141.055 42.345 141.855 ;
        RECT 42.525 141.135 42.855 141.645 ;
        RECT 41.625 140.835 41.805 140.875 ;
        RECT 38.050 140.075 39.700 140.595 ;
        RECT 39.890 140.295 40.220 140.545 ;
        RECT 32.510 139.305 32.890 139.705 ;
        RECT 33.060 139.525 33.230 139.875 ;
        RECT 33.400 139.305 33.730 139.705 ;
        RECT 33.930 139.525 34.100 139.875 ;
        RECT 34.300 139.305 34.630 139.805 ;
        RECT 34.810 139.305 35.100 140.030 ;
        RECT 36.190 139.305 39.700 140.075 ;
        RECT 39.910 139.305 40.140 140.125 ;
        RECT 40.390 140.105 40.640 140.705 ;
        RECT 41.540 140.665 41.805 140.835 ;
        RECT 40.310 139.475 40.640 140.105 ;
        RECT 40.810 139.305 41.020 140.125 ;
        RECT 41.625 140.015 41.805 140.665 ;
        RECT 42.525 140.545 42.775 141.135 ;
        RECT 43.125 140.985 43.295 141.595 ;
        RECT 43.465 141.165 43.795 141.855 ;
        RECT 44.025 141.305 44.265 141.595 ;
        RECT 44.465 141.475 44.885 141.855 ;
        RECT 45.065 141.385 45.695 141.635 ;
        RECT 46.165 141.475 46.495 141.855 ;
        RECT 45.065 141.305 45.235 141.385 ;
        RECT 46.665 141.305 46.835 141.595 ;
        RECT 47.015 141.475 47.395 141.855 ;
        RECT 47.635 141.470 48.465 141.640 ;
        RECT 44.025 141.135 45.235 141.305 ;
        RECT 41.975 140.215 42.775 140.545 ;
        RECT 41.625 139.485 41.880 140.015 ;
        RECT 42.060 139.305 42.345 139.765 ;
        RECT 42.525 139.565 42.775 140.215 ;
        RECT 42.975 140.965 43.295 140.985 ;
        RECT 42.975 140.795 44.895 140.965 ;
        RECT 42.975 139.900 43.165 140.795 ;
        RECT 45.065 140.625 45.235 141.135 ;
        RECT 45.405 140.875 45.925 141.185 ;
        RECT 43.335 140.455 45.235 140.625 ;
        RECT 43.335 140.395 43.665 140.455 ;
        RECT 43.815 140.225 44.145 140.285 ;
        RECT 43.485 139.955 44.145 140.225 ;
        RECT 42.975 139.570 43.295 139.900 ;
        RECT 43.475 139.305 44.135 139.785 ;
        RECT 44.335 139.695 44.505 140.455 ;
        RECT 45.405 140.285 45.585 140.695 ;
        RECT 44.675 140.115 45.005 140.235 ;
        RECT 45.755 140.115 45.925 140.875 ;
        RECT 44.675 139.945 45.925 140.115 ;
        RECT 46.095 141.055 47.465 141.305 ;
        RECT 46.095 140.285 46.285 141.055 ;
        RECT 47.215 140.795 47.465 141.055 ;
        RECT 46.455 140.625 46.705 140.785 ;
        RECT 47.635 140.625 47.805 141.470 ;
        RECT 48.700 141.185 48.870 141.685 ;
        RECT 49.040 141.355 49.370 141.855 ;
        RECT 47.975 140.795 48.475 141.175 ;
        RECT 48.700 141.015 49.395 141.185 ;
        RECT 46.455 140.455 47.805 140.625 ;
        RECT 47.385 140.415 47.805 140.455 ;
        RECT 46.095 139.945 46.515 140.285 ;
        RECT 46.805 139.955 47.215 140.285 ;
        RECT 44.335 139.525 45.185 139.695 ;
        RECT 45.745 139.305 46.065 139.765 ;
        RECT 46.265 139.515 46.515 139.945 ;
        RECT 46.805 139.305 47.215 139.745 ;
        RECT 47.385 139.685 47.555 140.415 ;
        RECT 47.725 139.865 48.075 140.235 ;
        RECT 48.255 139.925 48.475 140.795 ;
        RECT 48.645 140.225 49.055 140.845 ;
        RECT 49.225 140.045 49.395 141.015 ;
        RECT 48.700 139.855 49.395 140.045 ;
        RECT 47.385 139.485 48.400 139.685 ;
        RECT 48.700 139.525 48.870 139.855 ;
        RECT 49.040 139.305 49.370 139.685 ;
        RECT 49.585 139.565 49.810 141.685 ;
        RECT 49.980 141.355 50.310 141.855 ;
        RECT 50.480 141.185 50.650 141.685 ;
        RECT 49.985 141.015 50.650 141.185 ;
        RECT 49.985 140.025 50.215 141.015 ;
        RECT 50.385 140.195 50.735 140.845 ;
        RECT 50.910 140.715 51.180 141.685 ;
        RECT 51.390 141.055 51.670 141.855 ;
        RECT 51.840 141.345 53.495 141.635 ;
        RECT 51.905 141.005 53.495 141.175 ;
        RECT 51.905 140.885 52.075 141.005 ;
        RECT 51.350 140.715 52.075 140.885 ;
        RECT 49.985 139.855 50.650 140.025 ;
        RECT 49.980 139.305 50.310 139.685 ;
        RECT 50.480 139.565 50.650 139.855 ;
        RECT 50.910 139.980 51.080 140.715 ;
        RECT 51.350 140.545 51.520 140.715 ;
        RECT 51.250 140.215 51.520 140.545 ;
        RECT 51.690 140.215 52.095 140.545 ;
        RECT 52.265 140.215 52.975 140.835 ;
        RECT 53.175 140.715 53.495 141.005 ;
        RECT 53.670 140.765 56.260 141.855 ;
        RECT 51.350 140.045 51.520 140.215 ;
        RECT 50.910 139.635 51.180 139.980 ;
        RECT 51.350 139.875 52.960 140.045 ;
        RECT 53.145 139.975 53.495 140.545 ;
        RECT 53.670 140.245 54.880 140.765 ;
        RECT 56.430 140.715 56.770 141.685 ;
        RECT 56.940 140.715 57.110 141.855 ;
        RECT 57.380 141.055 57.630 141.855 ;
        RECT 58.275 140.885 58.605 141.685 ;
        RECT 58.905 141.055 59.235 141.855 ;
        RECT 59.405 140.885 59.735 141.685 ;
        RECT 57.300 140.715 59.735 140.885 ;
        RECT 55.050 140.075 56.260 140.595 ;
        RECT 51.370 139.305 51.750 139.705 ;
        RECT 51.920 139.525 52.090 139.875 ;
        RECT 52.260 139.305 52.590 139.705 ;
        RECT 52.790 139.525 52.960 139.875 ;
        RECT 53.160 139.305 53.490 139.805 ;
        RECT 53.670 139.305 56.260 140.075 ;
        RECT 56.430 140.155 56.605 140.715 ;
        RECT 57.300 140.465 57.470 140.715 ;
        RECT 56.775 140.295 57.470 140.465 ;
        RECT 57.645 140.295 58.065 140.495 ;
        RECT 58.235 140.295 58.565 140.495 ;
        RECT 58.735 140.295 59.065 140.495 ;
        RECT 56.430 140.105 56.660 140.155 ;
        RECT 56.430 139.475 56.770 140.105 ;
        RECT 56.940 139.305 57.190 140.105 ;
        RECT 57.380 139.955 58.605 140.125 ;
        RECT 57.380 139.475 57.710 139.955 ;
        RECT 57.880 139.305 58.105 139.765 ;
        RECT 58.275 139.475 58.605 139.955 ;
        RECT 59.235 140.085 59.405 140.715 ;
        RECT 60.570 140.690 60.860 141.855 ;
        RECT 61.405 140.875 61.660 141.545 ;
        RECT 61.840 141.055 62.125 141.855 ;
        RECT 62.305 141.135 62.635 141.645 ;
        RECT 59.590 140.295 59.940 140.545 ;
        RECT 59.235 139.475 59.735 140.085 ;
        RECT 60.570 139.305 60.860 140.030 ;
        RECT 61.405 140.015 61.585 140.875 ;
        RECT 62.305 140.545 62.555 141.135 ;
        RECT 62.905 140.985 63.075 141.595 ;
        RECT 63.245 141.165 63.575 141.855 ;
        RECT 63.805 141.305 64.045 141.595 ;
        RECT 64.245 141.475 64.665 141.855 ;
        RECT 64.845 141.385 65.475 141.635 ;
        RECT 65.945 141.475 66.275 141.855 ;
        RECT 64.845 141.305 65.015 141.385 ;
        RECT 66.445 141.305 66.615 141.595 ;
        RECT 66.795 141.475 67.175 141.855 ;
        RECT 67.415 141.470 68.245 141.640 ;
        RECT 63.805 141.135 65.015 141.305 ;
        RECT 61.755 140.215 62.555 140.545 ;
        RECT 61.405 139.815 61.660 140.015 ;
        RECT 61.320 139.645 61.660 139.815 ;
        RECT 61.405 139.485 61.660 139.645 ;
        RECT 61.840 139.305 62.125 139.765 ;
        RECT 62.305 139.565 62.555 140.215 ;
        RECT 62.755 140.965 63.075 140.985 ;
        RECT 62.755 140.795 64.675 140.965 ;
        RECT 62.755 139.900 62.945 140.795 ;
        RECT 64.845 140.625 65.015 141.135 ;
        RECT 65.185 140.875 65.705 141.185 ;
        RECT 63.115 140.455 65.015 140.625 ;
        RECT 63.115 140.395 63.445 140.455 ;
        RECT 63.595 140.225 63.925 140.285 ;
        RECT 63.265 139.955 63.925 140.225 ;
        RECT 62.755 139.570 63.075 139.900 ;
        RECT 63.255 139.305 63.915 139.785 ;
        RECT 64.115 139.695 64.285 140.455 ;
        RECT 65.185 140.285 65.365 140.695 ;
        RECT 64.455 140.115 64.785 140.235 ;
        RECT 65.535 140.115 65.705 140.875 ;
        RECT 64.455 139.945 65.705 140.115 ;
        RECT 65.875 141.055 67.245 141.305 ;
        RECT 65.875 140.285 66.065 141.055 ;
        RECT 66.995 140.795 67.245 141.055 ;
        RECT 66.235 140.625 66.485 140.785 ;
        RECT 67.415 140.625 67.585 141.470 ;
        RECT 68.480 141.185 68.650 141.685 ;
        RECT 68.820 141.355 69.150 141.855 ;
        RECT 67.755 140.795 68.255 141.175 ;
        RECT 68.480 141.015 69.175 141.185 ;
        RECT 66.235 140.455 67.585 140.625 ;
        RECT 67.165 140.415 67.585 140.455 ;
        RECT 65.875 139.945 66.295 140.285 ;
        RECT 66.585 139.955 66.995 140.285 ;
        RECT 64.115 139.525 64.965 139.695 ;
        RECT 65.525 139.305 65.845 139.765 ;
        RECT 66.045 139.515 66.295 139.945 ;
        RECT 66.585 139.305 66.995 139.745 ;
        RECT 67.165 139.685 67.335 140.415 ;
        RECT 67.505 139.865 67.855 140.235 ;
        RECT 68.035 139.925 68.255 140.795 ;
        RECT 68.425 140.225 68.835 140.845 ;
        RECT 69.005 140.045 69.175 141.015 ;
        RECT 68.480 139.855 69.175 140.045 ;
        RECT 67.165 139.485 68.180 139.685 ;
        RECT 68.480 139.525 68.650 139.855 ;
        RECT 68.820 139.305 69.150 139.685 ;
        RECT 69.365 139.565 69.590 141.685 ;
        RECT 69.760 141.355 70.090 141.855 ;
        RECT 70.260 141.185 70.430 141.685 ;
        RECT 69.765 141.015 70.430 141.185 ;
        RECT 69.765 140.025 69.995 141.015 ;
        RECT 70.165 140.195 70.515 140.845 ;
        RECT 71.150 140.765 72.820 141.855 ;
        RECT 71.150 140.245 71.900 140.765 ;
        RECT 72.990 140.715 73.330 141.685 ;
        RECT 73.500 140.715 73.670 141.855 ;
        RECT 73.940 141.055 74.190 141.855 ;
        RECT 74.835 140.885 75.165 141.685 ;
        RECT 75.465 141.055 75.795 141.855 ;
        RECT 75.965 140.885 76.295 141.685 ;
        RECT 77.045 141.175 77.300 141.545 ;
        RECT 76.960 141.005 77.300 141.175 ;
        RECT 77.480 141.055 77.765 141.855 ;
        RECT 77.945 141.135 78.275 141.645 ;
        RECT 73.860 140.715 76.295 140.885 ;
        RECT 77.045 140.875 77.300 141.005 ;
        RECT 72.070 140.075 72.820 140.595 ;
        RECT 69.765 139.855 70.430 140.025 ;
        RECT 69.760 139.305 70.090 139.685 ;
        RECT 70.260 139.565 70.430 139.855 ;
        RECT 71.150 139.305 72.820 140.075 ;
        RECT 72.990 140.105 73.165 140.715 ;
        RECT 73.860 140.465 74.030 140.715 ;
        RECT 73.335 140.295 74.030 140.465 ;
        RECT 74.205 140.295 74.625 140.495 ;
        RECT 74.795 140.295 75.125 140.495 ;
        RECT 75.295 140.295 75.625 140.495 ;
        RECT 72.990 139.475 73.330 140.105 ;
        RECT 73.500 139.305 73.750 140.105 ;
        RECT 73.940 139.955 75.165 140.125 ;
        RECT 73.940 139.475 74.270 139.955 ;
        RECT 74.440 139.305 74.665 139.765 ;
        RECT 74.835 139.475 75.165 139.955 ;
        RECT 75.795 140.085 75.965 140.715 ;
        RECT 76.150 140.295 76.500 140.545 ;
        RECT 75.795 139.475 76.295 140.085 ;
        RECT 77.045 140.015 77.225 140.875 ;
        RECT 77.945 140.545 78.195 141.135 ;
        RECT 78.545 140.985 78.715 141.595 ;
        RECT 78.885 141.165 79.215 141.855 ;
        RECT 79.445 141.305 79.685 141.595 ;
        RECT 79.885 141.475 80.305 141.855 ;
        RECT 80.485 141.385 81.115 141.635 ;
        RECT 81.585 141.475 81.915 141.855 ;
        RECT 80.485 141.305 80.655 141.385 ;
        RECT 82.085 141.305 82.255 141.595 ;
        RECT 82.435 141.475 82.815 141.855 ;
        RECT 83.055 141.470 83.885 141.640 ;
        RECT 79.445 141.135 80.655 141.305 ;
        RECT 77.395 140.215 78.195 140.545 ;
        RECT 77.045 139.485 77.300 140.015 ;
        RECT 77.480 139.305 77.765 139.765 ;
        RECT 77.945 139.565 78.195 140.215 ;
        RECT 78.395 140.965 78.715 140.985 ;
        RECT 78.395 140.795 80.315 140.965 ;
        RECT 78.395 139.900 78.585 140.795 ;
        RECT 80.485 140.625 80.655 141.135 ;
        RECT 80.825 140.875 81.345 141.185 ;
        RECT 78.755 140.455 80.655 140.625 ;
        RECT 78.755 140.395 79.085 140.455 ;
        RECT 79.235 140.225 79.565 140.285 ;
        RECT 78.905 139.955 79.565 140.225 ;
        RECT 78.395 139.570 78.715 139.900 ;
        RECT 78.895 139.305 79.555 139.785 ;
        RECT 79.755 139.695 79.925 140.455 ;
        RECT 80.825 140.285 81.005 140.695 ;
        RECT 80.095 140.115 80.425 140.235 ;
        RECT 81.175 140.115 81.345 140.875 ;
        RECT 80.095 139.945 81.345 140.115 ;
        RECT 81.515 141.055 82.885 141.305 ;
        RECT 81.515 140.285 81.705 141.055 ;
        RECT 82.635 140.795 82.885 141.055 ;
        RECT 81.875 140.625 82.125 140.785 ;
        RECT 83.055 140.625 83.225 141.470 ;
        RECT 84.120 141.185 84.290 141.685 ;
        RECT 84.460 141.355 84.790 141.855 ;
        RECT 83.395 140.795 83.895 141.175 ;
        RECT 84.120 141.015 84.815 141.185 ;
        RECT 81.875 140.455 83.225 140.625 ;
        RECT 82.805 140.415 83.225 140.455 ;
        RECT 81.515 139.945 81.935 140.285 ;
        RECT 82.225 139.955 82.635 140.285 ;
        RECT 79.755 139.525 80.605 139.695 ;
        RECT 81.165 139.305 81.485 139.765 ;
        RECT 81.685 139.515 81.935 139.945 ;
        RECT 82.225 139.305 82.635 139.745 ;
        RECT 82.805 139.685 82.975 140.415 ;
        RECT 83.145 139.865 83.495 140.235 ;
        RECT 83.675 139.925 83.895 140.795 ;
        RECT 84.065 140.225 84.475 140.845 ;
        RECT 84.645 140.045 84.815 141.015 ;
        RECT 84.120 139.855 84.815 140.045 ;
        RECT 82.805 139.485 83.820 139.685 ;
        RECT 84.120 139.525 84.290 139.855 ;
        RECT 84.460 139.305 84.790 139.685 ;
        RECT 85.005 139.565 85.230 141.685 ;
        RECT 85.400 141.355 85.730 141.855 ;
        RECT 85.900 141.185 86.070 141.685 ;
        RECT 85.405 141.015 86.070 141.185 ;
        RECT 85.405 140.025 85.635 141.015 ;
        RECT 85.805 140.195 86.155 140.845 ;
        RECT 86.330 140.690 86.620 141.855 ;
        RECT 86.850 140.715 87.060 141.855 ;
        RECT 87.230 140.705 87.560 141.685 ;
        RECT 87.730 140.715 87.960 141.855 ;
        RECT 88.170 140.765 90.760 141.855 ;
        RECT 85.405 139.855 86.070 140.025 ;
        RECT 85.400 139.305 85.730 139.685 ;
        RECT 85.900 139.565 86.070 139.855 ;
        RECT 86.330 139.305 86.620 140.030 ;
        RECT 86.850 139.305 87.060 140.125 ;
        RECT 87.230 140.105 87.480 140.705 ;
        RECT 87.650 140.295 87.980 140.545 ;
        RECT 88.170 140.245 89.380 140.765 ;
        RECT 90.930 140.715 91.200 141.685 ;
        RECT 91.410 141.055 91.690 141.855 ;
        RECT 91.860 141.345 93.515 141.635 ;
        RECT 91.925 141.005 93.515 141.175 ;
        RECT 91.925 140.885 92.095 141.005 ;
        RECT 91.370 140.715 92.095 140.885 ;
        RECT 87.230 139.475 87.560 140.105 ;
        RECT 87.730 139.305 87.960 140.125 ;
        RECT 89.550 140.075 90.760 140.595 ;
        RECT 88.170 139.305 90.760 140.075 ;
        RECT 90.930 139.980 91.100 140.715 ;
        RECT 91.370 140.545 91.540 140.715 ;
        RECT 92.285 140.665 93.000 140.835 ;
        RECT 93.195 140.715 93.515 141.005 ;
        RECT 93.690 140.715 94.030 141.685 ;
        RECT 94.200 140.715 94.370 141.855 ;
        RECT 94.640 141.055 94.890 141.855 ;
        RECT 95.535 140.885 95.865 141.685 ;
        RECT 96.165 141.055 96.495 141.855 ;
        RECT 96.665 140.885 96.995 141.685 ;
        RECT 94.560 140.715 96.995 140.885 ;
        RECT 97.370 141.095 97.885 141.505 ;
        RECT 98.120 141.095 98.290 141.855 ;
        RECT 98.460 141.515 100.490 141.685 ;
        RECT 91.270 140.215 91.540 140.545 ;
        RECT 91.710 140.215 92.115 140.545 ;
        RECT 92.285 140.215 92.995 140.665 ;
        RECT 91.370 140.045 91.540 140.215 ;
        RECT 90.930 139.635 91.200 139.980 ;
        RECT 91.370 139.875 92.980 140.045 ;
        RECT 93.165 139.975 93.515 140.545 ;
        RECT 93.690 140.155 93.865 140.715 ;
        RECT 94.560 140.465 94.730 140.715 ;
        RECT 94.035 140.295 94.730 140.465 ;
        RECT 94.905 140.295 95.325 140.495 ;
        RECT 95.495 140.295 95.825 140.495 ;
        RECT 95.995 140.295 96.325 140.495 ;
        RECT 93.690 140.105 93.920 140.155 ;
        RECT 91.390 139.305 91.770 139.705 ;
        RECT 91.940 139.525 92.110 139.875 ;
        RECT 92.280 139.305 92.610 139.705 ;
        RECT 92.810 139.525 92.980 139.875 ;
        RECT 93.180 139.305 93.510 139.805 ;
        RECT 93.690 139.475 94.030 140.105 ;
        RECT 94.200 139.305 94.450 140.105 ;
        RECT 94.640 139.955 95.865 140.125 ;
        RECT 94.640 139.475 94.970 139.955 ;
        RECT 95.140 139.305 95.365 139.765 ;
        RECT 95.535 139.475 95.865 139.955 ;
        RECT 96.495 140.085 96.665 140.715 ;
        RECT 96.850 140.295 97.200 140.545 ;
        RECT 97.370 140.285 97.710 141.095 ;
        RECT 98.460 140.850 98.630 141.515 ;
        RECT 99.025 141.175 100.150 141.345 ;
        RECT 97.880 140.660 98.630 140.850 ;
        RECT 98.800 140.835 99.810 141.005 ;
        RECT 97.370 140.115 98.600 140.285 ;
        RECT 96.495 139.475 96.995 140.085 ;
        RECT 97.645 139.510 97.890 140.115 ;
        RECT 98.110 139.305 98.620 139.840 ;
        RECT 98.800 139.475 98.990 140.835 ;
        RECT 99.160 140.495 99.435 140.635 ;
        RECT 99.160 140.325 99.440 140.495 ;
        RECT 99.160 139.475 99.435 140.325 ;
        RECT 99.640 140.035 99.810 140.835 ;
        RECT 99.980 140.045 100.150 141.175 ;
        RECT 100.320 140.545 100.490 141.515 ;
        RECT 100.660 140.715 100.830 141.855 ;
        RECT 101.000 140.715 101.335 141.685 ;
        RECT 100.320 140.215 100.515 140.545 ;
        RECT 100.740 140.215 100.995 140.545 ;
        RECT 100.740 140.045 100.910 140.215 ;
        RECT 101.165 140.045 101.335 140.715 ;
        RECT 101.885 140.875 102.140 141.545 ;
        RECT 102.320 141.055 102.605 141.855 ;
        RECT 102.785 141.135 103.115 141.645 ;
        RECT 101.885 140.155 102.065 140.875 ;
        RECT 102.785 140.545 103.035 141.135 ;
        RECT 103.385 140.985 103.555 141.595 ;
        RECT 103.725 141.165 104.055 141.855 ;
        RECT 104.285 141.305 104.525 141.595 ;
        RECT 104.725 141.475 105.145 141.855 ;
        RECT 105.325 141.385 105.955 141.635 ;
        RECT 106.425 141.475 106.755 141.855 ;
        RECT 105.325 141.305 105.495 141.385 ;
        RECT 106.925 141.305 107.095 141.595 ;
        RECT 107.275 141.475 107.655 141.855 ;
        RECT 107.895 141.470 108.725 141.640 ;
        RECT 104.285 141.135 105.495 141.305 ;
        RECT 102.235 140.215 103.035 140.545 ;
        RECT 99.980 139.875 100.910 140.045 ;
        RECT 99.980 139.840 100.155 139.875 ;
        RECT 99.625 139.475 100.155 139.840 ;
        RECT 100.580 139.305 100.910 139.705 ;
        RECT 101.080 139.475 101.335 140.045 ;
        RECT 101.800 140.015 102.065 140.155 ;
        RECT 101.800 139.985 102.140 140.015 ;
        RECT 101.885 139.485 102.140 139.985 ;
        RECT 102.320 139.305 102.605 139.765 ;
        RECT 102.785 139.565 103.035 140.215 ;
        RECT 103.235 140.965 103.555 140.985 ;
        RECT 103.235 140.795 105.155 140.965 ;
        RECT 103.235 139.900 103.425 140.795 ;
        RECT 105.325 140.625 105.495 141.135 ;
        RECT 105.665 140.875 106.185 141.185 ;
        RECT 103.595 140.455 105.495 140.625 ;
        RECT 103.595 140.395 103.925 140.455 ;
        RECT 104.075 140.225 104.405 140.285 ;
        RECT 103.745 139.955 104.405 140.225 ;
        RECT 103.235 139.570 103.555 139.900 ;
        RECT 103.735 139.305 104.395 139.785 ;
        RECT 104.595 139.695 104.765 140.455 ;
        RECT 105.665 140.285 105.845 140.695 ;
        RECT 104.935 140.115 105.265 140.235 ;
        RECT 106.015 140.115 106.185 140.875 ;
        RECT 104.935 139.945 106.185 140.115 ;
        RECT 106.355 141.055 107.725 141.305 ;
        RECT 106.355 140.285 106.545 141.055 ;
        RECT 107.475 140.795 107.725 141.055 ;
        RECT 106.715 140.625 106.965 140.785 ;
        RECT 107.895 140.625 108.065 141.470 ;
        RECT 108.960 141.185 109.130 141.685 ;
        RECT 109.300 141.355 109.630 141.855 ;
        RECT 108.235 140.795 108.735 141.175 ;
        RECT 108.960 141.015 109.655 141.185 ;
        RECT 106.715 140.455 108.065 140.625 ;
        RECT 107.645 140.415 108.065 140.455 ;
        RECT 106.355 139.945 106.775 140.285 ;
        RECT 107.065 139.955 107.475 140.285 ;
        RECT 104.595 139.525 105.445 139.695 ;
        RECT 106.005 139.305 106.325 139.765 ;
        RECT 106.525 139.515 106.775 139.945 ;
        RECT 107.065 139.305 107.475 139.745 ;
        RECT 107.645 139.685 107.815 140.415 ;
        RECT 107.985 139.865 108.335 140.235 ;
        RECT 108.515 139.925 108.735 140.795 ;
        RECT 108.905 140.225 109.315 140.845 ;
        RECT 109.485 140.045 109.655 141.015 ;
        RECT 108.960 139.855 109.655 140.045 ;
        RECT 107.645 139.485 108.660 139.685 ;
        RECT 108.960 139.525 109.130 139.855 ;
        RECT 109.300 139.305 109.630 139.685 ;
        RECT 109.845 139.565 110.070 141.685 ;
        RECT 110.240 141.355 110.570 141.855 ;
        RECT 110.740 141.185 110.910 141.685 ;
        RECT 110.245 141.015 110.910 141.185 ;
        RECT 110.245 140.025 110.475 141.015 ;
        RECT 110.645 140.195 110.995 140.845 ;
        RECT 111.170 140.765 112.380 141.855 ;
        RECT 111.170 140.225 111.690 140.765 ;
        RECT 111.860 140.055 112.380 140.595 ;
        RECT 110.245 139.855 110.910 140.025 ;
        RECT 110.240 139.305 110.570 139.685 ;
        RECT 110.740 139.565 110.910 139.855 ;
        RECT 111.170 139.305 112.380 140.055 ;
        RECT 18.165 139.135 112.465 139.305 ;
        RECT 18.250 138.385 19.460 139.135 ;
        RECT 18.250 137.845 18.770 138.385 ;
        RECT 20.090 138.365 21.760 139.135 ;
        RECT 21.930 138.410 22.220 139.135 ;
        RECT 23.310 138.365 26.820 139.135 ;
        RECT 26.995 138.590 32.340 139.135 ;
        RECT 32.520 138.635 32.850 139.135 ;
        RECT 18.940 137.675 19.460 138.215 ;
        RECT 18.250 136.585 19.460 137.675 ;
        RECT 20.090 137.675 20.840 138.195 ;
        RECT 21.010 137.845 21.760 138.365 ;
        RECT 20.090 136.585 21.760 137.675 ;
        RECT 21.930 136.585 22.220 137.750 ;
        RECT 23.310 137.675 25.000 138.195 ;
        RECT 25.170 137.845 26.820 138.365 ;
        RECT 23.310 136.585 26.820 137.675 ;
        RECT 28.585 137.020 28.935 138.270 ;
        RECT 30.415 137.760 30.755 138.590 ;
        RECT 33.050 138.565 33.220 138.915 ;
        RECT 33.420 138.735 33.750 139.135 ;
        RECT 33.920 138.565 34.090 138.915 ;
        RECT 34.260 138.735 34.640 139.135 ;
        RECT 32.515 137.895 32.865 138.465 ;
        RECT 33.050 138.395 34.660 138.565 ;
        RECT 34.830 138.460 35.100 138.805 ;
        RECT 34.490 138.225 34.660 138.395 ;
        RECT 32.515 137.435 32.835 137.725 ;
        RECT 33.035 137.605 33.745 138.225 ;
        RECT 33.915 137.895 34.320 138.225 ;
        RECT 34.490 137.895 34.760 138.225 ;
        RECT 34.490 137.725 34.660 137.895 ;
        RECT 34.930 137.725 35.100 138.460 ;
        RECT 35.270 138.365 37.860 139.135 ;
        RECT 33.935 137.555 34.660 137.725 ;
        RECT 33.935 137.435 34.105 137.555 ;
        RECT 32.515 137.265 34.105 137.435 ;
        RECT 26.995 136.585 32.340 137.020 ;
        RECT 32.515 136.805 34.170 137.095 ;
        RECT 34.340 136.585 34.620 137.385 ;
        RECT 34.830 136.755 35.100 137.725 ;
        RECT 35.270 137.675 36.480 138.195 ;
        RECT 36.650 137.845 37.860 138.365 ;
        RECT 38.030 138.335 38.370 138.965 ;
        RECT 38.540 138.335 38.790 139.135 ;
        RECT 38.980 138.485 39.310 138.965 ;
        RECT 39.480 138.675 39.705 139.135 ;
        RECT 39.875 138.485 40.205 138.965 ;
        RECT 38.030 138.285 38.260 138.335 ;
        RECT 38.980 138.315 40.205 138.485 ;
        RECT 40.835 138.355 41.335 138.965 ;
        RECT 41.710 138.365 43.380 139.135 ;
        RECT 43.640 138.585 43.810 138.965 ;
        RECT 43.990 138.755 44.320 139.135 ;
        RECT 43.640 138.415 44.305 138.585 ;
        RECT 44.500 138.460 44.760 138.965 ;
        RECT 38.030 137.725 38.205 138.285 ;
        RECT 38.375 137.975 39.070 138.145 ;
        RECT 38.900 137.725 39.070 137.975 ;
        RECT 39.245 137.945 39.665 138.145 ;
        RECT 39.835 137.945 40.165 138.145 ;
        RECT 40.335 137.945 40.665 138.145 ;
        RECT 40.835 137.725 41.005 138.355 ;
        RECT 41.190 137.895 41.540 138.145 ;
        RECT 35.270 136.585 37.860 137.675 ;
        RECT 38.030 136.755 38.370 137.725 ;
        RECT 38.540 136.585 38.710 137.725 ;
        RECT 38.900 137.555 41.335 137.725 ;
        RECT 38.980 136.585 39.230 137.385 ;
        RECT 39.875 136.755 40.205 137.555 ;
        RECT 40.505 136.585 40.835 137.385 ;
        RECT 41.005 136.755 41.335 137.555 ;
        RECT 41.710 137.675 42.460 138.195 ;
        RECT 42.630 137.845 43.380 138.365 ;
        RECT 43.570 137.865 43.900 138.235 ;
        RECT 44.135 138.160 44.305 138.415 ;
        RECT 44.135 137.830 44.420 138.160 ;
        RECT 44.135 137.685 44.305 137.830 ;
        RECT 41.710 136.585 43.380 137.675 ;
        RECT 43.640 137.515 44.305 137.685 ;
        RECT 44.590 137.660 44.760 138.460 ;
        RECT 43.640 136.755 43.810 137.515 ;
        RECT 43.990 136.585 44.320 137.345 ;
        RECT 44.490 136.755 44.760 137.660 ;
        RECT 44.930 138.460 45.200 138.805 ;
        RECT 45.390 138.735 45.770 139.135 ;
        RECT 45.940 138.565 46.110 138.915 ;
        RECT 46.280 138.735 46.610 139.135 ;
        RECT 46.810 138.565 46.980 138.915 ;
        RECT 47.180 138.635 47.510 139.135 ;
        RECT 44.930 137.725 45.100 138.460 ;
        RECT 45.370 138.395 46.980 138.565 ;
        RECT 45.370 138.225 45.540 138.395 ;
        RECT 45.270 137.895 45.540 138.225 ;
        RECT 45.710 137.895 46.115 138.225 ;
        RECT 45.370 137.725 45.540 137.895 ;
        RECT 46.285 137.775 46.995 138.225 ;
        RECT 47.165 137.895 47.515 138.465 ;
        RECT 47.690 138.410 47.980 139.135 ;
        RECT 48.150 138.365 50.740 139.135 ;
        RECT 50.915 138.590 56.260 139.135 ;
        RECT 44.930 136.755 45.200 137.725 ;
        RECT 45.370 137.555 46.095 137.725 ;
        RECT 46.285 137.605 47.000 137.775 ;
        RECT 45.925 137.435 46.095 137.555 ;
        RECT 47.195 137.435 47.515 137.725 ;
        RECT 45.410 136.585 45.690 137.385 ;
        RECT 45.925 137.265 47.515 137.435 ;
        RECT 45.860 136.805 47.515 137.095 ;
        RECT 47.690 136.585 47.980 137.750 ;
        RECT 48.150 137.675 49.360 138.195 ;
        RECT 49.530 137.845 50.740 138.365 ;
        RECT 48.150 136.585 50.740 137.675 ;
        RECT 52.505 137.020 52.855 138.270 ;
        RECT 54.335 137.760 54.675 138.590 ;
        RECT 56.430 138.335 56.770 138.965 ;
        RECT 56.940 138.335 57.190 139.135 ;
        RECT 57.380 138.485 57.710 138.965 ;
        RECT 57.880 138.675 58.105 139.135 ;
        RECT 58.275 138.485 58.605 138.965 ;
        RECT 56.430 138.285 56.660 138.335 ;
        RECT 57.380 138.315 58.605 138.485 ;
        RECT 59.235 138.355 59.735 138.965 ;
        RECT 56.430 137.725 56.605 138.285 ;
        RECT 56.775 137.975 57.470 138.145 ;
        RECT 57.300 137.725 57.470 137.975 ;
        RECT 57.645 137.945 58.065 138.145 ;
        RECT 58.235 137.945 58.565 138.145 ;
        RECT 58.735 137.945 59.065 138.145 ;
        RECT 59.235 137.725 59.405 138.355 ;
        RECT 61.305 138.325 61.550 138.930 ;
        RECT 61.770 138.600 62.280 139.135 ;
        RECT 61.030 138.155 62.260 138.325 ;
        RECT 59.590 137.895 59.940 138.145 ;
        RECT 50.915 136.585 56.260 137.020 ;
        RECT 56.430 136.755 56.770 137.725 ;
        RECT 56.940 136.585 57.110 137.725 ;
        RECT 57.300 137.555 59.735 137.725 ;
        RECT 57.380 136.585 57.630 137.385 ;
        RECT 58.275 136.755 58.605 137.555 ;
        RECT 58.905 136.585 59.235 137.385 ;
        RECT 59.405 136.755 59.735 137.555 ;
        RECT 61.030 137.345 61.370 138.155 ;
        RECT 61.540 137.590 62.290 137.780 ;
        RECT 61.030 136.935 61.545 137.345 ;
        RECT 61.780 136.585 61.950 137.345 ;
        RECT 62.120 136.925 62.290 137.590 ;
        RECT 62.460 137.605 62.650 138.965 ;
        RECT 62.820 138.455 63.095 138.965 ;
        RECT 63.285 138.600 63.815 138.965 ;
        RECT 64.240 138.735 64.570 139.135 ;
        RECT 63.640 138.565 63.815 138.600 ;
        RECT 62.820 138.285 63.100 138.455 ;
        RECT 62.820 137.805 63.095 138.285 ;
        RECT 63.300 137.605 63.470 138.405 ;
        RECT 62.460 137.435 63.470 137.605 ;
        RECT 63.640 138.395 64.570 138.565 ;
        RECT 64.740 138.395 64.995 138.965 ;
        RECT 63.640 137.265 63.810 138.395 ;
        RECT 64.400 138.225 64.570 138.395 ;
        RECT 62.685 137.095 63.810 137.265 ;
        RECT 63.980 137.895 64.175 138.225 ;
        RECT 64.400 137.895 64.655 138.225 ;
        RECT 63.980 136.925 64.150 137.895 ;
        RECT 64.825 137.725 64.995 138.395 ;
        RECT 62.120 136.755 64.150 136.925 ;
        RECT 64.320 136.585 64.490 137.725 ;
        RECT 64.660 136.755 64.995 137.725 ;
        RECT 65.170 138.460 65.430 138.965 ;
        RECT 65.610 138.755 65.940 139.135 ;
        RECT 66.120 138.585 66.290 138.965 ;
        RECT 65.170 137.660 65.350 138.460 ;
        RECT 65.625 138.415 66.290 138.585 ;
        RECT 65.625 138.160 65.795 138.415 ;
        RECT 66.610 138.315 66.820 139.135 ;
        RECT 66.990 138.335 67.320 138.965 ;
        RECT 65.520 137.830 65.795 138.160 ;
        RECT 66.020 137.865 66.360 138.235 ;
        RECT 65.625 137.685 65.795 137.830 ;
        RECT 66.990 137.735 67.240 138.335 ;
        RECT 67.490 138.315 67.720 139.135 ;
        RECT 68.020 138.585 68.190 138.965 ;
        RECT 68.370 138.755 68.700 139.135 ;
        RECT 68.020 138.415 68.685 138.585 ;
        RECT 68.880 138.460 69.140 138.965 ;
        RECT 67.410 137.895 67.740 138.145 ;
        RECT 67.950 137.865 68.280 138.235 ;
        RECT 68.515 138.160 68.685 138.415 ;
        RECT 68.515 137.830 68.800 138.160 ;
        RECT 65.170 136.755 65.440 137.660 ;
        RECT 65.625 137.515 66.300 137.685 ;
        RECT 65.610 136.585 65.940 137.345 ;
        RECT 66.120 136.755 66.300 137.515 ;
        RECT 66.610 136.585 66.820 137.725 ;
        RECT 66.990 136.755 67.320 137.735 ;
        RECT 67.490 136.585 67.720 137.725 ;
        RECT 68.515 137.685 68.685 137.830 ;
        RECT 68.020 137.515 68.685 137.685 ;
        RECT 68.970 137.660 69.140 138.460 ;
        RECT 69.310 138.385 70.520 139.135 ;
        RECT 68.020 136.755 68.190 137.515 ;
        RECT 68.370 136.585 68.700 137.345 ;
        RECT 68.870 136.755 69.140 137.660 ;
        RECT 69.310 137.675 69.830 138.215 ;
        RECT 70.000 137.845 70.520 138.385 ;
        RECT 70.690 138.460 70.960 138.805 ;
        RECT 71.150 138.735 71.530 139.135 ;
        RECT 71.700 138.565 71.870 138.915 ;
        RECT 72.040 138.735 72.370 139.135 ;
        RECT 72.570 138.565 72.740 138.915 ;
        RECT 72.940 138.635 73.270 139.135 ;
        RECT 70.690 137.725 70.860 138.460 ;
        RECT 71.130 138.395 72.740 138.565 ;
        RECT 71.130 138.225 71.300 138.395 ;
        RECT 71.030 137.895 71.300 138.225 ;
        RECT 71.470 137.895 71.875 138.225 ;
        RECT 71.130 137.725 71.300 137.895 ;
        RECT 72.045 137.775 72.755 138.225 ;
        RECT 72.925 137.895 73.275 138.465 ;
        RECT 73.450 138.410 73.740 139.135 ;
        RECT 74.830 138.365 78.340 139.135 ;
        RECT 69.310 136.585 70.520 137.675 ;
        RECT 70.690 136.755 70.960 137.725 ;
        RECT 71.130 137.555 71.855 137.725 ;
        RECT 72.045 137.605 72.760 137.775 ;
        RECT 71.685 137.435 71.855 137.555 ;
        RECT 72.955 137.435 73.275 137.725 ;
        RECT 71.170 136.585 71.450 137.385 ;
        RECT 71.685 137.265 73.275 137.435 ;
        RECT 71.620 136.805 73.275 137.095 ;
        RECT 73.450 136.585 73.740 137.750 ;
        RECT 74.830 137.675 76.520 138.195 ;
        RECT 76.690 137.845 78.340 138.365 ;
        RECT 78.785 138.325 79.030 138.930 ;
        RECT 79.250 138.600 79.760 139.135 ;
        RECT 78.510 138.155 79.740 138.325 ;
        RECT 74.830 136.585 78.340 137.675 ;
        RECT 78.510 137.345 78.850 138.155 ;
        RECT 79.020 137.590 79.770 137.780 ;
        RECT 78.510 136.935 79.025 137.345 ;
        RECT 79.260 136.585 79.430 137.345 ;
        RECT 79.600 136.925 79.770 137.590 ;
        RECT 79.940 137.605 80.130 138.965 ;
        RECT 80.300 138.115 80.575 138.965 ;
        RECT 80.765 138.600 81.295 138.965 ;
        RECT 81.720 138.735 82.050 139.135 ;
        RECT 81.120 138.565 81.295 138.600 ;
        RECT 80.300 137.945 80.580 138.115 ;
        RECT 80.300 137.805 80.575 137.945 ;
        RECT 80.780 137.605 80.950 138.405 ;
        RECT 79.940 137.435 80.950 137.605 ;
        RECT 81.120 138.395 82.050 138.565 ;
        RECT 82.220 138.395 82.475 138.965 ;
        RECT 82.740 138.585 82.910 138.965 ;
        RECT 83.090 138.755 83.420 139.135 ;
        RECT 82.740 138.415 83.405 138.585 ;
        RECT 83.600 138.460 83.860 138.965 ;
        RECT 81.120 137.265 81.290 138.395 ;
        RECT 81.880 138.225 82.050 138.395 ;
        RECT 80.165 137.095 81.290 137.265 ;
        RECT 81.460 137.895 81.655 138.225 ;
        RECT 81.880 137.895 82.135 138.225 ;
        RECT 81.460 136.925 81.630 137.895 ;
        RECT 82.305 137.725 82.475 138.395 ;
        RECT 82.670 137.865 83.000 138.235 ;
        RECT 83.235 138.160 83.405 138.415 ;
        RECT 79.600 136.755 81.630 136.925 ;
        RECT 81.800 136.585 81.970 137.725 ;
        RECT 82.140 136.755 82.475 137.725 ;
        RECT 83.235 137.830 83.520 138.160 ;
        RECT 83.235 137.685 83.405 137.830 ;
        RECT 82.740 137.515 83.405 137.685 ;
        RECT 83.690 137.660 83.860 138.460 ;
        RECT 82.740 136.755 82.910 137.515 ;
        RECT 83.090 136.585 83.420 137.345 ;
        RECT 83.590 136.755 83.860 137.660 ;
        RECT 84.030 138.460 84.300 138.805 ;
        RECT 84.490 138.735 84.870 139.135 ;
        RECT 85.040 138.565 85.210 138.915 ;
        RECT 85.380 138.735 85.710 139.135 ;
        RECT 85.910 138.565 86.080 138.915 ;
        RECT 86.280 138.635 86.610 139.135 ;
        RECT 84.030 137.725 84.200 138.460 ;
        RECT 84.470 138.395 86.080 138.565 ;
        RECT 84.470 138.225 84.640 138.395 ;
        RECT 84.370 137.895 84.640 138.225 ;
        RECT 84.810 137.895 85.215 138.225 ;
        RECT 84.470 137.725 84.640 137.895 ;
        RECT 85.385 137.775 86.095 138.225 ;
        RECT 86.265 137.895 86.615 138.465 ;
        RECT 86.995 138.355 87.495 138.965 ;
        RECT 86.790 137.895 87.140 138.145 ;
        RECT 84.030 136.755 84.300 137.725 ;
        RECT 84.470 137.555 85.195 137.725 ;
        RECT 85.385 137.605 86.100 137.775 ;
        RECT 87.325 137.725 87.495 138.355 ;
        RECT 88.125 138.485 88.455 138.965 ;
        RECT 88.625 138.675 88.850 139.135 ;
        RECT 89.020 138.485 89.350 138.965 ;
        RECT 88.125 138.315 89.350 138.485 ;
        RECT 89.540 138.335 89.790 139.135 ;
        RECT 89.960 138.335 90.300 138.965 ;
        RECT 87.665 137.945 87.995 138.145 ;
        RECT 88.165 137.945 88.495 138.145 ;
        RECT 88.665 137.945 89.085 138.145 ;
        RECT 89.260 137.975 89.955 138.145 ;
        RECT 89.260 137.725 89.430 137.975 ;
        RECT 90.125 137.725 90.300 138.335 ;
        RECT 85.025 137.435 85.195 137.555 ;
        RECT 86.295 137.435 86.615 137.725 ;
        RECT 84.510 136.585 84.790 137.385 ;
        RECT 85.025 137.265 86.615 137.435 ;
        RECT 86.995 137.555 89.430 137.725 ;
        RECT 84.960 136.805 86.615 137.095 ;
        RECT 86.995 136.755 87.325 137.555 ;
        RECT 87.495 136.585 87.825 137.385 ;
        RECT 88.125 136.755 88.455 137.555 ;
        RECT 89.100 136.585 89.350 137.385 ;
        RECT 89.620 136.585 89.790 137.725 ;
        RECT 89.960 136.755 90.300 137.725 ;
        RECT 90.470 138.335 90.810 138.965 ;
        RECT 90.980 138.335 91.230 139.135 ;
        RECT 91.420 138.485 91.750 138.965 ;
        RECT 91.920 138.675 92.145 139.135 ;
        RECT 92.315 138.485 92.645 138.965 ;
        RECT 90.470 138.285 90.700 138.335 ;
        RECT 91.420 138.315 92.645 138.485 ;
        RECT 93.275 138.355 93.775 138.965 ;
        RECT 90.470 137.725 90.645 138.285 ;
        RECT 90.815 137.975 91.510 138.145 ;
        RECT 91.340 137.725 91.510 137.975 ;
        RECT 91.685 137.945 92.105 138.145 ;
        RECT 92.275 137.945 92.605 138.145 ;
        RECT 92.775 137.945 93.105 138.145 ;
        RECT 93.275 137.725 93.445 138.355 ;
        RECT 95.345 138.325 95.590 138.930 ;
        RECT 95.810 138.600 96.320 139.135 ;
        RECT 95.070 138.155 96.300 138.325 ;
        RECT 93.630 137.895 93.980 138.145 ;
        RECT 90.470 136.755 90.810 137.725 ;
        RECT 90.980 136.585 91.150 137.725 ;
        RECT 91.340 137.555 93.775 137.725 ;
        RECT 91.420 136.585 91.670 137.385 ;
        RECT 92.315 136.755 92.645 137.555 ;
        RECT 92.945 136.585 93.275 137.385 ;
        RECT 93.445 136.755 93.775 137.555 ;
        RECT 95.070 137.345 95.410 138.155 ;
        RECT 95.580 137.590 96.330 137.780 ;
        RECT 95.070 136.935 95.585 137.345 ;
        RECT 95.820 136.585 95.990 137.345 ;
        RECT 96.160 136.925 96.330 137.590 ;
        RECT 96.500 137.605 96.690 138.965 ;
        RECT 96.860 138.795 97.135 138.965 ;
        RECT 96.860 138.625 97.140 138.795 ;
        RECT 96.860 137.805 97.135 138.625 ;
        RECT 97.325 138.600 97.855 138.965 ;
        RECT 98.280 138.735 98.610 139.135 ;
        RECT 97.680 138.565 97.855 138.600 ;
        RECT 97.340 137.605 97.510 138.405 ;
        RECT 96.500 137.435 97.510 137.605 ;
        RECT 97.680 138.395 98.610 138.565 ;
        RECT 98.780 138.395 99.035 138.965 ;
        RECT 99.210 138.410 99.500 139.135 ;
        RECT 97.680 137.265 97.850 138.395 ;
        RECT 98.440 138.225 98.610 138.395 ;
        RECT 96.725 137.095 97.850 137.265 ;
        RECT 98.020 137.895 98.215 138.225 ;
        RECT 98.440 137.895 98.695 138.225 ;
        RECT 98.020 136.925 98.190 137.895 ;
        RECT 98.865 137.725 99.035 138.395 ;
        RECT 100.170 138.315 100.400 139.135 ;
        RECT 100.570 138.335 100.900 138.965 ;
        RECT 100.150 137.895 100.480 138.145 ;
        RECT 96.160 136.755 98.190 136.925 ;
        RECT 98.360 136.585 98.530 137.725 ;
        RECT 98.700 136.755 99.035 137.725 ;
        RECT 99.210 136.585 99.500 137.750 ;
        RECT 100.650 137.735 100.900 138.335 ;
        RECT 101.070 138.315 101.280 139.135 ;
        RECT 101.885 138.425 102.140 138.955 ;
        RECT 102.320 138.675 102.605 139.135 ;
        RECT 100.170 136.585 100.400 137.725 ;
        RECT 100.570 136.755 100.900 137.735 ;
        RECT 101.070 136.585 101.280 137.725 ;
        RECT 101.885 137.565 102.065 138.425 ;
        RECT 102.785 138.225 103.035 138.875 ;
        RECT 102.235 137.895 103.035 138.225 ;
        RECT 101.885 137.435 102.140 137.565 ;
        RECT 101.800 137.265 102.140 137.435 ;
        RECT 101.885 136.895 102.140 137.265 ;
        RECT 102.320 136.585 102.605 137.385 ;
        RECT 102.785 137.305 103.035 137.895 ;
        RECT 103.235 138.540 103.555 138.870 ;
        RECT 103.735 138.655 104.395 139.135 ;
        RECT 104.595 138.745 105.445 138.915 ;
        RECT 103.235 137.645 103.425 138.540 ;
        RECT 103.745 138.215 104.405 138.485 ;
        RECT 104.075 138.155 104.405 138.215 ;
        RECT 103.595 137.985 103.925 138.045 ;
        RECT 104.595 137.985 104.765 138.745 ;
        RECT 106.005 138.675 106.325 139.135 ;
        RECT 106.525 138.495 106.775 138.925 ;
        RECT 107.065 138.695 107.475 139.135 ;
        RECT 107.645 138.755 108.660 138.955 ;
        RECT 104.935 138.325 106.185 138.495 ;
        RECT 104.935 138.205 105.265 138.325 ;
        RECT 103.595 137.815 105.495 137.985 ;
        RECT 103.235 137.475 105.155 137.645 ;
        RECT 103.235 137.455 103.555 137.475 ;
        RECT 102.785 136.795 103.115 137.305 ;
        RECT 103.385 136.845 103.555 137.455 ;
        RECT 105.325 137.305 105.495 137.815 ;
        RECT 105.665 137.745 105.845 138.155 ;
        RECT 106.015 137.565 106.185 138.325 ;
        RECT 103.725 136.585 104.055 137.275 ;
        RECT 104.285 137.135 105.495 137.305 ;
        RECT 105.665 137.255 106.185 137.565 ;
        RECT 106.355 138.155 106.775 138.495 ;
        RECT 107.065 138.155 107.475 138.485 ;
        RECT 106.355 137.385 106.545 138.155 ;
        RECT 107.645 138.025 107.815 138.755 ;
        RECT 108.960 138.585 109.130 138.915 ;
        RECT 109.300 138.755 109.630 139.135 ;
        RECT 107.985 138.205 108.335 138.575 ;
        RECT 107.645 137.985 108.065 138.025 ;
        RECT 106.715 137.815 108.065 137.985 ;
        RECT 106.715 137.655 106.965 137.815 ;
        RECT 107.475 137.385 107.725 137.645 ;
        RECT 106.355 137.135 107.725 137.385 ;
        RECT 104.285 136.845 104.525 137.135 ;
        RECT 105.325 137.055 105.495 137.135 ;
        RECT 104.725 136.585 105.145 136.965 ;
        RECT 105.325 136.805 105.955 137.055 ;
        RECT 106.425 136.585 106.755 136.965 ;
        RECT 106.925 136.845 107.095 137.135 ;
        RECT 107.895 136.970 108.065 137.815 ;
        RECT 108.515 137.645 108.735 138.515 ;
        RECT 108.960 138.395 109.655 138.585 ;
        RECT 108.235 137.265 108.735 137.645 ;
        RECT 108.905 137.595 109.315 138.215 ;
        RECT 109.485 137.425 109.655 138.395 ;
        RECT 108.960 137.255 109.655 137.425 ;
        RECT 107.275 136.585 107.655 136.965 ;
        RECT 107.895 136.800 108.725 136.970 ;
        RECT 108.960 136.755 109.130 137.255 ;
        RECT 109.300 136.585 109.630 137.085 ;
        RECT 109.845 136.755 110.070 138.875 ;
        RECT 110.240 138.755 110.570 139.135 ;
        RECT 110.740 138.585 110.910 138.875 ;
        RECT 110.245 138.415 110.910 138.585 ;
        RECT 110.245 137.425 110.475 138.415 ;
        RECT 111.170 138.385 112.380 139.135 ;
        RECT 110.645 137.595 110.995 138.245 ;
        RECT 111.170 137.675 111.690 138.215 ;
        RECT 111.860 137.845 112.380 138.385 ;
        RECT 110.245 137.255 110.910 137.425 ;
        RECT 110.240 136.585 110.570 137.085 ;
        RECT 110.740 136.755 110.910 137.255 ;
        RECT 111.170 136.585 112.380 137.675 ;
        RECT 18.165 136.415 112.465 136.585 ;
        RECT 18.250 135.325 19.460 136.415 ;
        RECT 18.250 134.615 18.770 135.155 ;
        RECT 18.940 134.785 19.460 135.325 ;
        RECT 19.630 135.325 20.840 136.415 ;
        RECT 21.015 135.980 26.360 136.415 ;
        RECT 26.535 135.980 31.880 136.415 ;
        RECT 19.630 134.785 20.150 135.325 ;
        RECT 20.320 134.615 20.840 135.155 ;
        RECT 22.605 134.730 22.955 135.980 ;
        RECT 18.250 133.865 19.460 134.615 ;
        RECT 19.630 133.865 20.840 134.615 ;
        RECT 24.435 134.410 24.775 135.240 ;
        RECT 28.125 134.730 28.475 135.980 ;
        RECT 32.055 135.905 33.710 136.195 ;
        RECT 32.055 135.565 33.645 135.735 ;
        RECT 33.880 135.615 34.160 136.415 ;
        RECT 32.055 135.275 32.375 135.565 ;
        RECT 33.475 135.445 33.645 135.565 ;
        RECT 29.955 134.410 30.295 135.240 ;
        RECT 32.055 134.535 32.405 135.105 ;
        RECT 32.575 134.775 33.285 135.395 ;
        RECT 33.475 135.275 34.200 135.445 ;
        RECT 34.370 135.275 34.640 136.245 ;
        RECT 34.030 135.105 34.200 135.275 ;
        RECT 33.455 134.775 33.860 135.105 ;
        RECT 34.030 134.775 34.300 135.105 ;
        RECT 34.030 134.605 34.200 134.775 ;
        RECT 32.590 134.435 34.200 134.605 ;
        RECT 34.470 134.540 34.640 135.275 ;
        RECT 34.810 135.250 35.100 136.415 ;
        RECT 35.730 135.325 37.400 136.415 ;
        RECT 35.730 134.805 36.480 135.325 ;
        RECT 37.610 135.275 37.840 136.415 ;
        RECT 38.010 135.265 38.340 136.245 ;
        RECT 38.510 135.275 38.720 136.415 ;
        RECT 38.950 135.275 39.290 136.245 ;
        RECT 39.460 135.275 39.630 136.415 ;
        RECT 39.900 135.615 40.150 136.415 ;
        RECT 40.795 135.445 41.125 136.245 ;
        RECT 41.425 135.615 41.755 136.415 ;
        RECT 41.925 135.445 42.255 136.245 ;
        RECT 39.820 135.275 42.255 135.445 ;
        RECT 43.090 135.325 45.680 136.415 ;
        RECT 46.225 135.435 46.480 136.105 ;
        RECT 46.660 135.615 46.945 136.415 ;
        RECT 47.125 135.695 47.455 136.205 ;
        RECT 46.225 135.395 46.405 135.435 ;
        RECT 36.650 134.635 37.400 135.155 ;
        RECT 37.590 134.855 37.920 135.105 ;
        RECT 21.015 133.865 26.360 134.410 ;
        RECT 26.535 133.865 31.880 134.410 ;
        RECT 32.060 133.865 32.390 134.365 ;
        RECT 32.590 134.085 32.760 134.435 ;
        RECT 32.960 133.865 33.290 134.265 ;
        RECT 33.460 134.085 33.630 134.435 ;
        RECT 33.800 133.865 34.180 134.265 ;
        RECT 34.370 134.195 34.640 134.540 ;
        RECT 34.810 133.865 35.100 134.590 ;
        RECT 35.730 133.865 37.400 134.635 ;
        RECT 37.610 133.865 37.840 134.685 ;
        RECT 38.090 134.665 38.340 135.265 ;
        RECT 38.950 134.715 39.125 135.275 ;
        RECT 39.820 135.025 39.990 135.275 ;
        RECT 39.295 134.855 39.990 135.025 ;
        RECT 40.165 134.855 40.585 135.055 ;
        RECT 40.755 134.855 41.085 135.055 ;
        RECT 41.255 134.855 41.585 135.055 ;
        RECT 38.010 134.035 38.340 134.665 ;
        RECT 38.510 133.865 38.720 134.685 ;
        RECT 38.950 134.665 39.180 134.715 ;
        RECT 38.950 134.035 39.290 134.665 ;
        RECT 39.460 133.865 39.710 134.665 ;
        RECT 39.900 134.515 41.125 134.685 ;
        RECT 39.900 134.035 40.230 134.515 ;
        RECT 40.400 133.865 40.625 134.325 ;
        RECT 40.795 134.035 41.125 134.515 ;
        RECT 41.755 134.645 41.925 135.275 ;
        RECT 42.110 134.855 42.460 135.105 ;
        RECT 43.090 134.805 44.300 135.325 ;
        RECT 46.140 135.225 46.405 135.395 ;
        RECT 41.755 134.035 42.255 134.645 ;
        RECT 44.470 134.635 45.680 135.155 ;
        RECT 43.090 133.865 45.680 134.635 ;
        RECT 46.225 134.575 46.405 135.225 ;
        RECT 47.125 135.105 47.375 135.695 ;
        RECT 47.725 135.545 47.895 136.155 ;
        RECT 48.065 135.725 48.395 136.415 ;
        RECT 48.625 135.865 48.865 136.155 ;
        RECT 49.065 136.035 49.485 136.415 ;
        RECT 49.665 135.945 50.295 136.195 ;
        RECT 50.765 136.035 51.095 136.415 ;
        RECT 49.665 135.865 49.835 135.945 ;
        RECT 51.265 135.865 51.435 136.155 ;
        RECT 51.615 136.035 51.995 136.415 ;
        RECT 52.235 136.030 53.065 136.200 ;
        RECT 48.625 135.695 49.835 135.865 ;
        RECT 46.575 134.775 47.375 135.105 ;
        RECT 46.225 134.045 46.480 134.575 ;
        RECT 46.660 133.865 46.945 134.325 ;
        RECT 47.125 134.125 47.375 134.775 ;
        RECT 47.575 135.525 47.895 135.545 ;
        RECT 47.575 135.355 49.495 135.525 ;
        RECT 47.575 134.460 47.765 135.355 ;
        RECT 49.665 135.185 49.835 135.695 ;
        RECT 50.005 135.435 50.525 135.745 ;
        RECT 47.935 135.015 49.835 135.185 ;
        RECT 47.935 134.955 48.265 135.015 ;
        RECT 48.415 134.785 48.745 134.845 ;
        RECT 48.085 134.515 48.745 134.785 ;
        RECT 47.575 134.130 47.895 134.460 ;
        RECT 48.075 133.865 48.735 134.345 ;
        RECT 48.935 134.255 49.105 135.015 ;
        RECT 50.005 134.845 50.185 135.255 ;
        RECT 49.275 134.675 49.605 134.795 ;
        RECT 50.355 134.675 50.525 135.435 ;
        RECT 49.275 134.505 50.525 134.675 ;
        RECT 50.695 135.615 52.065 135.865 ;
        RECT 50.695 134.845 50.885 135.615 ;
        RECT 51.815 135.355 52.065 135.615 ;
        RECT 51.055 135.185 51.305 135.345 ;
        RECT 52.235 135.185 52.405 136.030 ;
        RECT 53.300 135.745 53.470 136.245 ;
        RECT 53.640 135.915 53.970 136.415 ;
        RECT 52.575 135.355 53.075 135.735 ;
        RECT 53.300 135.575 53.995 135.745 ;
        RECT 51.055 135.015 52.405 135.185 ;
        RECT 51.985 134.975 52.405 135.015 ;
        RECT 50.695 134.505 51.115 134.845 ;
        RECT 51.405 134.515 51.815 134.845 ;
        RECT 48.935 134.085 49.785 134.255 ;
        RECT 50.345 133.865 50.665 134.325 ;
        RECT 50.865 134.075 51.115 134.505 ;
        RECT 51.405 133.865 51.815 134.305 ;
        RECT 51.985 134.245 52.155 134.975 ;
        RECT 52.325 134.425 52.675 134.795 ;
        RECT 52.855 134.485 53.075 135.355 ;
        RECT 53.245 134.785 53.655 135.405 ;
        RECT 53.825 134.605 53.995 135.575 ;
        RECT 53.300 134.415 53.995 134.605 ;
        RECT 51.985 134.045 53.000 134.245 ;
        RECT 53.300 134.085 53.470 134.415 ;
        RECT 53.640 133.865 53.970 134.245 ;
        RECT 54.185 134.125 54.410 136.245 ;
        RECT 54.580 135.915 54.910 136.415 ;
        RECT 55.080 135.745 55.250 136.245 ;
        RECT 54.585 135.575 55.250 135.745 ;
        RECT 56.430 135.655 56.945 136.065 ;
        RECT 57.180 135.655 57.350 136.415 ;
        RECT 57.520 136.075 59.550 136.245 ;
        RECT 54.585 134.585 54.815 135.575 ;
        RECT 54.985 134.755 55.335 135.405 ;
        RECT 56.430 134.845 56.770 135.655 ;
        RECT 57.520 135.410 57.690 136.075 ;
        RECT 58.085 135.735 59.210 135.905 ;
        RECT 56.940 135.220 57.690 135.410 ;
        RECT 57.860 135.395 58.870 135.565 ;
        RECT 56.430 134.675 57.660 134.845 ;
        RECT 54.585 134.415 55.250 134.585 ;
        RECT 54.580 133.865 54.910 134.245 ;
        RECT 55.080 134.125 55.250 134.415 ;
        RECT 56.705 134.070 56.950 134.675 ;
        RECT 57.170 133.865 57.680 134.400 ;
        RECT 57.860 134.035 58.050 135.395 ;
        RECT 58.220 134.375 58.495 135.195 ;
        RECT 58.700 134.595 58.870 135.395 ;
        RECT 59.040 134.605 59.210 135.735 ;
        RECT 59.380 135.105 59.550 136.075 ;
        RECT 59.720 135.275 59.890 136.415 ;
        RECT 60.060 135.275 60.395 136.245 ;
        RECT 59.380 134.775 59.575 135.105 ;
        RECT 59.800 134.775 60.055 135.105 ;
        RECT 59.800 134.605 59.970 134.775 ;
        RECT 60.225 134.605 60.395 135.275 ;
        RECT 60.570 135.250 60.860 136.415 ;
        RECT 61.405 135.435 61.660 136.105 ;
        RECT 61.840 135.615 62.125 136.415 ;
        RECT 62.305 135.695 62.635 136.205 ;
        RECT 61.405 135.395 61.585 135.435 ;
        RECT 61.320 135.225 61.585 135.395 ;
        RECT 59.040 134.435 59.970 134.605 ;
        RECT 59.040 134.400 59.215 134.435 ;
        RECT 58.220 134.205 58.500 134.375 ;
        RECT 58.220 134.035 58.495 134.205 ;
        RECT 58.685 134.035 59.215 134.400 ;
        RECT 59.640 133.865 59.970 134.265 ;
        RECT 60.140 134.035 60.395 134.605 ;
        RECT 60.570 133.865 60.860 134.590 ;
        RECT 61.405 134.575 61.585 135.225 ;
        RECT 62.305 135.105 62.555 135.695 ;
        RECT 62.905 135.545 63.075 136.155 ;
        RECT 63.245 135.725 63.575 136.415 ;
        RECT 63.805 135.865 64.045 136.155 ;
        RECT 64.245 136.035 64.665 136.415 ;
        RECT 64.845 135.945 65.475 136.195 ;
        RECT 65.945 136.035 66.275 136.415 ;
        RECT 64.845 135.865 65.015 135.945 ;
        RECT 66.445 135.865 66.615 136.155 ;
        RECT 66.795 136.035 67.175 136.415 ;
        RECT 67.415 136.030 68.245 136.200 ;
        RECT 63.805 135.695 65.015 135.865 ;
        RECT 61.755 134.775 62.555 135.105 ;
        RECT 61.405 134.045 61.660 134.575 ;
        RECT 61.840 133.865 62.125 134.325 ;
        RECT 62.305 134.125 62.555 134.775 ;
        RECT 62.755 135.525 63.075 135.545 ;
        RECT 62.755 135.355 64.675 135.525 ;
        RECT 62.755 134.460 62.945 135.355 ;
        RECT 64.845 135.185 65.015 135.695 ;
        RECT 65.185 135.435 65.705 135.745 ;
        RECT 63.115 135.015 65.015 135.185 ;
        RECT 63.115 134.955 63.445 135.015 ;
        RECT 63.595 134.785 63.925 134.845 ;
        RECT 63.265 134.515 63.925 134.785 ;
        RECT 62.755 134.130 63.075 134.460 ;
        RECT 63.255 133.865 63.915 134.345 ;
        RECT 64.115 134.255 64.285 135.015 ;
        RECT 65.185 134.845 65.365 135.255 ;
        RECT 64.455 134.675 64.785 134.795 ;
        RECT 65.535 134.675 65.705 135.435 ;
        RECT 64.455 134.505 65.705 134.675 ;
        RECT 65.875 135.615 67.245 135.865 ;
        RECT 65.875 134.845 66.065 135.615 ;
        RECT 66.995 135.355 67.245 135.615 ;
        RECT 66.235 135.185 66.485 135.345 ;
        RECT 67.415 135.185 67.585 136.030 ;
        RECT 68.480 135.745 68.650 136.245 ;
        RECT 68.820 135.915 69.150 136.415 ;
        RECT 67.755 135.355 68.255 135.735 ;
        RECT 68.480 135.575 69.175 135.745 ;
        RECT 66.235 135.015 67.585 135.185 ;
        RECT 67.165 134.975 67.585 135.015 ;
        RECT 65.875 134.505 66.295 134.845 ;
        RECT 66.585 134.515 66.995 134.845 ;
        RECT 64.115 134.085 64.965 134.255 ;
        RECT 65.525 133.865 65.845 134.325 ;
        RECT 66.045 134.075 66.295 134.505 ;
        RECT 66.585 133.865 66.995 134.305 ;
        RECT 67.165 134.245 67.335 134.975 ;
        RECT 67.505 134.425 67.855 134.795 ;
        RECT 68.035 134.485 68.255 135.355 ;
        RECT 68.425 134.785 68.835 135.405 ;
        RECT 69.005 134.605 69.175 135.575 ;
        RECT 68.480 134.415 69.175 134.605 ;
        RECT 67.165 134.045 68.180 134.245 ;
        RECT 68.480 134.085 68.650 134.415 ;
        RECT 68.820 133.865 69.150 134.245 ;
        RECT 69.365 134.125 69.590 136.245 ;
        RECT 69.760 135.915 70.090 136.415 ;
        RECT 70.260 135.745 70.430 136.245 ;
        RECT 69.765 135.575 70.430 135.745 ;
        RECT 69.765 134.585 69.995 135.575 ;
        RECT 70.165 134.755 70.515 135.405 ;
        RECT 71.150 135.325 73.740 136.415 ;
        RECT 71.150 134.805 72.360 135.325 ;
        RECT 73.910 135.275 74.250 136.245 ;
        RECT 74.420 135.275 74.590 136.415 ;
        RECT 74.860 135.615 75.110 136.415 ;
        RECT 75.755 135.445 76.085 136.245 ;
        RECT 76.385 135.615 76.715 136.415 ;
        RECT 76.885 135.445 77.215 136.245 ;
        RECT 74.780 135.275 77.215 135.445 ;
        RECT 77.590 135.325 79.260 136.415 ;
        RECT 79.430 135.655 79.945 136.065 ;
        RECT 80.180 135.655 80.350 136.415 ;
        RECT 80.520 136.075 82.550 136.245 ;
        RECT 72.530 134.635 73.740 135.155 ;
        RECT 69.765 134.415 70.430 134.585 ;
        RECT 69.760 133.865 70.090 134.245 ;
        RECT 70.260 134.125 70.430 134.415 ;
        RECT 71.150 133.865 73.740 134.635 ;
        RECT 73.910 134.665 74.085 135.275 ;
        RECT 74.780 135.025 74.950 135.275 ;
        RECT 74.255 134.855 74.950 135.025 ;
        RECT 75.125 134.855 75.545 135.055 ;
        RECT 75.715 134.855 76.045 135.055 ;
        RECT 76.215 134.855 76.545 135.055 ;
        RECT 73.910 134.035 74.250 134.665 ;
        RECT 74.420 133.865 74.670 134.665 ;
        RECT 74.860 134.515 76.085 134.685 ;
        RECT 74.860 134.035 75.190 134.515 ;
        RECT 75.360 133.865 75.585 134.325 ;
        RECT 75.755 134.035 76.085 134.515 ;
        RECT 76.715 134.645 76.885 135.275 ;
        RECT 77.070 134.855 77.420 135.105 ;
        RECT 77.590 134.805 78.340 135.325 ;
        RECT 76.715 134.035 77.215 134.645 ;
        RECT 78.510 134.635 79.260 135.155 ;
        RECT 79.430 134.845 79.770 135.655 ;
        RECT 80.520 135.410 80.690 136.075 ;
        RECT 81.085 135.735 82.210 135.905 ;
        RECT 79.940 135.220 80.690 135.410 ;
        RECT 80.860 135.395 81.870 135.565 ;
        RECT 79.430 134.675 80.660 134.845 ;
        RECT 77.590 133.865 79.260 134.635 ;
        RECT 79.705 134.070 79.950 134.675 ;
        RECT 80.170 133.865 80.680 134.400 ;
        RECT 80.860 134.035 81.050 135.395 ;
        RECT 81.220 134.375 81.495 135.195 ;
        RECT 81.700 134.595 81.870 135.395 ;
        RECT 82.040 134.605 82.210 135.735 ;
        RECT 82.380 135.105 82.550 136.075 ;
        RECT 82.720 135.275 82.890 136.415 ;
        RECT 83.060 135.275 83.395 136.245 ;
        RECT 83.660 135.485 83.830 136.245 ;
        RECT 84.010 135.655 84.340 136.415 ;
        RECT 83.660 135.315 84.325 135.485 ;
        RECT 84.510 135.340 84.780 136.245 ;
        RECT 82.380 134.775 82.575 135.105 ;
        RECT 82.800 134.775 83.055 135.105 ;
        RECT 82.800 134.605 82.970 134.775 ;
        RECT 83.225 134.605 83.395 135.275 ;
        RECT 84.155 135.170 84.325 135.315 ;
        RECT 83.590 134.765 83.920 135.135 ;
        RECT 84.155 134.840 84.440 135.170 ;
        RECT 82.040 134.435 82.970 134.605 ;
        RECT 82.040 134.400 82.215 134.435 ;
        RECT 81.220 134.205 81.500 134.375 ;
        RECT 81.220 134.035 81.495 134.205 ;
        RECT 81.685 134.035 82.215 134.400 ;
        RECT 82.640 133.865 82.970 134.265 ;
        RECT 83.140 134.035 83.395 134.605 ;
        RECT 84.155 134.585 84.325 134.840 ;
        RECT 83.660 134.415 84.325 134.585 ;
        RECT 84.610 134.540 84.780 135.340 ;
        RECT 84.950 135.325 86.160 136.415 ;
        RECT 84.950 134.785 85.470 135.325 ;
        RECT 86.330 135.250 86.620 136.415 ;
        RECT 87.250 135.325 89.840 136.415 ;
        RECT 90.010 135.655 90.525 136.065 ;
        RECT 90.760 135.655 90.930 136.415 ;
        RECT 91.100 136.075 93.130 136.245 ;
        RECT 85.640 134.615 86.160 135.155 ;
        RECT 87.250 134.805 88.460 135.325 ;
        RECT 88.630 134.635 89.840 135.155 ;
        RECT 90.010 134.845 90.350 135.655 ;
        RECT 91.100 135.410 91.270 136.075 ;
        RECT 91.665 135.735 92.790 135.905 ;
        RECT 90.520 135.220 91.270 135.410 ;
        RECT 91.440 135.395 92.450 135.565 ;
        RECT 90.010 134.675 91.240 134.845 ;
        RECT 83.660 134.035 83.830 134.415 ;
        RECT 84.010 133.865 84.340 134.245 ;
        RECT 84.520 134.035 84.780 134.540 ;
        RECT 84.950 133.865 86.160 134.615 ;
        RECT 86.330 133.865 86.620 134.590 ;
        RECT 87.250 133.865 89.840 134.635 ;
        RECT 90.285 134.070 90.530 134.675 ;
        RECT 90.750 133.865 91.260 134.400 ;
        RECT 91.440 134.035 91.630 135.395 ;
        RECT 91.800 135.055 92.075 135.195 ;
        RECT 91.800 134.885 92.080 135.055 ;
        RECT 91.800 134.035 92.075 134.885 ;
        RECT 92.280 134.595 92.450 135.395 ;
        RECT 92.620 134.605 92.790 135.735 ;
        RECT 92.960 135.105 93.130 136.075 ;
        RECT 93.300 135.275 93.470 136.415 ;
        RECT 93.640 135.275 93.975 136.245 ;
        RECT 92.960 134.775 93.155 135.105 ;
        RECT 93.380 134.775 93.635 135.105 ;
        RECT 93.380 134.605 93.550 134.775 ;
        RECT 93.805 134.605 93.975 135.275 ;
        RECT 92.620 134.435 93.550 134.605 ;
        RECT 92.620 134.400 92.795 134.435 ;
        RECT 92.265 134.035 92.795 134.400 ;
        RECT 93.220 133.865 93.550 134.265 ;
        RECT 93.720 134.035 93.975 134.605 ;
        RECT 94.150 135.275 94.420 136.245 ;
        RECT 94.630 135.615 94.910 136.415 ;
        RECT 95.080 135.905 96.735 136.195 ;
        RECT 97.285 136.075 97.540 136.105 ;
        RECT 97.200 135.905 97.540 136.075 ;
        RECT 95.145 135.565 96.735 135.735 ;
        RECT 95.145 135.445 95.315 135.565 ;
        RECT 94.590 135.275 95.315 135.445 ;
        RECT 94.150 134.540 94.320 135.275 ;
        RECT 94.590 135.105 94.760 135.275 ;
        RECT 95.505 135.225 96.220 135.395 ;
        RECT 96.415 135.275 96.735 135.565 ;
        RECT 97.285 135.435 97.540 135.905 ;
        RECT 97.720 135.615 98.005 136.415 ;
        RECT 98.185 135.695 98.515 136.205 ;
        RECT 94.490 134.775 94.760 135.105 ;
        RECT 94.930 134.775 95.335 135.105 ;
        RECT 95.505 134.775 96.215 135.225 ;
        RECT 94.590 134.605 94.760 134.775 ;
        RECT 94.150 134.195 94.420 134.540 ;
        RECT 94.590 134.435 96.200 134.605 ;
        RECT 96.385 134.535 96.735 135.105 ;
        RECT 97.285 134.575 97.465 135.435 ;
        RECT 98.185 135.105 98.435 135.695 ;
        RECT 98.785 135.545 98.955 136.155 ;
        RECT 99.125 135.725 99.455 136.415 ;
        RECT 99.685 135.865 99.925 136.155 ;
        RECT 100.125 136.035 100.545 136.415 ;
        RECT 100.725 135.945 101.355 136.195 ;
        RECT 101.825 136.035 102.155 136.415 ;
        RECT 100.725 135.865 100.895 135.945 ;
        RECT 102.325 135.865 102.495 136.155 ;
        RECT 102.675 136.035 103.055 136.415 ;
        RECT 103.295 136.030 104.125 136.200 ;
        RECT 99.685 135.695 100.895 135.865 ;
        RECT 97.635 134.775 98.435 135.105 ;
        RECT 94.610 133.865 94.990 134.265 ;
        RECT 95.160 134.085 95.330 134.435 ;
        RECT 95.500 133.865 95.830 134.265 ;
        RECT 96.030 134.085 96.200 134.435 ;
        RECT 96.400 133.865 96.730 134.365 ;
        RECT 97.285 134.045 97.540 134.575 ;
        RECT 97.720 133.865 98.005 134.325 ;
        RECT 98.185 134.125 98.435 134.775 ;
        RECT 98.635 135.525 98.955 135.545 ;
        RECT 98.635 135.355 100.555 135.525 ;
        RECT 98.635 134.460 98.825 135.355 ;
        RECT 100.725 135.185 100.895 135.695 ;
        RECT 101.065 135.435 101.585 135.745 ;
        RECT 98.995 135.015 100.895 135.185 ;
        RECT 98.995 134.955 99.325 135.015 ;
        RECT 99.475 134.785 99.805 134.845 ;
        RECT 99.145 134.515 99.805 134.785 ;
        RECT 98.635 134.130 98.955 134.460 ;
        RECT 99.135 133.865 99.795 134.345 ;
        RECT 99.995 134.255 100.165 135.015 ;
        RECT 101.065 134.845 101.245 135.255 ;
        RECT 100.335 134.675 100.665 134.795 ;
        RECT 101.415 134.675 101.585 135.435 ;
        RECT 100.335 134.505 101.585 134.675 ;
        RECT 101.755 135.615 103.125 135.865 ;
        RECT 101.755 134.845 101.945 135.615 ;
        RECT 102.875 135.355 103.125 135.615 ;
        RECT 102.115 135.185 102.365 135.345 ;
        RECT 103.295 135.185 103.465 136.030 ;
        RECT 104.360 135.745 104.530 136.245 ;
        RECT 104.700 135.915 105.030 136.415 ;
        RECT 103.635 135.355 104.135 135.735 ;
        RECT 104.360 135.575 105.055 135.745 ;
        RECT 102.115 135.015 103.465 135.185 ;
        RECT 103.045 134.975 103.465 135.015 ;
        RECT 101.755 134.505 102.175 134.845 ;
        RECT 102.465 134.515 102.875 134.845 ;
        RECT 99.995 134.085 100.845 134.255 ;
        RECT 101.405 133.865 101.725 134.325 ;
        RECT 101.925 134.075 102.175 134.505 ;
        RECT 102.465 133.865 102.875 134.305 ;
        RECT 103.045 134.245 103.215 134.975 ;
        RECT 103.385 134.425 103.735 134.795 ;
        RECT 103.915 134.485 104.135 135.355 ;
        RECT 104.305 134.785 104.715 135.405 ;
        RECT 104.885 134.605 105.055 135.575 ;
        RECT 104.360 134.415 105.055 134.605 ;
        RECT 103.045 134.045 104.060 134.245 ;
        RECT 104.360 134.085 104.530 134.415 ;
        RECT 104.700 133.865 105.030 134.245 ;
        RECT 105.245 134.125 105.470 136.245 ;
        RECT 105.640 135.915 105.970 136.415 ;
        RECT 106.140 135.745 106.310 136.245 ;
        RECT 105.645 135.575 106.310 135.745 ;
        RECT 105.645 134.585 105.875 135.575 ;
        RECT 106.660 135.485 106.830 136.245 ;
        RECT 107.010 135.655 107.340 136.415 ;
        RECT 106.045 134.755 106.395 135.405 ;
        RECT 106.660 135.315 107.325 135.485 ;
        RECT 107.510 135.340 107.780 136.245 ;
        RECT 107.155 135.170 107.325 135.315 ;
        RECT 106.590 134.765 106.920 135.135 ;
        RECT 107.155 134.840 107.440 135.170 ;
        RECT 107.155 134.585 107.325 134.840 ;
        RECT 105.645 134.415 106.310 134.585 ;
        RECT 105.640 133.865 105.970 134.245 ;
        RECT 106.140 134.125 106.310 134.415 ;
        RECT 106.660 134.415 107.325 134.585 ;
        RECT 107.610 134.540 107.780 135.340 ;
        RECT 108.410 135.325 111.000 136.415 ;
        RECT 111.170 135.325 112.380 136.415 ;
        RECT 108.410 134.805 109.620 135.325 ;
        RECT 109.790 134.635 111.000 135.155 ;
        RECT 111.170 134.785 111.690 135.325 ;
        RECT 106.660 134.035 106.830 134.415 ;
        RECT 107.010 133.865 107.340 134.245 ;
        RECT 107.520 134.035 107.780 134.540 ;
        RECT 108.410 133.865 111.000 134.635 ;
        RECT 111.860 134.615 112.380 135.155 ;
        RECT 111.170 133.865 112.380 134.615 ;
        RECT 18.165 133.695 112.465 133.865 ;
        RECT 18.250 132.945 19.460 133.695 ;
        RECT 18.250 132.405 18.770 132.945 ;
        RECT 20.090 132.925 21.760 133.695 ;
        RECT 21.930 132.970 22.220 133.695 ;
        RECT 18.940 132.235 19.460 132.775 ;
        RECT 18.250 131.145 19.460 132.235 ;
        RECT 20.090 132.235 20.840 132.755 ;
        RECT 21.010 132.405 21.760 132.925 ;
        RECT 22.890 132.875 23.120 133.695 ;
        RECT 23.290 132.895 23.620 133.525 ;
        RECT 22.870 132.455 23.200 132.705 ;
        RECT 20.090 131.145 21.760 132.235 ;
        RECT 21.930 131.145 22.220 132.310 ;
        RECT 23.370 132.295 23.620 132.895 ;
        RECT 23.790 132.875 24.000 133.695 ;
        RECT 25.155 132.955 25.410 133.525 ;
        RECT 25.580 133.295 25.910 133.695 ;
        RECT 26.335 133.160 26.865 133.525 ;
        RECT 26.335 133.125 26.510 133.160 ;
        RECT 25.580 132.955 26.510 133.125 ;
        RECT 22.890 131.145 23.120 132.285 ;
        RECT 23.290 131.315 23.620 132.295 ;
        RECT 25.155 132.285 25.325 132.955 ;
        RECT 25.580 132.785 25.750 132.955 ;
        RECT 25.495 132.455 25.750 132.785 ;
        RECT 25.975 132.455 26.170 132.785 ;
        RECT 23.790 131.145 24.000 132.285 ;
        RECT 25.155 131.315 25.490 132.285 ;
        RECT 25.660 131.145 25.830 132.285 ;
        RECT 26.000 131.485 26.170 132.455 ;
        RECT 26.340 131.825 26.510 132.955 ;
        RECT 26.680 132.165 26.850 132.965 ;
        RECT 27.055 132.675 27.330 133.525 ;
        RECT 27.050 132.505 27.330 132.675 ;
        RECT 27.055 132.365 27.330 132.505 ;
        RECT 27.500 132.165 27.690 133.525 ;
        RECT 27.870 133.160 28.380 133.695 ;
        RECT 28.600 132.885 28.845 133.490 ;
        RECT 29.290 132.945 30.500 133.695 ;
        RECT 27.890 132.715 29.120 132.885 ;
        RECT 26.680 131.995 27.690 132.165 ;
        RECT 27.860 132.150 28.610 132.340 ;
        RECT 26.340 131.655 27.465 131.825 ;
        RECT 27.860 131.485 28.030 132.150 ;
        RECT 28.780 131.905 29.120 132.715 ;
        RECT 26.000 131.315 28.030 131.485 ;
        RECT 28.200 131.145 28.370 131.905 ;
        RECT 28.605 131.495 29.120 131.905 ;
        RECT 29.290 132.235 29.810 132.775 ;
        RECT 29.980 132.405 30.500 132.945 ;
        RECT 30.670 133.020 30.940 133.365 ;
        RECT 31.130 133.295 31.510 133.695 ;
        RECT 31.680 133.125 31.850 133.475 ;
        RECT 32.020 133.295 32.350 133.695 ;
        RECT 32.550 133.125 32.720 133.475 ;
        RECT 32.920 133.195 33.250 133.695 ;
        RECT 33.430 133.235 33.990 133.525 ;
        RECT 34.160 133.235 34.410 133.695 ;
        RECT 30.670 132.285 30.840 133.020 ;
        RECT 31.110 132.955 32.720 133.125 ;
        RECT 31.110 132.785 31.280 132.955 ;
        RECT 31.010 132.455 31.280 132.785 ;
        RECT 31.450 132.455 31.855 132.785 ;
        RECT 31.110 132.285 31.280 132.455 ;
        RECT 29.290 131.145 30.500 132.235 ;
        RECT 30.670 131.315 30.940 132.285 ;
        RECT 31.110 132.115 31.835 132.285 ;
        RECT 32.025 132.165 32.735 132.785 ;
        RECT 32.905 132.455 33.255 133.025 ;
        RECT 31.665 131.995 31.835 132.115 ;
        RECT 32.935 131.995 33.255 132.285 ;
        RECT 31.150 131.145 31.430 131.945 ;
        RECT 31.665 131.825 33.255 131.995 ;
        RECT 33.430 131.865 33.680 133.235 ;
        RECT 35.030 133.065 35.360 133.425 ;
        RECT 33.970 132.875 35.360 133.065 ;
        RECT 35.730 132.895 36.070 133.525 ;
        RECT 36.240 132.895 36.490 133.695 ;
        RECT 36.680 133.045 37.010 133.525 ;
        RECT 37.180 133.235 37.405 133.695 ;
        RECT 37.575 133.045 37.905 133.525 ;
        RECT 33.970 132.785 34.140 132.875 ;
        RECT 33.850 132.455 34.140 132.785 ;
        RECT 35.730 132.845 35.960 132.895 ;
        RECT 36.680 132.875 37.905 133.045 ;
        RECT 38.535 132.915 39.035 133.525 ;
        RECT 34.310 132.455 34.650 132.705 ;
        RECT 34.870 132.455 35.545 132.705 ;
        RECT 33.970 132.205 34.140 132.455 ;
        RECT 33.970 132.035 34.910 132.205 ;
        RECT 35.280 132.095 35.545 132.455 ;
        RECT 35.730 132.285 35.905 132.845 ;
        RECT 36.075 132.535 36.770 132.705 ;
        RECT 36.600 132.285 36.770 132.535 ;
        RECT 36.945 132.505 37.365 132.705 ;
        RECT 37.535 132.505 37.865 132.705 ;
        RECT 38.035 132.505 38.365 132.705 ;
        RECT 38.535 132.285 38.705 132.915 ;
        RECT 39.685 132.885 39.930 133.490 ;
        RECT 40.150 133.160 40.660 133.695 ;
        RECT 39.410 132.715 40.640 132.885 ;
        RECT 38.890 132.455 39.240 132.705 ;
        RECT 31.600 131.365 33.255 131.655 ;
        RECT 33.430 131.315 33.890 131.865 ;
        RECT 34.080 131.145 34.410 131.865 ;
        RECT 34.610 131.485 34.910 132.035 ;
        RECT 35.080 131.145 35.360 131.815 ;
        RECT 35.730 131.315 36.070 132.285 ;
        RECT 36.240 131.145 36.410 132.285 ;
        RECT 36.600 132.115 39.035 132.285 ;
        RECT 36.680 131.145 36.930 131.945 ;
        RECT 37.575 131.315 37.905 132.115 ;
        RECT 38.205 131.145 38.535 131.945 ;
        RECT 38.705 131.315 39.035 132.115 ;
        RECT 39.410 131.905 39.750 132.715 ;
        RECT 39.920 132.150 40.670 132.340 ;
        RECT 39.410 131.495 39.925 131.905 ;
        RECT 40.160 131.145 40.330 131.905 ;
        RECT 40.500 131.485 40.670 132.150 ;
        RECT 40.840 132.165 41.030 133.525 ;
        RECT 41.200 133.355 41.475 133.525 ;
        RECT 41.200 133.185 41.480 133.355 ;
        RECT 41.200 132.365 41.475 133.185 ;
        RECT 41.665 133.160 42.195 133.525 ;
        RECT 42.620 133.295 42.950 133.695 ;
        RECT 42.020 133.125 42.195 133.160 ;
        RECT 41.680 132.165 41.850 132.965 ;
        RECT 40.840 131.995 41.850 132.165 ;
        RECT 42.020 132.955 42.950 133.125 ;
        RECT 43.120 132.955 43.375 133.525 ;
        RECT 42.020 131.825 42.190 132.955 ;
        RECT 42.780 132.785 42.950 132.955 ;
        RECT 41.065 131.655 42.190 131.825 ;
        RECT 42.360 132.455 42.555 132.785 ;
        RECT 42.780 132.455 43.035 132.785 ;
        RECT 42.360 131.485 42.530 132.455 ;
        RECT 43.205 132.285 43.375 132.955 ;
        RECT 43.825 132.885 44.070 133.490 ;
        RECT 44.290 133.160 44.800 133.695 ;
        RECT 40.500 131.315 42.530 131.485 ;
        RECT 42.700 131.145 42.870 132.285 ;
        RECT 43.040 131.315 43.375 132.285 ;
        RECT 43.550 132.715 44.780 132.885 ;
        RECT 43.550 131.905 43.890 132.715 ;
        RECT 44.060 132.150 44.810 132.340 ;
        RECT 43.550 131.495 44.065 131.905 ;
        RECT 44.300 131.145 44.470 131.905 ;
        RECT 44.640 131.485 44.810 132.150 ;
        RECT 44.980 132.165 45.170 133.525 ;
        RECT 45.340 133.015 45.615 133.525 ;
        RECT 45.805 133.160 46.335 133.525 ;
        RECT 46.760 133.295 47.090 133.695 ;
        RECT 46.160 133.125 46.335 133.160 ;
        RECT 45.340 132.845 45.620 133.015 ;
        RECT 45.340 132.365 45.615 132.845 ;
        RECT 45.820 132.165 45.990 132.965 ;
        RECT 44.980 131.995 45.990 132.165 ;
        RECT 46.160 132.955 47.090 133.125 ;
        RECT 47.260 132.955 47.515 133.525 ;
        RECT 47.690 132.970 47.980 133.695 ;
        RECT 46.160 131.825 46.330 132.955 ;
        RECT 46.920 132.785 47.090 132.955 ;
        RECT 45.205 131.655 46.330 131.825 ;
        RECT 46.500 132.455 46.695 132.785 ;
        RECT 46.920 132.455 47.175 132.785 ;
        RECT 46.500 131.485 46.670 132.455 ;
        RECT 47.345 132.285 47.515 132.955 ;
        RECT 49.110 132.875 49.340 133.695 ;
        RECT 49.510 132.895 49.840 133.525 ;
        RECT 49.090 132.455 49.420 132.705 ;
        RECT 44.640 131.315 46.670 131.485 ;
        RECT 46.840 131.145 47.010 132.285 ;
        RECT 47.180 131.315 47.515 132.285 ;
        RECT 47.690 131.145 47.980 132.310 ;
        RECT 49.590 132.295 49.840 132.895 ;
        RECT 50.010 132.875 50.220 133.695 ;
        RECT 50.540 133.145 50.710 133.525 ;
        RECT 50.890 133.315 51.220 133.695 ;
        RECT 50.540 132.975 51.205 133.145 ;
        RECT 51.400 133.020 51.660 133.525 ;
        RECT 50.470 132.425 50.800 132.795 ;
        RECT 51.035 132.720 51.205 132.975 ;
        RECT 49.110 131.145 49.340 132.285 ;
        RECT 49.510 131.315 49.840 132.295 ;
        RECT 51.035 132.390 51.320 132.720 ;
        RECT 50.010 131.145 50.220 132.285 ;
        RECT 51.035 132.245 51.205 132.390 ;
        RECT 50.540 132.075 51.205 132.245 ;
        RECT 51.490 132.220 51.660 133.020 ;
        RECT 50.540 131.315 50.710 132.075 ;
        RECT 50.890 131.145 51.220 131.905 ;
        RECT 51.390 131.315 51.660 132.220 ;
        RECT 51.830 132.895 52.170 133.525 ;
        RECT 52.340 132.895 52.590 133.695 ;
        RECT 52.780 133.045 53.110 133.525 ;
        RECT 53.280 133.235 53.505 133.695 ;
        RECT 53.675 133.045 54.005 133.525 ;
        RECT 51.830 132.285 52.005 132.895 ;
        RECT 52.780 132.875 54.005 133.045 ;
        RECT 54.635 132.915 55.135 133.525 ;
        RECT 55.885 132.985 56.140 133.515 ;
        RECT 56.320 133.235 56.605 133.695 ;
        RECT 52.175 132.535 52.870 132.705 ;
        RECT 52.700 132.285 52.870 132.535 ;
        RECT 53.045 132.505 53.465 132.705 ;
        RECT 53.635 132.505 53.965 132.705 ;
        RECT 54.135 132.505 54.465 132.705 ;
        RECT 54.635 132.285 54.805 132.915 ;
        RECT 54.990 132.455 55.340 132.705 ;
        RECT 51.830 131.315 52.170 132.285 ;
        RECT 52.340 131.145 52.510 132.285 ;
        RECT 52.700 132.115 55.135 132.285 ;
        RECT 52.780 131.145 53.030 131.945 ;
        RECT 53.675 131.315 54.005 132.115 ;
        RECT 54.305 131.145 54.635 131.945 ;
        RECT 54.805 131.315 55.135 132.115 ;
        RECT 55.885 132.125 56.065 132.985 ;
        RECT 56.785 132.785 57.035 133.435 ;
        RECT 56.235 132.455 57.035 132.785 ;
        RECT 55.885 131.655 56.140 132.125 ;
        RECT 55.800 131.485 56.140 131.655 ;
        RECT 55.885 131.455 56.140 131.485 ;
        RECT 56.320 131.145 56.605 131.945 ;
        RECT 56.785 131.865 57.035 132.455 ;
        RECT 57.235 133.100 57.555 133.430 ;
        RECT 57.735 133.215 58.395 133.695 ;
        RECT 58.595 133.305 59.445 133.475 ;
        RECT 57.235 132.205 57.425 133.100 ;
        RECT 57.745 132.775 58.405 133.045 ;
        RECT 58.075 132.715 58.405 132.775 ;
        RECT 57.595 132.545 57.925 132.605 ;
        RECT 58.595 132.545 58.765 133.305 ;
        RECT 60.005 133.235 60.325 133.695 ;
        RECT 60.525 133.055 60.775 133.485 ;
        RECT 61.065 133.255 61.475 133.695 ;
        RECT 61.645 133.315 62.660 133.515 ;
        RECT 58.935 132.885 60.185 133.055 ;
        RECT 58.935 132.765 59.265 132.885 ;
        RECT 57.595 132.375 59.495 132.545 ;
        RECT 57.235 132.035 59.155 132.205 ;
        RECT 57.235 132.015 57.555 132.035 ;
        RECT 56.785 131.355 57.115 131.865 ;
        RECT 57.385 131.405 57.555 132.015 ;
        RECT 59.325 131.865 59.495 132.375 ;
        RECT 59.665 132.305 59.845 132.715 ;
        RECT 60.015 132.125 60.185 132.885 ;
        RECT 57.725 131.145 58.055 131.835 ;
        RECT 58.285 131.695 59.495 131.865 ;
        RECT 59.665 131.815 60.185 132.125 ;
        RECT 60.355 132.715 60.775 133.055 ;
        RECT 61.065 132.715 61.475 133.045 ;
        RECT 60.355 131.945 60.545 132.715 ;
        RECT 61.645 132.585 61.815 133.315 ;
        RECT 62.960 133.145 63.130 133.475 ;
        RECT 63.300 133.315 63.630 133.695 ;
        RECT 61.985 132.765 62.335 133.135 ;
        RECT 61.645 132.545 62.065 132.585 ;
        RECT 60.715 132.375 62.065 132.545 ;
        RECT 60.715 132.215 60.965 132.375 ;
        RECT 61.475 131.945 61.725 132.205 ;
        RECT 60.355 131.695 61.725 131.945 ;
        RECT 58.285 131.405 58.525 131.695 ;
        RECT 59.325 131.615 59.495 131.695 ;
        RECT 58.725 131.145 59.145 131.525 ;
        RECT 59.325 131.365 59.955 131.615 ;
        RECT 60.425 131.145 60.755 131.525 ;
        RECT 60.925 131.405 61.095 131.695 ;
        RECT 61.895 131.530 62.065 132.375 ;
        RECT 62.515 132.205 62.735 133.075 ;
        RECT 62.960 132.955 63.655 133.145 ;
        RECT 62.235 131.825 62.735 132.205 ;
        RECT 62.905 132.155 63.315 132.775 ;
        RECT 63.485 131.985 63.655 132.955 ;
        RECT 62.960 131.815 63.655 131.985 ;
        RECT 61.275 131.145 61.655 131.525 ;
        RECT 61.895 131.360 62.725 131.530 ;
        RECT 62.960 131.315 63.130 131.815 ;
        RECT 63.300 131.145 63.630 131.645 ;
        RECT 63.845 131.315 64.070 133.435 ;
        RECT 64.240 133.315 64.570 133.695 ;
        RECT 64.740 133.145 64.910 133.435 ;
        RECT 64.245 132.975 64.910 133.145 ;
        RECT 64.245 131.985 64.475 132.975 ;
        RECT 65.230 132.875 65.440 133.695 ;
        RECT 65.610 132.895 65.940 133.525 ;
        RECT 64.645 132.155 64.995 132.805 ;
        RECT 65.610 132.295 65.860 132.895 ;
        RECT 66.110 132.875 66.340 133.695 ;
        RECT 66.640 133.145 66.810 133.525 ;
        RECT 66.990 133.315 67.320 133.695 ;
        RECT 66.640 132.975 67.305 133.145 ;
        RECT 67.500 133.020 67.760 133.525 ;
        RECT 66.030 132.455 66.360 132.705 ;
        RECT 66.570 132.425 66.900 132.795 ;
        RECT 67.135 132.720 67.305 132.975 ;
        RECT 67.135 132.390 67.420 132.720 ;
        RECT 64.245 131.815 64.910 131.985 ;
        RECT 64.240 131.145 64.570 131.645 ;
        RECT 64.740 131.315 64.910 131.815 ;
        RECT 65.230 131.145 65.440 132.285 ;
        RECT 65.610 131.315 65.940 132.295 ;
        RECT 66.110 131.145 66.340 132.285 ;
        RECT 67.135 132.245 67.305 132.390 ;
        RECT 66.640 132.075 67.305 132.245 ;
        RECT 67.590 132.220 67.760 133.020 ;
        RECT 67.930 132.925 70.520 133.695 ;
        RECT 66.640 131.315 66.810 132.075 ;
        RECT 66.990 131.145 67.320 131.905 ;
        RECT 67.490 131.315 67.760 132.220 ;
        RECT 67.930 132.235 69.140 132.755 ;
        RECT 69.310 132.405 70.520 132.925 ;
        RECT 70.690 133.020 70.960 133.365 ;
        RECT 71.150 133.295 71.530 133.695 ;
        RECT 71.700 133.125 71.870 133.475 ;
        RECT 72.040 133.295 72.370 133.695 ;
        RECT 72.570 133.125 72.740 133.475 ;
        RECT 72.940 133.195 73.270 133.695 ;
        RECT 70.690 132.285 70.860 133.020 ;
        RECT 71.130 132.955 72.740 133.125 ;
        RECT 71.130 132.785 71.300 132.955 ;
        RECT 71.030 132.455 71.300 132.785 ;
        RECT 71.470 132.455 71.875 132.785 ;
        RECT 71.130 132.285 71.300 132.455 ;
        RECT 72.045 132.335 72.755 132.785 ;
        RECT 72.925 132.455 73.275 133.025 ;
        RECT 73.450 132.970 73.740 133.695 ;
        RECT 73.910 132.895 74.250 133.525 ;
        RECT 74.420 132.895 74.670 133.695 ;
        RECT 74.860 133.045 75.190 133.525 ;
        RECT 75.360 133.235 75.585 133.695 ;
        RECT 75.755 133.045 76.085 133.525 ;
        RECT 67.930 131.145 70.520 132.235 ;
        RECT 70.690 131.315 70.960 132.285 ;
        RECT 71.130 132.115 71.855 132.285 ;
        RECT 72.045 132.165 72.760 132.335 ;
        RECT 71.685 131.995 71.855 132.115 ;
        RECT 72.955 131.995 73.275 132.285 ;
        RECT 71.170 131.145 71.450 131.945 ;
        RECT 71.685 131.825 73.275 131.995 ;
        RECT 71.620 131.365 73.275 131.655 ;
        RECT 73.450 131.145 73.740 132.310 ;
        RECT 73.910 132.285 74.085 132.895 ;
        RECT 74.860 132.875 76.085 133.045 ;
        RECT 76.715 132.915 77.215 133.525 ;
        RECT 77.965 133.355 78.220 133.515 ;
        RECT 77.880 133.185 78.220 133.355 ;
        RECT 78.400 133.235 78.685 133.695 ;
        RECT 77.965 132.985 78.220 133.185 ;
        RECT 74.255 132.535 74.950 132.705 ;
        RECT 74.780 132.285 74.950 132.535 ;
        RECT 75.125 132.505 75.545 132.705 ;
        RECT 75.715 132.505 76.045 132.705 ;
        RECT 76.215 132.505 76.545 132.705 ;
        RECT 76.715 132.285 76.885 132.915 ;
        RECT 77.070 132.455 77.420 132.705 ;
        RECT 73.910 131.315 74.250 132.285 ;
        RECT 74.420 131.145 74.590 132.285 ;
        RECT 74.780 132.115 77.215 132.285 ;
        RECT 74.860 131.145 75.110 131.945 ;
        RECT 75.755 131.315 76.085 132.115 ;
        RECT 76.385 131.145 76.715 131.945 ;
        RECT 76.885 131.315 77.215 132.115 ;
        RECT 77.965 132.125 78.145 132.985 ;
        RECT 78.865 132.785 79.115 133.435 ;
        RECT 78.315 132.455 79.115 132.785 ;
        RECT 77.965 131.455 78.220 132.125 ;
        RECT 78.400 131.145 78.685 131.945 ;
        RECT 78.865 131.865 79.115 132.455 ;
        RECT 79.315 133.100 79.635 133.430 ;
        RECT 79.815 133.215 80.475 133.695 ;
        RECT 80.675 133.305 81.525 133.475 ;
        RECT 79.315 132.205 79.505 133.100 ;
        RECT 79.825 132.775 80.485 133.045 ;
        RECT 80.155 132.715 80.485 132.775 ;
        RECT 79.675 132.545 80.005 132.605 ;
        RECT 80.675 132.545 80.845 133.305 ;
        RECT 82.085 133.235 82.405 133.695 ;
        RECT 82.605 133.055 82.855 133.485 ;
        RECT 83.145 133.255 83.555 133.695 ;
        RECT 83.725 133.315 84.740 133.515 ;
        RECT 81.015 132.885 82.265 133.055 ;
        RECT 81.015 132.765 81.345 132.885 ;
        RECT 79.675 132.375 81.575 132.545 ;
        RECT 79.315 132.035 81.235 132.205 ;
        RECT 79.315 132.015 79.635 132.035 ;
        RECT 78.865 131.355 79.195 131.865 ;
        RECT 79.465 131.405 79.635 132.015 ;
        RECT 81.405 131.865 81.575 132.375 ;
        RECT 81.745 132.305 81.925 132.715 ;
        RECT 82.095 132.125 82.265 132.885 ;
        RECT 79.805 131.145 80.135 131.835 ;
        RECT 80.365 131.695 81.575 131.865 ;
        RECT 81.745 131.815 82.265 132.125 ;
        RECT 82.435 132.715 82.855 133.055 ;
        RECT 83.145 132.715 83.555 133.045 ;
        RECT 82.435 131.945 82.625 132.715 ;
        RECT 83.725 132.585 83.895 133.315 ;
        RECT 85.040 133.145 85.210 133.475 ;
        RECT 85.380 133.315 85.710 133.695 ;
        RECT 84.065 132.765 84.415 133.135 ;
        RECT 83.725 132.545 84.145 132.585 ;
        RECT 82.795 132.375 84.145 132.545 ;
        RECT 82.795 132.215 83.045 132.375 ;
        RECT 83.555 131.945 83.805 132.205 ;
        RECT 82.435 131.695 83.805 131.945 ;
        RECT 80.365 131.405 80.605 131.695 ;
        RECT 81.405 131.615 81.575 131.695 ;
        RECT 80.805 131.145 81.225 131.525 ;
        RECT 81.405 131.365 82.035 131.615 ;
        RECT 82.505 131.145 82.835 131.525 ;
        RECT 83.005 131.405 83.175 131.695 ;
        RECT 83.975 131.530 84.145 132.375 ;
        RECT 84.595 132.205 84.815 133.075 ;
        RECT 85.040 132.955 85.735 133.145 ;
        RECT 84.315 131.825 84.815 132.205 ;
        RECT 84.985 132.155 85.395 132.775 ;
        RECT 85.565 131.985 85.735 132.955 ;
        RECT 85.040 131.815 85.735 131.985 ;
        RECT 83.355 131.145 83.735 131.525 ;
        RECT 83.975 131.360 84.805 131.530 ;
        RECT 85.040 131.315 85.210 131.815 ;
        RECT 85.380 131.145 85.710 131.645 ;
        RECT 85.925 131.315 86.150 133.435 ;
        RECT 86.320 133.315 86.650 133.695 ;
        RECT 86.820 133.145 86.990 133.435 ;
        RECT 87.625 133.355 87.880 133.515 ;
        RECT 87.540 133.185 87.880 133.355 ;
        RECT 88.060 133.235 88.345 133.695 ;
        RECT 86.325 132.975 86.990 133.145 ;
        RECT 87.625 132.985 87.880 133.185 ;
        RECT 86.325 131.985 86.555 132.975 ;
        RECT 86.725 132.155 87.075 132.805 ;
        RECT 87.625 132.125 87.805 132.985 ;
        RECT 88.525 132.785 88.775 133.435 ;
        RECT 87.975 132.455 88.775 132.785 ;
        RECT 86.325 131.815 86.990 131.985 ;
        RECT 86.320 131.145 86.650 131.645 ;
        RECT 86.820 131.315 86.990 131.815 ;
        RECT 87.625 131.455 87.880 132.125 ;
        RECT 88.060 131.145 88.345 131.945 ;
        RECT 88.525 131.865 88.775 132.455 ;
        RECT 88.975 133.100 89.295 133.430 ;
        RECT 89.475 133.215 90.135 133.695 ;
        RECT 90.335 133.305 91.185 133.475 ;
        RECT 88.975 132.205 89.165 133.100 ;
        RECT 89.485 132.775 90.145 133.045 ;
        RECT 89.815 132.715 90.145 132.775 ;
        RECT 89.335 132.545 89.665 132.605 ;
        RECT 90.335 132.545 90.505 133.305 ;
        RECT 91.745 133.235 92.065 133.695 ;
        RECT 92.265 133.055 92.515 133.485 ;
        RECT 92.805 133.255 93.215 133.695 ;
        RECT 93.385 133.315 94.400 133.515 ;
        RECT 90.675 132.885 91.925 133.055 ;
        RECT 90.675 132.765 91.005 132.885 ;
        RECT 89.335 132.375 91.235 132.545 ;
        RECT 88.975 132.035 90.895 132.205 ;
        RECT 88.975 132.015 89.295 132.035 ;
        RECT 88.525 131.355 88.855 131.865 ;
        RECT 89.125 131.405 89.295 132.015 ;
        RECT 91.065 131.865 91.235 132.375 ;
        RECT 91.405 132.305 91.585 132.715 ;
        RECT 91.755 132.125 91.925 132.885 ;
        RECT 89.465 131.145 89.795 131.835 ;
        RECT 90.025 131.695 91.235 131.865 ;
        RECT 91.405 131.815 91.925 132.125 ;
        RECT 92.095 132.715 92.515 133.055 ;
        RECT 92.805 132.715 93.215 133.045 ;
        RECT 92.095 131.945 92.285 132.715 ;
        RECT 93.385 132.585 93.555 133.315 ;
        RECT 94.700 133.145 94.870 133.475 ;
        RECT 95.040 133.315 95.370 133.695 ;
        RECT 93.725 132.765 94.075 133.135 ;
        RECT 93.385 132.545 93.805 132.585 ;
        RECT 92.455 132.375 93.805 132.545 ;
        RECT 92.455 132.215 92.705 132.375 ;
        RECT 93.215 131.945 93.465 132.205 ;
        RECT 92.095 131.695 93.465 131.945 ;
        RECT 90.025 131.405 90.265 131.695 ;
        RECT 91.065 131.615 91.235 131.695 ;
        RECT 90.465 131.145 90.885 131.525 ;
        RECT 91.065 131.365 91.695 131.615 ;
        RECT 92.165 131.145 92.495 131.525 ;
        RECT 92.665 131.405 92.835 131.695 ;
        RECT 93.635 131.530 93.805 132.375 ;
        RECT 94.255 132.205 94.475 133.075 ;
        RECT 94.700 132.955 95.395 133.145 ;
        RECT 93.975 131.825 94.475 132.205 ;
        RECT 94.645 132.155 95.055 132.775 ;
        RECT 95.225 131.985 95.395 132.955 ;
        RECT 94.700 131.815 95.395 131.985 ;
        RECT 93.015 131.145 93.395 131.525 ;
        RECT 93.635 131.360 94.465 131.530 ;
        RECT 94.700 131.315 94.870 131.815 ;
        RECT 95.040 131.145 95.370 131.645 ;
        RECT 95.585 131.315 95.810 133.435 ;
        RECT 95.980 133.315 96.310 133.695 ;
        RECT 96.480 133.145 96.650 133.435 ;
        RECT 95.985 132.975 96.650 133.145 ;
        RECT 95.985 131.985 96.215 132.975 ;
        RECT 97.870 132.875 98.100 133.695 ;
        RECT 98.270 132.895 98.600 133.525 ;
        RECT 96.385 132.155 96.735 132.805 ;
        RECT 97.850 132.455 98.180 132.705 ;
        RECT 98.350 132.295 98.600 132.895 ;
        RECT 98.770 132.875 98.980 133.695 ;
        RECT 99.210 132.970 99.500 133.695 ;
        RECT 99.945 132.885 100.190 133.490 ;
        RECT 100.410 133.160 100.920 133.695 ;
        RECT 99.670 132.715 100.900 132.885 ;
        RECT 95.985 131.815 96.650 131.985 ;
        RECT 95.980 131.145 96.310 131.645 ;
        RECT 96.480 131.315 96.650 131.815 ;
        RECT 97.870 131.145 98.100 132.285 ;
        RECT 98.270 131.315 98.600 132.295 ;
        RECT 98.770 131.145 98.980 132.285 ;
        RECT 99.210 131.145 99.500 132.310 ;
        RECT 99.670 131.905 100.010 132.715 ;
        RECT 100.180 132.150 100.930 132.340 ;
        RECT 99.670 131.495 100.185 131.905 ;
        RECT 100.420 131.145 100.590 131.905 ;
        RECT 100.760 131.485 100.930 132.150 ;
        RECT 101.100 132.165 101.290 133.525 ;
        RECT 101.460 133.355 101.735 133.525 ;
        RECT 101.460 133.185 101.740 133.355 ;
        RECT 101.460 132.365 101.735 133.185 ;
        RECT 101.925 133.160 102.455 133.525 ;
        RECT 102.880 133.295 103.210 133.695 ;
        RECT 102.280 133.125 102.455 133.160 ;
        RECT 101.940 132.165 102.110 132.965 ;
        RECT 101.100 131.995 102.110 132.165 ;
        RECT 102.280 132.955 103.210 133.125 ;
        RECT 103.380 132.955 103.635 133.525 ;
        RECT 103.900 133.145 104.070 133.525 ;
        RECT 104.250 133.315 104.580 133.695 ;
        RECT 103.900 132.975 104.565 133.145 ;
        RECT 104.760 133.020 105.020 133.525 ;
        RECT 105.655 133.150 111.000 133.695 ;
        RECT 102.280 131.825 102.450 132.955 ;
        RECT 103.040 132.785 103.210 132.955 ;
        RECT 101.325 131.655 102.450 131.825 ;
        RECT 102.620 132.455 102.815 132.785 ;
        RECT 103.040 132.455 103.295 132.785 ;
        RECT 102.620 131.485 102.790 132.455 ;
        RECT 103.465 132.285 103.635 132.955 ;
        RECT 103.830 132.425 104.160 132.795 ;
        RECT 104.395 132.720 104.565 132.975 ;
        RECT 100.760 131.315 102.790 131.485 ;
        RECT 102.960 131.145 103.130 132.285 ;
        RECT 103.300 131.315 103.635 132.285 ;
        RECT 104.395 132.390 104.680 132.720 ;
        RECT 104.395 132.245 104.565 132.390 ;
        RECT 103.900 132.075 104.565 132.245 ;
        RECT 104.850 132.220 105.020 133.020 ;
        RECT 103.900 131.315 104.070 132.075 ;
        RECT 104.250 131.145 104.580 131.905 ;
        RECT 104.750 131.315 105.020 132.220 ;
        RECT 107.245 131.580 107.595 132.830 ;
        RECT 109.075 132.320 109.415 133.150 ;
        RECT 111.170 132.945 112.380 133.695 ;
        RECT 111.170 132.235 111.690 132.775 ;
        RECT 111.860 132.405 112.380 132.945 ;
        RECT 105.655 131.145 111.000 131.580 ;
        RECT 111.170 131.145 112.380 132.235 ;
        RECT 18.165 130.975 112.465 131.145 ;
        RECT 18.250 129.885 19.460 130.975 ;
        RECT 18.250 129.175 18.770 129.715 ;
        RECT 18.940 129.345 19.460 129.885 ;
        RECT 20.005 129.995 20.260 130.665 ;
        RECT 20.440 130.175 20.725 130.975 ;
        RECT 20.905 130.255 21.235 130.765 ;
        RECT 18.250 128.425 19.460 129.175 ;
        RECT 20.005 129.135 20.185 129.995 ;
        RECT 20.905 129.665 21.155 130.255 ;
        RECT 21.505 130.105 21.675 130.715 ;
        RECT 21.845 130.285 22.175 130.975 ;
        RECT 22.405 130.425 22.645 130.715 ;
        RECT 22.845 130.595 23.265 130.975 ;
        RECT 23.445 130.505 24.075 130.755 ;
        RECT 24.545 130.595 24.875 130.975 ;
        RECT 23.445 130.425 23.615 130.505 ;
        RECT 25.045 130.425 25.215 130.715 ;
        RECT 25.395 130.595 25.775 130.975 ;
        RECT 26.015 130.590 26.845 130.760 ;
        RECT 22.405 130.255 23.615 130.425 ;
        RECT 20.355 129.335 21.155 129.665 ;
        RECT 20.005 128.935 20.260 129.135 ;
        RECT 19.920 128.765 20.260 128.935 ;
        RECT 20.005 128.605 20.260 128.765 ;
        RECT 20.440 128.425 20.725 128.885 ;
        RECT 20.905 128.685 21.155 129.335 ;
        RECT 21.355 130.085 21.675 130.105 ;
        RECT 21.355 129.915 23.275 130.085 ;
        RECT 21.355 129.020 21.545 129.915 ;
        RECT 23.445 129.745 23.615 130.255 ;
        RECT 23.785 129.995 24.305 130.305 ;
        RECT 21.715 129.575 23.615 129.745 ;
        RECT 21.715 129.515 22.045 129.575 ;
        RECT 22.195 129.345 22.525 129.405 ;
        RECT 21.865 129.075 22.525 129.345 ;
        RECT 21.355 128.690 21.675 129.020 ;
        RECT 21.855 128.425 22.515 128.905 ;
        RECT 22.715 128.815 22.885 129.575 ;
        RECT 23.785 129.405 23.965 129.815 ;
        RECT 23.055 129.235 23.385 129.355 ;
        RECT 24.135 129.235 24.305 129.995 ;
        RECT 23.055 129.065 24.305 129.235 ;
        RECT 24.475 130.175 25.845 130.425 ;
        RECT 24.475 129.405 24.665 130.175 ;
        RECT 25.595 129.915 25.845 130.175 ;
        RECT 24.835 129.745 25.085 129.905 ;
        RECT 26.015 129.745 26.185 130.590 ;
        RECT 27.080 130.305 27.250 130.805 ;
        RECT 27.420 130.475 27.750 130.975 ;
        RECT 26.355 129.915 26.855 130.295 ;
        RECT 27.080 130.135 27.775 130.305 ;
        RECT 24.835 129.575 26.185 129.745 ;
        RECT 25.765 129.535 26.185 129.575 ;
        RECT 24.475 129.065 24.895 129.405 ;
        RECT 25.185 129.075 25.595 129.405 ;
        RECT 22.715 128.645 23.565 128.815 ;
        RECT 24.125 128.425 24.445 128.885 ;
        RECT 24.645 128.635 24.895 129.065 ;
        RECT 25.185 128.425 25.595 128.865 ;
        RECT 25.765 128.805 25.935 129.535 ;
        RECT 26.105 128.985 26.455 129.355 ;
        RECT 26.635 129.045 26.855 129.915 ;
        RECT 27.025 129.345 27.435 129.965 ;
        RECT 27.605 129.165 27.775 130.135 ;
        RECT 27.080 128.975 27.775 129.165 ;
        RECT 25.765 128.605 26.780 128.805 ;
        RECT 27.080 128.645 27.250 128.975 ;
        RECT 27.420 128.425 27.750 128.805 ;
        RECT 27.965 128.685 28.190 130.805 ;
        RECT 28.360 130.475 28.690 130.975 ;
        RECT 28.860 130.305 29.030 130.805 ;
        RECT 28.365 130.135 29.030 130.305 ;
        RECT 28.365 129.145 28.595 130.135 ;
        RECT 28.765 129.315 29.115 129.965 ;
        RECT 29.790 129.835 30.020 130.975 ;
        RECT 30.190 129.825 30.520 130.805 ;
        RECT 30.690 129.835 30.900 130.975 ;
        RECT 31.330 130.305 31.610 130.975 ;
        RECT 31.780 130.085 32.080 130.635 ;
        RECT 32.280 130.255 32.610 130.975 ;
        RECT 32.800 130.255 33.260 130.805 ;
        RECT 29.770 129.415 30.100 129.665 ;
        RECT 28.365 128.975 29.030 129.145 ;
        RECT 28.360 128.425 28.690 128.805 ;
        RECT 28.860 128.685 29.030 128.975 ;
        RECT 29.790 128.425 30.020 129.245 ;
        RECT 30.270 129.225 30.520 129.825 ;
        RECT 31.145 129.665 31.410 130.025 ;
        RECT 31.780 129.915 32.720 130.085 ;
        RECT 32.550 129.665 32.720 129.915 ;
        RECT 31.145 129.415 31.820 129.665 ;
        RECT 32.040 129.415 32.380 129.665 ;
        RECT 32.550 129.335 32.840 129.665 ;
        RECT 32.550 129.245 32.720 129.335 ;
        RECT 30.190 128.595 30.520 129.225 ;
        RECT 30.690 128.425 30.900 129.245 ;
        RECT 31.330 129.055 32.720 129.245 ;
        RECT 31.330 128.695 31.660 129.055 ;
        RECT 33.010 128.885 33.260 130.255 ;
        RECT 33.430 129.885 34.640 130.975 ;
        RECT 33.430 129.345 33.950 129.885 ;
        RECT 34.810 129.810 35.100 130.975 ;
        RECT 35.730 130.255 36.190 130.805 ;
        RECT 36.380 130.255 36.710 130.975 ;
        RECT 34.120 129.175 34.640 129.715 ;
        RECT 32.280 128.425 32.530 128.885 ;
        RECT 32.700 128.595 33.260 128.885 ;
        RECT 33.430 128.425 34.640 129.175 ;
        RECT 34.810 128.425 35.100 129.150 ;
        RECT 35.730 128.885 35.980 130.255 ;
        RECT 36.910 130.085 37.210 130.635 ;
        RECT 37.380 130.305 37.660 130.975 ;
        RECT 38.405 130.635 38.660 130.665 ;
        RECT 38.320 130.465 38.660 130.635 ;
        RECT 36.270 129.915 37.210 130.085 ;
        RECT 36.270 129.665 36.440 129.915 ;
        RECT 37.580 129.665 37.845 130.025 ;
        RECT 36.150 129.335 36.440 129.665 ;
        RECT 36.610 129.415 36.950 129.665 ;
        RECT 37.170 129.415 37.845 129.665 ;
        RECT 38.405 129.995 38.660 130.465 ;
        RECT 38.840 130.175 39.125 130.975 ;
        RECT 39.305 130.255 39.635 130.765 ;
        RECT 36.270 129.245 36.440 129.335 ;
        RECT 36.270 129.055 37.660 129.245 ;
        RECT 35.730 128.595 36.290 128.885 ;
        RECT 36.460 128.425 36.710 128.885 ;
        RECT 37.330 128.695 37.660 129.055 ;
        RECT 38.405 129.135 38.585 129.995 ;
        RECT 39.305 129.665 39.555 130.255 ;
        RECT 39.905 130.105 40.075 130.715 ;
        RECT 40.245 130.285 40.575 130.975 ;
        RECT 40.805 130.425 41.045 130.715 ;
        RECT 41.245 130.595 41.665 130.975 ;
        RECT 41.845 130.505 42.475 130.755 ;
        RECT 42.945 130.595 43.275 130.975 ;
        RECT 41.845 130.425 42.015 130.505 ;
        RECT 43.445 130.425 43.615 130.715 ;
        RECT 43.795 130.595 44.175 130.975 ;
        RECT 44.415 130.590 45.245 130.760 ;
        RECT 40.805 130.255 42.015 130.425 ;
        RECT 38.755 129.335 39.555 129.665 ;
        RECT 38.405 128.605 38.660 129.135 ;
        RECT 38.840 128.425 39.125 128.885 ;
        RECT 39.305 128.685 39.555 129.335 ;
        RECT 39.755 130.085 40.075 130.105 ;
        RECT 39.755 129.915 41.675 130.085 ;
        RECT 39.755 129.020 39.945 129.915 ;
        RECT 41.845 129.745 42.015 130.255 ;
        RECT 42.185 129.995 42.705 130.305 ;
        RECT 40.115 129.575 42.015 129.745 ;
        RECT 40.115 129.515 40.445 129.575 ;
        RECT 40.595 129.345 40.925 129.405 ;
        RECT 40.265 129.075 40.925 129.345 ;
        RECT 39.755 128.690 40.075 129.020 ;
        RECT 40.255 128.425 40.915 128.905 ;
        RECT 41.115 128.815 41.285 129.575 ;
        RECT 42.185 129.405 42.365 129.815 ;
        RECT 41.455 129.235 41.785 129.355 ;
        RECT 42.535 129.235 42.705 129.995 ;
        RECT 41.455 129.065 42.705 129.235 ;
        RECT 42.875 130.175 44.245 130.425 ;
        RECT 42.875 129.405 43.065 130.175 ;
        RECT 43.995 129.915 44.245 130.175 ;
        RECT 43.235 129.745 43.485 129.905 ;
        RECT 44.415 129.745 44.585 130.590 ;
        RECT 45.480 130.305 45.650 130.805 ;
        RECT 45.820 130.475 46.150 130.975 ;
        RECT 44.755 129.915 45.255 130.295 ;
        RECT 45.480 130.135 46.175 130.305 ;
        RECT 43.235 129.575 44.585 129.745 ;
        RECT 44.165 129.535 44.585 129.575 ;
        RECT 42.875 129.065 43.295 129.405 ;
        RECT 43.585 129.075 43.995 129.405 ;
        RECT 41.115 128.645 41.965 128.815 ;
        RECT 42.525 128.425 42.845 128.885 ;
        RECT 43.045 128.635 43.295 129.065 ;
        RECT 43.585 128.425 43.995 128.865 ;
        RECT 44.165 128.805 44.335 129.535 ;
        RECT 44.505 128.985 44.855 129.355 ;
        RECT 45.035 129.045 45.255 129.915 ;
        RECT 45.425 129.345 45.835 129.965 ;
        RECT 46.005 129.165 46.175 130.135 ;
        RECT 45.480 128.975 46.175 129.165 ;
        RECT 44.165 128.605 45.180 128.805 ;
        RECT 45.480 128.645 45.650 128.975 ;
        RECT 45.820 128.425 46.150 128.805 ;
        RECT 46.365 128.685 46.590 130.805 ;
        RECT 46.760 130.475 47.090 130.975 ;
        RECT 47.260 130.305 47.430 130.805 ;
        RECT 46.765 130.135 47.430 130.305 ;
        RECT 46.765 129.145 46.995 130.135 ;
        RECT 47.165 129.315 47.515 129.965 ;
        RECT 47.690 129.835 47.960 130.805 ;
        RECT 48.170 130.175 48.450 130.975 ;
        RECT 48.620 130.465 50.275 130.755 ;
        RECT 50.455 130.540 55.800 130.975 ;
        RECT 48.685 130.125 50.275 130.295 ;
        RECT 48.685 130.005 48.855 130.125 ;
        RECT 48.130 129.835 48.855 130.005 ;
        RECT 46.765 128.975 47.430 129.145 ;
        RECT 46.760 128.425 47.090 128.805 ;
        RECT 47.260 128.685 47.430 128.975 ;
        RECT 47.690 129.100 47.860 129.835 ;
        RECT 48.130 129.665 48.300 129.835 ;
        RECT 48.030 129.335 48.300 129.665 ;
        RECT 48.470 129.335 48.875 129.665 ;
        RECT 49.045 129.335 49.755 129.955 ;
        RECT 49.955 129.835 50.275 130.125 ;
        RECT 48.130 129.165 48.300 129.335 ;
        RECT 47.690 128.755 47.960 129.100 ;
        RECT 48.130 128.995 49.740 129.165 ;
        RECT 49.925 129.095 50.275 129.665 ;
        RECT 52.045 129.290 52.395 130.540 ;
        RECT 55.970 130.215 56.485 130.625 ;
        RECT 56.720 130.215 56.890 130.975 ;
        RECT 57.060 130.635 59.090 130.805 ;
        RECT 48.150 128.425 48.530 128.825 ;
        RECT 48.700 128.645 48.870 128.995 ;
        RECT 49.040 128.425 49.370 128.825 ;
        RECT 49.570 128.645 49.740 128.995 ;
        RECT 53.875 128.970 54.215 129.800 ;
        RECT 55.970 129.405 56.310 130.215 ;
        RECT 57.060 129.970 57.230 130.635 ;
        RECT 57.625 130.295 58.750 130.465 ;
        RECT 56.480 129.780 57.230 129.970 ;
        RECT 57.400 129.955 58.410 130.125 ;
        RECT 55.970 129.235 57.200 129.405 ;
        RECT 49.940 128.425 50.270 128.925 ;
        RECT 50.455 128.425 55.800 128.970 ;
        RECT 56.245 128.630 56.490 129.235 ;
        RECT 56.710 128.425 57.220 128.960 ;
        RECT 57.400 128.595 57.590 129.955 ;
        RECT 57.760 129.615 58.035 129.755 ;
        RECT 57.760 129.445 58.040 129.615 ;
        RECT 57.760 128.595 58.035 129.445 ;
        RECT 58.240 129.155 58.410 129.955 ;
        RECT 58.580 129.165 58.750 130.295 ;
        RECT 58.920 129.665 59.090 130.635 ;
        RECT 59.260 129.835 59.430 130.975 ;
        RECT 59.600 129.835 59.935 130.805 ;
        RECT 58.920 129.335 59.115 129.665 ;
        RECT 59.340 129.335 59.595 129.665 ;
        RECT 59.340 129.165 59.510 129.335 ;
        RECT 59.765 129.165 59.935 129.835 ;
        RECT 60.570 129.810 60.860 130.975 ;
        RECT 61.120 130.045 61.290 130.805 ;
        RECT 61.470 130.215 61.800 130.975 ;
        RECT 61.120 129.875 61.785 130.045 ;
        RECT 61.970 129.900 62.240 130.805 ;
        RECT 61.615 129.730 61.785 129.875 ;
        RECT 61.050 129.325 61.380 129.695 ;
        RECT 61.615 129.400 61.900 129.730 ;
        RECT 58.580 128.995 59.510 129.165 ;
        RECT 58.580 128.960 58.755 128.995 ;
        RECT 58.225 128.595 58.755 128.960 ;
        RECT 59.180 128.425 59.510 128.825 ;
        RECT 59.680 128.595 59.935 129.165 ;
        RECT 60.570 128.425 60.860 129.150 ;
        RECT 61.615 129.145 61.785 129.400 ;
        RECT 61.120 128.975 61.785 129.145 ;
        RECT 62.070 129.100 62.240 129.900 ;
        RECT 62.470 129.835 62.680 130.975 ;
        RECT 62.850 129.825 63.180 130.805 ;
        RECT 63.350 129.835 63.580 130.975 ;
        RECT 64.710 129.885 68.220 130.975 ;
        RECT 68.590 130.305 68.870 130.975 ;
        RECT 69.040 130.085 69.340 130.635 ;
        RECT 69.540 130.255 69.870 130.975 ;
        RECT 70.060 130.255 70.520 130.805 ;
        RECT 61.120 128.595 61.290 128.975 ;
        RECT 61.470 128.425 61.800 128.805 ;
        RECT 61.980 128.595 62.240 129.100 ;
        RECT 62.470 128.425 62.680 129.245 ;
        RECT 62.850 129.225 63.100 129.825 ;
        RECT 63.270 129.415 63.600 129.665 ;
        RECT 64.710 129.365 66.400 129.885 ;
        RECT 62.850 128.595 63.180 129.225 ;
        RECT 63.350 128.425 63.580 129.245 ;
        RECT 66.570 129.195 68.220 129.715 ;
        RECT 68.405 129.665 68.670 130.025 ;
        RECT 69.040 129.915 69.980 130.085 ;
        RECT 69.810 129.665 69.980 129.915 ;
        RECT 68.405 129.415 69.080 129.665 ;
        RECT 69.300 129.415 69.640 129.665 ;
        RECT 69.810 129.335 70.100 129.665 ;
        RECT 69.810 129.245 69.980 129.335 ;
        RECT 64.710 128.425 68.220 129.195 ;
        RECT 68.590 129.055 69.980 129.245 ;
        RECT 68.590 128.695 68.920 129.055 ;
        RECT 70.270 128.885 70.520 130.255 ;
        RECT 70.780 130.230 71.050 130.975 ;
        RECT 71.680 130.970 77.955 130.975 ;
        RECT 71.220 130.060 71.510 130.800 ;
        RECT 71.680 130.245 71.935 130.970 ;
        RECT 72.120 130.075 72.380 130.800 ;
        RECT 72.550 130.245 72.795 130.970 ;
        RECT 72.980 130.075 73.240 130.800 ;
        RECT 73.410 130.245 73.655 130.970 ;
        RECT 73.840 130.075 74.100 130.800 ;
        RECT 74.270 130.245 74.515 130.970 ;
        RECT 74.685 130.075 74.945 130.800 ;
        RECT 75.115 130.245 75.375 130.970 ;
        RECT 75.545 130.075 75.805 130.800 ;
        RECT 75.975 130.245 76.235 130.970 ;
        RECT 76.405 130.075 76.665 130.800 ;
        RECT 76.835 130.245 77.095 130.970 ;
        RECT 77.265 130.075 77.525 130.800 ;
        RECT 77.695 130.175 77.955 130.970 ;
        RECT 72.120 130.060 77.525 130.075 ;
        RECT 70.780 129.835 77.525 130.060 ;
        RECT 70.780 129.245 71.945 129.835 ;
        RECT 78.125 129.665 78.375 130.800 ;
        RECT 78.555 130.165 78.815 130.975 ;
        RECT 78.990 129.665 79.235 130.805 ;
        RECT 79.415 130.165 79.710 130.975 ;
        RECT 80.350 129.885 82.020 130.975 ;
        RECT 72.115 129.415 79.235 129.665 ;
        RECT 70.780 129.075 77.525 129.245 ;
        RECT 69.540 128.425 69.790 128.885 ;
        RECT 69.960 128.595 70.520 128.885 ;
        RECT 70.780 128.425 71.080 128.905 ;
        RECT 71.250 128.620 71.510 129.075 ;
        RECT 71.680 128.425 71.940 128.905 ;
        RECT 72.120 128.620 72.380 129.075 ;
        RECT 72.550 128.425 72.800 128.905 ;
        RECT 72.980 128.620 73.240 129.075 ;
        RECT 73.410 128.425 73.660 128.905 ;
        RECT 73.840 128.620 74.100 129.075 ;
        RECT 74.270 128.425 74.515 128.905 ;
        RECT 74.685 128.620 74.960 129.075 ;
        RECT 75.130 128.425 75.375 128.905 ;
        RECT 75.545 128.620 75.805 129.075 ;
        RECT 75.975 128.425 76.235 128.905 ;
        RECT 76.405 128.620 76.665 129.075 ;
        RECT 76.835 128.425 77.095 128.905 ;
        RECT 77.265 128.620 77.525 129.075 ;
        RECT 77.695 128.425 77.955 128.985 ;
        RECT 78.125 128.605 78.375 129.415 ;
        RECT 78.555 128.425 78.815 128.950 ;
        RECT 78.985 128.605 79.235 129.415 ;
        RECT 79.405 129.105 79.720 129.665 ;
        RECT 80.350 129.365 81.100 129.885 ;
        RECT 82.250 129.835 82.460 130.975 ;
        RECT 82.630 129.825 82.960 130.805 ;
        RECT 83.130 129.835 83.360 130.975 ;
        RECT 83.570 129.885 84.780 130.975 ;
        RECT 81.270 129.195 82.020 129.715 ;
        RECT 79.415 128.425 79.720 128.935 ;
        RECT 80.350 128.425 82.020 129.195 ;
        RECT 82.250 128.425 82.460 129.245 ;
        RECT 82.630 129.225 82.880 129.825 ;
        RECT 83.050 129.415 83.380 129.665 ;
        RECT 83.570 129.345 84.090 129.885 ;
        RECT 84.990 129.835 85.220 130.975 ;
        RECT 85.390 129.825 85.720 130.805 ;
        RECT 85.890 129.835 86.100 130.975 ;
        RECT 82.630 128.595 82.960 129.225 ;
        RECT 83.130 128.425 83.360 129.245 ;
        RECT 84.260 129.175 84.780 129.715 ;
        RECT 84.970 129.415 85.300 129.665 ;
        RECT 83.570 128.425 84.780 129.175 ;
        RECT 84.990 128.425 85.220 129.245 ;
        RECT 85.470 129.225 85.720 129.825 ;
        RECT 86.330 129.810 86.620 130.975 ;
        RECT 86.800 130.165 87.095 130.975 ;
        RECT 87.275 129.665 87.520 130.805 ;
        RECT 87.695 130.165 87.955 130.975 ;
        RECT 88.555 130.970 94.830 130.975 ;
        RECT 88.135 129.665 88.385 130.800 ;
        RECT 88.555 130.175 88.815 130.970 ;
        RECT 88.985 130.075 89.245 130.800 ;
        RECT 89.415 130.245 89.675 130.970 ;
        RECT 89.845 130.075 90.105 130.800 ;
        RECT 90.275 130.245 90.535 130.970 ;
        RECT 90.705 130.075 90.965 130.800 ;
        RECT 91.135 130.245 91.395 130.970 ;
        RECT 91.565 130.075 91.825 130.800 ;
        RECT 91.995 130.245 92.240 130.970 ;
        RECT 92.410 130.075 92.670 130.800 ;
        RECT 92.855 130.245 93.100 130.970 ;
        RECT 93.270 130.075 93.530 130.800 ;
        RECT 93.715 130.245 93.960 130.970 ;
        RECT 94.130 130.075 94.390 130.800 ;
        RECT 94.575 130.245 94.830 130.970 ;
        RECT 88.985 130.060 94.390 130.075 ;
        RECT 95.000 130.060 95.290 130.800 ;
        RECT 95.460 130.230 95.730 130.975 ;
        RECT 88.985 129.835 95.730 130.060 ;
        RECT 85.390 128.595 85.720 129.225 ;
        RECT 85.890 128.425 86.100 129.245 ;
        RECT 86.330 128.425 86.620 129.150 ;
        RECT 86.790 129.105 87.105 129.665 ;
        RECT 87.275 129.415 94.395 129.665 ;
        RECT 86.790 128.425 87.095 128.935 ;
        RECT 87.275 128.605 87.525 129.415 ;
        RECT 87.695 128.425 87.955 128.950 ;
        RECT 88.135 128.605 88.385 129.415 ;
        RECT 94.565 129.245 95.730 129.835 ;
        RECT 88.985 129.075 95.730 129.245 ;
        RECT 95.990 129.900 96.260 130.805 ;
        RECT 96.430 130.215 96.760 130.975 ;
        RECT 96.940 130.045 97.110 130.805 ;
        RECT 95.990 129.100 96.160 129.900 ;
        RECT 96.445 129.875 97.110 130.045 ;
        RECT 97.370 129.885 99.960 130.975 ;
        RECT 100.135 130.540 105.480 130.975 ;
        RECT 105.655 130.540 111.000 130.975 ;
        RECT 96.445 129.730 96.615 129.875 ;
        RECT 96.330 129.400 96.615 129.730 ;
        RECT 96.445 129.145 96.615 129.400 ;
        RECT 96.850 129.325 97.180 129.695 ;
        RECT 97.370 129.365 98.580 129.885 ;
        RECT 98.750 129.195 99.960 129.715 ;
        RECT 101.725 129.290 102.075 130.540 ;
        RECT 88.555 128.425 88.815 128.985 ;
        RECT 88.985 128.620 89.245 129.075 ;
        RECT 89.415 128.425 89.675 128.905 ;
        RECT 89.845 128.620 90.105 129.075 ;
        RECT 90.275 128.425 90.535 128.905 ;
        RECT 90.705 128.620 90.965 129.075 ;
        RECT 91.135 128.425 91.380 128.905 ;
        RECT 91.550 128.620 91.825 129.075 ;
        RECT 91.995 128.425 92.240 128.905 ;
        RECT 92.410 128.620 92.670 129.075 ;
        RECT 92.850 128.425 93.100 128.905 ;
        RECT 93.270 128.620 93.530 129.075 ;
        RECT 93.710 128.425 93.960 128.905 ;
        RECT 94.130 128.620 94.390 129.075 ;
        RECT 94.570 128.425 94.830 128.905 ;
        RECT 95.000 128.620 95.260 129.075 ;
        RECT 95.430 128.425 95.730 128.905 ;
        RECT 95.990 128.595 96.250 129.100 ;
        RECT 96.445 128.975 97.110 129.145 ;
        RECT 96.430 128.425 96.760 128.805 ;
        RECT 96.940 128.595 97.110 128.975 ;
        RECT 97.370 128.425 99.960 129.195 ;
        RECT 103.555 128.970 103.895 129.800 ;
        RECT 107.245 129.290 107.595 130.540 ;
        RECT 111.170 129.885 112.380 130.975 ;
        RECT 109.075 128.970 109.415 129.800 ;
        RECT 111.170 129.345 111.690 129.885 ;
        RECT 111.860 129.175 112.380 129.715 ;
        RECT 100.135 128.425 105.480 128.970 ;
        RECT 105.655 128.425 111.000 128.970 ;
        RECT 111.170 128.425 112.380 129.175 ;
        RECT 18.165 128.255 112.465 128.425 ;
        RECT 18.250 127.505 19.460 128.255 ;
        RECT 20.640 127.705 20.810 128.085 ;
        RECT 20.990 127.875 21.320 128.255 ;
        RECT 20.640 127.535 21.305 127.705 ;
        RECT 21.500 127.580 21.760 128.085 ;
        RECT 18.250 126.965 18.770 127.505 ;
        RECT 18.940 126.795 19.460 127.335 ;
        RECT 20.570 126.985 20.900 127.355 ;
        RECT 21.135 127.280 21.305 127.535 ;
        RECT 21.135 126.950 21.420 127.280 ;
        RECT 21.135 126.805 21.305 126.950 ;
        RECT 18.250 125.705 19.460 126.795 ;
        RECT 20.640 126.635 21.305 126.805 ;
        RECT 21.590 126.780 21.760 127.580 ;
        RECT 21.930 127.530 22.220 128.255 ;
        RECT 22.395 127.515 22.650 128.085 ;
        RECT 22.820 127.855 23.150 128.255 ;
        RECT 23.575 127.720 24.105 128.085 ;
        RECT 23.575 127.685 23.750 127.720 ;
        RECT 22.820 127.515 23.750 127.685 ;
        RECT 20.640 125.875 20.810 126.635 ;
        RECT 20.990 125.705 21.320 126.465 ;
        RECT 21.490 125.875 21.760 126.780 ;
        RECT 21.930 125.705 22.220 126.870 ;
        RECT 22.395 126.845 22.565 127.515 ;
        RECT 22.820 127.345 22.990 127.515 ;
        RECT 22.735 127.015 22.990 127.345 ;
        RECT 23.215 127.015 23.410 127.345 ;
        RECT 22.395 125.875 22.730 126.845 ;
        RECT 22.900 125.705 23.070 126.845 ;
        RECT 23.240 126.045 23.410 127.015 ;
        RECT 23.580 126.385 23.750 127.515 ;
        RECT 23.920 126.725 24.090 127.525 ;
        RECT 24.295 127.235 24.570 128.085 ;
        RECT 24.290 127.065 24.570 127.235 ;
        RECT 24.295 126.925 24.570 127.065 ;
        RECT 24.740 126.725 24.930 128.085 ;
        RECT 25.110 127.720 25.620 128.255 ;
        RECT 25.840 127.445 26.085 128.050 ;
        RECT 26.620 127.705 26.790 128.085 ;
        RECT 26.970 127.875 27.300 128.255 ;
        RECT 26.620 127.535 27.285 127.705 ;
        RECT 27.480 127.580 27.740 128.085 ;
        RECT 28.285 127.915 28.540 128.075 ;
        RECT 28.200 127.745 28.540 127.915 ;
        RECT 28.720 127.795 29.005 128.255 ;
        RECT 25.130 127.275 26.360 127.445 ;
        RECT 23.920 126.555 24.930 126.725 ;
        RECT 25.100 126.710 25.850 126.900 ;
        RECT 23.580 126.215 24.705 126.385 ;
        RECT 25.100 126.045 25.270 126.710 ;
        RECT 26.020 126.465 26.360 127.275 ;
        RECT 26.550 126.985 26.880 127.355 ;
        RECT 27.115 127.280 27.285 127.535 ;
        RECT 27.115 126.950 27.400 127.280 ;
        RECT 27.115 126.805 27.285 126.950 ;
        RECT 23.240 125.875 25.270 126.045 ;
        RECT 25.440 125.705 25.610 126.465 ;
        RECT 25.845 126.055 26.360 126.465 ;
        RECT 26.620 126.635 27.285 126.805 ;
        RECT 27.570 126.780 27.740 127.580 ;
        RECT 26.620 125.875 26.790 126.635 ;
        RECT 26.970 125.705 27.300 126.465 ;
        RECT 27.470 125.875 27.740 126.780 ;
        RECT 28.285 127.545 28.540 127.745 ;
        RECT 28.285 126.685 28.465 127.545 ;
        RECT 29.185 127.345 29.435 127.995 ;
        RECT 28.635 127.015 29.435 127.345 ;
        RECT 28.285 126.015 28.540 126.685 ;
        RECT 28.720 125.705 29.005 126.505 ;
        RECT 29.185 126.425 29.435 127.015 ;
        RECT 29.635 127.660 29.955 127.990 ;
        RECT 30.135 127.775 30.795 128.255 ;
        RECT 30.995 127.865 31.845 128.035 ;
        RECT 29.635 126.765 29.825 127.660 ;
        RECT 30.145 127.335 30.805 127.605 ;
        RECT 30.475 127.275 30.805 127.335 ;
        RECT 29.995 127.105 30.325 127.165 ;
        RECT 30.995 127.105 31.165 127.865 ;
        RECT 32.405 127.795 32.725 128.255 ;
        RECT 32.925 127.615 33.175 128.045 ;
        RECT 33.465 127.815 33.875 128.255 ;
        RECT 34.045 127.875 35.060 128.075 ;
        RECT 31.335 127.445 32.585 127.615 ;
        RECT 31.335 127.325 31.665 127.445 ;
        RECT 29.995 126.935 31.895 127.105 ;
        RECT 29.635 126.595 31.555 126.765 ;
        RECT 29.635 126.575 29.955 126.595 ;
        RECT 29.185 125.915 29.515 126.425 ;
        RECT 29.785 125.965 29.955 126.575 ;
        RECT 31.725 126.425 31.895 126.935 ;
        RECT 32.065 126.865 32.245 127.275 ;
        RECT 32.415 126.685 32.585 127.445 ;
        RECT 30.125 125.705 30.455 126.395 ;
        RECT 30.685 126.255 31.895 126.425 ;
        RECT 32.065 126.375 32.585 126.685 ;
        RECT 32.755 127.275 33.175 127.615 ;
        RECT 33.465 127.275 33.875 127.605 ;
        RECT 32.755 126.505 32.945 127.275 ;
        RECT 34.045 127.145 34.215 127.875 ;
        RECT 35.360 127.705 35.530 128.035 ;
        RECT 35.700 127.875 36.030 128.255 ;
        RECT 34.385 127.325 34.735 127.695 ;
        RECT 34.045 127.105 34.465 127.145 ;
        RECT 33.115 126.935 34.465 127.105 ;
        RECT 33.115 126.775 33.365 126.935 ;
        RECT 33.875 126.505 34.125 126.765 ;
        RECT 32.755 126.255 34.125 126.505 ;
        RECT 30.685 125.965 30.925 126.255 ;
        RECT 31.725 126.175 31.895 126.255 ;
        RECT 31.125 125.705 31.545 126.085 ;
        RECT 31.725 125.925 32.355 126.175 ;
        RECT 32.825 125.705 33.155 126.085 ;
        RECT 33.325 125.965 33.495 126.255 ;
        RECT 34.295 126.090 34.465 126.935 ;
        RECT 34.915 126.765 35.135 127.635 ;
        RECT 35.360 127.515 36.055 127.705 ;
        RECT 34.635 126.385 35.135 126.765 ;
        RECT 35.305 126.715 35.715 127.335 ;
        RECT 35.885 126.545 36.055 127.515 ;
        RECT 35.360 126.375 36.055 126.545 ;
        RECT 33.675 125.705 34.055 126.085 ;
        RECT 34.295 125.920 35.125 126.090 ;
        RECT 35.360 125.875 35.530 126.375 ;
        RECT 35.700 125.705 36.030 126.205 ;
        RECT 36.245 125.875 36.470 127.995 ;
        RECT 36.640 127.875 36.970 128.255 ;
        RECT 37.140 127.705 37.310 127.995 ;
        RECT 36.645 127.535 37.310 127.705 ;
        RECT 36.645 126.545 36.875 127.535 ;
        RECT 37.575 127.515 37.830 128.085 ;
        RECT 38.000 127.855 38.330 128.255 ;
        RECT 38.755 127.720 39.285 128.085 ;
        RECT 39.475 127.915 39.750 128.085 ;
        RECT 39.470 127.745 39.750 127.915 ;
        RECT 38.755 127.685 38.930 127.720 ;
        RECT 38.000 127.515 38.930 127.685 ;
        RECT 37.045 126.715 37.395 127.365 ;
        RECT 37.575 126.845 37.745 127.515 ;
        RECT 38.000 127.345 38.170 127.515 ;
        RECT 37.915 127.015 38.170 127.345 ;
        RECT 38.395 127.015 38.590 127.345 ;
        RECT 36.645 126.375 37.310 126.545 ;
        RECT 36.640 125.705 36.970 126.205 ;
        RECT 37.140 125.875 37.310 126.375 ;
        RECT 37.575 125.875 37.910 126.845 ;
        RECT 38.080 125.705 38.250 126.845 ;
        RECT 38.420 126.045 38.590 127.015 ;
        RECT 38.760 126.385 38.930 127.515 ;
        RECT 39.100 126.725 39.270 127.525 ;
        RECT 39.475 126.925 39.750 127.745 ;
        RECT 39.920 126.725 40.110 128.085 ;
        RECT 40.290 127.720 40.800 128.255 ;
        RECT 41.020 127.445 41.265 128.050 ;
        RECT 41.800 127.705 41.970 128.085 ;
        RECT 42.150 127.875 42.480 128.255 ;
        RECT 41.800 127.535 42.465 127.705 ;
        RECT 42.660 127.580 42.920 128.085 ;
        RECT 40.310 127.275 41.540 127.445 ;
        RECT 39.100 126.555 40.110 126.725 ;
        RECT 40.280 126.710 41.030 126.900 ;
        RECT 38.760 126.215 39.885 126.385 ;
        RECT 40.280 126.045 40.450 126.710 ;
        RECT 41.200 126.465 41.540 127.275 ;
        RECT 41.730 126.985 42.060 127.355 ;
        RECT 42.295 127.280 42.465 127.535 ;
        RECT 42.295 126.950 42.580 127.280 ;
        RECT 42.295 126.805 42.465 126.950 ;
        RECT 38.420 125.875 40.450 126.045 ;
        RECT 40.620 125.705 40.790 126.465 ;
        RECT 41.025 126.055 41.540 126.465 ;
        RECT 41.800 126.635 42.465 126.805 ;
        RECT 42.750 126.780 42.920 127.580 ;
        RECT 43.290 127.625 43.620 127.985 ;
        RECT 44.240 127.795 44.490 128.255 ;
        RECT 44.660 127.795 45.220 128.085 ;
        RECT 43.290 127.435 44.680 127.625 ;
        RECT 44.510 127.345 44.680 127.435 ;
        RECT 41.800 125.875 41.970 126.635 ;
        RECT 42.150 125.705 42.480 126.465 ;
        RECT 42.650 125.875 42.920 126.780 ;
        RECT 43.105 127.015 43.780 127.265 ;
        RECT 44.000 127.015 44.340 127.265 ;
        RECT 44.510 127.015 44.800 127.345 ;
        RECT 43.105 126.655 43.370 127.015 ;
        RECT 44.510 126.765 44.680 127.015 ;
        RECT 43.740 126.595 44.680 126.765 ;
        RECT 43.290 125.705 43.570 126.375 ;
        RECT 43.740 126.045 44.040 126.595 ;
        RECT 44.970 126.425 45.220 127.795 ;
        RECT 45.590 127.625 45.920 127.985 ;
        RECT 46.540 127.795 46.790 128.255 ;
        RECT 46.960 127.795 47.520 128.085 ;
        RECT 45.590 127.435 46.980 127.625 ;
        RECT 46.810 127.345 46.980 127.435 ;
        RECT 45.405 127.015 46.080 127.265 ;
        RECT 46.300 127.015 46.640 127.265 ;
        RECT 46.810 127.015 47.100 127.345 ;
        RECT 45.405 126.655 45.670 127.015 ;
        RECT 46.810 126.765 46.980 127.015 ;
        RECT 44.240 125.705 44.570 126.425 ;
        RECT 44.760 125.875 45.220 126.425 ;
        RECT 46.040 126.595 46.980 126.765 ;
        RECT 45.590 125.705 45.870 126.375 ;
        RECT 46.040 126.045 46.340 126.595 ;
        RECT 47.270 126.425 47.520 127.795 ;
        RECT 47.690 127.530 47.980 128.255 ;
        RECT 48.610 127.795 49.170 128.085 ;
        RECT 49.340 127.795 49.590 128.255 ;
        RECT 46.540 125.705 46.870 126.425 ;
        RECT 47.060 125.875 47.520 126.425 ;
        RECT 47.690 125.705 47.980 126.870 ;
        RECT 48.610 126.425 48.860 127.795 ;
        RECT 50.210 127.625 50.540 127.985 ;
        RECT 49.150 127.435 50.540 127.625 ;
        RECT 50.910 127.505 52.120 128.255 ;
        RECT 52.810 127.785 53.110 128.255 ;
        RECT 53.280 127.615 53.535 128.060 ;
        RECT 53.705 127.785 53.965 128.255 ;
        RECT 54.135 127.615 54.395 128.060 ;
        RECT 54.565 127.785 54.860 128.255 ;
        RECT 49.150 127.345 49.320 127.435 ;
        RECT 49.030 127.015 49.320 127.345 ;
        RECT 49.490 127.015 49.830 127.265 ;
        RECT 50.050 127.015 50.725 127.265 ;
        RECT 49.150 126.765 49.320 127.015 ;
        RECT 49.150 126.595 50.090 126.765 ;
        RECT 50.460 126.655 50.725 127.015 ;
        RECT 50.910 126.795 51.430 127.335 ;
        RECT 51.600 126.965 52.120 127.505 ;
        RECT 52.290 127.445 55.320 127.615 ;
        RECT 55.510 127.485 57.180 128.255 ;
        RECT 57.440 127.705 57.610 128.085 ;
        RECT 57.790 127.875 58.120 128.255 ;
        RECT 57.440 127.535 58.105 127.705 ;
        RECT 58.300 127.580 58.560 128.085 ;
        RECT 52.290 126.880 52.590 127.445 ;
        RECT 52.765 127.050 54.980 127.275 ;
        RECT 55.150 126.880 55.320 127.445 ;
        RECT 48.610 125.875 49.070 126.425 ;
        RECT 49.260 125.705 49.590 126.425 ;
        RECT 49.790 126.045 50.090 126.595 ;
        RECT 50.260 125.705 50.540 126.375 ;
        RECT 50.910 125.705 52.120 126.795 ;
        RECT 52.290 126.710 55.320 126.880 ;
        RECT 55.510 126.795 56.260 127.315 ;
        RECT 56.430 126.965 57.180 127.485 ;
        RECT 57.370 126.985 57.700 127.355 ;
        RECT 57.935 127.280 58.105 127.535 ;
        RECT 57.935 126.950 58.220 127.280 ;
        RECT 57.935 126.805 58.105 126.950 ;
        RECT 52.290 125.705 52.675 126.540 ;
        RECT 52.845 125.905 53.105 126.710 ;
        RECT 53.275 125.705 53.535 126.540 ;
        RECT 53.705 125.905 53.960 126.710 ;
        RECT 54.135 125.705 54.395 126.540 ;
        RECT 54.565 125.905 54.820 126.710 ;
        RECT 54.995 125.705 55.340 126.540 ;
        RECT 55.510 125.705 57.180 126.795 ;
        RECT 57.440 126.635 58.105 126.805 ;
        RECT 58.390 126.780 58.560 127.580 ;
        RECT 57.440 125.875 57.610 126.635 ;
        RECT 57.790 125.705 58.120 126.465 ;
        RECT 58.290 125.875 58.560 126.780 ;
        RECT 58.730 127.755 58.990 128.085 ;
        RECT 59.200 127.775 59.475 128.255 ;
        RECT 58.730 126.845 58.900 127.755 ;
        RECT 59.685 127.685 59.890 128.085 ;
        RECT 60.060 127.855 60.395 128.255 ;
        RECT 60.575 127.855 60.910 128.255 ;
        RECT 61.080 127.685 61.285 128.085 ;
        RECT 61.495 127.775 61.770 128.255 ;
        RECT 61.980 127.755 62.240 128.085 ;
        RECT 59.070 127.015 59.430 127.595 ;
        RECT 59.685 127.515 60.370 127.685 ;
        RECT 59.610 126.845 59.860 127.345 ;
        RECT 58.730 126.675 59.860 126.845 ;
        RECT 58.730 125.905 59.000 126.675 ;
        RECT 60.030 126.485 60.370 127.515 ;
        RECT 59.170 125.705 59.500 126.485 ;
        RECT 59.705 126.310 60.370 126.485 ;
        RECT 60.600 127.515 61.285 127.685 ;
        RECT 60.600 126.485 60.940 127.515 ;
        RECT 61.110 126.845 61.360 127.345 ;
        RECT 61.540 127.015 61.900 127.595 ;
        RECT 62.070 126.845 62.240 127.755 ;
        RECT 61.110 126.675 62.240 126.845 ;
        RECT 60.600 126.310 61.265 126.485 ;
        RECT 59.705 125.905 59.890 126.310 ;
        RECT 60.060 125.705 60.395 126.130 ;
        RECT 60.575 125.705 60.910 126.130 ;
        RECT 61.080 125.905 61.265 126.310 ;
        RECT 61.470 125.705 61.800 126.485 ;
        RECT 61.970 125.905 62.240 126.675 ;
        RECT 62.410 127.795 62.970 128.085 ;
        RECT 63.140 127.795 63.390 128.255 ;
        RECT 62.410 126.425 62.660 127.795 ;
        RECT 64.010 127.625 64.340 127.985 ;
        RECT 62.950 127.435 64.340 127.625 ;
        RECT 64.710 127.485 68.220 128.255 ;
        RECT 62.950 127.345 63.120 127.435 ;
        RECT 62.830 127.015 63.120 127.345 ;
        RECT 63.290 127.015 63.630 127.265 ;
        RECT 63.850 127.015 64.525 127.265 ;
        RECT 62.950 126.765 63.120 127.015 ;
        RECT 62.950 126.595 63.890 126.765 ;
        RECT 64.260 126.655 64.525 127.015 ;
        RECT 64.710 126.795 66.400 127.315 ;
        RECT 66.570 126.965 68.220 127.485 ;
        RECT 68.590 127.625 68.920 127.985 ;
        RECT 69.540 127.795 69.790 128.255 ;
        RECT 69.960 127.795 70.520 128.085 ;
        RECT 68.590 127.435 69.980 127.625 ;
        RECT 69.810 127.345 69.980 127.435 ;
        RECT 68.405 127.015 69.080 127.265 ;
        RECT 69.300 127.015 69.640 127.265 ;
        RECT 69.810 127.015 70.100 127.345 ;
        RECT 62.410 125.875 62.870 126.425 ;
        RECT 63.060 125.705 63.390 126.425 ;
        RECT 63.590 126.045 63.890 126.595 ;
        RECT 64.060 125.705 64.340 126.375 ;
        RECT 64.710 125.705 68.220 126.795 ;
        RECT 68.405 126.655 68.670 127.015 ;
        RECT 69.810 126.765 69.980 127.015 ;
        RECT 69.040 126.595 69.980 126.765 ;
        RECT 68.590 125.705 68.870 126.375 ;
        RECT 69.040 126.045 69.340 126.595 ;
        RECT 70.270 126.425 70.520 127.795 ;
        RECT 69.540 125.705 69.870 126.425 ;
        RECT 70.060 125.875 70.520 126.425 ;
        RECT 70.690 127.580 70.960 127.925 ;
        RECT 71.150 127.855 71.530 128.255 ;
        RECT 71.700 127.685 71.870 128.035 ;
        RECT 72.040 127.855 72.370 128.255 ;
        RECT 72.570 127.685 72.740 128.035 ;
        RECT 72.940 127.755 73.270 128.255 ;
        RECT 70.690 126.845 70.860 127.580 ;
        RECT 71.130 127.515 72.740 127.685 ;
        RECT 71.130 127.345 71.300 127.515 ;
        RECT 71.030 127.015 71.300 127.345 ;
        RECT 71.470 127.015 71.875 127.345 ;
        RECT 71.130 126.845 71.300 127.015 ;
        RECT 70.690 125.875 70.960 126.845 ;
        RECT 71.130 126.675 71.855 126.845 ;
        RECT 72.045 126.725 72.755 127.345 ;
        RECT 72.925 127.015 73.275 127.585 ;
        RECT 73.450 127.530 73.740 128.255 ;
        RECT 74.645 127.445 74.890 128.050 ;
        RECT 75.110 127.720 75.620 128.255 ;
        RECT 74.370 127.275 75.600 127.445 ;
        RECT 71.685 126.555 71.855 126.675 ;
        RECT 72.955 126.555 73.275 126.845 ;
        RECT 71.170 125.705 71.450 126.505 ;
        RECT 71.685 126.385 73.275 126.555 ;
        RECT 71.620 125.925 73.275 126.215 ;
        RECT 73.450 125.705 73.740 126.870 ;
        RECT 74.370 126.465 74.710 127.275 ;
        RECT 74.880 126.710 75.630 126.900 ;
        RECT 74.370 126.055 74.885 126.465 ;
        RECT 75.120 125.705 75.290 126.465 ;
        RECT 75.460 126.045 75.630 126.710 ;
        RECT 75.800 126.725 75.990 128.085 ;
        RECT 76.160 127.915 76.435 128.085 ;
        RECT 76.160 127.745 76.440 127.915 ;
        RECT 76.160 126.925 76.435 127.745 ;
        RECT 76.625 127.720 77.155 128.085 ;
        RECT 77.580 127.855 77.910 128.255 ;
        RECT 76.980 127.685 77.155 127.720 ;
        RECT 76.640 126.725 76.810 127.525 ;
        RECT 75.800 126.555 76.810 126.725 ;
        RECT 76.980 127.515 77.910 127.685 ;
        RECT 78.080 127.515 78.335 128.085 ;
        RECT 79.180 127.565 79.510 128.255 ;
        RECT 79.970 127.660 80.590 128.085 ;
        RECT 80.760 127.765 81.090 128.255 ;
        RECT 76.980 126.385 77.150 127.515 ;
        RECT 77.740 127.345 77.910 127.515 ;
        RECT 76.025 126.215 77.150 126.385 ;
        RECT 77.320 127.015 77.515 127.345 ;
        RECT 77.740 127.015 77.995 127.345 ;
        RECT 77.320 126.045 77.490 127.015 ;
        RECT 78.165 126.845 78.335 127.515 ;
        RECT 80.230 127.325 80.590 127.660 ;
        RECT 79.170 127.045 80.590 127.325 ;
        RECT 75.460 125.875 77.490 126.045 ;
        RECT 77.660 125.705 77.830 126.845 ;
        RECT 78.000 125.875 78.335 126.845 ;
        RECT 78.640 125.705 78.970 126.875 ;
        RECT 79.170 125.875 79.500 127.045 ;
        RECT 79.700 125.705 80.030 126.875 ;
        RECT 80.230 125.875 80.590 127.045 ;
        RECT 80.760 127.015 81.100 127.595 ;
        RECT 81.330 127.435 81.540 128.255 ;
        RECT 81.710 127.455 82.040 128.085 ;
        RECT 81.710 126.855 81.960 127.455 ;
        RECT 82.210 127.435 82.440 128.255 ;
        RECT 83.200 127.705 83.370 127.995 ;
        RECT 83.540 127.875 83.870 128.255 ;
        RECT 83.200 127.535 83.865 127.705 ;
        RECT 82.130 127.015 82.460 127.265 ;
        RECT 80.760 125.705 81.090 126.845 ;
        RECT 81.330 125.705 81.540 126.845 ;
        RECT 81.710 125.875 82.040 126.855 ;
        RECT 82.210 125.705 82.440 126.845 ;
        RECT 83.115 126.715 83.465 127.365 ;
        RECT 83.635 126.545 83.865 127.535 ;
        RECT 83.200 126.375 83.865 126.545 ;
        RECT 83.200 125.875 83.370 126.375 ;
        RECT 83.540 125.705 83.870 126.205 ;
        RECT 84.040 125.875 84.265 127.995 ;
        RECT 84.480 127.875 84.810 128.255 ;
        RECT 84.980 127.705 85.150 128.035 ;
        RECT 85.450 127.875 86.465 128.075 ;
        RECT 84.455 127.515 85.150 127.705 ;
        RECT 84.455 126.545 84.625 127.515 ;
        RECT 84.795 126.715 85.205 127.335 ;
        RECT 85.375 126.765 85.595 127.635 ;
        RECT 85.775 127.325 86.125 127.695 ;
        RECT 86.295 127.145 86.465 127.875 ;
        RECT 86.635 127.815 87.045 128.255 ;
        RECT 87.335 127.615 87.585 128.045 ;
        RECT 87.785 127.795 88.105 128.255 ;
        RECT 88.665 127.865 89.515 128.035 ;
        RECT 86.635 127.275 87.045 127.605 ;
        RECT 87.335 127.275 87.755 127.615 ;
        RECT 86.045 127.105 86.465 127.145 ;
        RECT 86.045 126.935 87.395 127.105 ;
        RECT 84.455 126.375 85.150 126.545 ;
        RECT 85.375 126.385 85.875 126.765 ;
        RECT 84.480 125.705 84.810 126.205 ;
        RECT 84.980 125.875 85.150 126.375 ;
        RECT 86.045 126.090 86.215 126.935 ;
        RECT 87.145 126.775 87.395 126.935 ;
        RECT 86.385 126.505 86.635 126.765 ;
        RECT 87.565 126.505 87.755 127.275 ;
        RECT 86.385 126.255 87.755 126.505 ;
        RECT 87.925 127.445 89.175 127.615 ;
        RECT 87.925 126.685 88.095 127.445 ;
        RECT 88.845 127.325 89.175 127.445 ;
        RECT 88.265 126.865 88.445 127.275 ;
        RECT 89.345 127.105 89.515 127.865 ;
        RECT 89.715 127.775 90.375 128.255 ;
        RECT 90.555 127.660 90.875 127.990 ;
        RECT 89.705 127.335 90.365 127.605 ;
        RECT 89.705 127.275 90.035 127.335 ;
        RECT 90.185 127.105 90.515 127.165 ;
        RECT 88.615 126.935 90.515 127.105 ;
        RECT 87.925 126.375 88.445 126.685 ;
        RECT 88.615 126.425 88.785 126.935 ;
        RECT 90.685 126.765 90.875 127.660 ;
        RECT 88.955 126.595 90.875 126.765 ;
        RECT 90.555 126.575 90.875 126.595 ;
        RECT 91.075 127.345 91.325 127.995 ;
        RECT 91.505 127.795 91.790 128.255 ;
        RECT 91.970 127.545 92.225 128.075 ;
        RECT 91.075 127.015 91.875 127.345 ;
        RECT 88.615 126.255 89.825 126.425 ;
        RECT 85.385 125.920 86.215 126.090 ;
        RECT 86.455 125.705 86.835 126.085 ;
        RECT 87.015 125.965 87.185 126.255 ;
        RECT 88.615 126.175 88.785 126.255 ;
        RECT 87.355 125.705 87.685 126.085 ;
        RECT 88.155 125.925 88.785 126.175 ;
        RECT 88.965 125.705 89.385 126.085 ;
        RECT 89.585 125.965 89.825 126.255 ;
        RECT 90.055 125.705 90.385 126.395 ;
        RECT 90.555 125.965 90.725 126.575 ;
        RECT 91.075 126.425 91.325 127.015 ;
        RECT 92.045 126.685 92.225 127.545 ;
        RECT 90.995 125.915 91.325 126.425 ;
        RECT 91.505 125.705 91.790 126.505 ;
        RECT 91.970 126.215 92.225 126.685 ;
        RECT 93.690 127.795 94.250 128.085 ;
        RECT 94.420 127.795 94.670 128.255 ;
        RECT 93.690 126.425 93.940 127.795 ;
        RECT 95.290 127.625 95.620 127.985 ;
        RECT 94.230 127.435 95.620 127.625 ;
        RECT 96.910 127.795 97.470 128.085 ;
        RECT 97.640 127.795 97.890 128.255 ;
        RECT 94.230 127.345 94.400 127.435 ;
        RECT 94.110 127.015 94.400 127.345 ;
        RECT 94.570 127.015 94.910 127.265 ;
        RECT 95.130 127.015 95.805 127.265 ;
        RECT 94.230 126.765 94.400 127.015 ;
        RECT 94.230 126.595 95.170 126.765 ;
        RECT 95.540 126.655 95.805 127.015 ;
        RECT 91.970 126.045 92.310 126.215 ;
        RECT 91.970 126.015 92.225 126.045 ;
        RECT 93.690 125.875 94.150 126.425 ;
        RECT 94.340 125.705 94.670 126.425 ;
        RECT 94.870 126.045 95.170 126.595 ;
        RECT 96.910 126.425 97.160 127.795 ;
        RECT 98.510 127.625 98.840 127.985 ;
        RECT 97.450 127.435 98.840 127.625 ;
        RECT 99.210 127.530 99.500 128.255 ;
        RECT 100.170 127.435 100.400 128.255 ;
        RECT 100.570 127.455 100.900 128.085 ;
        RECT 97.450 127.345 97.620 127.435 ;
        RECT 97.330 127.015 97.620 127.345 ;
        RECT 97.790 127.015 98.130 127.265 ;
        RECT 98.350 127.015 99.025 127.265 ;
        RECT 100.150 127.015 100.480 127.265 ;
        RECT 97.450 126.765 97.620 127.015 ;
        RECT 97.450 126.595 98.390 126.765 ;
        RECT 98.760 126.655 99.025 127.015 ;
        RECT 95.340 125.705 95.620 126.375 ;
        RECT 96.910 125.875 97.370 126.425 ;
        RECT 97.560 125.705 97.890 126.425 ;
        RECT 98.090 126.045 98.390 126.595 ;
        RECT 98.560 125.705 98.840 126.375 ;
        RECT 99.210 125.705 99.500 126.870 ;
        RECT 100.650 126.855 100.900 127.455 ;
        RECT 101.070 127.435 101.280 128.255 ;
        RECT 101.885 127.545 102.140 128.075 ;
        RECT 102.320 127.795 102.605 128.255 ;
        RECT 101.885 126.895 102.065 127.545 ;
        RECT 102.785 127.345 103.035 127.995 ;
        RECT 102.235 127.015 103.035 127.345 ;
        RECT 100.170 125.705 100.400 126.845 ;
        RECT 100.570 125.875 100.900 126.855 ;
        RECT 101.070 125.705 101.280 126.845 ;
        RECT 101.800 126.725 102.065 126.895 ;
        RECT 101.885 126.685 102.065 126.725 ;
        RECT 101.885 126.015 102.140 126.685 ;
        RECT 102.320 125.705 102.605 126.505 ;
        RECT 102.785 126.425 103.035 127.015 ;
        RECT 103.235 127.660 103.555 127.990 ;
        RECT 103.735 127.775 104.395 128.255 ;
        RECT 104.595 127.865 105.445 128.035 ;
        RECT 103.235 126.765 103.425 127.660 ;
        RECT 103.745 127.335 104.405 127.605 ;
        RECT 104.075 127.275 104.405 127.335 ;
        RECT 103.595 127.105 103.925 127.165 ;
        RECT 104.595 127.105 104.765 127.865 ;
        RECT 106.005 127.795 106.325 128.255 ;
        RECT 106.525 127.615 106.775 128.045 ;
        RECT 107.065 127.815 107.475 128.255 ;
        RECT 107.645 127.875 108.660 128.075 ;
        RECT 104.935 127.445 106.185 127.615 ;
        RECT 104.935 127.325 105.265 127.445 ;
        RECT 103.595 126.935 105.495 127.105 ;
        RECT 103.235 126.595 105.155 126.765 ;
        RECT 103.235 126.575 103.555 126.595 ;
        RECT 102.785 125.915 103.115 126.425 ;
        RECT 103.385 125.965 103.555 126.575 ;
        RECT 105.325 126.425 105.495 126.935 ;
        RECT 105.665 126.865 105.845 127.275 ;
        RECT 106.015 126.685 106.185 127.445 ;
        RECT 103.725 125.705 104.055 126.395 ;
        RECT 104.285 126.255 105.495 126.425 ;
        RECT 105.665 126.375 106.185 126.685 ;
        RECT 106.355 127.275 106.775 127.615 ;
        RECT 107.065 127.275 107.475 127.605 ;
        RECT 106.355 126.505 106.545 127.275 ;
        RECT 107.645 127.145 107.815 127.875 ;
        RECT 108.960 127.705 109.130 128.035 ;
        RECT 109.300 127.875 109.630 128.255 ;
        RECT 107.985 127.325 108.335 127.695 ;
        RECT 107.645 127.105 108.065 127.145 ;
        RECT 106.715 126.935 108.065 127.105 ;
        RECT 106.715 126.775 106.965 126.935 ;
        RECT 107.475 126.505 107.725 126.765 ;
        RECT 106.355 126.255 107.725 126.505 ;
        RECT 104.285 125.965 104.525 126.255 ;
        RECT 105.325 126.175 105.495 126.255 ;
        RECT 104.725 125.705 105.145 126.085 ;
        RECT 105.325 125.925 105.955 126.175 ;
        RECT 106.425 125.705 106.755 126.085 ;
        RECT 106.925 125.965 107.095 126.255 ;
        RECT 107.895 126.090 108.065 126.935 ;
        RECT 108.515 126.765 108.735 127.635 ;
        RECT 108.960 127.515 109.655 127.705 ;
        RECT 108.235 126.385 108.735 126.765 ;
        RECT 108.905 126.715 109.315 127.335 ;
        RECT 109.485 126.545 109.655 127.515 ;
        RECT 108.960 126.375 109.655 126.545 ;
        RECT 107.275 125.705 107.655 126.085 ;
        RECT 107.895 125.920 108.725 126.090 ;
        RECT 108.960 125.875 109.130 126.375 ;
        RECT 109.300 125.705 109.630 126.205 ;
        RECT 109.845 125.875 110.070 127.995 ;
        RECT 110.240 127.875 110.570 128.255 ;
        RECT 110.740 127.705 110.910 127.995 ;
        RECT 110.245 127.535 110.910 127.705 ;
        RECT 110.245 126.545 110.475 127.535 ;
        RECT 111.170 127.505 112.380 128.255 ;
        RECT 110.645 126.715 110.995 127.365 ;
        RECT 111.170 126.795 111.690 127.335 ;
        RECT 111.860 126.965 112.380 127.505 ;
        RECT 110.245 126.375 110.910 126.545 ;
        RECT 110.240 125.705 110.570 126.205 ;
        RECT 110.740 125.875 110.910 126.375 ;
        RECT 111.170 125.705 112.380 126.795 ;
        RECT 18.165 125.535 112.465 125.705 ;
        RECT 18.250 124.445 19.460 125.535 ;
        RECT 20.005 125.195 20.260 125.225 ;
        RECT 19.920 125.025 20.260 125.195 ;
        RECT 18.250 123.735 18.770 124.275 ;
        RECT 18.940 123.905 19.460 124.445 ;
        RECT 20.005 124.555 20.260 125.025 ;
        RECT 20.440 124.735 20.725 125.535 ;
        RECT 20.905 124.815 21.235 125.325 ;
        RECT 18.250 122.985 19.460 123.735 ;
        RECT 20.005 123.695 20.185 124.555 ;
        RECT 20.905 124.225 21.155 124.815 ;
        RECT 21.505 124.665 21.675 125.275 ;
        RECT 21.845 124.845 22.175 125.535 ;
        RECT 22.405 124.985 22.645 125.275 ;
        RECT 22.845 125.155 23.265 125.535 ;
        RECT 23.445 125.065 24.075 125.315 ;
        RECT 24.545 125.155 24.875 125.535 ;
        RECT 23.445 124.985 23.615 125.065 ;
        RECT 25.045 124.985 25.215 125.275 ;
        RECT 25.395 125.155 25.775 125.535 ;
        RECT 26.015 125.150 26.845 125.320 ;
        RECT 22.405 124.815 23.615 124.985 ;
        RECT 20.355 123.895 21.155 124.225 ;
        RECT 20.005 123.165 20.260 123.695 ;
        RECT 20.440 122.985 20.725 123.445 ;
        RECT 20.905 123.245 21.155 123.895 ;
        RECT 21.355 124.645 21.675 124.665 ;
        RECT 21.355 124.475 23.275 124.645 ;
        RECT 21.355 123.580 21.545 124.475 ;
        RECT 23.445 124.305 23.615 124.815 ;
        RECT 23.785 124.555 24.305 124.865 ;
        RECT 21.715 124.135 23.615 124.305 ;
        RECT 21.715 124.075 22.045 124.135 ;
        RECT 22.195 123.905 22.525 123.965 ;
        RECT 21.865 123.635 22.525 123.905 ;
        RECT 21.355 123.250 21.675 123.580 ;
        RECT 21.855 122.985 22.515 123.465 ;
        RECT 22.715 123.375 22.885 124.135 ;
        RECT 23.785 123.965 23.965 124.375 ;
        RECT 23.055 123.795 23.385 123.915 ;
        RECT 24.135 123.795 24.305 124.555 ;
        RECT 23.055 123.625 24.305 123.795 ;
        RECT 24.475 124.735 25.845 124.985 ;
        RECT 24.475 123.965 24.665 124.735 ;
        RECT 25.595 124.475 25.845 124.735 ;
        RECT 24.835 124.305 25.085 124.465 ;
        RECT 26.015 124.305 26.185 125.150 ;
        RECT 27.080 124.865 27.250 125.365 ;
        RECT 27.420 125.035 27.750 125.535 ;
        RECT 26.355 124.475 26.855 124.855 ;
        RECT 27.080 124.695 27.775 124.865 ;
        RECT 24.835 124.135 26.185 124.305 ;
        RECT 25.765 124.095 26.185 124.135 ;
        RECT 24.475 123.625 24.895 123.965 ;
        RECT 25.185 123.635 25.595 123.965 ;
        RECT 22.715 123.205 23.565 123.375 ;
        RECT 24.125 122.985 24.445 123.445 ;
        RECT 24.645 123.195 24.895 123.625 ;
        RECT 25.185 122.985 25.595 123.425 ;
        RECT 25.765 123.365 25.935 124.095 ;
        RECT 26.105 123.545 26.455 123.915 ;
        RECT 26.635 123.605 26.855 124.475 ;
        RECT 27.025 123.905 27.435 124.525 ;
        RECT 27.605 123.725 27.775 124.695 ;
        RECT 27.080 123.535 27.775 123.725 ;
        RECT 25.765 123.165 26.780 123.365 ;
        RECT 27.080 123.205 27.250 123.535 ;
        RECT 27.420 122.985 27.750 123.365 ;
        RECT 27.965 123.245 28.190 125.365 ;
        RECT 28.360 125.035 28.690 125.535 ;
        RECT 28.860 124.865 29.030 125.365 ;
        RECT 29.950 124.865 30.230 125.535 ;
        RECT 28.365 124.695 29.030 124.865 ;
        RECT 28.365 123.705 28.595 124.695 ;
        RECT 30.400 124.645 30.700 125.195 ;
        RECT 30.900 124.815 31.230 125.535 ;
        RECT 31.420 124.815 31.880 125.365 ;
        RECT 28.765 123.875 29.115 124.525 ;
        RECT 29.765 124.225 30.030 124.585 ;
        RECT 30.400 124.475 31.340 124.645 ;
        RECT 31.170 124.225 31.340 124.475 ;
        RECT 29.765 123.975 30.440 124.225 ;
        RECT 30.660 123.975 31.000 124.225 ;
        RECT 31.170 123.895 31.460 124.225 ;
        RECT 31.170 123.805 31.340 123.895 ;
        RECT 28.365 123.535 29.030 123.705 ;
        RECT 28.360 122.985 28.690 123.365 ;
        RECT 28.860 123.245 29.030 123.535 ;
        RECT 29.950 123.615 31.340 123.805 ;
        RECT 29.950 123.255 30.280 123.615 ;
        RECT 31.630 123.445 31.880 124.815 ;
        RECT 30.900 122.985 31.150 123.445 ;
        RECT 31.320 123.155 31.880 123.445 ;
        RECT 32.050 124.815 32.510 125.365 ;
        RECT 32.700 124.815 33.030 125.535 ;
        RECT 32.050 123.445 32.300 124.815 ;
        RECT 33.230 124.645 33.530 125.195 ;
        RECT 33.700 124.865 33.980 125.535 ;
        RECT 32.590 124.475 33.530 124.645 ;
        RECT 32.590 124.225 32.760 124.475 ;
        RECT 33.900 124.225 34.165 124.585 ;
        RECT 34.810 124.370 35.100 125.535 ;
        RECT 35.360 124.790 35.630 125.535 ;
        RECT 36.260 125.530 42.535 125.535 ;
        RECT 35.800 124.620 36.090 125.360 ;
        RECT 36.260 124.805 36.515 125.530 ;
        RECT 36.700 124.635 36.960 125.360 ;
        RECT 37.130 124.805 37.375 125.530 ;
        RECT 37.560 124.635 37.820 125.360 ;
        RECT 37.990 124.805 38.235 125.530 ;
        RECT 38.420 124.635 38.680 125.360 ;
        RECT 38.850 124.805 39.095 125.530 ;
        RECT 39.265 124.635 39.525 125.360 ;
        RECT 39.695 124.805 39.955 125.530 ;
        RECT 40.125 124.635 40.385 125.360 ;
        RECT 40.555 124.805 40.815 125.530 ;
        RECT 40.985 124.635 41.245 125.360 ;
        RECT 41.415 124.805 41.675 125.530 ;
        RECT 41.845 124.635 42.105 125.360 ;
        RECT 42.275 124.735 42.535 125.530 ;
        RECT 36.700 124.620 42.105 124.635 ;
        RECT 35.360 124.395 42.105 124.620 ;
        RECT 32.470 123.895 32.760 124.225 ;
        RECT 32.930 123.975 33.270 124.225 ;
        RECT 33.490 123.975 34.165 124.225 ;
        RECT 32.590 123.805 32.760 123.895 ;
        RECT 35.360 123.805 36.525 124.395 ;
        RECT 42.705 124.225 42.955 125.360 ;
        RECT 43.135 124.725 43.395 125.535 ;
        RECT 43.570 124.225 43.815 125.365 ;
        RECT 43.995 124.725 44.290 125.535 ;
        RECT 45.020 124.605 45.190 125.365 ;
        RECT 45.370 124.775 45.700 125.535 ;
        RECT 45.020 124.435 45.685 124.605 ;
        RECT 45.870 124.460 46.140 125.365 ;
        RECT 46.320 124.725 46.615 125.535 ;
        RECT 45.515 124.290 45.685 124.435 ;
        RECT 36.695 123.975 43.815 124.225 ;
        RECT 32.590 123.615 33.980 123.805 ;
        RECT 32.050 123.155 32.610 123.445 ;
        RECT 32.780 122.985 33.030 123.445 ;
        RECT 33.650 123.255 33.980 123.615 ;
        RECT 34.810 122.985 35.100 123.710 ;
        RECT 35.360 123.635 42.105 123.805 ;
        RECT 35.360 122.985 35.660 123.465 ;
        RECT 35.830 123.180 36.090 123.635 ;
        RECT 36.260 122.985 36.520 123.465 ;
        RECT 36.700 123.180 36.960 123.635 ;
        RECT 37.130 122.985 37.380 123.465 ;
        RECT 37.560 123.180 37.820 123.635 ;
        RECT 37.990 122.985 38.240 123.465 ;
        RECT 38.420 123.180 38.680 123.635 ;
        RECT 38.850 122.985 39.095 123.465 ;
        RECT 39.265 123.180 39.540 123.635 ;
        RECT 39.710 122.985 39.955 123.465 ;
        RECT 40.125 123.180 40.385 123.635 ;
        RECT 40.555 122.985 40.815 123.465 ;
        RECT 40.985 123.180 41.245 123.635 ;
        RECT 41.415 122.985 41.675 123.465 ;
        RECT 41.845 123.180 42.105 123.635 ;
        RECT 42.275 122.985 42.535 123.545 ;
        RECT 42.705 123.165 42.955 123.975 ;
        RECT 43.135 122.985 43.395 123.510 ;
        RECT 43.565 123.165 43.815 123.975 ;
        RECT 43.985 123.665 44.300 124.225 ;
        RECT 44.950 123.885 45.280 124.255 ;
        RECT 45.515 123.960 45.800 124.290 ;
        RECT 45.515 123.705 45.685 123.960 ;
        RECT 45.020 123.535 45.685 123.705 ;
        RECT 45.970 123.660 46.140 124.460 ;
        RECT 46.795 124.225 47.040 125.365 ;
        RECT 47.215 124.725 47.475 125.535 ;
        RECT 48.075 125.530 54.350 125.535 ;
        RECT 47.655 124.225 47.905 125.360 ;
        RECT 48.075 124.735 48.335 125.530 ;
        RECT 48.505 124.635 48.765 125.360 ;
        RECT 48.935 124.805 49.195 125.530 ;
        RECT 49.365 124.635 49.625 125.360 ;
        RECT 49.795 124.805 50.055 125.530 ;
        RECT 50.225 124.635 50.485 125.360 ;
        RECT 50.655 124.805 50.915 125.530 ;
        RECT 51.085 124.635 51.345 125.360 ;
        RECT 51.515 124.805 51.760 125.530 ;
        RECT 51.930 124.635 52.190 125.360 ;
        RECT 52.375 124.805 52.620 125.530 ;
        RECT 52.790 124.635 53.050 125.360 ;
        RECT 53.235 124.805 53.480 125.530 ;
        RECT 53.650 124.635 53.910 125.360 ;
        RECT 54.095 124.805 54.350 125.530 ;
        RECT 48.505 124.620 53.910 124.635 ;
        RECT 54.520 124.620 54.810 125.360 ;
        RECT 54.980 124.790 55.250 125.535 ;
        RECT 48.505 124.395 55.250 124.620 ;
        RECT 46.310 123.665 46.625 124.225 ;
        RECT 46.795 123.975 53.915 124.225 ;
        RECT 43.995 122.985 44.300 123.495 ;
        RECT 45.020 123.155 45.190 123.535 ;
        RECT 45.370 122.985 45.700 123.365 ;
        RECT 45.880 123.155 46.140 123.660 ;
        RECT 46.310 122.985 46.615 123.495 ;
        RECT 46.795 123.165 47.045 123.975 ;
        RECT 47.215 122.985 47.475 123.510 ;
        RECT 47.655 123.165 47.905 123.975 ;
        RECT 54.085 123.805 55.250 124.395 ;
        RECT 55.510 124.445 56.720 125.535 ;
        RECT 56.945 124.665 57.230 125.535 ;
        RECT 57.400 124.905 57.660 125.365 ;
        RECT 57.835 125.075 58.090 125.535 ;
        RECT 58.260 124.905 58.520 125.365 ;
        RECT 57.400 124.735 58.520 124.905 ;
        RECT 58.690 124.735 59.000 125.535 ;
        RECT 57.400 124.485 57.660 124.735 ;
        RECT 59.170 124.565 59.480 125.365 ;
        RECT 55.510 123.905 56.030 124.445 ;
        RECT 56.905 124.315 57.660 124.485 ;
        RECT 58.450 124.395 59.480 124.565 ;
        RECT 48.505 123.635 55.250 123.805 ;
        RECT 56.200 123.735 56.720 124.275 ;
        RECT 48.075 122.985 48.335 123.545 ;
        RECT 48.505 123.180 48.765 123.635 ;
        RECT 48.935 122.985 49.195 123.465 ;
        RECT 49.365 123.180 49.625 123.635 ;
        RECT 49.795 122.985 50.055 123.465 ;
        RECT 50.225 123.180 50.485 123.635 ;
        RECT 50.655 122.985 50.900 123.465 ;
        RECT 51.070 123.180 51.345 123.635 ;
        RECT 51.515 122.985 51.760 123.465 ;
        RECT 51.930 123.180 52.190 123.635 ;
        RECT 52.370 122.985 52.620 123.465 ;
        RECT 52.790 123.180 53.050 123.635 ;
        RECT 53.230 122.985 53.480 123.465 ;
        RECT 53.650 123.180 53.910 123.635 ;
        RECT 54.090 122.985 54.350 123.465 ;
        RECT 54.520 123.180 54.780 123.635 ;
        RECT 54.950 122.985 55.250 123.465 ;
        RECT 55.510 122.985 56.720 123.735 ;
        RECT 56.905 123.805 57.310 124.315 ;
        RECT 58.450 124.145 58.620 124.395 ;
        RECT 57.480 123.975 58.620 124.145 ;
        RECT 56.905 123.635 58.555 123.805 ;
        RECT 58.790 123.655 59.140 124.225 ;
        RECT 56.950 122.985 57.230 123.465 ;
        RECT 57.400 123.245 57.660 123.635 ;
        RECT 57.835 122.985 58.090 123.465 ;
        RECT 58.260 123.245 58.555 123.635 ;
        RECT 59.310 123.485 59.480 124.395 ;
        RECT 60.570 124.370 60.860 125.535 ;
        RECT 61.030 124.445 62.700 125.535 ;
        RECT 62.870 124.565 63.180 125.365 ;
        RECT 63.350 124.735 63.660 125.535 ;
        RECT 63.830 124.905 64.090 125.365 ;
        RECT 64.260 125.075 64.515 125.535 ;
        RECT 64.690 124.905 64.950 125.365 ;
        RECT 63.830 124.735 64.950 124.905 ;
        RECT 61.030 123.925 61.780 124.445 ;
        RECT 62.870 124.395 63.900 124.565 ;
        RECT 61.950 123.755 62.700 124.275 ;
        RECT 58.735 122.985 59.010 123.465 ;
        RECT 59.180 123.155 59.480 123.485 ;
        RECT 60.570 122.985 60.860 123.710 ;
        RECT 61.030 122.985 62.700 123.755 ;
        RECT 62.870 123.485 63.040 124.395 ;
        RECT 63.210 123.655 63.560 124.225 ;
        RECT 63.730 124.145 63.900 124.395 ;
        RECT 64.690 124.485 64.950 124.735 ;
        RECT 65.120 124.665 65.405 125.535 ;
        RECT 64.690 124.315 65.445 124.485 ;
        RECT 63.730 123.975 64.870 124.145 ;
        RECT 65.040 123.805 65.445 124.315 ;
        RECT 65.630 124.445 67.300 125.535 ;
        RECT 65.630 123.925 66.380 124.445 ;
        RECT 67.510 124.395 67.740 125.535 ;
        RECT 67.910 124.385 68.240 125.365 ;
        RECT 68.410 124.395 68.620 125.535 ;
        RECT 69.050 124.865 69.330 125.535 ;
        RECT 69.500 124.645 69.800 125.195 ;
        RECT 70.000 124.815 70.330 125.535 ;
        RECT 70.520 124.815 70.980 125.365 ;
        RECT 71.350 124.865 71.630 125.535 ;
        RECT 63.795 123.635 65.445 123.805 ;
        RECT 66.550 123.755 67.300 124.275 ;
        RECT 67.490 123.975 67.820 124.225 ;
        RECT 62.870 123.155 63.170 123.485 ;
        RECT 63.340 122.985 63.615 123.465 ;
        RECT 63.795 123.245 64.090 123.635 ;
        RECT 64.260 122.985 64.515 123.465 ;
        RECT 64.690 123.245 64.950 123.635 ;
        RECT 65.120 122.985 65.400 123.465 ;
        RECT 65.630 122.985 67.300 123.755 ;
        RECT 67.510 122.985 67.740 123.805 ;
        RECT 67.990 123.785 68.240 124.385 ;
        RECT 68.865 124.225 69.130 124.585 ;
        RECT 69.500 124.475 70.440 124.645 ;
        RECT 70.270 124.225 70.440 124.475 ;
        RECT 68.865 123.975 69.540 124.225 ;
        RECT 69.760 123.975 70.100 124.225 ;
        RECT 70.270 123.895 70.560 124.225 ;
        RECT 70.270 123.805 70.440 123.895 ;
        RECT 67.910 123.155 68.240 123.785 ;
        RECT 68.410 122.985 68.620 123.805 ;
        RECT 69.050 123.615 70.440 123.805 ;
        RECT 69.050 123.255 69.380 123.615 ;
        RECT 70.730 123.445 70.980 124.815 ;
        RECT 71.800 124.645 72.100 125.195 ;
        RECT 72.300 124.815 72.630 125.535 ;
        RECT 72.820 124.815 73.280 125.365 ;
        RECT 71.165 124.225 71.430 124.585 ;
        RECT 71.800 124.475 72.740 124.645 ;
        RECT 72.570 124.225 72.740 124.475 ;
        RECT 71.165 123.975 71.840 124.225 ;
        RECT 72.060 123.975 72.400 124.225 ;
        RECT 72.570 123.895 72.860 124.225 ;
        RECT 72.570 123.805 72.740 123.895 ;
        RECT 70.000 122.985 70.250 123.445 ;
        RECT 70.420 123.155 70.980 123.445 ;
        RECT 71.350 123.615 72.740 123.805 ;
        RECT 71.350 123.255 71.680 123.615 ;
        RECT 73.030 123.445 73.280 124.815 ;
        RECT 74.285 124.555 74.540 125.225 ;
        RECT 74.720 124.735 75.005 125.535 ;
        RECT 75.185 124.815 75.515 125.325 ;
        RECT 74.285 123.695 74.465 124.555 ;
        RECT 75.185 124.225 75.435 124.815 ;
        RECT 75.785 124.665 75.955 125.275 ;
        RECT 76.125 124.845 76.455 125.535 ;
        RECT 76.685 124.985 76.925 125.275 ;
        RECT 77.125 125.155 77.545 125.535 ;
        RECT 77.725 125.065 78.355 125.315 ;
        RECT 78.825 125.155 79.155 125.535 ;
        RECT 77.725 124.985 77.895 125.065 ;
        RECT 79.325 124.985 79.495 125.275 ;
        RECT 79.675 125.155 80.055 125.535 ;
        RECT 80.295 125.150 81.125 125.320 ;
        RECT 76.685 124.815 77.895 124.985 ;
        RECT 74.635 123.895 75.435 124.225 ;
        RECT 74.285 123.495 74.540 123.695 ;
        RECT 72.300 122.985 72.550 123.445 ;
        RECT 72.720 123.155 73.280 123.445 ;
        RECT 74.200 123.325 74.540 123.495 ;
        RECT 74.285 123.165 74.540 123.325 ;
        RECT 74.720 122.985 75.005 123.445 ;
        RECT 75.185 123.245 75.435 123.895 ;
        RECT 75.635 124.645 75.955 124.665 ;
        RECT 75.635 124.475 77.555 124.645 ;
        RECT 75.635 123.580 75.825 124.475 ;
        RECT 77.725 124.305 77.895 124.815 ;
        RECT 78.065 124.555 78.585 124.865 ;
        RECT 75.995 124.135 77.895 124.305 ;
        RECT 75.995 124.075 76.325 124.135 ;
        RECT 76.475 123.905 76.805 123.965 ;
        RECT 76.145 123.635 76.805 123.905 ;
        RECT 75.635 123.250 75.955 123.580 ;
        RECT 76.135 122.985 76.795 123.465 ;
        RECT 76.995 123.375 77.165 124.135 ;
        RECT 78.065 123.965 78.245 124.375 ;
        RECT 77.335 123.795 77.665 123.915 ;
        RECT 78.415 123.795 78.585 124.555 ;
        RECT 77.335 123.625 78.585 123.795 ;
        RECT 78.755 124.735 80.125 124.985 ;
        RECT 78.755 123.965 78.945 124.735 ;
        RECT 79.875 124.475 80.125 124.735 ;
        RECT 79.115 124.305 79.365 124.465 ;
        RECT 80.295 124.305 80.465 125.150 ;
        RECT 81.360 124.865 81.530 125.365 ;
        RECT 81.700 125.035 82.030 125.535 ;
        RECT 80.635 124.475 81.135 124.855 ;
        RECT 81.360 124.695 82.055 124.865 ;
        RECT 79.115 124.135 80.465 124.305 ;
        RECT 80.045 124.095 80.465 124.135 ;
        RECT 78.755 123.625 79.175 123.965 ;
        RECT 79.465 123.635 79.875 123.965 ;
        RECT 76.995 123.205 77.845 123.375 ;
        RECT 78.405 122.985 78.725 123.445 ;
        RECT 78.925 123.195 79.175 123.625 ;
        RECT 79.465 122.985 79.875 123.425 ;
        RECT 80.045 123.365 80.215 124.095 ;
        RECT 80.385 123.545 80.735 123.915 ;
        RECT 80.915 123.605 81.135 124.475 ;
        RECT 81.305 123.905 81.715 124.525 ;
        RECT 81.885 123.725 82.055 124.695 ;
        RECT 81.360 123.535 82.055 123.725 ;
        RECT 80.045 123.165 81.060 123.365 ;
        RECT 81.360 123.205 81.530 123.535 ;
        RECT 81.700 122.985 82.030 123.365 ;
        RECT 82.245 123.245 82.470 125.365 ;
        RECT 82.640 125.035 82.970 125.535 ;
        RECT 83.140 124.865 83.310 125.365 ;
        RECT 82.645 124.695 83.310 124.865 ;
        RECT 82.645 123.705 82.875 124.695 ;
        RECT 83.045 123.875 83.395 124.525 ;
        RECT 83.570 124.445 84.780 125.535 ;
        RECT 83.570 123.905 84.090 124.445 ;
        RECT 84.990 124.395 85.220 125.535 ;
        RECT 85.390 124.385 85.720 125.365 ;
        RECT 85.890 124.395 86.100 125.535 ;
        RECT 84.260 123.735 84.780 124.275 ;
        RECT 84.970 123.975 85.300 124.225 ;
        RECT 82.645 123.535 83.310 123.705 ;
        RECT 82.640 122.985 82.970 123.365 ;
        RECT 83.140 123.245 83.310 123.535 ;
        RECT 83.570 122.985 84.780 123.735 ;
        RECT 84.990 122.985 85.220 123.805 ;
        RECT 85.470 123.785 85.720 124.385 ;
        RECT 86.330 124.370 86.620 125.535 ;
        RECT 86.790 124.460 87.060 125.365 ;
        RECT 87.230 124.775 87.560 125.535 ;
        RECT 87.740 124.605 87.910 125.365 ;
        RECT 85.390 123.155 85.720 123.785 ;
        RECT 85.890 122.985 86.100 123.805 ;
        RECT 86.330 122.985 86.620 123.710 ;
        RECT 86.790 123.660 86.960 124.460 ;
        RECT 87.245 124.435 87.910 124.605 ;
        RECT 88.170 124.815 88.630 125.365 ;
        RECT 88.820 124.815 89.150 125.535 ;
        RECT 87.245 124.290 87.415 124.435 ;
        RECT 87.130 123.960 87.415 124.290 ;
        RECT 87.245 123.705 87.415 123.960 ;
        RECT 87.650 123.885 87.980 124.255 ;
        RECT 86.790 123.155 87.050 123.660 ;
        RECT 87.245 123.535 87.910 123.705 ;
        RECT 87.230 122.985 87.560 123.365 ;
        RECT 87.740 123.155 87.910 123.535 ;
        RECT 88.170 123.445 88.420 124.815 ;
        RECT 89.350 124.645 89.650 125.195 ;
        RECT 89.820 124.865 90.100 125.535 ;
        RECT 88.710 124.475 89.650 124.645 ;
        RECT 88.710 124.225 88.880 124.475 ;
        RECT 90.020 124.225 90.285 124.585 ;
        RECT 88.590 123.895 88.880 124.225 ;
        RECT 89.050 123.975 89.390 124.225 ;
        RECT 89.610 123.975 90.285 124.225 ;
        RECT 90.930 124.445 94.440 125.535 ;
        RECT 94.610 124.815 95.070 125.365 ;
        RECT 95.260 124.815 95.590 125.535 ;
        RECT 90.930 123.925 92.620 124.445 ;
        RECT 88.710 123.805 88.880 123.895 ;
        RECT 88.710 123.615 90.100 123.805 ;
        RECT 92.790 123.755 94.440 124.275 ;
        RECT 88.170 123.155 88.730 123.445 ;
        RECT 88.900 122.985 89.150 123.445 ;
        RECT 89.770 123.255 90.100 123.615 ;
        RECT 90.930 122.985 94.440 123.755 ;
        RECT 94.610 123.445 94.860 124.815 ;
        RECT 95.790 124.645 96.090 125.195 ;
        RECT 96.260 124.865 96.540 125.535 ;
        RECT 95.150 124.475 96.090 124.645 ;
        RECT 96.910 124.815 97.370 125.365 ;
        RECT 97.560 124.815 97.890 125.535 ;
        RECT 95.150 124.225 95.320 124.475 ;
        RECT 96.460 124.225 96.725 124.585 ;
        RECT 95.030 123.895 95.320 124.225 ;
        RECT 95.490 123.975 95.830 124.225 ;
        RECT 96.050 123.975 96.725 124.225 ;
        RECT 95.150 123.805 95.320 123.895 ;
        RECT 95.150 123.615 96.540 123.805 ;
        RECT 94.610 123.155 95.170 123.445 ;
        RECT 95.340 122.985 95.590 123.445 ;
        RECT 96.210 123.255 96.540 123.615 ;
        RECT 96.910 123.445 97.160 124.815 ;
        RECT 98.090 124.645 98.390 125.195 ;
        RECT 98.560 124.865 98.840 125.535 ;
        RECT 97.450 124.475 98.390 124.645 ;
        RECT 99.210 124.775 99.725 125.185 ;
        RECT 99.960 124.775 100.130 125.535 ;
        RECT 100.300 125.195 102.330 125.365 ;
        RECT 97.450 124.225 97.620 124.475 ;
        RECT 98.760 124.225 99.025 124.585 ;
        RECT 97.330 123.895 97.620 124.225 ;
        RECT 97.790 123.975 98.130 124.225 ;
        RECT 98.350 123.975 99.025 124.225 ;
        RECT 97.450 123.805 97.620 123.895 ;
        RECT 99.210 123.965 99.550 124.775 ;
        RECT 100.300 124.530 100.470 125.195 ;
        RECT 100.865 124.855 101.990 125.025 ;
        RECT 99.720 124.340 100.470 124.530 ;
        RECT 100.640 124.515 101.650 124.685 ;
        RECT 97.450 123.615 98.840 123.805 ;
        RECT 99.210 123.795 100.440 123.965 ;
        RECT 96.910 123.155 97.470 123.445 ;
        RECT 97.640 122.985 97.890 123.445 ;
        RECT 98.510 123.255 98.840 123.615 ;
        RECT 99.485 123.190 99.730 123.795 ;
        RECT 99.950 122.985 100.460 123.520 ;
        RECT 100.640 123.155 100.830 124.515 ;
        RECT 101.000 123.495 101.275 124.315 ;
        RECT 101.480 123.715 101.650 124.515 ;
        RECT 101.820 123.725 101.990 124.855 ;
        RECT 102.160 124.225 102.330 125.195 ;
        RECT 102.500 124.395 102.670 125.535 ;
        RECT 102.840 124.395 103.175 125.365 ;
        RECT 104.360 124.605 104.530 125.365 ;
        RECT 104.710 124.775 105.040 125.535 ;
        RECT 104.360 124.435 105.025 124.605 ;
        RECT 105.210 124.460 105.480 125.365 ;
        RECT 102.160 123.895 102.355 124.225 ;
        RECT 102.580 123.895 102.835 124.225 ;
        RECT 102.580 123.725 102.750 123.895 ;
        RECT 103.005 123.725 103.175 124.395 ;
        RECT 104.855 124.290 105.025 124.435 ;
        RECT 104.290 123.885 104.620 124.255 ;
        RECT 104.855 123.960 105.140 124.290 ;
        RECT 101.820 123.555 102.750 123.725 ;
        RECT 101.820 123.520 101.995 123.555 ;
        RECT 101.000 123.325 101.280 123.495 ;
        RECT 101.000 123.155 101.275 123.325 ;
        RECT 101.465 123.155 101.995 123.520 ;
        RECT 102.420 122.985 102.750 123.385 ;
        RECT 102.920 123.155 103.175 123.725 ;
        RECT 104.855 123.705 105.025 123.960 ;
        RECT 104.360 123.535 105.025 123.705 ;
        RECT 105.310 123.660 105.480 124.460 ;
        RECT 106.200 124.605 106.370 125.365 ;
        RECT 106.550 124.775 106.880 125.535 ;
        RECT 106.200 124.435 106.865 124.605 ;
        RECT 107.050 124.460 107.320 125.365 ;
        RECT 106.695 124.290 106.865 124.435 ;
        RECT 106.130 123.885 106.460 124.255 ;
        RECT 106.695 123.960 106.980 124.290 ;
        RECT 106.695 123.705 106.865 123.960 ;
        RECT 104.360 123.155 104.530 123.535 ;
        RECT 104.710 122.985 105.040 123.365 ;
        RECT 105.220 123.155 105.480 123.660 ;
        RECT 106.200 123.535 106.865 123.705 ;
        RECT 107.150 123.660 107.320 124.460 ;
        RECT 107.490 124.445 111.000 125.535 ;
        RECT 111.170 124.445 112.380 125.535 ;
        RECT 107.490 123.925 109.180 124.445 ;
        RECT 109.350 123.755 111.000 124.275 ;
        RECT 111.170 123.905 111.690 124.445 ;
        RECT 106.200 123.155 106.370 123.535 ;
        RECT 106.550 122.985 106.880 123.365 ;
        RECT 107.060 123.155 107.320 123.660 ;
        RECT 107.490 122.985 111.000 123.755 ;
        RECT 111.860 123.735 112.380 124.275 ;
        RECT 111.170 122.985 112.380 123.735 ;
        RECT 18.165 122.815 112.465 122.985 ;
        RECT 18.250 122.065 19.460 122.815 ;
        RECT 18.250 121.525 18.770 122.065 ;
        RECT 20.610 121.995 20.820 122.815 ;
        RECT 20.990 122.015 21.320 122.645 ;
        RECT 18.940 121.355 19.460 121.895 ;
        RECT 20.990 121.415 21.240 122.015 ;
        RECT 21.490 121.995 21.720 122.815 ;
        RECT 21.930 122.090 22.220 122.815 ;
        RECT 22.765 122.475 23.020 122.635 ;
        RECT 22.680 122.305 23.020 122.475 ;
        RECT 23.200 122.355 23.485 122.815 ;
        RECT 22.765 122.105 23.020 122.305 ;
        RECT 21.410 121.575 21.740 121.825 ;
        RECT 18.250 120.265 19.460 121.355 ;
        RECT 20.610 120.265 20.820 121.405 ;
        RECT 20.990 120.435 21.320 121.415 ;
        RECT 21.490 120.265 21.720 121.405 ;
        RECT 21.930 120.265 22.220 121.430 ;
        RECT 22.765 121.245 22.945 122.105 ;
        RECT 23.665 121.905 23.915 122.555 ;
        RECT 23.115 121.575 23.915 121.905 ;
        RECT 22.765 120.575 23.020 121.245 ;
        RECT 23.200 120.265 23.485 121.065 ;
        RECT 23.665 120.985 23.915 121.575 ;
        RECT 24.115 122.220 24.435 122.550 ;
        RECT 24.615 122.335 25.275 122.815 ;
        RECT 25.475 122.425 26.325 122.595 ;
        RECT 24.115 121.325 24.305 122.220 ;
        RECT 24.625 121.895 25.285 122.165 ;
        RECT 24.955 121.835 25.285 121.895 ;
        RECT 24.475 121.665 24.805 121.725 ;
        RECT 25.475 121.665 25.645 122.425 ;
        RECT 26.885 122.355 27.205 122.815 ;
        RECT 27.405 122.175 27.655 122.605 ;
        RECT 27.945 122.375 28.355 122.815 ;
        RECT 28.525 122.435 29.540 122.635 ;
        RECT 25.815 122.005 27.065 122.175 ;
        RECT 25.815 121.885 26.145 122.005 ;
        RECT 24.475 121.495 26.375 121.665 ;
        RECT 24.115 121.155 26.035 121.325 ;
        RECT 24.115 121.135 24.435 121.155 ;
        RECT 23.665 120.475 23.995 120.985 ;
        RECT 24.265 120.525 24.435 121.135 ;
        RECT 26.205 120.985 26.375 121.495 ;
        RECT 26.545 121.425 26.725 121.835 ;
        RECT 26.895 121.245 27.065 122.005 ;
        RECT 24.605 120.265 24.935 120.955 ;
        RECT 25.165 120.815 26.375 120.985 ;
        RECT 26.545 120.935 27.065 121.245 ;
        RECT 27.235 121.835 27.655 122.175 ;
        RECT 27.945 121.835 28.355 122.165 ;
        RECT 27.235 121.065 27.425 121.835 ;
        RECT 28.525 121.705 28.695 122.435 ;
        RECT 29.840 122.265 30.010 122.595 ;
        RECT 30.180 122.435 30.510 122.815 ;
        RECT 28.865 121.885 29.215 122.255 ;
        RECT 28.525 121.665 28.945 121.705 ;
        RECT 27.595 121.495 28.945 121.665 ;
        RECT 27.595 121.335 27.845 121.495 ;
        RECT 28.355 121.065 28.605 121.325 ;
        RECT 27.235 120.815 28.605 121.065 ;
        RECT 25.165 120.525 25.405 120.815 ;
        RECT 26.205 120.735 26.375 120.815 ;
        RECT 25.605 120.265 26.025 120.645 ;
        RECT 26.205 120.485 26.835 120.735 ;
        RECT 27.305 120.265 27.635 120.645 ;
        RECT 27.805 120.525 27.975 120.815 ;
        RECT 28.775 120.650 28.945 121.495 ;
        RECT 29.395 121.325 29.615 122.195 ;
        RECT 29.840 122.075 30.535 122.265 ;
        RECT 29.115 120.945 29.615 121.325 ;
        RECT 29.785 121.275 30.195 121.895 ;
        RECT 30.365 121.105 30.535 122.075 ;
        RECT 29.840 120.935 30.535 121.105 ;
        RECT 28.155 120.265 28.535 120.645 ;
        RECT 28.775 120.480 29.605 120.650 ;
        RECT 29.840 120.435 30.010 120.935 ;
        RECT 30.180 120.265 30.510 120.765 ;
        RECT 30.725 120.435 30.950 122.555 ;
        RECT 31.120 122.435 31.450 122.815 ;
        RECT 31.620 122.265 31.790 122.555 ;
        RECT 31.125 122.095 31.790 122.265 ;
        RECT 31.125 121.105 31.355 122.095 ;
        RECT 32.055 122.075 32.310 122.645 ;
        RECT 32.480 122.415 32.810 122.815 ;
        RECT 33.235 122.280 33.765 122.645 ;
        RECT 33.955 122.475 34.230 122.645 ;
        RECT 33.950 122.305 34.230 122.475 ;
        RECT 33.235 122.245 33.410 122.280 ;
        RECT 32.480 122.075 33.410 122.245 ;
        RECT 31.525 121.275 31.875 121.925 ;
        RECT 32.055 121.405 32.225 122.075 ;
        RECT 32.480 121.905 32.650 122.075 ;
        RECT 32.395 121.575 32.650 121.905 ;
        RECT 32.875 121.575 33.070 121.905 ;
        RECT 31.125 120.935 31.790 121.105 ;
        RECT 31.120 120.265 31.450 120.765 ;
        RECT 31.620 120.435 31.790 120.935 ;
        RECT 32.055 120.435 32.390 121.405 ;
        RECT 32.560 120.265 32.730 121.405 ;
        RECT 32.900 120.605 33.070 121.575 ;
        RECT 33.240 120.945 33.410 122.075 ;
        RECT 33.580 121.285 33.750 122.085 ;
        RECT 33.955 121.485 34.230 122.305 ;
        RECT 34.400 121.285 34.590 122.645 ;
        RECT 34.770 122.280 35.280 122.815 ;
        RECT 35.500 122.005 35.745 122.610 ;
        RECT 36.190 122.140 36.450 122.645 ;
        RECT 36.630 122.435 36.960 122.815 ;
        RECT 37.140 122.265 37.310 122.645 ;
        RECT 34.790 121.835 36.020 122.005 ;
        RECT 33.580 121.115 34.590 121.285 ;
        RECT 34.760 121.270 35.510 121.460 ;
        RECT 33.240 120.775 34.365 120.945 ;
        RECT 34.760 120.605 34.930 121.270 ;
        RECT 35.680 121.025 36.020 121.835 ;
        RECT 32.900 120.435 34.930 120.605 ;
        RECT 35.100 120.265 35.270 121.025 ;
        RECT 35.505 120.615 36.020 121.025 ;
        RECT 36.190 121.340 36.360 122.140 ;
        RECT 36.645 122.095 37.310 122.265 ;
        RECT 36.645 121.840 36.815 122.095 ;
        RECT 38.530 121.995 38.760 122.815 ;
        RECT 38.930 122.015 39.260 122.645 ;
        RECT 36.530 121.510 36.815 121.840 ;
        RECT 37.050 121.545 37.380 121.915 ;
        RECT 38.510 121.575 38.840 121.825 ;
        RECT 36.645 121.365 36.815 121.510 ;
        RECT 39.010 121.415 39.260 122.015 ;
        RECT 39.430 121.995 39.640 122.815 ;
        RECT 39.870 122.310 40.155 122.815 ;
        RECT 40.325 122.140 40.650 122.645 ;
        RECT 39.870 121.610 40.650 122.140 ;
        RECT 36.190 120.435 36.460 121.340 ;
        RECT 36.645 121.195 37.310 121.365 ;
        RECT 36.630 120.265 36.960 121.025 ;
        RECT 37.140 120.435 37.310 121.195 ;
        RECT 38.530 120.265 38.760 121.405 ;
        RECT 38.930 120.435 39.260 121.415 ;
        RECT 39.430 120.265 39.640 121.405 ;
        RECT 39.870 120.265 40.150 121.235 ;
        RECT 40.320 120.435 40.650 121.610 ;
        RECT 40.840 121.575 41.080 122.525 ;
        RECT 41.450 122.185 41.780 122.545 ;
        RECT 42.400 122.355 42.650 122.815 ;
        RECT 42.820 122.355 43.380 122.645 ;
        RECT 41.450 121.995 42.840 122.185 ;
        RECT 42.670 121.905 42.840 121.995 ;
        RECT 41.265 121.575 41.940 121.825 ;
        RECT 42.160 121.575 42.500 121.825 ;
        RECT 42.670 121.575 42.960 121.905 ;
        RECT 40.820 120.265 41.080 121.235 ;
        RECT 41.265 121.215 41.530 121.575 ;
        RECT 42.670 121.325 42.840 121.575 ;
        RECT 41.900 121.155 42.840 121.325 ;
        RECT 41.450 120.265 41.730 120.935 ;
        RECT 41.900 120.605 42.200 121.155 ;
        RECT 43.130 120.985 43.380 122.355 ;
        RECT 42.400 120.265 42.730 120.985 ;
        RECT 42.920 120.435 43.380 120.985 ;
        RECT 43.555 122.075 43.810 122.645 ;
        RECT 43.980 122.415 44.310 122.815 ;
        RECT 44.735 122.280 45.265 122.645 ;
        RECT 44.735 122.245 44.910 122.280 ;
        RECT 43.980 122.075 44.910 122.245 ;
        RECT 43.555 121.405 43.725 122.075 ;
        RECT 43.980 121.905 44.150 122.075 ;
        RECT 43.895 121.575 44.150 121.905 ;
        RECT 44.375 121.575 44.570 121.905 ;
        RECT 43.555 120.435 43.890 121.405 ;
        RECT 44.060 120.265 44.230 121.405 ;
        RECT 44.400 120.605 44.570 121.575 ;
        RECT 44.740 120.945 44.910 122.075 ;
        RECT 45.080 121.285 45.250 122.085 ;
        RECT 45.455 121.795 45.730 122.645 ;
        RECT 45.450 121.625 45.730 121.795 ;
        RECT 45.455 121.485 45.730 121.625 ;
        RECT 45.900 121.285 46.090 122.645 ;
        RECT 46.270 122.280 46.780 122.815 ;
        RECT 47.000 122.005 47.245 122.610 ;
        RECT 47.690 122.090 47.980 122.815 ;
        RECT 46.290 121.835 47.520 122.005 ;
        RECT 49.110 121.995 49.340 122.815 ;
        RECT 49.510 122.015 49.840 122.645 ;
        RECT 45.080 121.115 46.090 121.285 ;
        RECT 46.260 121.270 47.010 121.460 ;
        RECT 44.740 120.775 45.865 120.945 ;
        RECT 46.260 120.605 46.430 121.270 ;
        RECT 47.180 121.025 47.520 121.835 ;
        RECT 49.090 121.575 49.420 121.825 ;
        RECT 44.400 120.435 46.430 120.605 ;
        RECT 46.600 120.265 46.770 121.025 ;
        RECT 47.005 120.615 47.520 121.025 ;
        RECT 47.690 120.265 47.980 121.430 ;
        RECT 49.590 121.415 49.840 122.015 ;
        RECT 50.010 121.995 50.220 122.815 ;
        RECT 50.650 122.185 50.980 122.545 ;
        RECT 51.600 122.355 51.850 122.815 ;
        RECT 52.020 122.355 52.580 122.645 ;
        RECT 50.650 121.995 52.040 122.185 ;
        RECT 51.870 121.905 52.040 121.995 ;
        RECT 49.110 120.265 49.340 121.405 ;
        RECT 49.510 120.435 49.840 121.415 ;
        RECT 50.465 121.575 51.140 121.825 ;
        RECT 51.360 121.575 51.700 121.825 ;
        RECT 51.870 121.575 52.160 121.905 ;
        RECT 50.010 120.265 50.220 121.405 ;
        RECT 50.465 121.215 50.730 121.575 ;
        RECT 51.870 121.325 52.040 121.575 ;
        RECT 51.100 121.155 52.040 121.325 ;
        RECT 50.650 120.265 50.930 120.935 ;
        RECT 51.100 120.605 51.400 121.155 ;
        RECT 52.330 120.985 52.580 122.355 ;
        RECT 53.025 122.005 53.270 122.610 ;
        RECT 53.490 122.280 54.000 122.815 ;
        RECT 51.600 120.265 51.930 120.985 ;
        RECT 52.120 120.435 52.580 120.985 ;
        RECT 52.750 121.835 53.980 122.005 ;
        RECT 52.750 121.025 53.090 121.835 ;
        RECT 53.260 121.270 54.010 121.460 ;
        RECT 52.750 120.615 53.265 121.025 ;
        RECT 53.500 120.265 53.670 121.025 ;
        RECT 53.840 120.605 54.010 121.270 ;
        RECT 54.180 121.285 54.370 122.645 ;
        RECT 54.540 122.135 54.815 122.645 ;
        RECT 55.005 122.280 55.535 122.645 ;
        RECT 55.960 122.415 56.290 122.815 ;
        RECT 55.360 122.245 55.535 122.280 ;
        RECT 54.540 121.965 54.820 122.135 ;
        RECT 54.540 121.485 54.815 121.965 ;
        RECT 55.020 121.285 55.190 122.085 ;
        RECT 54.180 121.115 55.190 121.285 ;
        RECT 55.360 122.075 56.290 122.245 ;
        RECT 56.460 122.075 56.715 122.645 ;
        RECT 55.360 120.945 55.530 122.075 ;
        RECT 56.120 121.905 56.290 122.075 ;
        RECT 54.405 120.775 55.530 120.945 ;
        RECT 55.700 121.575 55.895 121.905 ;
        RECT 56.120 121.575 56.375 121.905 ;
        RECT 55.700 120.605 55.870 121.575 ;
        RECT 56.545 121.405 56.715 122.075 ;
        RECT 57.040 122.015 57.370 122.815 ;
        RECT 57.540 122.165 57.710 122.645 ;
        RECT 57.880 122.335 58.210 122.815 ;
        RECT 58.380 122.165 58.550 122.645 ;
        RECT 58.800 122.335 59.040 122.815 ;
        RECT 59.220 122.165 59.390 122.645 ;
        RECT 57.540 121.995 58.550 122.165 ;
        RECT 58.755 121.995 59.390 122.165 ;
        RECT 60.110 122.045 63.620 122.815 ;
        RECT 63.880 122.265 64.050 122.555 ;
        RECT 64.220 122.435 64.550 122.815 ;
        RECT 63.880 122.095 64.545 122.265 ;
        RECT 57.540 121.965 58.040 121.995 ;
        RECT 57.540 121.455 58.035 121.965 ;
        RECT 58.755 121.825 58.925 121.995 ;
        RECT 58.425 121.655 58.925 121.825 ;
        RECT 53.840 120.435 55.870 120.605 ;
        RECT 56.040 120.265 56.210 121.405 ;
        RECT 56.380 120.435 56.715 121.405 ;
        RECT 57.040 120.265 57.370 121.415 ;
        RECT 57.540 121.285 58.550 121.455 ;
        RECT 57.540 120.435 57.710 121.285 ;
        RECT 57.880 120.265 58.210 121.065 ;
        RECT 58.380 120.435 58.550 121.285 ;
        RECT 58.755 121.415 58.925 121.655 ;
        RECT 59.095 121.585 59.475 121.825 ;
        RECT 58.755 121.245 59.470 121.415 ;
        RECT 58.730 120.265 58.970 121.065 ;
        RECT 59.140 120.435 59.470 121.245 ;
        RECT 60.110 121.355 61.800 121.875 ;
        RECT 61.970 121.525 63.620 122.045 ;
        RECT 60.110 120.265 63.620 121.355 ;
        RECT 63.795 121.275 64.145 121.925 ;
        RECT 64.315 121.105 64.545 122.095 ;
        RECT 63.880 120.935 64.545 121.105 ;
        RECT 63.880 120.435 64.050 120.935 ;
        RECT 64.220 120.265 64.550 120.765 ;
        RECT 64.720 120.435 64.945 122.555 ;
        RECT 65.160 122.435 65.490 122.815 ;
        RECT 65.660 122.265 65.830 122.595 ;
        RECT 66.130 122.435 67.145 122.635 ;
        RECT 65.135 122.075 65.830 122.265 ;
        RECT 65.135 121.105 65.305 122.075 ;
        RECT 65.475 121.275 65.885 121.895 ;
        RECT 66.055 121.325 66.275 122.195 ;
        RECT 66.455 121.885 66.805 122.255 ;
        RECT 66.975 121.705 67.145 122.435 ;
        RECT 67.315 122.375 67.725 122.815 ;
        RECT 68.015 122.175 68.265 122.605 ;
        RECT 68.465 122.355 68.785 122.815 ;
        RECT 69.345 122.425 70.195 122.595 ;
        RECT 67.315 121.835 67.725 122.165 ;
        RECT 68.015 121.835 68.435 122.175 ;
        RECT 66.725 121.665 67.145 121.705 ;
        RECT 66.725 121.495 68.075 121.665 ;
        RECT 65.135 120.935 65.830 121.105 ;
        RECT 66.055 120.945 66.555 121.325 ;
        RECT 65.160 120.265 65.490 120.765 ;
        RECT 65.660 120.435 65.830 120.935 ;
        RECT 66.725 120.650 66.895 121.495 ;
        RECT 67.825 121.335 68.075 121.495 ;
        RECT 67.065 121.065 67.315 121.325 ;
        RECT 68.245 121.065 68.435 121.835 ;
        RECT 67.065 120.815 68.435 121.065 ;
        RECT 68.605 122.005 69.855 122.175 ;
        RECT 68.605 121.245 68.775 122.005 ;
        RECT 69.525 121.885 69.855 122.005 ;
        RECT 68.945 121.425 69.125 121.835 ;
        RECT 70.025 121.665 70.195 122.425 ;
        RECT 70.395 122.335 71.055 122.815 ;
        RECT 71.235 122.220 71.555 122.550 ;
        RECT 70.385 121.895 71.045 122.165 ;
        RECT 70.385 121.835 70.715 121.895 ;
        RECT 70.865 121.665 71.195 121.725 ;
        RECT 69.295 121.495 71.195 121.665 ;
        RECT 68.605 120.935 69.125 121.245 ;
        RECT 69.295 120.985 69.465 121.495 ;
        RECT 71.365 121.325 71.555 122.220 ;
        RECT 69.635 121.155 71.555 121.325 ;
        RECT 71.235 121.135 71.555 121.155 ;
        RECT 71.755 121.905 72.005 122.555 ;
        RECT 72.185 122.355 72.470 122.815 ;
        RECT 72.650 122.105 72.905 122.635 ;
        RECT 71.755 121.575 72.555 121.905 ;
        RECT 69.295 120.815 70.505 120.985 ;
        RECT 66.065 120.480 66.895 120.650 ;
        RECT 67.135 120.265 67.515 120.645 ;
        RECT 67.695 120.525 67.865 120.815 ;
        RECT 69.295 120.735 69.465 120.815 ;
        RECT 68.035 120.265 68.365 120.645 ;
        RECT 68.835 120.485 69.465 120.735 ;
        RECT 69.645 120.265 70.065 120.645 ;
        RECT 70.265 120.525 70.505 120.815 ;
        RECT 70.735 120.265 71.065 120.955 ;
        RECT 71.235 120.525 71.405 121.135 ;
        RECT 71.755 120.985 72.005 121.575 ;
        RECT 72.725 121.245 72.905 122.105 ;
        RECT 73.450 122.090 73.740 122.815 ;
        RECT 74.370 122.140 74.630 122.645 ;
        RECT 74.810 122.435 75.140 122.815 ;
        RECT 75.320 122.265 75.490 122.645 ;
        RECT 71.675 120.475 72.005 120.985 ;
        RECT 72.185 120.265 72.470 121.065 ;
        RECT 72.650 120.775 72.905 121.245 ;
        RECT 72.650 120.605 72.990 120.775 ;
        RECT 72.650 120.575 72.905 120.605 ;
        RECT 73.450 120.265 73.740 121.430 ;
        RECT 74.370 121.340 74.540 122.140 ;
        RECT 74.825 122.095 75.490 122.265 ;
        RECT 74.825 121.840 74.995 122.095 ;
        RECT 76.210 122.045 78.800 122.815 ;
        RECT 79.060 122.265 79.230 122.645 ;
        RECT 79.410 122.435 79.740 122.815 ;
        RECT 79.060 122.095 79.725 122.265 ;
        RECT 79.920 122.140 80.180 122.645 ;
        RECT 74.710 121.510 74.995 121.840 ;
        RECT 75.230 121.545 75.560 121.915 ;
        RECT 74.825 121.365 74.995 121.510 ;
        RECT 74.370 120.435 74.640 121.340 ;
        RECT 74.825 121.195 75.490 121.365 ;
        RECT 74.810 120.265 75.140 121.025 ;
        RECT 75.320 120.435 75.490 121.195 ;
        RECT 76.210 121.355 77.420 121.875 ;
        RECT 77.590 121.525 78.800 122.045 ;
        RECT 78.990 121.545 79.320 121.915 ;
        RECT 79.555 121.840 79.725 122.095 ;
        RECT 79.555 121.510 79.840 121.840 ;
        RECT 79.555 121.365 79.725 121.510 ;
        RECT 76.210 120.265 78.800 121.355 ;
        RECT 79.060 121.195 79.725 121.365 ;
        RECT 80.010 121.340 80.180 122.140 ;
        RECT 80.810 122.045 83.400 122.815 ;
        RECT 79.060 120.435 79.230 121.195 ;
        RECT 79.410 120.265 79.740 121.025 ;
        RECT 79.910 120.435 80.180 121.340 ;
        RECT 80.810 121.355 82.020 121.875 ;
        RECT 82.190 121.525 83.400 122.045 ;
        RECT 83.845 122.005 84.090 122.610 ;
        RECT 84.310 122.280 84.820 122.815 ;
        RECT 83.570 121.835 84.800 122.005 ;
        RECT 80.810 120.265 83.400 121.355 ;
        RECT 83.570 121.025 83.910 121.835 ;
        RECT 84.080 121.270 84.830 121.460 ;
        RECT 83.570 120.615 84.085 121.025 ;
        RECT 84.320 120.265 84.490 121.025 ;
        RECT 84.660 120.605 84.830 121.270 ;
        RECT 85.000 121.285 85.190 122.645 ;
        RECT 85.360 122.475 85.635 122.645 ;
        RECT 85.360 122.305 85.640 122.475 ;
        RECT 85.360 121.485 85.635 122.305 ;
        RECT 85.825 122.280 86.355 122.645 ;
        RECT 86.780 122.415 87.110 122.815 ;
        RECT 86.180 122.245 86.355 122.280 ;
        RECT 85.840 121.285 86.010 122.085 ;
        RECT 85.000 121.115 86.010 121.285 ;
        RECT 86.180 122.075 87.110 122.245 ;
        RECT 87.280 122.075 87.535 122.645 ;
        RECT 86.180 120.945 86.350 122.075 ;
        RECT 86.940 121.905 87.110 122.075 ;
        RECT 85.225 120.775 86.350 120.945 ;
        RECT 86.520 121.575 86.715 121.905 ;
        RECT 86.940 121.575 87.195 121.905 ;
        RECT 86.520 120.605 86.690 121.575 ;
        RECT 87.365 121.405 87.535 122.075 ;
        RECT 84.660 120.435 86.690 120.605 ;
        RECT 86.860 120.265 87.030 121.405 ;
        RECT 87.200 120.435 87.535 121.405 ;
        RECT 87.715 122.075 87.970 122.645 ;
        RECT 88.140 122.415 88.470 122.815 ;
        RECT 88.895 122.280 89.425 122.645 ;
        RECT 88.895 122.245 89.070 122.280 ;
        RECT 88.140 122.075 89.070 122.245 ;
        RECT 87.715 121.405 87.885 122.075 ;
        RECT 88.140 121.905 88.310 122.075 ;
        RECT 88.055 121.575 88.310 121.905 ;
        RECT 88.535 121.575 88.730 121.905 ;
        RECT 87.715 120.435 88.050 121.405 ;
        RECT 88.220 120.265 88.390 121.405 ;
        RECT 88.560 120.605 88.730 121.575 ;
        RECT 88.900 120.945 89.070 122.075 ;
        RECT 89.240 121.285 89.410 122.085 ;
        RECT 89.615 121.795 89.890 122.645 ;
        RECT 89.610 121.625 89.890 121.795 ;
        RECT 89.615 121.485 89.890 121.625 ;
        RECT 90.060 121.285 90.250 122.645 ;
        RECT 90.430 122.280 90.940 122.815 ;
        RECT 91.160 122.005 91.405 122.610 ;
        RECT 92.050 122.185 92.380 122.545 ;
        RECT 93.000 122.355 93.250 122.815 ;
        RECT 93.420 122.355 93.980 122.645 ;
        RECT 90.450 121.835 91.680 122.005 ;
        RECT 92.050 121.995 93.440 122.185 ;
        RECT 89.240 121.115 90.250 121.285 ;
        RECT 90.420 121.270 91.170 121.460 ;
        RECT 88.900 120.775 90.025 120.945 ;
        RECT 90.420 120.605 90.590 121.270 ;
        RECT 91.340 121.025 91.680 121.835 ;
        RECT 93.270 121.905 93.440 121.995 ;
        RECT 91.865 121.575 92.540 121.825 ;
        RECT 92.760 121.575 93.100 121.825 ;
        RECT 93.270 121.575 93.560 121.905 ;
        RECT 91.865 121.215 92.130 121.575 ;
        RECT 93.270 121.325 93.440 121.575 ;
        RECT 88.560 120.435 90.590 120.605 ;
        RECT 90.760 120.265 90.930 121.025 ;
        RECT 91.165 120.615 91.680 121.025 ;
        RECT 92.500 121.155 93.440 121.325 ;
        RECT 92.050 120.265 92.330 120.935 ;
        RECT 92.500 120.605 92.800 121.155 ;
        RECT 93.730 120.985 93.980 122.355 ;
        RECT 94.425 122.005 94.670 122.610 ;
        RECT 94.890 122.280 95.400 122.815 ;
        RECT 93.000 120.265 93.330 120.985 ;
        RECT 93.520 120.435 93.980 120.985 ;
        RECT 94.150 121.835 95.380 122.005 ;
        RECT 94.150 121.025 94.490 121.835 ;
        RECT 94.660 121.270 95.410 121.460 ;
        RECT 94.150 120.615 94.665 121.025 ;
        RECT 94.900 120.265 95.070 121.025 ;
        RECT 95.240 120.605 95.410 121.270 ;
        RECT 95.580 121.285 95.770 122.645 ;
        RECT 95.940 122.135 96.215 122.645 ;
        RECT 96.405 122.280 96.935 122.645 ;
        RECT 97.360 122.415 97.690 122.815 ;
        RECT 96.760 122.245 96.935 122.280 ;
        RECT 95.940 121.965 96.220 122.135 ;
        RECT 95.940 121.485 96.215 121.965 ;
        RECT 96.420 121.285 96.590 122.085 ;
        RECT 95.580 121.115 96.590 121.285 ;
        RECT 96.760 122.075 97.690 122.245 ;
        RECT 97.860 122.075 98.115 122.645 ;
        RECT 99.210 122.090 99.500 122.815 ;
        RECT 96.760 120.945 96.930 122.075 ;
        RECT 97.520 121.905 97.690 122.075 ;
        RECT 95.805 120.775 96.930 120.945 ;
        RECT 97.100 121.575 97.295 121.905 ;
        RECT 97.520 121.575 97.775 121.905 ;
        RECT 97.100 120.605 97.270 121.575 ;
        RECT 97.945 121.405 98.115 122.075 ;
        RECT 100.865 122.005 101.110 122.610 ;
        RECT 101.330 122.280 101.840 122.815 ;
        RECT 100.590 121.835 101.820 122.005 ;
        RECT 95.240 120.435 97.270 120.605 ;
        RECT 97.440 120.265 97.610 121.405 ;
        RECT 97.780 120.435 98.115 121.405 ;
        RECT 99.210 120.265 99.500 121.430 ;
        RECT 100.590 121.025 100.930 121.835 ;
        RECT 101.100 121.270 101.850 121.460 ;
        RECT 100.590 120.615 101.105 121.025 ;
        RECT 101.340 120.265 101.510 121.025 ;
        RECT 101.680 120.605 101.850 121.270 ;
        RECT 102.020 121.285 102.210 122.645 ;
        RECT 102.380 121.795 102.655 122.645 ;
        RECT 102.845 122.280 103.375 122.645 ;
        RECT 103.800 122.415 104.130 122.815 ;
        RECT 103.200 122.245 103.375 122.280 ;
        RECT 102.380 121.625 102.660 121.795 ;
        RECT 102.380 121.485 102.655 121.625 ;
        RECT 102.860 121.285 103.030 122.085 ;
        RECT 102.020 121.115 103.030 121.285 ;
        RECT 103.200 122.075 104.130 122.245 ;
        RECT 104.300 122.075 104.555 122.645 ;
        RECT 103.200 120.945 103.370 122.075 ;
        RECT 103.960 121.905 104.130 122.075 ;
        RECT 102.245 120.775 103.370 120.945 ;
        RECT 103.540 121.575 103.735 121.905 ;
        RECT 103.960 121.575 104.215 121.905 ;
        RECT 103.540 120.605 103.710 121.575 ;
        RECT 104.385 121.405 104.555 122.075 ;
        RECT 104.770 121.995 105.000 122.815 ;
        RECT 105.170 122.015 105.500 122.645 ;
        RECT 104.750 121.575 105.080 121.825 ;
        RECT 105.250 121.415 105.500 122.015 ;
        RECT 105.670 121.995 105.880 122.815 ;
        RECT 106.660 122.265 106.830 122.645 ;
        RECT 107.010 122.435 107.340 122.815 ;
        RECT 106.660 122.095 107.325 122.265 ;
        RECT 107.520 122.140 107.780 122.645 ;
        RECT 106.590 121.545 106.920 121.915 ;
        RECT 107.155 121.840 107.325 122.095 ;
        RECT 101.680 120.435 103.710 120.605 ;
        RECT 103.880 120.265 104.050 121.405 ;
        RECT 104.220 120.435 104.555 121.405 ;
        RECT 104.770 120.265 105.000 121.405 ;
        RECT 105.170 120.435 105.500 121.415 ;
        RECT 107.155 121.510 107.440 121.840 ;
        RECT 105.670 120.265 105.880 121.405 ;
        RECT 107.155 121.365 107.325 121.510 ;
        RECT 106.660 121.195 107.325 121.365 ;
        RECT 107.610 121.340 107.780 122.140 ;
        RECT 108.410 122.045 111.000 122.815 ;
        RECT 111.170 122.065 112.380 122.815 ;
        RECT 106.660 120.435 106.830 121.195 ;
        RECT 107.010 120.265 107.340 121.025 ;
        RECT 107.510 120.435 107.780 121.340 ;
        RECT 108.410 121.355 109.620 121.875 ;
        RECT 109.790 121.525 111.000 122.045 ;
        RECT 111.170 121.355 111.690 121.895 ;
        RECT 111.860 121.525 112.380 122.065 ;
        RECT 108.410 120.265 111.000 121.355 ;
        RECT 111.170 120.265 112.380 121.355 ;
        RECT 18.165 120.095 112.465 120.265 ;
        RECT 18.250 119.005 19.460 120.095 ;
        RECT 18.250 118.295 18.770 118.835 ;
        RECT 18.940 118.465 19.460 119.005 ;
        RECT 19.630 119.005 20.840 120.095 ;
        RECT 21.010 119.335 21.525 119.745 ;
        RECT 21.760 119.335 21.930 120.095 ;
        RECT 22.100 119.755 24.130 119.925 ;
        RECT 19.630 118.465 20.150 119.005 ;
        RECT 20.320 118.295 20.840 118.835 ;
        RECT 21.010 118.525 21.350 119.335 ;
        RECT 22.100 119.090 22.270 119.755 ;
        RECT 22.665 119.415 23.790 119.585 ;
        RECT 21.520 118.900 22.270 119.090 ;
        RECT 22.440 119.075 23.450 119.245 ;
        RECT 21.010 118.355 22.240 118.525 ;
        RECT 18.250 117.545 19.460 118.295 ;
        RECT 19.630 117.545 20.840 118.295 ;
        RECT 21.285 117.750 21.530 118.355 ;
        RECT 21.750 117.545 22.260 118.080 ;
        RECT 22.440 117.715 22.630 119.075 ;
        RECT 22.800 118.735 23.075 118.875 ;
        RECT 22.800 118.565 23.080 118.735 ;
        RECT 22.800 117.715 23.075 118.565 ;
        RECT 23.280 118.275 23.450 119.075 ;
        RECT 23.620 118.285 23.790 119.415 ;
        RECT 23.960 118.785 24.130 119.755 ;
        RECT 24.300 118.955 24.470 120.095 ;
        RECT 24.640 118.955 24.975 119.925 ;
        RECT 25.525 119.115 25.780 119.785 ;
        RECT 25.960 119.295 26.245 120.095 ;
        RECT 26.425 119.375 26.755 119.885 ;
        RECT 25.525 119.075 25.705 119.115 ;
        RECT 23.960 118.455 24.155 118.785 ;
        RECT 24.380 118.455 24.635 118.785 ;
        RECT 24.380 118.285 24.550 118.455 ;
        RECT 24.805 118.285 24.975 118.955 ;
        RECT 25.440 118.905 25.705 119.075 ;
        RECT 23.620 118.115 24.550 118.285 ;
        RECT 23.620 118.080 23.795 118.115 ;
        RECT 23.265 117.715 23.795 118.080 ;
        RECT 24.220 117.545 24.550 117.945 ;
        RECT 24.720 117.715 24.975 118.285 ;
        RECT 25.525 118.255 25.705 118.905 ;
        RECT 26.425 118.785 26.675 119.375 ;
        RECT 27.025 119.225 27.195 119.835 ;
        RECT 27.365 119.405 27.695 120.095 ;
        RECT 27.925 119.545 28.165 119.835 ;
        RECT 28.365 119.715 28.785 120.095 ;
        RECT 28.965 119.625 29.595 119.875 ;
        RECT 30.065 119.715 30.395 120.095 ;
        RECT 28.965 119.545 29.135 119.625 ;
        RECT 30.565 119.545 30.735 119.835 ;
        RECT 30.915 119.715 31.295 120.095 ;
        RECT 31.535 119.710 32.365 119.880 ;
        RECT 27.925 119.375 29.135 119.545 ;
        RECT 25.875 118.455 26.675 118.785 ;
        RECT 25.525 117.725 25.780 118.255 ;
        RECT 25.960 117.545 26.245 118.005 ;
        RECT 26.425 117.805 26.675 118.455 ;
        RECT 26.875 119.205 27.195 119.225 ;
        RECT 26.875 119.035 28.795 119.205 ;
        RECT 26.875 118.140 27.065 119.035 ;
        RECT 28.965 118.865 29.135 119.375 ;
        RECT 29.305 119.115 29.825 119.425 ;
        RECT 27.235 118.695 29.135 118.865 ;
        RECT 27.235 118.635 27.565 118.695 ;
        RECT 27.715 118.465 28.045 118.525 ;
        RECT 27.385 118.195 28.045 118.465 ;
        RECT 26.875 117.810 27.195 118.140 ;
        RECT 27.375 117.545 28.035 118.025 ;
        RECT 28.235 117.935 28.405 118.695 ;
        RECT 29.305 118.525 29.485 118.935 ;
        RECT 28.575 118.355 28.905 118.475 ;
        RECT 29.655 118.355 29.825 119.115 ;
        RECT 28.575 118.185 29.825 118.355 ;
        RECT 29.995 119.295 31.365 119.545 ;
        RECT 29.995 118.525 30.185 119.295 ;
        RECT 31.115 119.035 31.365 119.295 ;
        RECT 30.355 118.865 30.605 119.025 ;
        RECT 31.535 118.865 31.705 119.710 ;
        RECT 32.600 119.425 32.770 119.925 ;
        RECT 32.940 119.595 33.270 120.095 ;
        RECT 31.875 119.035 32.375 119.415 ;
        RECT 32.600 119.255 33.295 119.425 ;
        RECT 30.355 118.695 31.705 118.865 ;
        RECT 31.285 118.655 31.705 118.695 ;
        RECT 29.995 118.185 30.415 118.525 ;
        RECT 30.705 118.195 31.115 118.525 ;
        RECT 28.235 117.765 29.085 117.935 ;
        RECT 29.645 117.545 29.965 118.005 ;
        RECT 30.165 117.755 30.415 118.185 ;
        RECT 30.705 117.545 31.115 117.985 ;
        RECT 31.285 117.925 31.455 118.655 ;
        RECT 31.625 118.105 31.975 118.475 ;
        RECT 32.155 118.165 32.375 119.035 ;
        RECT 32.545 118.465 32.955 119.085 ;
        RECT 33.125 118.285 33.295 119.255 ;
        RECT 32.600 118.095 33.295 118.285 ;
        RECT 31.285 117.725 32.300 117.925 ;
        RECT 32.600 117.765 32.770 118.095 ;
        RECT 32.940 117.545 33.270 117.925 ;
        RECT 33.485 117.805 33.710 119.925 ;
        RECT 33.880 119.595 34.210 120.095 ;
        RECT 34.380 119.425 34.550 119.925 ;
        RECT 33.885 119.255 34.550 119.425 ;
        RECT 33.885 118.265 34.115 119.255 ;
        RECT 34.285 118.435 34.635 119.085 ;
        RECT 34.810 118.930 35.100 120.095 ;
        RECT 35.790 118.955 36.000 120.095 ;
        RECT 36.170 118.945 36.500 119.925 ;
        RECT 36.670 118.955 36.900 120.095 ;
        RECT 37.115 118.955 37.450 119.925 ;
        RECT 37.620 118.955 37.790 120.095 ;
        RECT 37.960 119.755 39.990 119.925 ;
        RECT 33.885 118.095 34.550 118.265 ;
        RECT 33.880 117.545 34.210 117.925 ;
        RECT 34.380 117.805 34.550 118.095 ;
        RECT 34.810 117.545 35.100 118.270 ;
        RECT 35.790 117.545 36.000 118.365 ;
        RECT 36.170 118.345 36.420 118.945 ;
        RECT 36.590 118.535 36.920 118.785 ;
        RECT 36.170 117.715 36.500 118.345 ;
        RECT 36.670 117.545 36.900 118.365 ;
        RECT 37.115 118.285 37.285 118.955 ;
        RECT 37.960 118.785 38.130 119.755 ;
        RECT 37.455 118.455 37.710 118.785 ;
        RECT 37.935 118.455 38.130 118.785 ;
        RECT 38.300 119.415 39.425 119.585 ;
        RECT 37.540 118.285 37.710 118.455 ;
        RECT 38.300 118.285 38.470 119.415 ;
        RECT 37.115 117.715 37.370 118.285 ;
        RECT 37.540 118.115 38.470 118.285 ;
        RECT 38.640 119.075 39.650 119.245 ;
        RECT 38.640 118.275 38.810 119.075 ;
        RECT 38.295 118.080 38.470 118.115 ;
        RECT 37.540 117.545 37.870 117.945 ;
        RECT 38.295 117.715 38.825 118.080 ;
        RECT 39.015 118.055 39.290 118.875 ;
        RECT 39.010 117.885 39.290 118.055 ;
        RECT 39.015 117.715 39.290 117.885 ;
        RECT 39.460 117.715 39.650 119.075 ;
        RECT 39.820 119.090 39.990 119.755 ;
        RECT 40.160 119.335 40.330 120.095 ;
        RECT 40.565 119.335 41.080 119.745 ;
        RECT 39.820 118.900 40.570 119.090 ;
        RECT 40.740 118.525 41.080 119.335 ;
        RECT 41.625 119.115 41.880 119.785 ;
        RECT 42.060 119.295 42.345 120.095 ;
        RECT 42.525 119.375 42.855 119.885 ;
        RECT 41.625 118.735 41.805 119.115 ;
        RECT 42.525 118.785 42.775 119.375 ;
        RECT 43.125 119.225 43.295 119.835 ;
        RECT 43.465 119.405 43.795 120.095 ;
        RECT 44.025 119.545 44.265 119.835 ;
        RECT 44.465 119.715 44.885 120.095 ;
        RECT 45.065 119.625 45.695 119.875 ;
        RECT 46.165 119.715 46.495 120.095 ;
        RECT 45.065 119.545 45.235 119.625 ;
        RECT 46.665 119.545 46.835 119.835 ;
        RECT 47.015 119.715 47.395 120.095 ;
        RECT 47.635 119.710 48.465 119.880 ;
        RECT 44.025 119.375 45.235 119.545 ;
        RECT 41.540 118.565 41.805 118.735 ;
        RECT 39.850 118.355 41.080 118.525 ;
        RECT 39.830 117.545 40.340 118.080 ;
        RECT 40.560 117.750 40.805 118.355 ;
        RECT 41.625 118.255 41.805 118.565 ;
        RECT 41.975 118.455 42.775 118.785 ;
        RECT 41.625 117.725 41.880 118.255 ;
        RECT 42.060 117.545 42.345 118.005 ;
        RECT 42.525 117.805 42.775 118.455 ;
        RECT 42.975 119.205 43.295 119.225 ;
        RECT 42.975 119.035 44.895 119.205 ;
        RECT 42.975 118.140 43.165 119.035 ;
        RECT 45.065 118.865 45.235 119.375 ;
        RECT 45.405 119.115 45.925 119.425 ;
        RECT 43.335 118.695 45.235 118.865 ;
        RECT 43.335 118.635 43.665 118.695 ;
        RECT 43.815 118.465 44.145 118.525 ;
        RECT 43.485 118.195 44.145 118.465 ;
        RECT 42.975 117.810 43.295 118.140 ;
        RECT 43.475 117.545 44.135 118.025 ;
        RECT 44.335 117.935 44.505 118.695 ;
        RECT 45.405 118.525 45.585 118.935 ;
        RECT 44.675 118.355 45.005 118.475 ;
        RECT 45.755 118.355 45.925 119.115 ;
        RECT 44.675 118.185 45.925 118.355 ;
        RECT 46.095 119.295 47.465 119.545 ;
        RECT 46.095 118.525 46.285 119.295 ;
        RECT 47.215 119.035 47.465 119.295 ;
        RECT 46.455 118.865 46.705 119.025 ;
        RECT 47.635 118.865 47.805 119.710 ;
        RECT 48.700 119.425 48.870 119.925 ;
        RECT 49.040 119.595 49.370 120.095 ;
        RECT 47.975 119.035 48.475 119.415 ;
        RECT 48.700 119.255 49.395 119.425 ;
        RECT 46.455 118.695 47.805 118.865 ;
        RECT 47.385 118.655 47.805 118.695 ;
        RECT 46.095 118.185 46.515 118.525 ;
        RECT 46.805 118.195 47.215 118.525 ;
        RECT 44.335 117.765 45.185 117.935 ;
        RECT 45.745 117.545 46.065 118.005 ;
        RECT 46.265 117.755 46.515 118.185 ;
        RECT 46.805 117.545 47.215 117.985 ;
        RECT 47.385 117.925 47.555 118.655 ;
        RECT 47.725 118.105 48.075 118.475 ;
        RECT 48.255 118.165 48.475 119.035 ;
        RECT 48.645 118.465 49.055 119.085 ;
        RECT 49.225 118.285 49.395 119.255 ;
        RECT 48.700 118.095 49.395 118.285 ;
        RECT 47.385 117.725 48.400 117.925 ;
        RECT 48.700 117.765 48.870 118.095 ;
        RECT 49.040 117.545 49.370 117.925 ;
        RECT 49.585 117.805 49.810 119.925 ;
        RECT 49.980 119.595 50.310 120.095 ;
        RECT 50.480 119.425 50.650 119.925 ;
        RECT 51.285 119.755 51.540 119.785 ;
        RECT 51.200 119.585 51.540 119.755 ;
        RECT 49.985 119.255 50.650 119.425 ;
        RECT 49.985 118.265 50.215 119.255 ;
        RECT 51.285 119.115 51.540 119.585 ;
        RECT 51.720 119.295 52.005 120.095 ;
        RECT 52.185 119.375 52.515 119.885 ;
        RECT 50.385 118.435 50.735 119.085 ;
        RECT 49.985 118.095 50.650 118.265 ;
        RECT 49.980 117.545 50.310 117.925 ;
        RECT 50.480 117.805 50.650 118.095 ;
        RECT 51.285 118.255 51.465 119.115 ;
        RECT 52.185 118.785 52.435 119.375 ;
        RECT 52.785 119.225 52.955 119.835 ;
        RECT 53.125 119.405 53.455 120.095 ;
        RECT 53.685 119.545 53.925 119.835 ;
        RECT 54.125 119.715 54.545 120.095 ;
        RECT 54.725 119.625 55.355 119.875 ;
        RECT 55.825 119.715 56.155 120.095 ;
        RECT 54.725 119.545 54.895 119.625 ;
        RECT 56.325 119.545 56.495 119.835 ;
        RECT 56.675 119.715 57.055 120.095 ;
        RECT 57.295 119.710 58.125 119.880 ;
        RECT 53.685 119.375 54.895 119.545 ;
        RECT 51.635 118.455 52.435 118.785 ;
        RECT 51.285 117.725 51.540 118.255 ;
        RECT 51.720 117.545 52.005 118.005 ;
        RECT 52.185 117.805 52.435 118.455 ;
        RECT 52.635 119.205 52.955 119.225 ;
        RECT 52.635 119.035 54.555 119.205 ;
        RECT 52.635 118.140 52.825 119.035 ;
        RECT 54.725 118.865 54.895 119.375 ;
        RECT 55.065 119.115 55.585 119.425 ;
        RECT 52.995 118.695 54.895 118.865 ;
        RECT 52.995 118.635 53.325 118.695 ;
        RECT 53.475 118.465 53.805 118.525 ;
        RECT 53.145 118.195 53.805 118.465 ;
        RECT 52.635 117.810 52.955 118.140 ;
        RECT 53.135 117.545 53.795 118.025 ;
        RECT 53.995 117.935 54.165 118.695 ;
        RECT 55.065 118.525 55.245 118.935 ;
        RECT 54.335 118.355 54.665 118.475 ;
        RECT 55.415 118.355 55.585 119.115 ;
        RECT 54.335 118.185 55.585 118.355 ;
        RECT 55.755 119.295 57.125 119.545 ;
        RECT 55.755 118.525 55.945 119.295 ;
        RECT 56.875 119.035 57.125 119.295 ;
        RECT 56.115 118.865 56.365 119.025 ;
        RECT 57.295 118.865 57.465 119.710 ;
        RECT 58.360 119.425 58.530 119.925 ;
        RECT 58.700 119.595 59.030 120.095 ;
        RECT 57.635 119.035 58.135 119.415 ;
        RECT 58.360 119.255 59.055 119.425 ;
        RECT 56.115 118.695 57.465 118.865 ;
        RECT 57.045 118.655 57.465 118.695 ;
        RECT 55.755 118.185 56.175 118.525 ;
        RECT 56.465 118.195 56.875 118.525 ;
        RECT 53.995 117.765 54.845 117.935 ;
        RECT 55.405 117.545 55.725 118.005 ;
        RECT 55.925 117.755 56.175 118.185 ;
        RECT 56.465 117.545 56.875 117.985 ;
        RECT 57.045 117.925 57.215 118.655 ;
        RECT 57.385 118.105 57.735 118.475 ;
        RECT 57.915 118.165 58.135 119.035 ;
        RECT 58.305 118.465 58.715 119.085 ;
        RECT 58.885 118.285 59.055 119.255 ;
        RECT 58.360 118.095 59.055 118.285 ;
        RECT 57.045 117.725 58.060 117.925 ;
        RECT 58.360 117.765 58.530 118.095 ;
        RECT 58.700 117.545 59.030 117.925 ;
        RECT 59.245 117.805 59.470 119.925 ;
        RECT 59.640 119.595 59.970 120.095 ;
        RECT 60.140 119.425 60.310 119.925 ;
        RECT 59.645 119.255 60.310 119.425 ;
        RECT 59.645 118.265 59.875 119.255 ;
        RECT 60.045 118.435 60.395 119.085 ;
        RECT 60.570 118.930 60.860 120.095 ;
        RECT 61.030 119.020 61.300 119.925 ;
        RECT 61.470 119.335 61.800 120.095 ;
        RECT 61.980 119.165 62.150 119.925 ;
        RECT 63.705 119.755 63.960 119.785 ;
        RECT 63.620 119.585 63.960 119.755 ;
        RECT 59.645 118.095 60.310 118.265 ;
        RECT 59.640 117.545 59.970 117.925 ;
        RECT 60.140 117.805 60.310 118.095 ;
        RECT 60.570 117.545 60.860 118.270 ;
        RECT 61.030 118.220 61.200 119.020 ;
        RECT 61.485 118.995 62.150 119.165 ;
        RECT 63.705 119.115 63.960 119.585 ;
        RECT 64.140 119.295 64.425 120.095 ;
        RECT 64.605 119.375 64.935 119.885 ;
        RECT 61.485 118.850 61.655 118.995 ;
        RECT 61.370 118.520 61.655 118.850 ;
        RECT 61.485 118.265 61.655 118.520 ;
        RECT 61.890 118.445 62.220 118.815 ;
        RECT 61.030 117.715 61.290 118.220 ;
        RECT 61.485 118.095 62.150 118.265 ;
        RECT 61.470 117.545 61.800 117.925 ;
        RECT 61.980 117.715 62.150 118.095 ;
        RECT 63.705 118.255 63.885 119.115 ;
        RECT 64.605 118.785 64.855 119.375 ;
        RECT 65.205 119.225 65.375 119.835 ;
        RECT 65.545 119.405 65.875 120.095 ;
        RECT 66.105 119.545 66.345 119.835 ;
        RECT 66.545 119.715 66.965 120.095 ;
        RECT 67.145 119.625 67.775 119.875 ;
        RECT 68.245 119.715 68.575 120.095 ;
        RECT 67.145 119.545 67.315 119.625 ;
        RECT 68.745 119.545 68.915 119.835 ;
        RECT 69.095 119.715 69.475 120.095 ;
        RECT 69.715 119.710 70.545 119.880 ;
        RECT 66.105 119.375 67.315 119.545 ;
        RECT 64.055 118.455 64.855 118.785 ;
        RECT 63.705 117.725 63.960 118.255 ;
        RECT 64.140 117.545 64.425 118.005 ;
        RECT 64.605 117.805 64.855 118.455 ;
        RECT 65.055 119.205 65.375 119.225 ;
        RECT 65.055 119.035 66.975 119.205 ;
        RECT 65.055 118.140 65.245 119.035 ;
        RECT 67.145 118.865 67.315 119.375 ;
        RECT 67.485 119.115 68.005 119.425 ;
        RECT 65.415 118.695 67.315 118.865 ;
        RECT 65.415 118.635 65.745 118.695 ;
        RECT 65.895 118.465 66.225 118.525 ;
        RECT 65.565 118.195 66.225 118.465 ;
        RECT 65.055 117.810 65.375 118.140 ;
        RECT 65.555 117.545 66.215 118.025 ;
        RECT 66.415 117.935 66.585 118.695 ;
        RECT 67.485 118.525 67.665 118.935 ;
        RECT 66.755 118.355 67.085 118.475 ;
        RECT 67.835 118.355 68.005 119.115 ;
        RECT 66.755 118.185 68.005 118.355 ;
        RECT 68.175 119.295 69.545 119.545 ;
        RECT 68.175 118.525 68.365 119.295 ;
        RECT 69.295 119.035 69.545 119.295 ;
        RECT 68.535 118.865 68.785 119.025 ;
        RECT 69.715 118.865 69.885 119.710 ;
        RECT 70.780 119.425 70.950 119.925 ;
        RECT 71.120 119.595 71.450 120.095 ;
        RECT 70.055 119.035 70.555 119.415 ;
        RECT 70.780 119.255 71.475 119.425 ;
        RECT 68.535 118.695 69.885 118.865 ;
        RECT 69.465 118.655 69.885 118.695 ;
        RECT 68.175 118.185 68.595 118.525 ;
        RECT 68.885 118.195 69.295 118.525 ;
        RECT 66.415 117.765 67.265 117.935 ;
        RECT 67.825 117.545 68.145 118.005 ;
        RECT 68.345 117.755 68.595 118.185 ;
        RECT 68.885 117.545 69.295 117.985 ;
        RECT 69.465 117.925 69.635 118.655 ;
        RECT 69.805 118.105 70.155 118.475 ;
        RECT 70.335 118.165 70.555 119.035 ;
        RECT 70.725 118.465 71.135 119.085 ;
        RECT 71.305 118.285 71.475 119.255 ;
        RECT 70.780 118.095 71.475 118.285 ;
        RECT 69.465 117.725 70.480 117.925 ;
        RECT 70.780 117.765 70.950 118.095 ;
        RECT 71.120 117.545 71.450 117.925 ;
        RECT 71.665 117.805 71.890 119.925 ;
        RECT 72.060 119.595 72.390 120.095 ;
        RECT 72.560 119.425 72.730 119.925 ;
        RECT 72.065 119.255 72.730 119.425 ;
        RECT 72.065 118.265 72.295 119.255 ;
        RECT 72.465 118.435 72.815 119.085 ;
        RECT 72.995 118.955 73.330 119.925 ;
        RECT 73.500 118.955 73.670 120.095 ;
        RECT 73.840 119.755 75.870 119.925 ;
        RECT 72.995 118.285 73.165 118.955 ;
        RECT 73.840 118.785 74.010 119.755 ;
        RECT 73.335 118.455 73.590 118.785 ;
        RECT 73.815 118.455 74.010 118.785 ;
        RECT 74.180 119.415 75.305 119.585 ;
        RECT 73.420 118.285 73.590 118.455 ;
        RECT 74.180 118.285 74.350 119.415 ;
        RECT 72.065 118.095 72.730 118.265 ;
        RECT 72.060 117.545 72.390 117.925 ;
        RECT 72.560 117.805 72.730 118.095 ;
        RECT 72.995 117.715 73.250 118.285 ;
        RECT 73.420 118.115 74.350 118.285 ;
        RECT 74.520 119.075 75.530 119.245 ;
        RECT 74.520 118.275 74.690 119.075 ;
        RECT 74.175 118.080 74.350 118.115 ;
        RECT 73.420 117.545 73.750 117.945 ;
        RECT 74.175 117.715 74.705 118.080 ;
        RECT 74.895 118.055 75.170 118.875 ;
        RECT 74.890 117.885 75.170 118.055 ;
        RECT 74.895 117.715 75.170 117.885 ;
        RECT 75.340 117.715 75.530 119.075 ;
        RECT 75.700 119.090 75.870 119.755 ;
        RECT 76.040 119.335 76.210 120.095 ;
        RECT 76.445 119.335 76.960 119.745 ;
        RECT 75.700 118.900 76.450 119.090 ;
        RECT 76.620 118.525 76.960 119.335 ;
        RECT 75.730 118.355 76.960 118.525 ;
        RECT 77.130 119.005 78.340 120.095 ;
        RECT 77.130 118.465 77.650 119.005 ;
        RECT 78.515 118.955 78.850 119.925 ;
        RECT 79.020 118.955 79.190 120.095 ;
        RECT 79.360 119.755 81.390 119.925 ;
        RECT 75.710 117.545 76.220 118.080 ;
        RECT 76.440 117.750 76.685 118.355 ;
        RECT 77.820 118.295 78.340 118.835 ;
        RECT 77.130 117.545 78.340 118.295 ;
        RECT 78.515 118.285 78.685 118.955 ;
        RECT 79.360 118.785 79.530 119.755 ;
        RECT 78.855 118.455 79.110 118.785 ;
        RECT 79.335 118.455 79.530 118.785 ;
        RECT 79.700 119.415 80.825 119.585 ;
        RECT 78.940 118.285 79.110 118.455 ;
        RECT 79.700 118.285 79.870 119.415 ;
        RECT 78.515 117.715 78.770 118.285 ;
        RECT 78.940 118.115 79.870 118.285 ;
        RECT 80.040 119.075 81.050 119.245 ;
        RECT 80.040 118.275 80.210 119.075 ;
        RECT 80.415 118.735 80.690 118.875 ;
        RECT 80.410 118.565 80.690 118.735 ;
        RECT 79.695 118.080 79.870 118.115 ;
        RECT 78.940 117.545 79.270 117.945 ;
        RECT 79.695 117.715 80.225 118.080 ;
        RECT 80.415 117.715 80.690 118.565 ;
        RECT 80.860 117.715 81.050 119.075 ;
        RECT 81.220 119.090 81.390 119.755 ;
        RECT 81.560 119.335 81.730 120.095 ;
        RECT 81.965 119.335 82.480 119.745 ;
        RECT 81.220 118.900 81.970 119.090 ;
        RECT 82.140 118.525 82.480 119.335 ;
        RECT 81.250 118.355 82.480 118.525 ;
        RECT 82.650 119.005 86.160 120.095 ;
        RECT 82.650 118.485 84.340 119.005 ;
        RECT 86.330 118.930 86.620 120.095 ;
        RECT 86.790 119.005 88.000 120.095 ;
        RECT 81.230 117.545 81.740 118.080 ;
        RECT 81.960 117.750 82.205 118.355 ;
        RECT 84.510 118.315 86.160 118.835 ;
        RECT 86.790 118.465 87.310 119.005 ;
        RECT 88.210 118.955 88.440 120.095 ;
        RECT 88.610 118.945 88.940 119.925 ;
        RECT 89.110 118.955 89.320 120.095 ;
        RECT 89.925 119.755 90.180 119.785 ;
        RECT 89.840 119.585 90.180 119.755 ;
        RECT 89.925 119.115 90.180 119.585 ;
        RECT 90.360 119.295 90.645 120.095 ;
        RECT 90.825 119.375 91.155 119.885 ;
        RECT 82.650 117.545 86.160 118.315 ;
        RECT 87.480 118.295 88.000 118.835 ;
        RECT 88.190 118.535 88.520 118.785 ;
        RECT 86.330 117.545 86.620 118.270 ;
        RECT 86.790 117.545 88.000 118.295 ;
        RECT 88.210 117.545 88.440 118.365 ;
        RECT 88.690 118.345 88.940 118.945 ;
        RECT 88.610 117.715 88.940 118.345 ;
        RECT 89.110 117.545 89.320 118.365 ;
        RECT 89.925 118.255 90.105 119.115 ;
        RECT 90.825 118.785 91.075 119.375 ;
        RECT 91.425 119.225 91.595 119.835 ;
        RECT 91.765 119.405 92.095 120.095 ;
        RECT 92.325 119.545 92.565 119.835 ;
        RECT 92.765 119.715 93.185 120.095 ;
        RECT 93.365 119.625 93.995 119.875 ;
        RECT 94.465 119.715 94.795 120.095 ;
        RECT 93.365 119.545 93.535 119.625 ;
        RECT 94.965 119.545 95.135 119.835 ;
        RECT 95.315 119.715 95.695 120.095 ;
        RECT 95.935 119.710 96.765 119.880 ;
        RECT 92.325 119.375 93.535 119.545 ;
        RECT 90.275 118.455 91.075 118.785 ;
        RECT 89.925 117.725 90.180 118.255 ;
        RECT 90.360 117.545 90.645 118.005 ;
        RECT 90.825 117.805 91.075 118.455 ;
        RECT 91.275 119.205 91.595 119.225 ;
        RECT 91.275 119.035 93.195 119.205 ;
        RECT 91.275 118.140 91.465 119.035 ;
        RECT 93.365 118.865 93.535 119.375 ;
        RECT 93.705 119.115 94.225 119.425 ;
        RECT 91.635 118.695 93.535 118.865 ;
        RECT 91.635 118.635 91.965 118.695 ;
        RECT 92.115 118.465 92.445 118.525 ;
        RECT 91.785 118.195 92.445 118.465 ;
        RECT 91.275 117.810 91.595 118.140 ;
        RECT 91.775 117.545 92.435 118.025 ;
        RECT 92.635 117.935 92.805 118.695 ;
        RECT 93.705 118.525 93.885 118.935 ;
        RECT 92.975 118.355 93.305 118.475 ;
        RECT 94.055 118.355 94.225 119.115 ;
        RECT 92.975 118.185 94.225 118.355 ;
        RECT 94.395 119.295 95.765 119.545 ;
        RECT 94.395 118.525 94.585 119.295 ;
        RECT 95.515 119.035 95.765 119.295 ;
        RECT 94.755 118.865 95.005 119.025 ;
        RECT 95.935 118.865 96.105 119.710 ;
        RECT 97.000 119.425 97.170 119.925 ;
        RECT 97.340 119.595 97.670 120.095 ;
        RECT 96.275 119.035 96.775 119.415 ;
        RECT 97.000 119.255 97.695 119.425 ;
        RECT 94.755 118.695 96.105 118.865 ;
        RECT 95.685 118.655 96.105 118.695 ;
        RECT 94.395 118.185 94.815 118.525 ;
        RECT 95.105 118.195 95.515 118.525 ;
        RECT 92.635 117.765 93.485 117.935 ;
        RECT 94.045 117.545 94.365 118.005 ;
        RECT 94.565 117.755 94.815 118.185 ;
        RECT 95.105 117.545 95.515 117.985 ;
        RECT 95.685 117.925 95.855 118.655 ;
        RECT 96.025 118.105 96.375 118.475 ;
        RECT 96.555 118.165 96.775 119.035 ;
        RECT 96.945 118.465 97.355 119.085 ;
        RECT 97.525 118.285 97.695 119.255 ;
        RECT 97.000 118.095 97.695 118.285 ;
        RECT 95.685 117.725 96.700 117.925 ;
        RECT 97.000 117.765 97.170 118.095 ;
        RECT 97.340 117.545 97.670 117.925 ;
        RECT 97.885 117.805 98.110 119.925 ;
        RECT 98.280 119.595 98.610 120.095 ;
        RECT 98.780 119.425 98.950 119.925 ;
        RECT 98.285 119.255 98.950 119.425 ;
        RECT 98.285 118.265 98.515 119.255 ;
        RECT 98.685 118.435 99.035 119.085 ;
        RECT 100.170 118.955 100.400 120.095 ;
        RECT 100.570 118.945 100.900 119.925 ;
        RECT 101.070 118.955 101.280 120.095 ;
        RECT 101.885 119.755 102.140 119.785 ;
        RECT 101.800 119.585 102.140 119.755 ;
        RECT 101.885 119.115 102.140 119.585 ;
        RECT 102.320 119.295 102.605 120.095 ;
        RECT 102.785 119.375 103.115 119.885 ;
        RECT 100.150 118.535 100.480 118.785 ;
        RECT 98.285 118.095 98.950 118.265 ;
        RECT 98.280 117.545 98.610 117.925 ;
        RECT 98.780 117.805 98.950 118.095 ;
        RECT 100.170 117.545 100.400 118.365 ;
        RECT 100.650 118.345 100.900 118.945 ;
        RECT 100.570 117.715 100.900 118.345 ;
        RECT 101.070 117.545 101.280 118.365 ;
        RECT 101.885 118.255 102.065 119.115 ;
        RECT 102.785 118.785 103.035 119.375 ;
        RECT 103.385 119.225 103.555 119.835 ;
        RECT 103.725 119.405 104.055 120.095 ;
        RECT 104.285 119.545 104.525 119.835 ;
        RECT 104.725 119.715 105.145 120.095 ;
        RECT 105.325 119.625 105.955 119.875 ;
        RECT 106.425 119.715 106.755 120.095 ;
        RECT 105.325 119.545 105.495 119.625 ;
        RECT 106.925 119.545 107.095 119.835 ;
        RECT 107.275 119.715 107.655 120.095 ;
        RECT 107.895 119.710 108.725 119.880 ;
        RECT 104.285 119.375 105.495 119.545 ;
        RECT 102.235 118.455 103.035 118.785 ;
        RECT 101.885 117.725 102.140 118.255 ;
        RECT 102.320 117.545 102.605 118.005 ;
        RECT 102.785 117.805 103.035 118.455 ;
        RECT 103.235 119.205 103.555 119.225 ;
        RECT 103.235 119.035 105.155 119.205 ;
        RECT 103.235 118.140 103.425 119.035 ;
        RECT 105.325 118.865 105.495 119.375 ;
        RECT 105.665 119.115 106.185 119.425 ;
        RECT 103.595 118.695 105.495 118.865 ;
        RECT 103.595 118.635 103.925 118.695 ;
        RECT 104.075 118.465 104.405 118.525 ;
        RECT 103.745 118.195 104.405 118.465 ;
        RECT 103.235 117.810 103.555 118.140 ;
        RECT 103.735 117.545 104.395 118.025 ;
        RECT 104.595 117.935 104.765 118.695 ;
        RECT 105.665 118.525 105.845 118.935 ;
        RECT 104.935 118.355 105.265 118.475 ;
        RECT 106.015 118.355 106.185 119.115 ;
        RECT 104.935 118.185 106.185 118.355 ;
        RECT 106.355 119.295 107.725 119.545 ;
        RECT 106.355 118.525 106.545 119.295 ;
        RECT 107.475 119.035 107.725 119.295 ;
        RECT 106.715 118.865 106.965 119.025 ;
        RECT 107.895 118.865 108.065 119.710 ;
        RECT 108.960 119.425 109.130 119.925 ;
        RECT 109.300 119.595 109.630 120.095 ;
        RECT 108.235 119.035 108.735 119.415 ;
        RECT 108.960 119.255 109.655 119.425 ;
        RECT 106.715 118.695 108.065 118.865 ;
        RECT 107.645 118.655 108.065 118.695 ;
        RECT 106.355 118.185 106.775 118.525 ;
        RECT 107.065 118.195 107.475 118.525 ;
        RECT 104.595 117.765 105.445 117.935 ;
        RECT 106.005 117.545 106.325 118.005 ;
        RECT 106.525 117.755 106.775 118.185 ;
        RECT 107.065 117.545 107.475 117.985 ;
        RECT 107.645 117.925 107.815 118.655 ;
        RECT 107.985 118.105 108.335 118.475 ;
        RECT 108.515 118.165 108.735 119.035 ;
        RECT 108.905 118.465 109.315 119.085 ;
        RECT 109.485 118.285 109.655 119.255 ;
        RECT 108.960 118.095 109.655 118.285 ;
        RECT 107.645 117.725 108.660 117.925 ;
        RECT 108.960 117.765 109.130 118.095 ;
        RECT 109.300 117.545 109.630 117.925 ;
        RECT 109.845 117.805 110.070 119.925 ;
        RECT 110.240 119.595 110.570 120.095 ;
        RECT 110.740 119.425 110.910 119.925 ;
        RECT 110.245 119.255 110.910 119.425 ;
        RECT 110.245 118.265 110.475 119.255 ;
        RECT 110.645 118.435 110.995 119.085 ;
        RECT 111.170 119.005 112.380 120.095 ;
        RECT 111.170 118.465 111.690 119.005 ;
        RECT 111.860 118.295 112.380 118.835 ;
        RECT 110.245 118.095 110.910 118.265 ;
        RECT 110.240 117.545 110.570 117.925 ;
        RECT 110.740 117.805 110.910 118.095 ;
        RECT 111.170 117.545 112.380 118.295 ;
        RECT 18.165 117.375 112.465 117.545 ;
        RECT 18.250 116.625 19.460 117.375 ;
        RECT 18.250 116.085 18.770 116.625 ;
        RECT 20.090 116.605 21.760 117.375 ;
        RECT 21.930 116.650 22.220 117.375 ;
        RECT 18.940 115.915 19.460 116.455 ;
        RECT 18.250 114.825 19.460 115.915 ;
        RECT 20.090 115.915 20.840 116.435 ;
        RECT 21.010 116.085 21.760 116.605 ;
        RECT 23.350 116.555 23.580 117.375 ;
        RECT 23.750 116.575 24.080 117.205 ;
        RECT 23.330 116.135 23.660 116.385 ;
        RECT 20.090 114.825 21.760 115.915 ;
        RECT 21.930 114.825 22.220 115.990 ;
        RECT 23.830 115.975 24.080 116.575 ;
        RECT 24.250 116.555 24.460 117.375 ;
        RECT 25.700 116.825 25.870 117.205 ;
        RECT 26.050 116.995 26.380 117.375 ;
        RECT 25.700 116.655 26.365 116.825 ;
        RECT 26.560 116.700 26.820 117.205 ;
        RECT 25.630 116.105 25.960 116.475 ;
        RECT 26.195 116.400 26.365 116.655 ;
        RECT 23.350 114.825 23.580 115.965 ;
        RECT 23.750 114.995 24.080 115.975 ;
        RECT 26.195 116.070 26.480 116.400 ;
        RECT 24.250 114.825 24.460 115.965 ;
        RECT 26.195 115.925 26.365 116.070 ;
        RECT 25.700 115.755 26.365 115.925 ;
        RECT 26.650 115.900 26.820 116.700 ;
        RECT 27.030 116.555 27.260 117.375 ;
        RECT 27.430 116.575 27.760 117.205 ;
        RECT 27.010 116.135 27.340 116.385 ;
        RECT 27.510 115.975 27.760 116.575 ;
        RECT 27.930 116.555 28.140 117.375 ;
        RECT 28.460 116.825 28.630 117.115 ;
        RECT 28.800 116.995 29.130 117.375 ;
        RECT 28.460 116.655 29.125 116.825 ;
        RECT 25.700 114.995 25.870 115.755 ;
        RECT 26.050 114.825 26.380 115.585 ;
        RECT 26.550 114.995 26.820 115.900 ;
        RECT 27.030 114.825 27.260 115.965 ;
        RECT 27.430 114.995 27.760 115.975 ;
        RECT 27.930 114.825 28.140 115.965 ;
        RECT 28.375 115.835 28.725 116.485 ;
        RECT 28.895 115.665 29.125 116.655 ;
        RECT 28.460 115.495 29.125 115.665 ;
        RECT 28.460 114.995 28.630 115.495 ;
        RECT 28.800 114.825 29.130 115.325 ;
        RECT 29.300 114.995 29.525 117.115 ;
        RECT 29.740 116.995 30.070 117.375 ;
        RECT 30.240 116.825 30.410 117.155 ;
        RECT 30.710 116.995 31.725 117.195 ;
        RECT 29.715 116.635 30.410 116.825 ;
        RECT 29.715 115.665 29.885 116.635 ;
        RECT 30.055 115.835 30.465 116.455 ;
        RECT 30.635 115.885 30.855 116.755 ;
        RECT 31.035 116.445 31.385 116.815 ;
        RECT 31.555 116.265 31.725 116.995 ;
        RECT 31.895 116.935 32.305 117.375 ;
        RECT 32.595 116.735 32.845 117.165 ;
        RECT 33.045 116.915 33.365 117.375 ;
        RECT 33.925 116.985 34.775 117.155 ;
        RECT 31.895 116.395 32.305 116.725 ;
        RECT 32.595 116.395 33.015 116.735 ;
        RECT 31.305 116.225 31.725 116.265 ;
        RECT 31.305 116.055 32.655 116.225 ;
        RECT 29.715 115.495 30.410 115.665 ;
        RECT 30.635 115.505 31.135 115.885 ;
        RECT 29.740 114.825 30.070 115.325 ;
        RECT 30.240 114.995 30.410 115.495 ;
        RECT 31.305 115.210 31.475 116.055 ;
        RECT 32.405 115.895 32.655 116.055 ;
        RECT 31.645 115.625 31.895 115.885 ;
        RECT 32.825 115.625 33.015 116.395 ;
        RECT 31.645 115.375 33.015 115.625 ;
        RECT 33.185 116.565 34.435 116.735 ;
        RECT 33.185 115.805 33.355 116.565 ;
        RECT 34.105 116.445 34.435 116.565 ;
        RECT 33.525 115.985 33.705 116.395 ;
        RECT 34.605 116.225 34.775 116.985 ;
        RECT 34.975 116.895 35.635 117.375 ;
        RECT 35.815 116.780 36.135 117.110 ;
        RECT 34.965 116.455 35.625 116.725 ;
        RECT 34.965 116.395 35.295 116.455 ;
        RECT 35.445 116.225 35.775 116.285 ;
        RECT 33.875 116.055 35.775 116.225 ;
        RECT 33.185 115.495 33.705 115.805 ;
        RECT 33.875 115.545 34.045 116.055 ;
        RECT 35.945 115.885 36.135 116.780 ;
        RECT 34.215 115.715 36.135 115.885 ;
        RECT 35.815 115.695 36.135 115.715 ;
        RECT 36.335 116.465 36.585 117.115 ;
        RECT 36.765 116.915 37.050 117.375 ;
        RECT 37.230 117.035 37.485 117.195 ;
        RECT 38.405 117.035 38.660 117.195 ;
        RECT 37.230 116.865 37.570 117.035 ;
        RECT 38.320 116.865 38.660 117.035 ;
        RECT 38.840 116.915 39.125 117.375 ;
        RECT 37.230 116.665 37.485 116.865 ;
        RECT 36.335 116.135 37.135 116.465 ;
        RECT 33.875 115.375 35.085 115.545 ;
        RECT 30.645 115.040 31.475 115.210 ;
        RECT 31.715 114.825 32.095 115.205 ;
        RECT 32.275 115.085 32.445 115.375 ;
        RECT 33.875 115.295 34.045 115.375 ;
        RECT 32.615 114.825 32.945 115.205 ;
        RECT 33.415 115.045 34.045 115.295 ;
        RECT 34.225 114.825 34.645 115.205 ;
        RECT 34.845 115.085 35.085 115.375 ;
        RECT 35.315 114.825 35.645 115.515 ;
        RECT 35.815 115.085 35.985 115.695 ;
        RECT 36.335 115.545 36.585 116.135 ;
        RECT 37.305 115.805 37.485 116.665 ;
        RECT 36.255 115.035 36.585 115.545 ;
        RECT 36.765 114.825 37.050 115.625 ;
        RECT 37.230 115.135 37.485 115.805 ;
        RECT 38.405 116.665 38.660 116.865 ;
        RECT 38.405 115.805 38.585 116.665 ;
        RECT 39.305 116.465 39.555 117.115 ;
        RECT 38.755 116.135 39.555 116.465 ;
        RECT 38.405 115.135 38.660 115.805 ;
        RECT 38.840 114.825 39.125 115.625 ;
        RECT 39.305 115.545 39.555 116.135 ;
        RECT 39.755 116.780 40.075 117.110 ;
        RECT 40.255 116.895 40.915 117.375 ;
        RECT 41.115 116.985 41.965 117.155 ;
        RECT 39.755 115.885 39.945 116.780 ;
        RECT 40.265 116.455 40.925 116.725 ;
        RECT 40.595 116.395 40.925 116.455 ;
        RECT 40.115 116.225 40.445 116.285 ;
        RECT 41.115 116.225 41.285 116.985 ;
        RECT 42.525 116.915 42.845 117.375 ;
        RECT 43.045 116.735 43.295 117.165 ;
        RECT 43.585 116.935 43.995 117.375 ;
        RECT 44.165 116.995 45.180 117.195 ;
        RECT 41.455 116.565 42.705 116.735 ;
        RECT 41.455 116.445 41.785 116.565 ;
        RECT 40.115 116.055 42.015 116.225 ;
        RECT 39.755 115.715 41.675 115.885 ;
        RECT 39.755 115.695 40.075 115.715 ;
        RECT 39.305 115.035 39.635 115.545 ;
        RECT 39.905 115.085 40.075 115.695 ;
        RECT 41.845 115.545 42.015 116.055 ;
        RECT 42.185 115.985 42.365 116.395 ;
        RECT 42.535 115.805 42.705 116.565 ;
        RECT 40.245 114.825 40.575 115.515 ;
        RECT 40.805 115.375 42.015 115.545 ;
        RECT 42.185 115.495 42.705 115.805 ;
        RECT 42.875 116.395 43.295 116.735 ;
        RECT 43.585 116.395 43.995 116.725 ;
        RECT 42.875 115.625 43.065 116.395 ;
        RECT 44.165 116.265 44.335 116.995 ;
        RECT 45.480 116.825 45.650 117.155 ;
        RECT 45.820 116.995 46.150 117.375 ;
        RECT 44.505 116.445 44.855 116.815 ;
        RECT 44.165 116.225 44.585 116.265 ;
        RECT 43.235 116.055 44.585 116.225 ;
        RECT 43.235 115.895 43.485 116.055 ;
        RECT 43.995 115.625 44.245 115.885 ;
        RECT 42.875 115.375 44.245 115.625 ;
        RECT 40.805 115.085 41.045 115.375 ;
        RECT 41.845 115.295 42.015 115.375 ;
        RECT 41.245 114.825 41.665 115.205 ;
        RECT 41.845 115.045 42.475 115.295 ;
        RECT 42.945 114.825 43.275 115.205 ;
        RECT 43.445 115.085 43.615 115.375 ;
        RECT 44.415 115.210 44.585 116.055 ;
        RECT 45.035 115.885 45.255 116.755 ;
        RECT 45.480 116.635 46.175 116.825 ;
        RECT 44.755 115.505 45.255 115.885 ;
        RECT 45.425 115.835 45.835 116.455 ;
        RECT 46.005 115.665 46.175 116.635 ;
        RECT 45.480 115.495 46.175 115.665 ;
        RECT 43.795 114.825 44.175 115.205 ;
        RECT 44.415 115.040 45.245 115.210 ;
        RECT 45.480 114.995 45.650 115.495 ;
        RECT 45.820 114.825 46.150 115.325 ;
        RECT 46.365 114.995 46.590 117.115 ;
        RECT 46.760 116.995 47.090 117.375 ;
        RECT 47.260 116.825 47.430 117.115 ;
        RECT 46.765 116.655 47.430 116.825 ;
        RECT 46.765 115.665 46.995 116.655 ;
        RECT 47.690 116.650 47.980 117.375 ;
        RECT 49.345 116.565 49.590 117.170 ;
        RECT 49.810 116.840 50.320 117.375 ;
        RECT 47.165 115.835 47.515 116.485 ;
        RECT 49.070 116.395 50.300 116.565 ;
        RECT 46.765 115.495 47.430 115.665 ;
        RECT 46.760 114.825 47.090 115.325 ;
        RECT 47.260 114.995 47.430 115.495 ;
        RECT 47.690 114.825 47.980 115.990 ;
        RECT 49.070 115.585 49.410 116.395 ;
        RECT 49.580 115.830 50.330 116.020 ;
        RECT 49.070 115.175 49.585 115.585 ;
        RECT 49.820 114.825 49.990 115.585 ;
        RECT 50.160 115.165 50.330 115.830 ;
        RECT 50.500 115.845 50.690 117.205 ;
        RECT 50.860 117.035 51.135 117.205 ;
        RECT 50.860 116.865 51.140 117.035 ;
        RECT 50.860 116.045 51.135 116.865 ;
        RECT 51.325 116.840 51.855 117.205 ;
        RECT 52.280 116.975 52.610 117.375 ;
        RECT 51.680 116.805 51.855 116.840 ;
        RECT 51.340 115.845 51.510 116.645 ;
        RECT 50.500 115.675 51.510 115.845 ;
        RECT 51.680 116.635 52.610 116.805 ;
        RECT 52.780 116.635 53.035 117.205 ;
        RECT 53.585 117.035 53.840 117.195 ;
        RECT 53.500 116.865 53.840 117.035 ;
        RECT 54.020 116.915 54.305 117.375 ;
        RECT 51.680 115.505 51.850 116.635 ;
        RECT 52.440 116.465 52.610 116.635 ;
        RECT 50.725 115.335 51.850 115.505 ;
        RECT 52.020 116.135 52.215 116.465 ;
        RECT 52.440 116.135 52.695 116.465 ;
        RECT 52.020 115.165 52.190 116.135 ;
        RECT 52.865 115.965 53.035 116.635 ;
        RECT 50.160 114.995 52.190 115.165 ;
        RECT 52.360 114.825 52.530 115.965 ;
        RECT 52.700 114.995 53.035 115.965 ;
        RECT 53.585 116.665 53.840 116.865 ;
        RECT 53.585 115.805 53.765 116.665 ;
        RECT 54.485 116.465 54.735 117.115 ;
        RECT 53.935 116.135 54.735 116.465 ;
        RECT 53.585 115.135 53.840 115.805 ;
        RECT 54.020 114.825 54.305 115.625 ;
        RECT 54.485 115.545 54.735 116.135 ;
        RECT 54.935 116.780 55.255 117.110 ;
        RECT 55.435 116.895 56.095 117.375 ;
        RECT 56.295 116.985 57.145 117.155 ;
        RECT 54.935 115.885 55.125 116.780 ;
        RECT 55.445 116.455 56.105 116.725 ;
        RECT 55.775 116.395 56.105 116.455 ;
        RECT 55.295 116.225 55.625 116.285 ;
        RECT 56.295 116.225 56.465 116.985 ;
        RECT 57.705 116.915 58.025 117.375 ;
        RECT 58.225 116.735 58.475 117.165 ;
        RECT 58.765 116.935 59.175 117.375 ;
        RECT 59.345 116.995 60.360 117.195 ;
        RECT 56.635 116.565 57.885 116.735 ;
        RECT 56.635 116.445 56.965 116.565 ;
        RECT 55.295 116.055 57.195 116.225 ;
        RECT 54.935 115.715 56.855 115.885 ;
        RECT 54.935 115.695 55.255 115.715 ;
        RECT 54.485 115.035 54.815 115.545 ;
        RECT 55.085 115.085 55.255 115.695 ;
        RECT 57.025 115.545 57.195 116.055 ;
        RECT 57.365 115.985 57.545 116.395 ;
        RECT 57.715 115.805 57.885 116.565 ;
        RECT 55.425 114.825 55.755 115.515 ;
        RECT 55.985 115.375 57.195 115.545 ;
        RECT 57.365 115.495 57.885 115.805 ;
        RECT 58.055 116.395 58.475 116.735 ;
        RECT 58.765 116.395 59.175 116.725 ;
        RECT 58.055 115.625 58.245 116.395 ;
        RECT 59.345 116.265 59.515 116.995 ;
        RECT 60.660 116.825 60.830 117.155 ;
        RECT 61.000 116.995 61.330 117.375 ;
        RECT 59.685 116.445 60.035 116.815 ;
        RECT 59.345 116.225 59.765 116.265 ;
        RECT 58.415 116.055 59.765 116.225 ;
        RECT 58.415 115.895 58.665 116.055 ;
        RECT 59.175 115.625 59.425 115.885 ;
        RECT 58.055 115.375 59.425 115.625 ;
        RECT 55.985 115.085 56.225 115.375 ;
        RECT 57.025 115.295 57.195 115.375 ;
        RECT 56.425 114.825 56.845 115.205 ;
        RECT 57.025 115.045 57.655 115.295 ;
        RECT 58.125 114.825 58.455 115.205 ;
        RECT 58.625 115.085 58.795 115.375 ;
        RECT 59.595 115.210 59.765 116.055 ;
        RECT 60.215 115.885 60.435 116.755 ;
        RECT 60.660 116.635 61.355 116.825 ;
        RECT 59.935 115.505 60.435 115.885 ;
        RECT 60.605 115.835 61.015 116.455 ;
        RECT 61.185 115.665 61.355 116.635 ;
        RECT 60.660 115.495 61.355 115.665 ;
        RECT 58.975 114.825 59.355 115.205 ;
        RECT 59.595 115.040 60.425 115.210 ;
        RECT 60.660 114.995 60.830 115.495 ;
        RECT 61.000 114.825 61.330 115.325 ;
        RECT 61.545 114.995 61.770 117.115 ;
        RECT 61.940 116.995 62.270 117.375 ;
        RECT 62.440 116.825 62.610 117.115 ;
        RECT 61.945 116.655 62.610 116.825 ;
        RECT 61.945 115.665 62.175 116.655 ;
        RECT 63.330 116.605 65.920 117.375 ;
        RECT 62.345 115.835 62.695 116.485 ;
        RECT 63.330 115.915 64.540 116.435 ;
        RECT 64.710 116.085 65.920 116.605 ;
        RECT 66.130 116.555 66.360 117.375 ;
        RECT 66.530 116.575 66.860 117.205 ;
        RECT 66.110 116.135 66.440 116.385 ;
        RECT 66.610 115.975 66.860 116.575 ;
        RECT 67.030 116.555 67.240 117.375 ;
        RECT 67.745 116.565 67.990 117.170 ;
        RECT 68.210 116.840 68.720 117.375 ;
        RECT 61.945 115.495 62.610 115.665 ;
        RECT 61.940 114.825 62.270 115.325 ;
        RECT 62.440 114.995 62.610 115.495 ;
        RECT 63.330 114.825 65.920 115.915 ;
        RECT 66.130 114.825 66.360 115.965 ;
        RECT 66.530 114.995 66.860 115.975 ;
        RECT 67.470 116.395 68.700 116.565 ;
        RECT 67.030 114.825 67.240 115.965 ;
        RECT 67.470 115.585 67.810 116.395 ;
        RECT 67.980 115.830 68.730 116.020 ;
        RECT 67.470 115.175 67.985 115.585 ;
        RECT 68.220 114.825 68.390 115.585 ;
        RECT 68.560 115.165 68.730 115.830 ;
        RECT 68.900 115.845 69.090 117.205 ;
        RECT 69.260 117.035 69.535 117.205 ;
        RECT 69.260 116.865 69.540 117.035 ;
        RECT 69.260 116.045 69.535 116.865 ;
        RECT 69.725 116.840 70.255 117.205 ;
        RECT 70.680 116.975 71.010 117.375 ;
        RECT 70.080 116.805 70.255 116.840 ;
        RECT 69.740 115.845 69.910 116.645 ;
        RECT 68.900 115.675 69.910 115.845 ;
        RECT 70.080 116.635 71.010 116.805 ;
        RECT 71.180 116.635 71.435 117.205 ;
        RECT 70.080 115.505 70.250 116.635 ;
        RECT 70.840 116.465 71.010 116.635 ;
        RECT 69.125 115.335 70.250 115.505 ;
        RECT 70.420 116.135 70.615 116.465 ;
        RECT 70.840 116.135 71.095 116.465 ;
        RECT 70.420 115.165 70.590 116.135 ;
        RECT 71.265 115.965 71.435 116.635 ;
        RECT 68.560 114.995 70.590 115.165 ;
        RECT 70.760 114.825 70.930 115.965 ;
        RECT 71.100 114.995 71.435 115.965 ;
        RECT 71.610 116.700 71.870 117.205 ;
        RECT 72.050 116.995 72.380 117.375 ;
        RECT 72.560 116.825 72.730 117.205 ;
        RECT 71.610 115.900 71.780 116.700 ;
        RECT 72.065 116.655 72.730 116.825 ;
        RECT 72.065 116.400 72.235 116.655 ;
        RECT 73.450 116.650 73.740 117.375 ;
        RECT 75.205 117.035 75.460 117.195 ;
        RECT 75.120 116.865 75.460 117.035 ;
        RECT 75.640 116.915 75.925 117.375 ;
        RECT 75.205 116.665 75.460 116.865 ;
        RECT 71.950 116.070 72.235 116.400 ;
        RECT 72.470 116.105 72.800 116.475 ;
        RECT 72.065 115.925 72.235 116.070 ;
        RECT 71.610 114.995 71.880 115.900 ;
        RECT 72.065 115.755 72.730 115.925 ;
        RECT 72.050 114.825 72.380 115.585 ;
        RECT 72.560 114.995 72.730 115.755 ;
        RECT 73.450 114.825 73.740 115.990 ;
        RECT 75.205 115.805 75.385 116.665 ;
        RECT 76.105 116.465 76.355 117.115 ;
        RECT 75.555 116.135 76.355 116.465 ;
        RECT 75.205 115.135 75.460 115.805 ;
        RECT 75.640 114.825 75.925 115.625 ;
        RECT 76.105 115.545 76.355 116.135 ;
        RECT 76.555 116.780 76.875 117.110 ;
        RECT 77.055 116.895 77.715 117.375 ;
        RECT 77.915 116.985 78.765 117.155 ;
        RECT 76.555 115.885 76.745 116.780 ;
        RECT 77.065 116.455 77.725 116.725 ;
        RECT 77.395 116.395 77.725 116.455 ;
        RECT 76.915 116.225 77.245 116.285 ;
        RECT 77.915 116.225 78.085 116.985 ;
        RECT 79.325 116.915 79.645 117.375 ;
        RECT 79.845 116.735 80.095 117.165 ;
        RECT 80.385 116.935 80.795 117.375 ;
        RECT 80.965 116.995 81.980 117.195 ;
        RECT 78.255 116.565 79.505 116.735 ;
        RECT 78.255 116.445 78.585 116.565 ;
        RECT 76.915 116.055 78.815 116.225 ;
        RECT 76.555 115.715 78.475 115.885 ;
        RECT 76.555 115.695 76.875 115.715 ;
        RECT 76.105 115.035 76.435 115.545 ;
        RECT 76.705 115.085 76.875 115.695 ;
        RECT 78.645 115.545 78.815 116.055 ;
        RECT 78.985 115.985 79.165 116.395 ;
        RECT 79.335 115.805 79.505 116.565 ;
        RECT 77.045 114.825 77.375 115.515 ;
        RECT 77.605 115.375 78.815 115.545 ;
        RECT 78.985 115.495 79.505 115.805 ;
        RECT 79.675 116.395 80.095 116.735 ;
        RECT 80.385 116.395 80.795 116.725 ;
        RECT 79.675 115.625 79.865 116.395 ;
        RECT 80.965 116.265 81.135 116.995 ;
        RECT 82.280 116.825 82.450 117.155 ;
        RECT 82.620 116.995 82.950 117.375 ;
        RECT 81.305 116.445 81.655 116.815 ;
        RECT 80.965 116.225 81.385 116.265 ;
        RECT 80.035 116.055 81.385 116.225 ;
        RECT 80.035 115.895 80.285 116.055 ;
        RECT 80.795 115.625 81.045 115.885 ;
        RECT 79.675 115.375 81.045 115.625 ;
        RECT 77.605 115.085 77.845 115.375 ;
        RECT 78.645 115.295 78.815 115.375 ;
        RECT 78.045 114.825 78.465 115.205 ;
        RECT 78.645 115.045 79.275 115.295 ;
        RECT 79.745 114.825 80.075 115.205 ;
        RECT 80.245 115.085 80.415 115.375 ;
        RECT 81.215 115.210 81.385 116.055 ;
        RECT 81.835 115.885 82.055 116.755 ;
        RECT 82.280 116.635 82.975 116.825 ;
        RECT 81.555 115.505 82.055 115.885 ;
        RECT 82.225 115.835 82.635 116.455 ;
        RECT 82.805 115.665 82.975 116.635 ;
        RECT 82.280 115.495 82.975 115.665 ;
        RECT 80.595 114.825 80.975 115.205 ;
        RECT 81.215 115.040 82.045 115.210 ;
        RECT 82.280 114.995 82.450 115.495 ;
        RECT 82.620 114.825 82.950 115.325 ;
        RECT 83.165 114.995 83.390 117.115 ;
        RECT 83.560 116.995 83.890 117.375 ;
        RECT 84.060 116.825 84.230 117.115 ;
        RECT 84.865 117.035 85.120 117.195 ;
        RECT 84.780 116.865 85.120 117.035 ;
        RECT 85.300 116.915 85.585 117.375 ;
        RECT 83.565 116.655 84.230 116.825 ;
        RECT 84.865 116.665 85.120 116.865 ;
        RECT 83.565 115.665 83.795 116.655 ;
        RECT 83.965 115.835 84.315 116.485 ;
        RECT 84.865 115.805 85.045 116.665 ;
        RECT 85.765 116.465 86.015 117.115 ;
        RECT 85.215 116.135 86.015 116.465 ;
        RECT 83.565 115.495 84.230 115.665 ;
        RECT 83.560 114.825 83.890 115.325 ;
        RECT 84.060 114.995 84.230 115.495 ;
        RECT 84.865 115.135 85.120 115.805 ;
        RECT 85.300 114.825 85.585 115.625 ;
        RECT 85.765 115.545 86.015 116.135 ;
        RECT 86.215 116.780 86.535 117.110 ;
        RECT 86.715 116.895 87.375 117.375 ;
        RECT 87.575 116.985 88.425 117.155 ;
        RECT 86.215 115.885 86.405 116.780 ;
        RECT 86.725 116.455 87.385 116.725 ;
        RECT 87.055 116.395 87.385 116.455 ;
        RECT 86.575 116.225 86.905 116.285 ;
        RECT 87.575 116.225 87.745 116.985 ;
        RECT 88.985 116.915 89.305 117.375 ;
        RECT 89.505 116.735 89.755 117.165 ;
        RECT 90.045 116.935 90.455 117.375 ;
        RECT 90.625 116.995 91.640 117.195 ;
        RECT 87.915 116.565 89.165 116.735 ;
        RECT 87.915 116.445 88.245 116.565 ;
        RECT 86.575 116.055 88.475 116.225 ;
        RECT 86.215 115.715 88.135 115.885 ;
        RECT 86.215 115.695 86.535 115.715 ;
        RECT 85.765 115.035 86.095 115.545 ;
        RECT 86.365 115.085 86.535 115.695 ;
        RECT 88.305 115.545 88.475 116.055 ;
        RECT 88.645 115.985 88.825 116.395 ;
        RECT 88.995 115.805 89.165 116.565 ;
        RECT 86.705 114.825 87.035 115.515 ;
        RECT 87.265 115.375 88.475 115.545 ;
        RECT 88.645 115.495 89.165 115.805 ;
        RECT 89.335 116.395 89.755 116.735 ;
        RECT 90.045 116.395 90.455 116.725 ;
        RECT 89.335 115.625 89.525 116.395 ;
        RECT 90.625 116.265 90.795 116.995 ;
        RECT 91.940 116.825 92.110 117.155 ;
        RECT 92.280 116.995 92.610 117.375 ;
        RECT 90.965 116.445 91.315 116.815 ;
        RECT 90.625 116.225 91.045 116.265 ;
        RECT 89.695 116.055 91.045 116.225 ;
        RECT 89.695 115.895 89.945 116.055 ;
        RECT 90.455 115.625 90.705 115.885 ;
        RECT 89.335 115.375 90.705 115.625 ;
        RECT 87.265 115.085 87.505 115.375 ;
        RECT 88.305 115.295 88.475 115.375 ;
        RECT 87.705 114.825 88.125 115.205 ;
        RECT 88.305 115.045 88.935 115.295 ;
        RECT 89.405 114.825 89.735 115.205 ;
        RECT 89.905 115.085 90.075 115.375 ;
        RECT 90.875 115.210 91.045 116.055 ;
        RECT 91.495 115.885 91.715 116.755 ;
        RECT 91.940 116.635 92.635 116.825 ;
        RECT 91.215 115.505 91.715 115.885 ;
        RECT 91.885 115.835 92.295 116.455 ;
        RECT 92.465 115.665 92.635 116.635 ;
        RECT 91.940 115.495 92.635 115.665 ;
        RECT 90.255 114.825 90.635 115.205 ;
        RECT 90.875 115.040 91.705 115.210 ;
        RECT 91.940 114.995 92.110 115.495 ;
        RECT 92.280 114.825 92.610 115.325 ;
        RECT 92.825 114.995 93.050 117.115 ;
        RECT 93.220 116.995 93.550 117.375 ;
        RECT 93.720 116.825 93.890 117.115 ;
        RECT 93.225 116.655 93.890 116.825 ;
        RECT 93.225 115.665 93.455 116.655 ;
        RECT 95.345 116.565 95.590 117.170 ;
        RECT 95.810 116.840 96.320 117.375 ;
        RECT 93.625 115.835 93.975 116.485 ;
        RECT 95.070 116.395 96.300 116.565 ;
        RECT 93.225 115.495 93.890 115.665 ;
        RECT 93.220 114.825 93.550 115.325 ;
        RECT 93.720 114.995 93.890 115.495 ;
        RECT 95.070 115.585 95.410 116.395 ;
        RECT 95.580 115.830 96.330 116.020 ;
        RECT 95.070 115.175 95.585 115.585 ;
        RECT 95.820 114.825 95.990 115.585 ;
        RECT 96.160 115.165 96.330 115.830 ;
        RECT 96.500 115.845 96.690 117.205 ;
        RECT 96.860 117.035 97.135 117.205 ;
        RECT 96.860 116.865 97.140 117.035 ;
        RECT 96.860 116.045 97.135 116.865 ;
        RECT 97.325 116.840 97.855 117.205 ;
        RECT 98.280 116.975 98.610 117.375 ;
        RECT 97.680 116.805 97.855 116.840 ;
        RECT 97.340 115.845 97.510 116.645 ;
        RECT 96.500 115.675 97.510 115.845 ;
        RECT 97.680 116.635 98.610 116.805 ;
        RECT 98.780 116.635 99.035 117.205 ;
        RECT 99.210 116.650 99.500 117.375 ;
        RECT 100.045 116.695 100.300 117.195 ;
        RECT 100.480 116.915 100.765 117.375 ;
        RECT 99.960 116.665 100.300 116.695 ;
        RECT 97.680 115.505 97.850 116.635 ;
        RECT 98.440 116.465 98.610 116.635 ;
        RECT 96.725 115.335 97.850 115.505 ;
        RECT 98.020 116.135 98.215 116.465 ;
        RECT 98.440 116.135 98.695 116.465 ;
        RECT 98.020 115.165 98.190 116.135 ;
        RECT 98.865 115.965 99.035 116.635 ;
        RECT 99.960 116.525 100.225 116.665 ;
        RECT 96.160 114.995 98.190 115.165 ;
        RECT 98.360 114.825 98.530 115.965 ;
        RECT 98.700 114.995 99.035 115.965 ;
        RECT 99.210 114.825 99.500 115.990 ;
        RECT 100.045 115.805 100.225 116.525 ;
        RECT 100.945 116.465 101.195 117.115 ;
        RECT 100.395 116.135 101.195 116.465 ;
        RECT 100.045 115.135 100.300 115.805 ;
        RECT 100.480 114.825 100.765 115.625 ;
        RECT 100.945 115.545 101.195 116.135 ;
        RECT 101.395 116.780 101.715 117.110 ;
        RECT 101.895 116.895 102.555 117.375 ;
        RECT 102.755 116.985 103.605 117.155 ;
        RECT 101.395 115.885 101.585 116.780 ;
        RECT 101.905 116.455 102.565 116.725 ;
        RECT 102.235 116.395 102.565 116.455 ;
        RECT 101.755 116.225 102.085 116.285 ;
        RECT 102.755 116.225 102.925 116.985 ;
        RECT 104.165 116.915 104.485 117.375 ;
        RECT 104.685 116.735 104.935 117.165 ;
        RECT 105.225 116.935 105.635 117.375 ;
        RECT 105.805 116.995 106.820 117.195 ;
        RECT 103.095 116.565 104.345 116.735 ;
        RECT 103.095 116.445 103.425 116.565 ;
        RECT 101.755 116.055 103.655 116.225 ;
        RECT 101.395 115.715 103.315 115.885 ;
        RECT 101.395 115.695 101.715 115.715 ;
        RECT 100.945 115.035 101.275 115.545 ;
        RECT 101.545 115.085 101.715 115.695 ;
        RECT 103.485 115.545 103.655 116.055 ;
        RECT 103.825 115.985 104.005 116.395 ;
        RECT 104.175 115.805 104.345 116.565 ;
        RECT 101.885 114.825 102.215 115.515 ;
        RECT 102.445 115.375 103.655 115.545 ;
        RECT 103.825 115.495 104.345 115.805 ;
        RECT 104.515 116.395 104.935 116.735 ;
        RECT 105.225 116.395 105.635 116.725 ;
        RECT 104.515 115.625 104.705 116.395 ;
        RECT 105.805 116.265 105.975 116.995 ;
        RECT 107.120 116.825 107.290 117.155 ;
        RECT 107.460 116.995 107.790 117.375 ;
        RECT 106.145 116.445 106.495 116.815 ;
        RECT 105.805 116.225 106.225 116.265 ;
        RECT 104.875 116.055 106.225 116.225 ;
        RECT 104.875 115.895 105.125 116.055 ;
        RECT 105.635 115.625 105.885 115.885 ;
        RECT 104.515 115.375 105.885 115.625 ;
        RECT 102.445 115.085 102.685 115.375 ;
        RECT 103.485 115.295 103.655 115.375 ;
        RECT 102.885 114.825 103.305 115.205 ;
        RECT 103.485 115.045 104.115 115.295 ;
        RECT 104.585 114.825 104.915 115.205 ;
        RECT 105.085 115.085 105.255 115.375 ;
        RECT 106.055 115.210 106.225 116.055 ;
        RECT 106.675 115.885 106.895 116.755 ;
        RECT 107.120 116.635 107.815 116.825 ;
        RECT 106.395 115.505 106.895 115.885 ;
        RECT 107.065 115.835 107.475 116.455 ;
        RECT 107.645 115.665 107.815 116.635 ;
        RECT 107.120 115.495 107.815 115.665 ;
        RECT 105.435 114.825 105.815 115.205 ;
        RECT 106.055 115.040 106.885 115.210 ;
        RECT 107.120 114.995 107.290 115.495 ;
        RECT 107.460 114.825 107.790 115.325 ;
        RECT 108.005 114.995 108.230 117.115 ;
        RECT 108.400 116.995 108.730 117.375 ;
        RECT 108.900 116.825 109.070 117.115 ;
        RECT 108.405 116.655 109.070 116.825 ;
        RECT 108.405 115.665 108.635 116.655 ;
        RECT 109.330 116.605 111.000 117.375 ;
        RECT 111.170 116.625 112.380 117.375 ;
        RECT 108.805 115.835 109.155 116.485 ;
        RECT 109.330 115.915 110.080 116.435 ;
        RECT 110.250 116.085 111.000 116.605 ;
        RECT 111.170 115.915 111.690 116.455 ;
        RECT 111.860 116.085 112.380 116.625 ;
        RECT 108.405 115.495 109.070 115.665 ;
        RECT 108.400 114.825 108.730 115.325 ;
        RECT 108.900 114.995 109.070 115.495 ;
        RECT 109.330 114.825 111.000 115.915 ;
        RECT 111.170 114.825 112.380 115.915 ;
        RECT 18.165 114.655 112.465 114.825 ;
        RECT 18.250 113.565 19.460 114.655 ;
        RECT 19.940 113.815 20.110 114.655 ;
        RECT 20.320 113.645 20.570 114.485 ;
        RECT 20.780 113.815 20.950 114.655 ;
        RECT 21.120 113.645 21.410 114.485 ;
        RECT 18.250 112.855 18.770 113.395 ;
        RECT 18.940 113.025 19.460 113.565 ;
        RECT 19.685 113.475 21.410 113.645 ;
        RECT 21.620 113.595 21.790 114.655 ;
        RECT 22.085 114.275 22.415 114.655 ;
        RECT 22.595 114.105 22.765 114.395 ;
        RECT 22.935 114.195 23.185 114.655 ;
        RECT 21.965 113.935 22.765 114.105 ;
        RECT 23.355 114.145 24.225 114.485 ;
        RECT 19.685 112.925 20.095 113.475 ;
        RECT 21.965 113.315 22.135 113.935 ;
        RECT 23.355 113.765 23.525 114.145 ;
        RECT 24.460 114.025 24.630 114.485 ;
        RECT 24.800 114.195 25.170 114.655 ;
        RECT 25.465 114.055 25.635 114.395 ;
        RECT 25.805 114.225 26.135 114.655 ;
        RECT 26.370 114.055 26.540 114.395 ;
        RECT 22.305 113.595 23.525 113.765 ;
        RECT 23.695 113.685 24.155 113.975 ;
        RECT 24.460 113.855 25.020 114.025 ;
        RECT 25.465 113.885 26.540 114.055 ;
        RECT 26.710 114.155 27.390 114.485 ;
        RECT 27.605 114.155 27.855 114.485 ;
        RECT 28.025 114.195 28.275 114.655 ;
        RECT 24.850 113.715 25.020 113.855 ;
        RECT 23.695 113.675 24.660 113.685 ;
        RECT 23.355 113.505 23.525 113.595 ;
        RECT 23.985 113.515 24.660 113.675 ;
        RECT 21.965 113.305 22.310 113.315 ;
        RECT 20.280 113.095 22.310 113.305 ;
        RECT 18.250 112.105 19.460 112.855 ;
        RECT 19.685 112.755 21.450 112.925 ;
        RECT 19.940 112.105 20.110 112.575 ;
        RECT 20.280 112.275 20.610 112.755 ;
        RECT 20.780 112.105 20.950 112.575 ;
        RECT 21.120 112.275 21.450 112.755 ;
        RECT 21.620 112.105 21.790 112.915 ;
        RECT 21.985 112.840 22.310 113.095 ;
        RECT 21.990 112.485 22.310 112.840 ;
        RECT 22.480 113.055 23.020 113.425 ;
        RECT 23.355 113.335 23.760 113.505 ;
        RECT 22.480 112.655 22.720 113.055 ;
        RECT 23.200 112.885 23.420 113.165 ;
        RECT 22.890 112.715 23.420 112.885 ;
        RECT 22.890 112.485 23.060 112.715 ;
        RECT 23.590 112.555 23.760 113.335 ;
        RECT 23.930 112.725 24.280 113.345 ;
        RECT 24.450 112.725 24.660 113.515 ;
        RECT 24.850 113.545 26.350 113.715 ;
        RECT 24.850 112.855 25.020 113.545 ;
        RECT 26.710 113.375 26.880 114.155 ;
        RECT 27.685 114.025 27.855 114.155 ;
        RECT 25.190 113.205 26.880 113.375 ;
        RECT 27.050 113.595 27.515 113.985 ;
        RECT 27.685 113.855 28.080 114.025 ;
        RECT 25.190 113.025 25.360 113.205 ;
        RECT 21.990 112.315 23.060 112.485 ;
        RECT 23.230 112.105 23.420 112.545 ;
        RECT 23.590 112.275 24.540 112.555 ;
        RECT 24.850 112.465 25.110 112.855 ;
        RECT 25.530 112.785 26.320 113.035 ;
        RECT 24.760 112.295 25.110 112.465 ;
        RECT 25.320 112.105 25.650 112.565 ;
        RECT 26.525 112.495 26.695 113.205 ;
        RECT 27.050 113.005 27.220 113.595 ;
        RECT 26.865 112.785 27.220 113.005 ;
        RECT 27.390 112.785 27.740 113.405 ;
        RECT 27.910 112.495 28.080 113.855 ;
        RECT 28.445 113.685 28.770 114.470 ;
        RECT 28.250 112.635 28.710 113.685 ;
        RECT 26.525 112.325 27.380 112.495 ;
        RECT 27.585 112.325 28.080 112.495 ;
        RECT 28.250 112.105 28.580 112.465 ;
        RECT 28.940 112.365 29.110 114.485 ;
        RECT 29.280 114.155 29.610 114.655 ;
        RECT 29.780 113.985 30.035 114.485 ;
        RECT 29.285 113.815 30.035 113.985 ;
        RECT 29.285 112.825 29.515 113.815 ;
        RECT 29.685 112.995 30.035 113.645 ;
        RECT 30.210 113.565 31.880 114.655 ;
        RECT 32.140 113.725 32.310 114.485 ;
        RECT 32.490 113.895 32.820 114.655 ;
        RECT 30.210 113.045 30.960 113.565 ;
        RECT 32.140 113.555 32.805 113.725 ;
        RECT 32.990 113.580 33.260 114.485 ;
        RECT 32.635 113.410 32.805 113.555 ;
        RECT 31.130 112.875 31.880 113.395 ;
        RECT 32.070 113.005 32.400 113.375 ;
        RECT 32.635 113.080 32.920 113.410 ;
        RECT 29.285 112.655 30.035 112.825 ;
        RECT 29.280 112.105 29.610 112.485 ;
        RECT 29.780 112.365 30.035 112.655 ;
        RECT 30.210 112.105 31.880 112.875 ;
        RECT 32.635 112.825 32.805 113.080 ;
        RECT 32.140 112.655 32.805 112.825 ;
        RECT 33.090 112.780 33.260 113.580 ;
        RECT 33.470 113.515 33.700 114.655 ;
        RECT 33.870 113.505 34.200 114.485 ;
        RECT 34.370 113.515 34.580 114.655 ;
        RECT 33.450 113.095 33.780 113.345 ;
        RECT 32.140 112.275 32.310 112.655 ;
        RECT 32.490 112.105 32.820 112.485 ;
        RECT 33.000 112.275 33.260 112.780 ;
        RECT 33.470 112.105 33.700 112.925 ;
        RECT 33.950 112.905 34.200 113.505 ;
        RECT 34.810 113.490 35.100 114.655 ;
        RECT 35.730 113.580 36.000 114.485 ;
        RECT 36.170 113.895 36.500 114.655 ;
        RECT 36.680 113.725 36.850 114.485 ;
        RECT 33.870 112.275 34.200 112.905 ;
        RECT 34.370 112.105 34.580 112.925 ;
        RECT 34.810 112.105 35.100 112.830 ;
        RECT 35.730 112.780 35.900 113.580 ;
        RECT 36.185 113.555 36.850 113.725 ;
        RECT 37.110 113.565 40.620 114.655 ;
        RECT 36.185 113.410 36.355 113.555 ;
        RECT 36.070 113.080 36.355 113.410 ;
        RECT 36.185 112.825 36.355 113.080 ;
        RECT 36.590 113.005 36.920 113.375 ;
        RECT 37.110 113.045 38.800 113.565 ;
        RECT 40.830 113.515 41.060 114.655 ;
        RECT 41.230 113.505 41.560 114.485 ;
        RECT 41.730 113.515 41.940 114.655 ;
        RECT 42.170 113.895 42.685 114.305 ;
        RECT 42.920 113.895 43.090 114.655 ;
        RECT 43.260 114.315 45.290 114.485 ;
        RECT 38.970 112.875 40.620 113.395 ;
        RECT 40.810 113.095 41.140 113.345 ;
        RECT 35.730 112.275 35.990 112.780 ;
        RECT 36.185 112.655 36.850 112.825 ;
        RECT 36.170 112.105 36.500 112.485 ;
        RECT 36.680 112.275 36.850 112.655 ;
        RECT 37.110 112.105 40.620 112.875 ;
        RECT 40.830 112.105 41.060 112.925 ;
        RECT 41.310 112.905 41.560 113.505 ;
        RECT 42.170 113.085 42.510 113.895 ;
        RECT 43.260 113.650 43.430 114.315 ;
        RECT 43.825 113.975 44.950 114.145 ;
        RECT 42.680 113.460 43.430 113.650 ;
        RECT 43.600 113.635 44.610 113.805 ;
        RECT 41.230 112.275 41.560 112.905 ;
        RECT 41.730 112.105 41.940 112.925 ;
        RECT 42.170 112.915 43.400 113.085 ;
        RECT 42.445 112.310 42.690 112.915 ;
        RECT 42.910 112.105 43.420 112.640 ;
        RECT 43.600 112.275 43.790 113.635 ;
        RECT 43.960 112.955 44.235 113.435 ;
        RECT 43.960 112.785 44.240 112.955 ;
        RECT 44.440 112.835 44.610 113.635 ;
        RECT 44.780 112.845 44.950 113.975 ;
        RECT 45.120 113.345 45.290 114.315 ;
        RECT 45.460 113.515 45.630 114.655 ;
        RECT 45.800 113.515 46.135 114.485 ;
        RECT 45.120 113.015 45.315 113.345 ;
        RECT 45.540 113.015 45.795 113.345 ;
        RECT 45.540 112.845 45.710 113.015 ;
        RECT 45.965 112.845 46.135 113.515 ;
        RECT 43.960 112.275 44.235 112.785 ;
        RECT 44.780 112.675 45.710 112.845 ;
        RECT 44.780 112.640 44.955 112.675 ;
        RECT 44.425 112.275 44.955 112.640 ;
        RECT 45.380 112.105 45.710 112.505 ;
        RECT 45.880 112.275 46.135 112.845 ;
        RECT 46.310 113.580 46.580 114.485 ;
        RECT 46.750 113.895 47.080 114.655 ;
        RECT 47.260 113.725 47.430 114.485 ;
        RECT 46.310 112.780 46.480 113.580 ;
        RECT 46.765 113.555 47.430 113.725 ;
        RECT 48.150 113.565 50.740 114.655 ;
        RECT 50.915 114.220 56.260 114.655 ;
        RECT 46.765 113.410 46.935 113.555 ;
        RECT 46.650 113.080 46.935 113.410 ;
        RECT 46.765 112.825 46.935 113.080 ;
        RECT 47.170 113.005 47.500 113.375 ;
        RECT 48.150 113.045 49.360 113.565 ;
        RECT 49.530 112.875 50.740 113.395 ;
        RECT 52.505 112.970 52.855 114.220 ;
        RECT 56.470 113.515 56.700 114.655 ;
        RECT 56.870 113.505 57.200 114.485 ;
        RECT 57.370 113.515 57.580 114.655 ;
        RECT 58.360 113.725 58.530 114.485 ;
        RECT 58.710 113.895 59.040 114.655 ;
        RECT 58.360 113.555 59.025 113.725 ;
        RECT 59.210 113.580 59.480 114.485 ;
        RECT 46.310 112.275 46.570 112.780 ;
        RECT 46.765 112.655 47.430 112.825 ;
        RECT 46.750 112.105 47.080 112.485 ;
        RECT 47.260 112.275 47.430 112.655 ;
        RECT 48.150 112.105 50.740 112.875 ;
        RECT 54.335 112.650 54.675 113.480 ;
        RECT 56.450 113.095 56.780 113.345 ;
        RECT 50.915 112.105 56.260 112.650 ;
        RECT 56.470 112.105 56.700 112.925 ;
        RECT 56.950 112.905 57.200 113.505 ;
        RECT 58.855 113.410 59.025 113.555 ;
        RECT 58.290 113.005 58.620 113.375 ;
        RECT 58.855 113.080 59.140 113.410 ;
        RECT 56.870 112.275 57.200 112.905 ;
        RECT 57.370 112.105 57.580 112.925 ;
        RECT 58.855 112.825 59.025 113.080 ;
        RECT 58.360 112.655 59.025 112.825 ;
        RECT 59.310 112.780 59.480 113.580 ;
        RECT 60.570 113.490 60.860 114.655 ;
        RECT 61.490 113.565 63.160 114.655 ;
        RECT 63.335 114.220 68.680 114.655 ;
        RECT 61.490 113.045 62.240 113.565 ;
        RECT 62.410 112.875 63.160 113.395 ;
        RECT 64.925 112.970 65.275 114.220 ;
        RECT 68.910 113.515 69.120 114.655 ;
        RECT 69.290 113.505 69.620 114.485 ;
        RECT 69.790 113.515 70.020 114.655 ;
        RECT 70.690 113.565 72.360 114.655 ;
        RECT 72.535 114.220 77.880 114.655 ;
        RECT 58.360 112.275 58.530 112.655 ;
        RECT 58.710 112.105 59.040 112.485 ;
        RECT 59.220 112.275 59.480 112.780 ;
        RECT 60.570 112.105 60.860 112.830 ;
        RECT 61.490 112.105 63.160 112.875 ;
        RECT 66.755 112.650 67.095 113.480 ;
        RECT 63.335 112.105 68.680 112.650 ;
        RECT 68.910 112.105 69.120 112.925 ;
        RECT 69.290 112.905 69.540 113.505 ;
        RECT 69.710 113.095 70.040 113.345 ;
        RECT 70.690 113.045 71.440 113.565 ;
        RECT 69.290 112.275 69.620 112.905 ;
        RECT 69.790 112.105 70.020 112.925 ;
        RECT 71.610 112.875 72.360 113.395 ;
        RECT 74.125 112.970 74.475 114.220 ;
        RECT 78.090 113.515 78.320 114.655 ;
        RECT 78.490 113.505 78.820 114.485 ;
        RECT 78.990 113.515 79.200 114.655 ;
        RECT 79.980 113.725 80.150 114.485 ;
        RECT 80.330 113.895 80.660 114.655 ;
        RECT 79.980 113.555 80.645 113.725 ;
        RECT 80.830 113.580 81.100 114.485 ;
        RECT 70.690 112.105 72.360 112.875 ;
        RECT 75.955 112.650 76.295 113.480 ;
        RECT 78.070 113.095 78.400 113.345 ;
        RECT 72.535 112.105 77.880 112.650 ;
        RECT 78.090 112.105 78.320 112.925 ;
        RECT 78.570 112.905 78.820 113.505 ;
        RECT 80.475 113.410 80.645 113.555 ;
        RECT 79.910 113.005 80.240 113.375 ;
        RECT 80.475 113.080 80.760 113.410 ;
        RECT 78.490 112.275 78.820 112.905 ;
        RECT 78.990 112.105 79.200 112.925 ;
        RECT 80.475 112.825 80.645 113.080 ;
        RECT 79.980 112.655 80.645 112.825 ;
        RECT 80.930 112.780 81.100 113.580 ;
        RECT 81.310 113.515 81.540 114.655 ;
        RECT 81.710 113.505 82.040 114.485 ;
        RECT 82.210 113.515 82.420 114.655 ;
        RECT 82.650 113.565 86.160 114.655 ;
        RECT 81.290 113.095 81.620 113.345 ;
        RECT 79.980 112.275 80.150 112.655 ;
        RECT 80.330 112.105 80.660 112.485 ;
        RECT 80.840 112.275 81.100 112.780 ;
        RECT 81.310 112.105 81.540 112.925 ;
        RECT 81.790 112.905 82.040 113.505 ;
        RECT 82.650 113.045 84.340 113.565 ;
        RECT 86.330 113.490 86.620 114.655 ;
        RECT 86.790 113.565 88.460 114.655 ;
        RECT 88.720 113.725 88.890 114.485 ;
        RECT 89.070 113.895 89.400 114.655 ;
        RECT 81.710 112.275 82.040 112.905 ;
        RECT 82.210 112.105 82.420 112.925 ;
        RECT 84.510 112.875 86.160 113.395 ;
        RECT 86.790 113.045 87.540 113.565 ;
        RECT 88.720 113.555 89.385 113.725 ;
        RECT 89.570 113.580 89.840 114.485 ;
        RECT 90.935 114.220 96.280 114.655 ;
        RECT 89.215 113.410 89.385 113.555 ;
        RECT 87.710 112.875 88.460 113.395 ;
        RECT 88.650 113.005 88.980 113.375 ;
        RECT 89.215 113.080 89.500 113.410 ;
        RECT 82.650 112.105 86.160 112.875 ;
        RECT 86.330 112.105 86.620 112.830 ;
        RECT 86.790 112.105 88.460 112.875 ;
        RECT 89.215 112.825 89.385 113.080 ;
        RECT 88.720 112.655 89.385 112.825 ;
        RECT 89.670 112.780 89.840 113.580 ;
        RECT 92.525 112.970 92.875 114.220 ;
        RECT 96.450 113.580 96.720 114.485 ;
        RECT 96.890 113.895 97.220 114.655 ;
        RECT 97.400 113.725 97.570 114.485 ;
        RECT 88.720 112.275 88.890 112.655 ;
        RECT 89.070 112.105 89.400 112.485 ;
        RECT 89.580 112.275 89.840 112.780 ;
        RECT 94.355 112.650 94.695 113.480 ;
        RECT 96.450 112.780 96.620 113.580 ;
        RECT 96.905 113.555 97.570 113.725 ;
        RECT 98.290 113.565 99.960 114.655 ;
        RECT 100.135 114.220 105.480 114.655 ;
        RECT 105.655 114.220 111.000 114.655 ;
        RECT 96.905 113.410 97.075 113.555 ;
        RECT 96.790 113.080 97.075 113.410 ;
        RECT 96.905 112.825 97.075 113.080 ;
        RECT 97.310 113.005 97.640 113.375 ;
        RECT 98.290 113.045 99.040 113.565 ;
        RECT 99.210 112.875 99.960 113.395 ;
        RECT 101.725 112.970 102.075 114.220 ;
        RECT 90.935 112.105 96.280 112.650 ;
        RECT 96.450 112.275 96.710 112.780 ;
        RECT 96.905 112.655 97.570 112.825 ;
        RECT 96.890 112.105 97.220 112.485 ;
        RECT 97.400 112.275 97.570 112.655 ;
        RECT 98.290 112.105 99.960 112.875 ;
        RECT 103.555 112.650 103.895 113.480 ;
        RECT 107.245 112.970 107.595 114.220 ;
        RECT 111.170 113.565 112.380 114.655 ;
        RECT 109.075 112.650 109.415 113.480 ;
        RECT 111.170 113.025 111.690 113.565 ;
        RECT 111.860 112.855 112.380 113.395 ;
        RECT 100.135 112.105 105.480 112.650 ;
        RECT 105.655 112.105 111.000 112.650 ;
        RECT 111.170 112.105 112.380 112.855 ;
        RECT 18.165 111.935 112.465 112.105 ;
        RECT 18.250 111.185 19.460 111.935 ;
        RECT 18.250 110.645 18.770 111.185 ;
        RECT 20.090 111.165 21.760 111.935 ;
        RECT 21.930 111.210 22.220 111.935 ;
        RECT 22.395 111.390 27.740 111.935 ;
        RECT 18.940 110.475 19.460 111.015 ;
        RECT 18.250 109.385 19.460 110.475 ;
        RECT 20.090 110.475 20.840 110.995 ;
        RECT 21.010 110.645 21.760 111.165 ;
        RECT 20.090 109.385 21.760 110.475 ;
        RECT 21.930 109.385 22.220 110.550 ;
        RECT 23.985 109.820 24.335 111.070 ;
        RECT 25.815 110.560 26.155 111.390 ;
        RECT 27.910 111.260 28.170 111.765 ;
        RECT 28.350 111.555 28.680 111.935 ;
        RECT 28.860 111.385 29.030 111.765 ;
        RECT 27.910 110.460 28.080 111.260 ;
        RECT 28.365 111.215 29.030 111.385 ;
        RECT 29.840 111.385 30.010 111.765 ;
        RECT 30.190 111.555 30.520 111.935 ;
        RECT 29.840 111.215 30.505 111.385 ;
        RECT 30.700 111.260 30.960 111.765 ;
        RECT 31.440 111.465 31.610 111.935 ;
        RECT 31.780 111.285 32.110 111.765 ;
        RECT 32.280 111.465 32.450 111.935 ;
        RECT 32.620 111.285 32.950 111.765 ;
        RECT 28.365 110.960 28.535 111.215 ;
        RECT 28.250 110.630 28.535 110.960 ;
        RECT 28.770 110.665 29.100 111.035 ;
        RECT 29.770 110.665 30.100 111.035 ;
        RECT 30.335 110.960 30.505 111.215 ;
        RECT 28.365 110.485 28.535 110.630 ;
        RECT 30.335 110.630 30.620 110.960 ;
        RECT 30.335 110.485 30.505 110.630 ;
        RECT 22.395 109.385 27.740 109.820 ;
        RECT 27.910 109.555 28.180 110.460 ;
        RECT 28.365 110.315 29.030 110.485 ;
        RECT 28.350 109.385 28.680 110.145 ;
        RECT 28.860 109.555 29.030 110.315 ;
        RECT 29.840 110.315 30.505 110.485 ;
        RECT 30.790 110.460 30.960 111.260 ;
        RECT 29.840 109.555 30.010 110.315 ;
        RECT 30.190 109.385 30.520 110.145 ;
        RECT 30.690 109.555 30.960 110.460 ;
        RECT 31.185 111.115 32.950 111.285 ;
        RECT 33.120 111.125 33.290 111.935 ;
        RECT 33.490 111.555 34.560 111.725 ;
        RECT 33.490 111.200 33.810 111.555 ;
        RECT 31.185 110.565 31.595 111.115 ;
        RECT 33.485 110.945 33.810 111.200 ;
        RECT 31.780 110.735 33.810 110.945 ;
        RECT 33.465 110.725 33.810 110.735 ;
        RECT 33.980 110.985 34.220 111.385 ;
        RECT 34.390 111.325 34.560 111.555 ;
        RECT 34.730 111.495 34.920 111.935 ;
        RECT 35.090 111.485 36.040 111.765 ;
        RECT 36.260 111.575 36.610 111.745 ;
        RECT 34.390 111.155 34.920 111.325 ;
        RECT 31.185 110.395 32.910 110.565 ;
        RECT 31.440 109.385 31.610 110.225 ;
        RECT 31.820 109.555 32.070 110.395 ;
        RECT 32.280 109.385 32.450 110.225 ;
        RECT 32.620 109.555 32.910 110.395 ;
        RECT 33.120 109.385 33.290 110.445 ;
        RECT 33.465 110.105 33.635 110.725 ;
        RECT 33.980 110.615 34.520 110.985 ;
        RECT 34.700 110.875 34.920 111.155 ;
        RECT 35.090 110.705 35.260 111.485 ;
        RECT 34.855 110.535 35.260 110.705 ;
        RECT 35.430 110.695 35.780 111.315 ;
        RECT 34.855 110.445 35.025 110.535 ;
        RECT 35.950 110.525 36.160 111.315 ;
        RECT 33.805 110.275 35.025 110.445 ;
        RECT 35.485 110.365 36.160 110.525 ;
        RECT 33.465 109.935 34.265 110.105 ;
        RECT 33.585 109.385 33.915 109.765 ;
        RECT 34.095 109.645 34.265 109.935 ;
        RECT 34.855 109.895 35.025 110.275 ;
        RECT 35.195 110.355 36.160 110.365 ;
        RECT 36.350 111.185 36.610 111.575 ;
        RECT 36.820 111.475 37.150 111.935 ;
        RECT 38.025 111.545 38.880 111.715 ;
        RECT 39.085 111.545 39.580 111.715 ;
        RECT 39.750 111.575 40.080 111.935 ;
        RECT 36.350 110.495 36.520 111.185 ;
        RECT 36.690 110.835 36.860 111.015 ;
        RECT 37.030 111.005 37.820 111.255 ;
        RECT 38.025 110.835 38.195 111.545 ;
        RECT 38.365 111.035 38.720 111.255 ;
        RECT 36.690 110.665 38.380 110.835 ;
        RECT 35.195 110.065 35.655 110.355 ;
        RECT 36.350 110.325 37.850 110.495 ;
        RECT 36.350 110.185 36.520 110.325 ;
        RECT 35.960 110.015 36.520 110.185 ;
        RECT 34.435 109.385 34.685 109.845 ;
        RECT 34.855 109.555 35.725 109.895 ;
        RECT 35.960 109.555 36.130 110.015 ;
        RECT 36.965 109.985 38.040 110.155 ;
        RECT 36.300 109.385 36.670 109.845 ;
        RECT 36.965 109.645 37.135 109.985 ;
        RECT 37.305 109.385 37.635 109.815 ;
        RECT 37.870 109.645 38.040 109.985 ;
        RECT 38.210 109.885 38.380 110.665 ;
        RECT 38.550 110.445 38.720 111.035 ;
        RECT 38.890 110.635 39.240 111.255 ;
        RECT 38.550 110.055 39.015 110.445 ;
        RECT 39.410 110.185 39.580 111.545 ;
        RECT 39.750 110.355 40.210 111.405 ;
        RECT 39.185 110.015 39.580 110.185 ;
        RECT 39.185 109.885 39.355 110.015 ;
        RECT 38.210 109.555 38.890 109.885 ;
        RECT 39.105 109.555 39.355 109.885 ;
        RECT 39.525 109.385 39.775 109.845 ;
        RECT 39.945 109.570 40.270 110.355 ;
        RECT 40.440 109.555 40.610 111.675 ;
        RECT 40.780 111.555 41.110 111.935 ;
        RECT 41.280 111.385 41.535 111.675 ;
        RECT 40.785 111.215 41.535 111.385 ;
        RECT 42.630 111.260 42.890 111.765 ;
        RECT 43.070 111.555 43.400 111.935 ;
        RECT 43.580 111.385 43.750 111.765 ;
        RECT 40.785 110.225 41.015 111.215 ;
        RECT 41.185 110.395 41.535 111.045 ;
        RECT 42.630 110.460 42.800 111.260 ;
        RECT 43.085 111.215 43.750 111.385 ;
        RECT 44.010 111.260 44.270 111.765 ;
        RECT 44.450 111.555 44.780 111.935 ;
        RECT 44.960 111.385 45.130 111.765 ;
        RECT 43.085 110.960 43.255 111.215 ;
        RECT 42.970 110.630 43.255 110.960 ;
        RECT 43.490 110.665 43.820 111.035 ;
        RECT 43.085 110.485 43.255 110.630 ;
        RECT 40.785 110.055 41.535 110.225 ;
        RECT 40.780 109.385 41.110 109.885 ;
        RECT 41.280 109.555 41.535 110.055 ;
        RECT 42.630 109.555 42.900 110.460 ;
        RECT 43.085 110.315 43.750 110.485 ;
        RECT 43.070 109.385 43.400 110.145 ;
        RECT 43.580 109.555 43.750 110.315 ;
        RECT 44.010 110.460 44.180 111.260 ;
        RECT 44.465 111.215 45.130 111.385 ;
        RECT 45.480 111.385 45.650 111.765 ;
        RECT 45.830 111.555 46.160 111.935 ;
        RECT 45.480 111.215 46.145 111.385 ;
        RECT 46.340 111.260 46.600 111.765 ;
        RECT 44.465 110.960 44.635 111.215 ;
        RECT 44.350 110.630 44.635 110.960 ;
        RECT 44.870 110.665 45.200 111.035 ;
        RECT 45.410 110.665 45.740 111.035 ;
        RECT 45.975 110.960 46.145 111.215 ;
        RECT 44.465 110.485 44.635 110.630 ;
        RECT 45.975 110.630 46.260 110.960 ;
        RECT 45.975 110.485 46.145 110.630 ;
        RECT 44.010 109.555 44.280 110.460 ;
        RECT 44.465 110.315 45.130 110.485 ;
        RECT 44.450 109.385 44.780 110.145 ;
        RECT 44.960 109.555 45.130 110.315 ;
        RECT 45.480 110.315 46.145 110.485 ;
        RECT 46.430 110.460 46.600 111.260 ;
        RECT 47.690 111.210 47.980 111.935 ;
        RECT 48.150 111.165 50.740 111.935 ;
        RECT 45.480 109.555 45.650 110.315 ;
        RECT 45.830 109.385 46.160 110.145 ;
        RECT 46.330 109.555 46.600 110.460 ;
        RECT 47.690 109.385 47.980 110.550 ;
        RECT 48.150 110.475 49.360 110.995 ;
        RECT 49.530 110.645 50.740 111.165 ;
        RECT 50.910 111.260 51.170 111.765 ;
        RECT 51.350 111.555 51.680 111.935 ;
        RECT 51.860 111.385 52.030 111.765 ;
        RECT 48.150 109.385 50.740 110.475 ;
        RECT 50.910 110.460 51.080 111.260 ;
        RECT 51.365 111.215 52.030 111.385 ;
        RECT 51.365 110.960 51.535 111.215 ;
        RECT 52.750 111.165 54.420 111.935 ;
        RECT 51.250 110.630 51.535 110.960 ;
        RECT 51.770 110.665 52.100 111.035 ;
        RECT 51.365 110.485 51.535 110.630 ;
        RECT 50.910 109.555 51.180 110.460 ;
        RECT 51.365 110.315 52.030 110.485 ;
        RECT 51.350 109.385 51.680 110.145 ;
        RECT 51.860 109.555 52.030 110.315 ;
        RECT 52.750 110.475 53.500 110.995 ;
        RECT 53.670 110.645 54.420 111.165 ;
        RECT 54.740 111.135 55.070 111.935 ;
        RECT 55.240 111.285 55.410 111.765 ;
        RECT 55.580 111.455 55.910 111.935 ;
        RECT 56.080 111.285 56.250 111.765 ;
        RECT 56.500 111.455 56.740 111.935 ;
        RECT 56.920 111.285 57.090 111.765 ;
        RECT 57.660 111.465 57.830 111.935 ;
        RECT 58.000 111.285 58.330 111.765 ;
        RECT 58.500 111.465 58.670 111.935 ;
        RECT 58.840 111.285 59.170 111.765 ;
        RECT 55.240 111.115 56.250 111.285 ;
        RECT 56.455 111.115 57.090 111.285 ;
        RECT 57.405 111.115 59.170 111.285 ;
        RECT 59.340 111.125 59.510 111.935 ;
        RECT 59.710 111.555 60.780 111.725 ;
        RECT 59.710 111.200 60.030 111.555 ;
        RECT 55.240 110.575 55.735 111.115 ;
        RECT 56.455 110.945 56.625 111.115 ;
        RECT 56.125 110.775 56.625 110.945 ;
        RECT 52.750 109.385 54.420 110.475 ;
        RECT 54.740 109.385 55.070 110.535 ;
        RECT 55.240 110.405 56.250 110.575 ;
        RECT 55.240 109.555 55.410 110.405 ;
        RECT 55.580 109.385 55.910 110.185 ;
        RECT 56.080 109.555 56.250 110.405 ;
        RECT 56.455 110.535 56.625 110.775 ;
        RECT 56.795 110.705 57.175 110.945 ;
        RECT 57.405 110.565 57.815 111.115 ;
        RECT 59.705 110.945 60.030 111.200 ;
        RECT 58.000 110.735 60.030 110.945 ;
        RECT 59.685 110.725 60.030 110.735 ;
        RECT 60.200 110.985 60.440 111.385 ;
        RECT 60.610 111.325 60.780 111.555 ;
        RECT 60.950 111.495 61.140 111.935 ;
        RECT 61.310 111.485 62.260 111.765 ;
        RECT 62.480 111.575 62.830 111.745 ;
        RECT 60.610 111.155 61.140 111.325 ;
        RECT 56.455 110.365 57.170 110.535 ;
        RECT 57.405 110.395 59.130 110.565 ;
        RECT 56.430 109.385 56.670 110.185 ;
        RECT 56.840 109.555 57.170 110.365 ;
        RECT 57.660 109.385 57.830 110.225 ;
        RECT 58.040 109.555 58.290 110.395 ;
        RECT 58.500 109.385 58.670 110.225 ;
        RECT 58.840 109.555 59.130 110.395 ;
        RECT 59.340 109.385 59.510 110.445 ;
        RECT 59.685 110.105 59.855 110.725 ;
        RECT 60.200 110.615 60.740 110.985 ;
        RECT 60.920 110.875 61.140 111.155 ;
        RECT 61.310 110.705 61.480 111.485 ;
        RECT 61.075 110.535 61.480 110.705 ;
        RECT 61.650 110.695 62.000 111.315 ;
        RECT 61.075 110.445 61.245 110.535 ;
        RECT 62.170 110.525 62.380 111.315 ;
        RECT 60.025 110.275 61.245 110.445 ;
        RECT 61.705 110.365 62.380 110.525 ;
        RECT 59.685 109.935 60.485 110.105 ;
        RECT 59.805 109.385 60.135 109.765 ;
        RECT 60.315 109.645 60.485 109.935 ;
        RECT 61.075 109.895 61.245 110.275 ;
        RECT 61.415 110.355 62.380 110.365 ;
        RECT 62.570 111.185 62.830 111.575 ;
        RECT 63.040 111.475 63.370 111.935 ;
        RECT 64.245 111.545 65.100 111.715 ;
        RECT 65.305 111.545 65.800 111.715 ;
        RECT 65.970 111.575 66.300 111.935 ;
        RECT 62.570 110.495 62.740 111.185 ;
        RECT 62.910 110.835 63.080 111.015 ;
        RECT 63.250 111.005 64.040 111.255 ;
        RECT 64.245 110.835 64.415 111.545 ;
        RECT 64.585 111.035 64.940 111.255 ;
        RECT 62.910 110.665 64.600 110.835 ;
        RECT 61.415 110.065 61.875 110.355 ;
        RECT 62.570 110.325 64.070 110.495 ;
        RECT 62.570 110.185 62.740 110.325 ;
        RECT 62.180 110.015 62.740 110.185 ;
        RECT 60.655 109.385 60.905 109.845 ;
        RECT 61.075 109.555 61.945 109.895 ;
        RECT 62.180 109.555 62.350 110.015 ;
        RECT 63.185 109.985 64.260 110.155 ;
        RECT 62.520 109.385 62.890 109.845 ;
        RECT 63.185 109.645 63.355 109.985 ;
        RECT 63.525 109.385 63.855 109.815 ;
        RECT 64.090 109.645 64.260 109.985 ;
        RECT 64.430 109.885 64.600 110.665 ;
        RECT 64.770 110.445 64.940 111.035 ;
        RECT 65.110 110.635 65.460 111.255 ;
        RECT 64.770 110.055 65.235 110.445 ;
        RECT 65.630 110.185 65.800 111.545 ;
        RECT 65.970 110.355 66.430 111.405 ;
        RECT 65.405 110.015 65.800 110.185 ;
        RECT 65.405 109.885 65.575 110.015 ;
        RECT 64.430 109.555 65.110 109.885 ;
        RECT 65.325 109.555 65.575 109.885 ;
        RECT 65.745 109.385 65.995 109.845 ;
        RECT 66.165 109.570 66.490 110.355 ;
        RECT 66.660 109.555 66.830 111.675 ;
        RECT 67.000 111.555 67.330 111.935 ;
        RECT 67.500 111.385 67.755 111.675 ;
        RECT 67.005 111.215 67.755 111.385 ;
        RECT 67.005 110.225 67.235 111.215 ;
        RECT 67.930 111.185 69.140 111.935 ;
        RECT 67.405 110.395 67.755 111.045 ;
        RECT 67.930 110.475 68.450 111.015 ;
        RECT 68.620 110.645 69.140 111.185 ;
        RECT 69.310 111.260 69.570 111.765 ;
        RECT 69.750 111.555 70.080 111.935 ;
        RECT 70.260 111.385 70.430 111.765 ;
        RECT 67.005 110.055 67.755 110.225 ;
        RECT 67.000 109.385 67.330 109.885 ;
        RECT 67.500 109.555 67.755 110.055 ;
        RECT 67.930 109.385 69.140 110.475 ;
        RECT 69.310 110.460 69.480 111.260 ;
        RECT 69.765 111.215 70.430 111.385 ;
        RECT 70.780 111.285 70.950 111.765 ;
        RECT 71.130 111.455 71.370 111.935 ;
        RECT 71.620 111.285 71.790 111.765 ;
        RECT 71.960 111.455 72.290 111.935 ;
        RECT 72.460 111.285 72.630 111.765 ;
        RECT 69.765 110.960 69.935 111.215 ;
        RECT 70.780 111.115 71.415 111.285 ;
        RECT 71.620 111.115 72.630 111.285 ;
        RECT 72.800 111.135 73.130 111.935 ;
        RECT 73.450 111.210 73.740 111.935 ;
        RECT 73.910 111.165 77.420 111.935 ;
        RECT 77.680 111.385 77.850 111.765 ;
        RECT 78.030 111.555 78.360 111.935 ;
        RECT 77.680 111.215 78.345 111.385 ;
        RECT 78.540 111.260 78.800 111.765 ;
        RECT 69.650 110.630 69.935 110.960 ;
        RECT 70.170 110.665 70.500 111.035 ;
        RECT 71.245 110.945 71.415 111.115 ;
        RECT 70.695 110.705 71.075 110.945 ;
        RECT 71.245 110.775 71.745 110.945 ;
        RECT 69.765 110.485 69.935 110.630 ;
        RECT 71.245 110.535 71.415 110.775 ;
        RECT 72.135 110.575 72.630 111.115 ;
        RECT 69.310 109.555 69.580 110.460 ;
        RECT 69.765 110.315 70.430 110.485 ;
        RECT 69.750 109.385 70.080 110.145 ;
        RECT 70.260 109.555 70.430 110.315 ;
        RECT 70.700 110.365 71.415 110.535 ;
        RECT 71.620 110.405 72.630 110.575 ;
        RECT 70.700 109.555 71.030 110.365 ;
        RECT 71.200 109.385 71.440 110.185 ;
        RECT 71.620 109.555 71.790 110.405 ;
        RECT 71.960 109.385 72.290 110.185 ;
        RECT 72.460 109.555 72.630 110.405 ;
        RECT 72.800 109.385 73.130 110.535 ;
        RECT 73.450 109.385 73.740 110.550 ;
        RECT 73.910 110.475 75.600 110.995 ;
        RECT 75.770 110.645 77.420 111.165 ;
        RECT 77.610 110.665 77.940 111.035 ;
        RECT 78.175 110.960 78.345 111.215 ;
        RECT 78.175 110.630 78.460 110.960 ;
        RECT 78.175 110.485 78.345 110.630 ;
        RECT 73.910 109.385 77.420 110.475 ;
        RECT 77.680 110.315 78.345 110.485 ;
        RECT 78.630 110.460 78.800 111.260 ;
        RECT 79.430 111.165 82.940 111.935 ;
        RECT 83.200 111.385 83.370 111.765 ;
        RECT 83.550 111.555 83.880 111.935 ;
        RECT 83.200 111.215 83.865 111.385 ;
        RECT 84.060 111.260 84.320 111.765 ;
        RECT 77.680 109.555 77.850 110.315 ;
        RECT 78.030 109.385 78.360 110.145 ;
        RECT 78.530 109.555 78.800 110.460 ;
        RECT 79.430 110.475 81.120 110.995 ;
        RECT 81.290 110.645 82.940 111.165 ;
        RECT 83.130 110.665 83.460 111.035 ;
        RECT 83.695 110.960 83.865 111.215 ;
        RECT 83.695 110.630 83.980 110.960 ;
        RECT 83.695 110.485 83.865 110.630 ;
        RECT 79.430 109.385 82.940 110.475 ;
        RECT 83.200 110.315 83.865 110.485 ;
        RECT 84.150 110.460 84.320 111.260 ;
        RECT 84.490 111.165 86.160 111.935 ;
        RECT 83.200 109.555 83.370 110.315 ;
        RECT 83.550 109.385 83.880 110.145 ;
        RECT 84.050 109.555 84.320 110.460 ;
        RECT 84.490 110.475 85.240 110.995 ;
        RECT 85.410 110.645 86.160 111.165 ;
        RECT 86.370 111.115 86.600 111.935 ;
        RECT 86.770 111.135 87.100 111.765 ;
        RECT 86.350 110.695 86.680 110.945 ;
        RECT 86.850 110.535 87.100 111.135 ;
        RECT 87.270 111.115 87.480 111.935 ;
        RECT 87.710 111.185 88.920 111.935 ;
        RECT 89.180 111.385 89.350 111.765 ;
        RECT 89.530 111.555 89.860 111.935 ;
        RECT 89.180 111.215 89.845 111.385 ;
        RECT 90.040 111.260 90.300 111.765 ;
        RECT 84.490 109.385 86.160 110.475 ;
        RECT 86.370 109.385 86.600 110.525 ;
        RECT 86.770 109.555 87.100 110.535 ;
        RECT 87.270 109.385 87.480 110.525 ;
        RECT 87.710 110.475 88.230 111.015 ;
        RECT 88.400 110.645 88.920 111.185 ;
        RECT 89.110 110.665 89.440 111.035 ;
        RECT 89.675 110.960 89.845 111.215 ;
        RECT 89.675 110.630 89.960 110.960 ;
        RECT 89.675 110.485 89.845 110.630 ;
        RECT 87.710 109.385 88.920 110.475 ;
        RECT 89.180 110.315 89.845 110.485 ;
        RECT 90.130 110.460 90.300 111.260 ;
        RECT 91.450 111.115 91.660 111.935 ;
        RECT 91.830 111.135 92.160 111.765 ;
        RECT 91.830 110.535 92.080 111.135 ;
        RECT 92.330 111.115 92.560 111.935 ;
        RECT 93.780 111.385 93.950 111.765 ;
        RECT 94.130 111.555 94.460 111.935 ;
        RECT 93.780 111.215 94.445 111.385 ;
        RECT 94.640 111.260 94.900 111.765 ;
        RECT 92.250 110.695 92.580 110.945 ;
        RECT 93.710 110.665 94.040 111.035 ;
        RECT 94.275 110.960 94.445 111.215 ;
        RECT 94.275 110.630 94.560 110.960 ;
        RECT 89.180 109.555 89.350 110.315 ;
        RECT 89.530 109.385 89.860 110.145 ;
        RECT 90.030 109.555 90.300 110.460 ;
        RECT 91.450 109.385 91.660 110.525 ;
        RECT 91.830 109.555 92.160 110.535 ;
        RECT 92.330 109.385 92.560 110.525 ;
        RECT 94.275 110.485 94.445 110.630 ;
        RECT 93.780 110.315 94.445 110.485 ;
        RECT 94.730 110.460 94.900 111.260 ;
        RECT 95.070 111.165 97.660 111.935 ;
        RECT 93.780 109.555 93.950 110.315 ;
        RECT 94.130 109.385 94.460 110.145 ;
        RECT 94.630 109.555 94.900 110.460 ;
        RECT 95.070 110.475 96.280 110.995 ;
        RECT 96.450 110.645 97.660 111.165 ;
        RECT 97.870 111.115 98.100 111.935 ;
        RECT 98.270 111.135 98.600 111.765 ;
        RECT 97.850 110.695 98.180 110.945 ;
        RECT 98.350 110.535 98.600 111.135 ;
        RECT 98.770 111.115 98.980 111.935 ;
        RECT 99.210 111.210 99.500 111.935 ;
        RECT 100.220 111.385 100.390 111.765 ;
        RECT 100.570 111.555 100.900 111.935 ;
        RECT 100.220 111.215 100.885 111.385 ;
        RECT 101.080 111.260 101.340 111.765 ;
        RECT 100.150 110.665 100.480 111.035 ;
        RECT 100.715 110.960 100.885 111.215 ;
        RECT 100.715 110.630 101.000 110.960 ;
        RECT 95.070 109.385 97.660 110.475 ;
        RECT 97.870 109.385 98.100 110.525 ;
        RECT 98.270 109.555 98.600 110.535 ;
        RECT 98.770 109.385 98.980 110.525 ;
        RECT 99.210 109.385 99.500 110.550 ;
        RECT 100.715 110.485 100.885 110.630 ;
        RECT 100.220 110.315 100.885 110.485 ;
        RECT 101.170 110.460 101.340 111.260 ;
        RECT 101.970 111.165 104.560 111.935 ;
        RECT 100.220 109.555 100.390 110.315 ;
        RECT 100.570 109.385 100.900 110.145 ;
        RECT 101.070 109.555 101.340 110.460 ;
        RECT 101.970 110.475 103.180 110.995 ;
        RECT 103.350 110.645 104.560 111.165 ;
        RECT 104.770 111.115 105.000 111.935 ;
        RECT 105.170 111.135 105.500 111.765 ;
        RECT 104.750 110.695 105.080 110.945 ;
        RECT 105.250 110.535 105.500 111.135 ;
        RECT 105.670 111.115 105.880 111.935 ;
        RECT 106.200 111.385 106.370 111.765 ;
        RECT 106.550 111.555 106.880 111.935 ;
        RECT 106.200 111.215 106.865 111.385 ;
        RECT 107.060 111.260 107.320 111.765 ;
        RECT 106.130 110.665 106.460 111.035 ;
        RECT 106.695 110.960 106.865 111.215 ;
        RECT 101.970 109.385 104.560 110.475 ;
        RECT 104.770 109.385 105.000 110.525 ;
        RECT 105.170 109.555 105.500 110.535 ;
        RECT 106.695 110.630 106.980 110.960 ;
        RECT 105.670 109.385 105.880 110.525 ;
        RECT 106.695 110.485 106.865 110.630 ;
        RECT 106.200 110.315 106.865 110.485 ;
        RECT 107.150 110.460 107.320 111.260 ;
        RECT 107.580 111.385 107.750 111.765 ;
        RECT 107.930 111.555 108.260 111.935 ;
        RECT 107.580 111.215 108.245 111.385 ;
        RECT 108.440 111.260 108.700 111.765 ;
        RECT 107.510 110.665 107.840 111.035 ;
        RECT 108.075 110.960 108.245 111.215 ;
        RECT 108.075 110.630 108.360 110.960 ;
        RECT 108.075 110.485 108.245 110.630 ;
        RECT 106.200 109.555 106.370 110.315 ;
        RECT 106.550 109.385 106.880 110.145 ;
        RECT 107.050 109.555 107.320 110.460 ;
        RECT 107.580 110.315 108.245 110.485 ;
        RECT 108.530 110.460 108.700 111.260 ;
        RECT 107.580 109.555 107.750 110.315 ;
        RECT 107.930 109.385 108.260 110.145 ;
        RECT 108.430 109.555 108.700 110.460 ;
        RECT 109.790 111.260 110.050 111.765 ;
        RECT 110.230 111.555 110.560 111.935 ;
        RECT 110.740 111.385 110.910 111.765 ;
        RECT 109.790 110.460 109.970 111.260 ;
        RECT 110.245 111.215 110.910 111.385 ;
        RECT 110.245 110.960 110.415 111.215 ;
        RECT 111.170 111.185 112.380 111.935 ;
        RECT 110.140 110.630 110.415 110.960 ;
        RECT 110.640 110.665 110.980 111.035 ;
        RECT 110.245 110.485 110.415 110.630 ;
        RECT 109.790 109.555 110.060 110.460 ;
        RECT 110.245 110.315 110.920 110.485 ;
        RECT 110.230 109.385 110.560 110.145 ;
        RECT 110.740 109.555 110.920 110.315 ;
        RECT 111.170 110.475 111.690 111.015 ;
        RECT 111.860 110.645 112.380 111.185 ;
        RECT 111.170 109.385 112.380 110.475 ;
        RECT 18.165 109.215 112.465 109.385 ;
        RECT 18.250 108.125 19.460 109.215 ;
        RECT 18.250 107.415 18.770 107.955 ;
        RECT 18.940 107.585 19.460 108.125 ;
        RECT 20.090 108.125 22.680 109.215 ;
        RECT 20.090 107.605 21.300 108.125 ;
        RECT 22.910 108.075 23.120 109.215 ;
        RECT 23.290 108.065 23.620 109.045 ;
        RECT 23.790 108.075 24.020 109.215 ;
        RECT 24.540 108.375 24.710 109.215 ;
        RECT 24.920 108.205 25.170 109.045 ;
        RECT 25.380 108.375 25.550 109.215 ;
        RECT 25.720 108.205 26.010 109.045 ;
        RECT 21.470 107.435 22.680 107.955 ;
        RECT 18.250 106.665 19.460 107.415 ;
        RECT 20.090 106.665 22.680 107.435 ;
        RECT 22.910 106.665 23.120 107.485 ;
        RECT 23.290 107.465 23.540 108.065 ;
        RECT 24.285 108.035 26.010 108.205 ;
        RECT 26.220 108.155 26.390 109.215 ;
        RECT 26.685 108.835 27.015 109.215 ;
        RECT 27.195 108.665 27.365 108.955 ;
        RECT 27.535 108.755 27.785 109.215 ;
        RECT 26.565 108.495 27.365 108.665 ;
        RECT 27.955 108.705 28.825 109.045 ;
        RECT 23.710 107.655 24.040 107.905 ;
        RECT 24.285 107.485 24.695 108.035 ;
        RECT 26.565 107.875 26.735 108.495 ;
        RECT 27.955 108.325 28.125 108.705 ;
        RECT 29.060 108.585 29.230 109.045 ;
        RECT 29.400 108.755 29.770 109.215 ;
        RECT 30.065 108.615 30.235 108.955 ;
        RECT 30.405 108.785 30.735 109.215 ;
        RECT 30.970 108.615 31.140 108.955 ;
        RECT 26.905 108.155 28.125 108.325 ;
        RECT 28.295 108.245 28.755 108.535 ;
        RECT 29.060 108.415 29.620 108.585 ;
        RECT 30.065 108.445 31.140 108.615 ;
        RECT 31.310 108.715 31.990 109.045 ;
        RECT 32.205 108.715 32.455 109.045 ;
        RECT 32.625 108.755 32.875 109.215 ;
        RECT 29.450 108.275 29.620 108.415 ;
        RECT 28.295 108.235 29.260 108.245 ;
        RECT 27.955 108.065 28.125 108.155 ;
        RECT 28.585 108.075 29.260 108.235 ;
        RECT 26.565 107.865 26.910 107.875 ;
        RECT 24.880 107.655 26.910 107.865 ;
        RECT 23.290 106.835 23.620 107.465 ;
        RECT 23.790 106.665 24.020 107.485 ;
        RECT 24.285 107.315 26.050 107.485 ;
        RECT 24.540 106.665 24.710 107.135 ;
        RECT 24.880 106.835 25.210 107.315 ;
        RECT 25.380 106.665 25.550 107.135 ;
        RECT 25.720 106.835 26.050 107.315 ;
        RECT 26.220 106.665 26.390 107.475 ;
        RECT 26.585 107.400 26.910 107.655 ;
        RECT 26.590 107.045 26.910 107.400 ;
        RECT 27.080 107.615 27.620 107.985 ;
        RECT 27.955 107.895 28.360 108.065 ;
        RECT 27.080 107.215 27.320 107.615 ;
        RECT 27.800 107.445 28.020 107.725 ;
        RECT 27.490 107.275 28.020 107.445 ;
        RECT 27.490 107.045 27.660 107.275 ;
        RECT 28.190 107.115 28.360 107.895 ;
        RECT 28.530 107.285 28.880 107.905 ;
        RECT 29.050 107.285 29.260 108.075 ;
        RECT 29.450 108.105 30.950 108.275 ;
        RECT 29.450 107.415 29.620 108.105 ;
        RECT 31.310 107.935 31.480 108.715 ;
        RECT 32.285 108.585 32.455 108.715 ;
        RECT 29.790 107.765 31.480 107.935 ;
        RECT 31.650 108.155 32.115 108.545 ;
        RECT 32.285 108.415 32.680 108.585 ;
        RECT 29.790 107.585 29.960 107.765 ;
        RECT 26.590 106.875 27.660 107.045 ;
        RECT 27.830 106.665 28.020 107.105 ;
        RECT 28.190 106.835 29.140 107.115 ;
        RECT 29.450 107.025 29.710 107.415 ;
        RECT 30.130 107.345 30.920 107.595 ;
        RECT 29.360 106.855 29.710 107.025 ;
        RECT 29.920 106.665 30.250 107.125 ;
        RECT 31.125 107.055 31.295 107.765 ;
        RECT 31.650 107.565 31.820 108.155 ;
        RECT 31.465 107.345 31.820 107.565 ;
        RECT 31.990 107.345 32.340 107.965 ;
        RECT 32.510 107.055 32.680 108.415 ;
        RECT 33.045 108.245 33.370 109.030 ;
        RECT 32.850 107.195 33.310 108.245 ;
        RECT 31.125 106.885 31.980 107.055 ;
        RECT 32.185 106.885 32.680 107.055 ;
        RECT 32.850 106.665 33.180 107.025 ;
        RECT 33.540 106.925 33.710 109.045 ;
        RECT 33.880 108.715 34.210 109.215 ;
        RECT 34.380 108.545 34.635 109.045 ;
        RECT 33.885 108.375 34.635 108.545 ;
        RECT 33.885 107.385 34.115 108.375 ;
        RECT 34.285 107.555 34.635 108.205 ;
        RECT 34.810 108.050 35.100 109.215 ;
        RECT 36.190 108.140 36.460 109.045 ;
        RECT 36.630 108.455 36.960 109.215 ;
        RECT 37.140 108.285 37.310 109.045 ;
        RECT 37.880 108.375 38.050 109.215 ;
        RECT 33.885 107.215 34.635 107.385 ;
        RECT 33.880 106.665 34.210 107.045 ;
        RECT 34.380 106.925 34.635 107.215 ;
        RECT 34.810 106.665 35.100 107.390 ;
        RECT 36.190 107.340 36.360 108.140 ;
        RECT 36.645 108.115 37.310 108.285 ;
        RECT 38.260 108.205 38.510 109.045 ;
        RECT 38.720 108.375 38.890 109.215 ;
        RECT 39.060 108.205 39.350 109.045 ;
        RECT 36.645 107.970 36.815 108.115 ;
        RECT 36.530 107.640 36.815 107.970 ;
        RECT 37.625 108.035 39.350 108.205 ;
        RECT 39.560 108.155 39.730 109.215 ;
        RECT 40.025 108.835 40.355 109.215 ;
        RECT 40.535 108.665 40.705 108.955 ;
        RECT 40.875 108.755 41.125 109.215 ;
        RECT 39.905 108.495 40.705 108.665 ;
        RECT 41.295 108.705 42.165 109.045 ;
        RECT 36.645 107.385 36.815 107.640 ;
        RECT 37.050 107.565 37.380 107.935 ;
        RECT 37.625 107.485 38.035 108.035 ;
        RECT 39.905 107.875 40.075 108.495 ;
        RECT 41.295 108.325 41.465 108.705 ;
        RECT 42.400 108.585 42.570 109.045 ;
        RECT 42.740 108.755 43.110 109.215 ;
        RECT 43.405 108.615 43.575 108.955 ;
        RECT 43.745 108.785 44.075 109.215 ;
        RECT 44.310 108.615 44.480 108.955 ;
        RECT 40.245 108.155 41.465 108.325 ;
        RECT 41.635 108.245 42.095 108.535 ;
        RECT 42.400 108.415 42.960 108.585 ;
        RECT 43.405 108.445 44.480 108.615 ;
        RECT 44.650 108.715 45.330 109.045 ;
        RECT 45.545 108.715 45.795 109.045 ;
        RECT 45.965 108.755 46.215 109.215 ;
        RECT 42.790 108.275 42.960 108.415 ;
        RECT 41.635 108.235 42.600 108.245 ;
        RECT 41.295 108.065 41.465 108.155 ;
        RECT 41.925 108.075 42.600 108.235 ;
        RECT 39.905 107.865 40.250 107.875 ;
        RECT 38.220 107.655 40.250 107.865 ;
        RECT 36.190 106.835 36.450 107.340 ;
        RECT 36.645 107.215 37.310 107.385 ;
        RECT 37.625 107.315 39.390 107.485 ;
        RECT 36.630 106.665 36.960 107.045 ;
        RECT 37.140 106.835 37.310 107.215 ;
        RECT 37.880 106.665 38.050 107.135 ;
        RECT 38.220 106.835 38.550 107.315 ;
        RECT 38.720 106.665 38.890 107.135 ;
        RECT 39.060 106.835 39.390 107.315 ;
        RECT 39.560 106.665 39.730 107.475 ;
        RECT 39.925 107.400 40.250 107.655 ;
        RECT 39.930 107.045 40.250 107.400 ;
        RECT 40.420 107.615 40.960 107.985 ;
        RECT 41.295 107.895 41.700 108.065 ;
        RECT 40.420 107.215 40.660 107.615 ;
        RECT 41.140 107.445 41.360 107.725 ;
        RECT 40.830 107.275 41.360 107.445 ;
        RECT 40.830 107.045 41.000 107.275 ;
        RECT 41.530 107.115 41.700 107.895 ;
        RECT 41.870 107.285 42.220 107.905 ;
        RECT 42.390 107.285 42.600 108.075 ;
        RECT 42.790 108.105 44.290 108.275 ;
        RECT 42.790 107.415 42.960 108.105 ;
        RECT 44.650 107.935 44.820 108.715 ;
        RECT 45.625 108.585 45.795 108.715 ;
        RECT 43.130 107.765 44.820 107.935 ;
        RECT 44.990 108.155 45.455 108.545 ;
        RECT 45.625 108.415 46.020 108.585 ;
        RECT 43.130 107.585 43.300 107.765 ;
        RECT 39.930 106.875 41.000 107.045 ;
        RECT 41.170 106.665 41.360 107.105 ;
        RECT 41.530 106.835 42.480 107.115 ;
        RECT 42.790 107.025 43.050 107.415 ;
        RECT 43.470 107.345 44.260 107.595 ;
        RECT 42.700 106.855 43.050 107.025 ;
        RECT 43.260 106.665 43.590 107.125 ;
        RECT 44.465 107.055 44.635 107.765 ;
        RECT 44.990 107.565 45.160 108.155 ;
        RECT 44.805 107.345 45.160 107.565 ;
        RECT 45.330 107.345 45.680 107.965 ;
        RECT 45.850 107.055 46.020 108.415 ;
        RECT 46.385 108.245 46.710 109.030 ;
        RECT 46.190 107.195 46.650 108.245 ;
        RECT 44.465 106.885 45.320 107.055 ;
        RECT 45.525 106.885 46.020 107.055 ;
        RECT 46.190 106.665 46.520 107.025 ;
        RECT 46.880 106.925 47.050 109.045 ;
        RECT 47.220 108.715 47.550 109.215 ;
        RECT 47.720 108.545 47.975 109.045 ;
        RECT 47.225 108.375 47.975 108.545 ;
        RECT 49.380 108.375 49.550 109.215 ;
        RECT 47.225 107.385 47.455 108.375 ;
        RECT 49.760 108.205 50.010 109.045 ;
        RECT 50.220 108.375 50.390 109.215 ;
        RECT 50.560 108.205 50.850 109.045 ;
        RECT 47.625 107.555 47.975 108.205 ;
        RECT 49.125 108.035 50.850 108.205 ;
        RECT 51.060 108.155 51.230 109.215 ;
        RECT 51.525 108.835 51.855 109.215 ;
        RECT 52.035 108.665 52.205 108.955 ;
        RECT 52.375 108.755 52.625 109.215 ;
        RECT 51.405 108.495 52.205 108.665 ;
        RECT 52.795 108.705 53.665 109.045 ;
        RECT 49.125 107.485 49.535 108.035 ;
        RECT 51.405 107.875 51.575 108.495 ;
        RECT 52.795 108.325 52.965 108.705 ;
        RECT 53.900 108.585 54.070 109.045 ;
        RECT 54.240 108.755 54.610 109.215 ;
        RECT 54.905 108.615 55.075 108.955 ;
        RECT 55.245 108.785 55.575 109.215 ;
        RECT 55.810 108.615 55.980 108.955 ;
        RECT 51.745 108.155 52.965 108.325 ;
        RECT 53.135 108.245 53.595 108.535 ;
        RECT 53.900 108.415 54.460 108.585 ;
        RECT 54.905 108.445 55.980 108.615 ;
        RECT 56.150 108.715 56.830 109.045 ;
        RECT 57.045 108.715 57.295 109.045 ;
        RECT 57.465 108.755 57.715 109.215 ;
        RECT 54.290 108.275 54.460 108.415 ;
        RECT 53.135 108.235 54.100 108.245 ;
        RECT 52.795 108.065 52.965 108.155 ;
        RECT 53.425 108.075 54.100 108.235 ;
        RECT 51.405 107.865 51.750 107.875 ;
        RECT 49.720 107.655 51.750 107.865 ;
        RECT 47.225 107.215 47.975 107.385 ;
        RECT 49.125 107.315 50.890 107.485 ;
        RECT 47.220 106.665 47.550 107.045 ;
        RECT 47.720 106.925 47.975 107.215 ;
        RECT 49.380 106.665 49.550 107.135 ;
        RECT 49.720 106.835 50.050 107.315 ;
        RECT 50.220 106.665 50.390 107.135 ;
        RECT 50.560 106.835 50.890 107.315 ;
        RECT 51.060 106.665 51.230 107.475 ;
        RECT 51.425 107.400 51.750 107.655 ;
        RECT 51.430 107.045 51.750 107.400 ;
        RECT 51.920 107.615 52.460 107.985 ;
        RECT 52.795 107.895 53.200 108.065 ;
        RECT 51.920 107.215 52.160 107.615 ;
        RECT 52.640 107.445 52.860 107.725 ;
        RECT 52.330 107.275 52.860 107.445 ;
        RECT 52.330 107.045 52.500 107.275 ;
        RECT 53.030 107.115 53.200 107.895 ;
        RECT 53.370 107.285 53.720 107.905 ;
        RECT 53.890 107.285 54.100 108.075 ;
        RECT 54.290 108.105 55.790 108.275 ;
        RECT 54.290 107.415 54.460 108.105 ;
        RECT 56.150 107.935 56.320 108.715 ;
        RECT 57.125 108.585 57.295 108.715 ;
        RECT 54.630 107.765 56.320 107.935 ;
        RECT 56.490 108.155 56.955 108.545 ;
        RECT 57.125 108.415 57.520 108.585 ;
        RECT 54.630 107.585 54.800 107.765 ;
        RECT 51.430 106.875 52.500 107.045 ;
        RECT 52.670 106.665 52.860 107.105 ;
        RECT 53.030 106.835 53.980 107.115 ;
        RECT 54.290 107.025 54.550 107.415 ;
        RECT 54.970 107.345 55.760 107.595 ;
        RECT 54.200 106.855 54.550 107.025 ;
        RECT 54.760 106.665 55.090 107.125 ;
        RECT 55.965 107.055 56.135 107.765 ;
        RECT 56.490 107.565 56.660 108.155 ;
        RECT 56.305 107.345 56.660 107.565 ;
        RECT 56.830 107.345 57.180 107.965 ;
        RECT 57.350 107.055 57.520 108.415 ;
        RECT 57.885 108.245 58.210 109.030 ;
        RECT 57.690 107.195 58.150 108.245 ;
        RECT 55.965 106.885 56.820 107.055 ;
        RECT 57.025 106.885 57.520 107.055 ;
        RECT 57.690 106.665 58.020 107.025 ;
        RECT 58.380 106.925 58.550 109.045 ;
        RECT 58.720 108.715 59.050 109.215 ;
        RECT 59.220 108.545 59.475 109.045 ;
        RECT 58.725 108.375 59.475 108.545 ;
        RECT 58.725 107.385 58.955 108.375 ;
        RECT 59.125 107.555 59.475 108.205 ;
        RECT 60.570 108.050 60.860 109.215 ;
        RECT 61.120 108.285 61.290 109.045 ;
        RECT 61.470 108.455 61.800 109.215 ;
        RECT 61.120 108.115 61.785 108.285 ;
        RECT 61.970 108.140 62.240 109.045 ;
        RECT 61.615 107.970 61.785 108.115 ;
        RECT 61.050 107.565 61.380 107.935 ;
        RECT 61.615 107.640 61.900 107.970 ;
        RECT 58.725 107.215 59.475 107.385 ;
        RECT 58.720 106.665 59.050 107.045 ;
        RECT 59.220 106.925 59.475 107.215 ;
        RECT 60.570 106.665 60.860 107.390 ;
        RECT 61.615 107.385 61.785 107.640 ;
        RECT 61.120 107.215 61.785 107.385 ;
        RECT 62.070 107.340 62.240 108.140 ;
        RECT 63.420 108.285 63.590 109.045 ;
        RECT 63.770 108.455 64.100 109.215 ;
        RECT 63.420 108.115 64.085 108.285 ;
        RECT 64.270 108.140 64.540 109.045 ;
        RECT 65.020 108.375 65.190 109.215 ;
        RECT 65.400 108.205 65.650 109.045 ;
        RECT 65.860 108.375 66.030 109.215 ;
        RECT 66.200 108.205 66.490 109.045 ;
        RECT 63.915 107.970 64.085 108.115 ;
        RECT 63.350 107.565 63.680 107.935 ;
        RECT 63.915 107.640 64.200 107.970 ;
        RECT 63.915 107.385 64.085 107.640 ;
        RECT 61.120 106.835 61.290 107.215 ;
        RECT 61.470 106.665 61.800 107.045 ;
        RECT 61.980 106.835 62.240 107.340 ;
        RECT 63.420 107.215 64.085 107.385 ;
        RECT 64.370 107.340 64.540 108.140 ;
        RECT 63.420 106.835 63.590 107.215 ;
        RECT 63.770 106.665 64.100 107.045 ;
        RECT 64.280 106.835 64.540 107.340 ;
        RECT 64.765 108.035 66.490 108.205 ;
        RECT 66.700 108.155 66.870 109.215 ;
        RECT 67.165 108.835 67.495 109.215 ;
        RECT 67.675 108.665 67.845 108.955 ;
        RECT 68.015 108.755 68.265 109.215 ;
        RECT 67.045 108.495 67.845 108.665 ;
        RECT 68.435 108.705 69.305 109.045 ;
        RECT 64.765 107.485 65.175 108.035 ;
        RECT 67.045 107.875 67.215 108.495 ;
        RECT 68.435 108.325 68.605 108.705 ;
        RECT 69.540 108.585 69.710 109.045 ;
        RECT 69.880 108.755 70.250 109.215 ;
        RECT 70.545 108.615 70.715 108.955 ;
        RECT 70.885 108.785 71.215 109.215 ;
        RECT 71.450 108.615 71.620 108.955 ;
        RECT 67.385 108.155 68.605 108.325 ;
        RECT 68.775 108.245 69.235 108.535 ;
        RECT 69.540 108.415 70.100 108.585 ;
        RECT 70.545 108.445 71.620 108.615 ;
        RECT 71.790 108.715 72.470 109.045 ;
        RECT 72.685 108.715 72.935 109.045 ;
        RECT 73.105 108.755 73.355 109.215 ;
        RECT 69.930 108.275 70.100 108.415 ;
        RECT 68.775 108.235 69.740 108.245 ;
        RECT 68.435 108.065 68.605 108.155 ;
        RECT 69.065 108.075 69.740 108.235 ;
        RECT 67.045 107.865 67.390 107.875 ;
        RECT 65.360 107.655 67.390 107.865 ;
        RECT 64.765 107.315 66.530 107.485 ;
        RECT 65.020 106.665 65.190 107.135 ;
        RECT 65.360 106.835 65.690 107.315 ;
        RECT 65.860 106.665 66.030 107.135 ;
        RECT 66.200 106.835 66.530 107.315 ;
        RECT 66.700 106.665 66.870 107.475 ;
        RECT 67.065 107.400 67.390 107.655 ;
        RECT 67.070 107.045 67.390 107.400 ;
        RECT 67.560 107.615 68.100 107.985 ;
        RECT 68.435 107.895 68.840 108.065 ;
        RECT 67.560 107.215 67.800 107.615 ;
        RECT 68.280 107.445 68.500 107.725 ;
        RECT 67.970 107.275 68.500 107.445 ;
        RECT 67.970 107.045 68.140 107.275 ;
        RECT 68.670 107.115 68.840 107.895 ;
        RECT 69.010 107.285 69.360 107.905 ;
        RECT 69.530 107.285 69.740 108.075 ;
        RECT 69.930 108.105 71.430 108.275 ;
        RECT 69.930 107.415 70.100 108.105 ;
        RECT 71.790 107.935 71.960 108.715 ;
        RECT 72.765 108.585 72.935 108.715 ;
        RECT 70.270 107.765 71.960 107.935 ;
        RECT 72.130 108.155 72.595 108.545 ;
        RECT 72.765 108.415 73.160 108.585 ;
        RECT 70.270 107.585 70.440 107.765 ;
        RECT 67.070 106.875 68.140 107.045 ;
        RECT 68.310 106.665 68.500 107.105 ;
        RECT 68.670 106.835 69.620 107.115 ;
        RECT 69.930 107.025 70.190 107.415 ;
        RECT 70.610 107.345 71.400 107.595 ;
        RECT 69.840 106.855 70.190 107.025 ;
        RECT 70.400 106.665 70.730 107.125 ;
        RECT 71.605 107.055 71.775 107.765 ;
        RECT 72.130 107.565 72.300 108.155 ;
        RECT 71.945 107.345 72.300 107.565 ;
        RECT 72.470 107.345 72.820 107.965 ;
        RECT 72.990 107.055 73.160 108.415 ;
        RECT 73.525 108.245 73.850 109.030 ;
        RECT 73.330 107.195 73.790 108.245 ;
        RECT 71.605 106.885 72.460 107.055 ;
        RECT 72.665 106.885 73.160 107.055 ;
        RECT 73.330 106.665 73.660 107.025 ;
        RECT 74.020 106.925 74.190 109.045 ;
        RECT 74.360 108.715 74.690 109.215 ;
        RECT 74.860 108.545 75.115 109.045 ;
        RECT 74.365 108.375 75.115 108.545 ;
        RECT 76.060 108.375 76.230 109.215 ;
        RECT 74.365 107.385 74.595 108.375 ;
        RECT 76.440 108.205 76.690 109.045 ;
        RECT 76.900 108.375 77.070 109.215 ;
        RECT 77.240 108.205 77.530 109.045 ;
        RECT 74.765 107.555 75.115 108.205 ;
        RECT 75.805 108.035 77.530 108.205 ;
        RECT 77.740 108.155 77.910 109.215 ;
        RECT 78.205 108.835 78.535 109.215 ;
        RECT 78.715 108.665 78.885 108.955 ;
        RECT 79.055 108.755 79.305 109.215 ;
        RECT 78.085 108.495 78.885 108.665 ;
        RECT 79.475 108.705 80.345 109.045 ;
        RECT 75.805 107.485 76.215 108.035 ;
        RECT 78.085 107.875 78.255 108.495 ;
        RECT 79.475 108.325 79.645 108.705 ;
        RECT 80.580 108.585 80.750 109.045 ;
        RECT 80.920 108.755 81.290 109.215 ;
        RECT 81.585 108.615 81.755 108.955 ;
        RECT 81.925 108.785 82.255 109.215 ;
        RECT 82.490 108.615 82.660 108.955 ;
        RECT 78.425 108.155 79.645 108.325 ;
        RECT 79.815 108.245 80.275 108.535 ;
        RECT 80.580 108.415 81.140 108.585 ;
        RECT 81.585 108.445 82.660 108.615 ;
        RECT 82.830 108.715 83.510 109.045 ;
        RECT 83.725 108.715 83.975 109.045 ;
        RECT 84.145 108.755 84.395 109.215 ;
        RECT 80.970 108.275 81.140 108.415 ;
        RECT 79.815 108.235 80.780 108.245 ;
        RECT 79.475 108.065 79.645 108.155 ;
        RECT 80.105 108.075 80.780 108.235 ;
        RECT 78.085 107.865 78.430 107.875 ;
        RECT 76.400 107.655 78.430 107.865 ;
        RECT 74.365 107.215 75.115 107.385 ;
        RECT 75.805 107.315 77.570 107.485 ;
        RECT 74.360 106.665 74.690 107.045 ;
        RECT 74.860 106.925 75.115 107.215 ;
        RECT 76.060 106.665 76.230 107.135 ;
        RECT 76.400 106.835 76.730 107.315 ;
        RECT 76.900 106.665 77.070 107.135 ;
        RECT 77.240 106.835 77.570 107.315 ;
        RECT 77.740 106.665 77.910 107.475 ;
        RECT 78.105 107.400 78.430 107.655 ;
        RECT 78.110 107.045 78.430 107.400 ;
        RECT 78.600 107.615 79.140 107.985 ;
        RECT 79.475 107.895 79.880 108.065 ;
        RECT 78.600 107.215 78.840 107.615 ;
        RECT 79.320 107.445 79.540 107.725 ;
        RECT 79.010 107.275 79.540 107.445 ;
        RECT 79.010 107.045 79.180 107.275 ;
        RECT 79.710 107.115 79.880 107.895 ;
        RECT 80.050 107.285 80.400 107.905 ;
        RECT 80.570 107.285 80.780 108.075 ;
        RECT 80.970 108.105 82.470 108.275 ;
        RECT 80.970 107.415 81.140 108.105 ;
        RECT 82.830 107.935 83.000 108.715 ;
        RECT 83.805 108.585 83.975 108.715 ;
        RECT 81.310 107.765 83.000 107.935 ;
        RECT 83.170 108.155 83.635 108.545 ;
        RECT 83.805 108.415 84.200 108.585 ;
        RECT 81.310 107.585 81.480 107.765 ;
        RECT 78.110 106.875 79.180 107.045 ;
        RECT 79.350 106.665 79.540 107.105 ;
        RECT 79.710 106.835 80.660 107.115 ;
        RECT 80.970 107.025 81.230 107.415 ;
        RECT 81.650 107.345 82.440 107.595 ;
        RECT 80.880 106.855 81.230 107.025 ;
        RECT 81.440 106.665 81.770 107.125 ;
        RECT 82.645 107.055 82.815 107.765 ;
        RECT 83.170 107.565 83.340 108.155 ;
        RECT 82.985 107.345 83.340 107.565 ;
        RECT 83.510 107.345 83.860 107.965 ;
        RECT 84.030 107.055 84.200 108.415 ;
        RECT 84.565 108.245 84.890 109.030 ;
        RECT 84.370 107.195 84.830 108.245 ;
        RECT 82.645 106.885 83.500 107.055 ;
        RECT 83.705 106.885 84.200 107.055 ;
        RECT 84.370 106.665 84.700 107.025 ;
        RECT 85.060 106.925 85.230 109.045 ;
        RECT 85.400 108.715 85.730 109.215 ;
        RECT 85.900 108.545 86.155 109.045 ;
        RECT 85.405 108.375 86.155 108.545 ;
        RECT 85.405 107.385 85.635 108.375 ;
        RECT 85.805 107.555 86.155 108.205 ;
        RECT 86.330 108.050 86.620 109.215 ;
        RECT 87.100 108.375 87.270 109.215 ;
        RECT 87.480 108.205 87.730 109.045 ;
        RECT 87.940 108.375 88.110 109.215 ;
        RECT 88.280 108.205 88.570 109.045 ;
        RECT 86.845 108.035 88.570 108.205 ;
        RECT 88.780 108.155 88.950 109.215 ;
        RECT 89.245 108.835 89.575 109.215 ;
        RECT 89.755 108.665 89.925 108.955 ;
        RECT 90.095 108.755 90.345 109.215 ;
        RECT 89.125 108.495 89.925 108.665 ;
        RECT 90.515 108.705 91.385 109.045 ;
        RECT 86.845 107.485 87.255 108.035 ;
        RECT 89.125 107.875 89.295 108.495 ;
        RECT 90.515 108.325 90.685 108.705 ;
        RECT 91.620 108.585 91.790 109.045 ;
        RECT 91.960 108.755 92.330 109.215 ;
        RECT 92.625 108.615 92.795 108.955 ;
        RECT 92.965 108.785 93.295 109.215 ;
        RECT 93.530 108.615 93.700 108.955 ;
        RECT 89.465 108.155 90.685 108.325 ;
        RECT 90.855 108.245 91.315 108.535 ;
        RECT 91.620 108.415 92.180 108.585 ;
        RECT 92.625 108.445 93.700 108.615 ;
        RECT 93.870 108.715 94.550 109.045 ;
        RECT 94.765 108.715 95.015 109.045 ;
        RECT 95.185 108.755 95.435 109.215 ;
        RECT 92.010 108.275 92.180 108.415 ;
        RECT 90.855 108.235 91.820 108.245 ;
        RECT 90.515 108.065 90.685 108.155 ;
        RECT 91.145 108.075 91.820 108.235 ;
        RECT 89.125 107.865 89.470 107.875 ;
        RECT 87.440 107.655 89.470 107.865 ;
        RECT 85.405 107.215 86.155 107.385 ;
        RECT 85.400 106.665 85.730 107.045 ;
        RECT 85.900 106.925 86.155 107.215 ;
        RECT 86.330 106.665 86.620 107.390 ;
        RECT 86.845 107.315 88.610 107.485 ;
        RECT 87.100 106.665 87.270 107.135 ;
        RECT 87.440 106.835 87.770 107.315 ;
        RECT 87.940 106.665 88.110 107.135 ;
        RECT 88.280 106.835 88.610 107.315 ;
        RECT 88.780 106.665 88.950 107.475 ;
        RECT 89.145 107.400 89.470 107.655 ;
        RECT 89.150 107.045 89.470 107.400 ;
        RECT 89.640 107.615 90.180 107.985 ;
        RECT 90.515 107.895 90.920 108.065 ;
        RECT 89.640 107.215 89.880 107.615 ;
        RECT 90.360 107.445 90.580 107.725 ;
        RECT 90.050 107.275 90.580 107.445 ;
        RECT 90.050 107.045 90.220 107.275 ;
        RECT 90.750 107.115 90.920 107.895 ;
        RECT 91.090 107.285 91.440 107.905 ;
        RECT 91.610 107.285 91.820 108.075 ;
        RECT 92.010 108.105 93.510 108.275 ;
        RECT 92.010 107.415 92.180 108.105 ;
        RECT 93.870 107.935 94.040 108.715 ;
        RECT 94.845 108.585 95.015 108.715 ;
        RECT 92.350 107.765 94.040 107.935 ;
        RECT 94.210 108.155 94.675 108.545 ;
        RECT 94.845 108.415 95.240 108.585 ;
        RECT 92.350 107.585 92.520 107.765 ;
        RECT 89.150 106.875 90.220 107.045 ;
        RECT 90.390 106.665 90.580 107.105 ;
        RECT 90.750 106.835 91.700 107.115 ;
        RECT 92.010 107.025 92.270 107.415 ;
        RECT 92.690 107.345 93.480 107.595 ;
        RECT 91.920 106.855 92.270 107.025 ;
        RECT 92.480 106.665 92.810 107.125 ;
        RECT 93.685 107.055 93.855 107.765 ;
        RECT 94.210 107.565 94.380 108.155 ;
        RECT 94.025 107.345 94.380 107.565 ;
        RECT 94.550 107.345 94.900 107.965 ;
        RECT 95.070 107.055 95.240 108.415 ;
        RECT 95.605 108.245 95.930 109.030 ;
        RECT 95.410 107.195 95.870 108.245 ;
        RECT 93.685 106.885 94.540 107.055 ;
        RECT 94.745 106.885 95.240 107.055 ;
        RECT 95.410 106.665 95.740 107.025 ;
        RECT 96.100 106.925 96.270 109.045 ;
        RECT 96.440 108.715 96.770 109.215 ;
        RECT 96.940 108.545 97.195 109.045 ;
        RECT 96.445 108.375 97.195 108.545 ;
        RECT 96.445 107.385 96.675 108.375 ;
        RECT 96.845 107.555 97.195 108.205 ;
        RECT 97.370 108.140 97.640 109.045 ;
        RECT 97.810 108.455 98.140 109.215 ;
        RECT 98.320 108.285 98.490 109.045 ;
        RECT 96.445 107.215 97.195 107.385 ;
        RECT 96.440 106.665 96.770 107.045 ;
        RECT 96.940 106.925 97.195 107.215 ;
        RECT 97.370 107.340 97.540 108.140 ;
        RECT 97.825 108.115 98.490 108.285 ;
        RECT 97.825 107.970 97.995 108.115 ;
        RECT 98.810 108.075 99.020 109.215 ;
        RECT 97.710 107.640 97.995 107.970 ;
        RECT 99.190 108.065 99.520 109.045 ;
        RECT 99.690 108.075 99.920 109.215 ;
        RECT 100.900 108.375 101.070 109.215 ;
        RECT 101.280 108.205 101.530 109.045 ;
        RECT 101.740 108.375 101.910 109.215 ;
        RECT 102.080 108.205 102.370 109.045 ;
        RECT 97.825 107.385 97.995 107.640 ;
        RECT 98.230 107.565 98.560 107.935 ;
        RECT 97.370 106.835 97.630 107.340 ;
        RECT 97.825 107.215 98.490 107.385 ;
        RECT 97.810 106.665 98.140 107.045 ;
        RECT 98.320 106.835 98.490 107.215 ;
        RECT 98.810 106.665 99.020 107.485 ;
        RECT 99.190 107.465 99.440 108.065 ;
        RECT 100.645 108.035 102.370 108.205 ;
        RECT 102.580 108.155 102.750 109.215 ;
        RECT 103.045 108.835 103.375 109.215 ;
        RECT 103.555 108.665 103.725 108.955 ;
        RECT 103.895 108.755 104.145 109.215 ;
        RECT 102.925 108.495 103.725 108.665 ;
        RECT 104.315 108.705 105.185 109.045 ;
        RECT 99.610 107.655 99.940 107.905 ;
        RECT 100.645 107.485 101.055 108.035 ;
        RECT 102.925 107.875 103.095 108.495 ;
        RECT 104.315 108.325 104.485 108.705 ;
        RECT 105.420 108.585 105.590 109.045 ;
        RECT 105.760 108.755 106.130 109.215 ;
        RECT 106.425 108.615 106.595 108.955 ;
        RECT 106.765 108.785 107.095 109.215 ;
        RECT 107.330 108.615 107.500 108.955 ;
        RECT 103.265 108.155 104.485 108.325 ;
        RECT 104.655 108.245 105.115 108.535 ;
        RECT 105.420 108.415 105.980 108.585 ;
        RECT 106.425 108.445 107.500 108.615 ;
        RECT 107.670 108.715 108.350 109.045 ;
        RECT 108.565 108.715 108.815 109.045 ;
        RECT 108.985 108.755 109.235 109.215 ;
        RECT 105.810 108.275 105.980 108.415 ;
        RECT 104.655 108.235 105.620 108.245 ;
        RECT 104.315 108.065 104.485 108.155 ;
        RECT 104.945 108.075 105.620 108.235 ;
        RECT 102.925 107.865 103.270 107.875 ;
        RECT 101.240 107.655 103.270 107.865 ;
        RECT 99.190 106.835 99.520 107.465 ;
        RECT 99.690 106.665 99.920 107.485 ;
        RECT 100.645 107.315 102.410 107.485 ;
        RECT 100.900 106.665 101.070 107.135 ;
        RECT 101.240 106.835 101.570 107.315 ;
        RECT 101.740 106.665 101.910 107.135 ;
        RECT 102.080 106.835 102.410 107.315 ;
        RECT 102.580 106.665 102.750 107.475 ;
        RECT 102.945 107.400 103.270 107.655 ;
        RECT 102.950 107.045 103.270 107.400 ;
        RECT 103.440 107.615 103.980 107.985 ;
        RECT 104.315 107.895 104.720 108.065 ;
        RECT 103.440 107.215 103.680 107.615 ;
        RECT 104.160 107.445 104.380 107.725 ;
        RECT 103.850 107.275 104.380 107.445 ;
        RECT 103.850 107.045 104.020 107.275 ;
        RECT 104.550 107.115 104.720 107.895 ;
        RECT 104.890 107.285 105.240 107.905 ;
        RECT 105.410 107.285 105.620 108.075 ;
        RECT 105.810 108.105 107.310 108.275 ;
        RECT 105.810 107.415 105.980 108.105 ;
        RECT 107.670 107.935 107.840 108.715 ;
        RECT 108.645 108.585 108.815 108.715 ;
        RECT 106.150 107.765 107.840 107.935 ;
        RECT 108.010 108.155 108.475 108.545 ;
        RECT 108.645 108.415 109.040 108.585 ;
        RECT 106.150 107.585 106.320 107.765 ;
        RECT 102.950 106.875 104.020 107.045 ;
        RECT 104.190 106.665 104.380 107.105 ;
        RECT 104.550 106.835 105.500 107.115 ;
        RECT 105.810 107.025 106.070 107.415 ;
        RECT 106.490 107.345 107.280 107.595 ;
        RECT 105.720 106.855 106.070 107.025 ;
        RECT 106.280 106.665 106.610 107.125 ;
        RECT 107.485 107.055 107.655 107.765 ;
        RECT 108.010 107.565 108.180 108.155 ;
        RECT 107.825 107.345 108.180 107.565 ;
        RECT 108.350 107.345 108.700 107.965 ;
        RECT 108.870 107.055 109.040 108.415 ;
        RECT 109.405 108.245 109.730 109.030 ;
        RECT 109.210 107.195 109.670 108.245 ;
        RECT 107.485 106.885 108.340 107.055 ;
        RECT 108.545 106.885 109.040 107.055 ;
        RECT 109.210 106.665 109.540 107.025 ;
        RECT 109.900 106.925 110.070 109.045 ;
        RECT 110.240 108.715 110.570 109.215 ;
        RECT 110.740 108.545 110.995 109.045 ;
        RECT 110.245 108.375 110.995 108.545 ;
        RECT 110.245 107.385 110.475 108.375 ;
        RECT 110.645 107.555 110.995 108.205 ;
        RECT 111.170 108.125 112.380 109.215 ;
        RECT 111.170 107.585 111.690 108.125 ;
        RECT 111.860 107.415 112.380 107.955 ;
        RECT 110.245 107.215 110.995 107.385 ;
        RECT 110.240 106.665 110.570 107.045 ;
        RECT 110.740 106.925 110.995 107.215 ;
        RECT 111.170 106.665 112.380 107.415 ;
        RECT 18.165 106.495 112.465 106.665 ;
        RECT 18.250 105.745 19.460 106.495 ;
        RECT 18.250 105.205 18.770 105.745 ;
        RECT 20.090 105.725 21.760 106.495 ;
        RECT 21.930 105.770 22.220 106.495 ;
        RECT 22.390 105.745 23.600 106.495 ;
        RECT 18.940 105.035 19.460 105.575 ;
        RECT 18.250 103.945 19.460 105.035 ;
        RECT 20.090 105.035 20.840 105.555 ;
        RECT 21.010 105.205 21.760 105.725 ;
        RECT 20.090 103.945 21.760 105.035 ;
        RECT 21.930 103.945 22.220 105.110 ;
        RECT 22.390 105.035 22.910 105.575 ;
        RECT 23.080 105.205 23.600 105.745 ;
        RECT 23.810 105.675 24.040 106.495 ;
        RECT 24.210 105.695 24.540 106.325 ;
        RECT 23.790 105.255 24.120 105.505 ;
        RECT 24.290 105.095 24.540 105.695 ;
        RECT 24.710 105.675 24.920 106.495 ;
        RECT 25.190 105.675 25.420 106.495 ;
        RECT 25.590 105.695 25.920 106.325 ;
        RECT 25.170 105.255 25.500 105.505 ;
        RECT 25.670 105.095 25.920 105.695 ;
        RECT 26.090 105.675 26.300 106.495 ;
        RECT 26.840 106.025 27.010 106.495 ;
        RECT 27.180 105.845 27.510 106.325 ;
        RECT 27.680 106.025 27.850 106.495 ;
        RECT 28.020 105.845 28.350 106.325 ;
        RECT 26.585 105.675 28.350 105.845 ;
        RECT 28.520 105.685 28.690 106.495 ;
        RECT 28.890 106.115 29.960 106.285 ;
        RECT 28.890 105.760 29.210 106.115 ;
        RECT 22.390 103.945 23.600 105.035 ;
        RECT 23.810 103.945 24.040 105.085 ;
        RECT 24.210 104.115 24.540 105.095 ;
        RECT 24.710 103.945 24.920 105.085 ;
        RECT 25.190 103.945 25.420 105.085 ;
        RECT 25.590 104.115 25.920 105.095 ;
        RECT 26.585 105.125 26.995 105.675 ;
        RECT 28.885 105.505 29.210 105.760 ;
        RECT 27.180 105.295 29.210 105.505 ;
        RECT 28.865 105.285 29.210 105.295 ;
        RECT 29.380 105.545 29.620 105.945 ;
        RECT 29.790 105.885 29.960 106.115 ;
        RECT 30.130 106.055 30.320 106.495 ;
        RECT 30.490 106.045 31.440 106.325 ;
        RECT 31.660 106.135 32.010 106.305 ;
        RECT 29.790 105.715 30.320 105.885 ;
        RECT 26.090 103.945 26.300 105.085 ;
        RECT 26.585 104.955 28.310 105.125 ;
        RECT 26.840 103.945 27.010 104.785 ;
        RECT 27.220 104.115 27.470 104.955 ;
        RECT 27.680 103.945 27.850 104.785 ;
        RECT 28.020 104.115 28.310 104.955 ;
        RECT 28.520 103.945 28.690 105.005 ;
        RECT 28.865 104.665 29.035 105.285 ;
        RECT 29.380 105.175 29.920 105.545 ;
        RECT 30.100 105.435 30.320 105.715 ;
        RECT 30.490 105.265 30.660 106.045 ;
        RECT 30.255 105.095 30.660 105.265 ;
        RECT 30.830 105.255 31.180 105.875 ;
        RECT 30.255 105.005 30.425 105.095 ;
        RECT 31.350 105.085 31.560 105.875 ;
        RECT 29.205 104.835 30.425 105.005 ;
        RECT 30.885 104.925 31.560 105.085 ;
        RECT 28.865 104.495 29.665 104.665 ;
        RECT 28.985 103.945 29.315 104.325 ;
        RECT 29.495 104.205 29.665 104.495 ;
        RECT 30.255 104.455 30.425 104.835 ;
        RECT 30.595 104.915 31.560 104.925 ;
        RECT 31.750 105.745 32.010 106.135 ;
        RECT 32.220 106.035 32.550 106.495 ;
        RECT 33.425 106.105 34.280 106.275 ;
        RECT 34.485 106.105 34.980 106.275 ;
        RECT 35.150 106.135 35.480 106.495 ;
        RECT 31.750 105.055 31.920 105.745 ;
        RECT 32.090 105.395 32.260 105.575 ;
        RECT 32.430 105.565 33.220 105.815 ;
        RECT 33.425 105.395 33.595 106.105 ;
        RECT 33.765 105.595 34.120 105.815 ;
        RECT 32.090 105.225 33.780 105.395 ;
        RECT 30.595 104.625 31.055 104.915 ;
        RECT 31.750 104.885 33.250 105.055 ;
        RECT 31.750 104.745 31.920 104.885 ;
        RECT 31.360 104.575 31.920 104.745 ;
        RECT 29.835 103.945 30.085 104.405 ;
        RECT 30.255 104.115 31.125 104.455 ;
        RECT 31.360 104.115 31.530 104.575 ;
        RECT 32.365 104.545 33.440 104.715 ;
        RECT 31.700 103.945 32.070 104.405 ;
        RECT 32.365 104.205 32.535 104.545 ;
        RECT 32.705 103.945 33.035 104.375 ;
        RECT 33.270 104.205 33.440 104.545 ;
        RECT 33.610 104.445 33.780 105.225 ;
        RECT 33.950 105.005 34.120 105.595 ;
        RECT 34.290 105.195 34.640 105.815 ;
        RECT 33.950 104.615 34.415 105.005 ;
        RECT 34.810 104.745 34.980 106.105 ;
        RECT 35.150 104.915 35.610 105.965 ;
        RECT 34.585 104.575 34.980 104.745 ;
        RECT 34.585 104.445 34.755 104.575 ;
        RECT 33.610 104.115 34.290 104.445 ;
        RECT 34.505 104.115 34.755 104.445 ;
        RECT 34.925 103.945 35.175 104.405 ;
        RECT 35.345 104.130 35.670 104.915 ;
        RECT 35.840 104.115 36.010 106.235 ;
        RECT 36.180 106.115 36.510 106.495 ;
        RECT 36.680 105.945 36.935 106.235 ;
        RECT 36.185 105.775 36.935 105.945 ;
        RECT 37.115 105.945 37.370 106.235 ;
        RECT 37.540 106.115 37.870 106.495 ;
        RECT 37.115 105.775 37.865 105.945 ;
        RECT 36.185 104.785 36.415 105.775 ;
        RECT 36.585 104.955 36.935 105.605 ;
        RECT 37.115 104.955 37.465 105.605 ;
        RECT 37.635 104.785 37.865 105.775 ;
        RECT 36.185 104.615 36.935 104.785 ;
        RECT 36.180 103.945 36.510 104.445 ;
        RECT 36.680 104.115 36.935 104.615 ;
        RECT 37.115 104.615 37.865 104.785 ;
        RECT 37.115 104.115 37.370 104.615 ;
        RECT 37.540 103.945 37.870 104.445 ;
        RECT 38.040 104.115 38.210 106.235 ;
        RECT 38.570 106.135 38.900 106.495 ;
        RECT 39.070 106.105 39.565 106.275 ;
        RECT 39.770 106.105 40.625 106.275 ;
        RECT 38.440 104.915 38.900 105.965 ;
        RECT 38.380 104.130 38.705 104.915 ;
        RECT 39.070 104.745 39.240 106.105 ;
        RECT 39.410 105.195 39.760 105.815 ;
        RECT 39.930 105.595 40.285 105.815 ;
        RECT 39.930 105.005 40.100 105.595 ;
        RECT 40.455 105.395 40.625 106.105 ;
        RECT 41.500 106.035 41.830 106.495 ;
        RECT 42.040 106.135 42.390 106.305 ;
        RECT 40.830 105.565 41.620 105.815 ;
        RECT 42.040 105.745 42.300 106.135 ;
        RECT 42.610 106.045 43.560 106.325 ;
        RECT 43.730 106.055 43.920 106.495 ;
        RECT 44.090 106.115 45.160 106.285 ;
        RECT 41.790 105.395 41.960 105.575 ;
        RECT 39.070 104.575 39.465 104.745 ;
        RECT 39.635 104.615 40.100 105.005 ;
        RECT 40.270 105.225 41.960 105.395 ;
        RECT 39.295 104.445 39.465 104.575 ;
        RECT 40.270 104.445 40.440 105.225 ;
        RECT 42.130 105.055 42.300 105.745 ;
        RECT 40.800 104.885 42.300 105.055 ;
        RECT 42.490 105.085 42.700 105.875 ;
        RECT 42.870 105.255 43.220 105.875 ;
        RECT 43.390 105.265 43.560 106.045 ;
        RECT 44.090 105.885 44.260 106.115 ;
        RECT 43.730 105.715 44.260 105.885 ;
        RECT 43.730 105.435 43.950 105.715 ;
        RECT 44.430 105.545 44.670 105.945 ;
        RECT 43.390 105.095 43.795 105.265 ;
        RECT 44.130 105.175 44.670 105.545 ;
        RECT 44.840 105.760 45.160 106.115 ;
        RECT 44.840 105.505 45.165 105.760 ;
        RECT 45.360 105.685 45.530 106.495 ;
        RECT 45.700 105.845 46.030 106.325 ;
        RECT 46.200 106.025 46.370 106.495 ;
        RECT 46.540 105.845 46.870 106.325 ;
        RECT 47.040 106.025 47.210 106.495 ;
        RECT 45.700 105.675 47.465 105.845 ;
        RECT 47.690 105.770 47.980 106.495 ;
        RECT 48.150 105.745 49.360 106.495 ;
        RECT 44.840 105.295 46.870 105.505 ;
        RECT 44.840 105.285 45.185 105.295 ;
        RECT 42.490 104.925 43.165 105.085 ;
        RECT 43.625 105.005 43.795 105.095 ;
        RECT 42.490 104.915 43.455 104.925 ;
        RECT 42.130 104.745 42.300 104.885 ;
        RECT 38.875 103.945 39.125 104.405 ;
        RECT 39.295 104.115 39.545 104.445 ;
        RECT 39.760 104.115 40.440 104.445 ;
        RECT 40.610 104.545 41.685 104.715 ;
        RECT 42.130 104.575 42.690 104.745 ;
        RECT 42.995 104.625 43.455 104.915 ;
        RECT 43.625 104.835 44.845 105.005 ;
        RECT 40.610 104.205 40.780 104.545 ;
        RECT 41.015 103.945 41.345 104.375 ;
        RECT 41.515 104.205 41.685 104.545 ;
        RECT 41.980 103.945 42.350 104.405 ;
        RECT 42.520 104.115 42.690 104.575 ;
        RECT 43.625 104.455 43.795 104.835 ;
        RECT 45.015 104.665 45.185 105.285 ;
        RECT 47.055 105.125 47.465 105.675 ;
        RECT 42.925 104.115 43.795 104.455 ;
        RECT 44.385 104.495 45.185 104.665 ;
        RECT 43.965 103.945 44.215 104.405 ;
        RECT 44.385 104.205 44.555 104.495 ;
        RECT 44.735 103.945 45.065 104.325 ;
        RECT 45.360 103.945 45.530 105.005 ;
        RECT 45.740 104.955 47.465 105.125 ;
        RECT 45.740 104.115 46.030 104.955 ;
        RECT 46.200 103.945 46.370 104.785 ;
        RECT 46.580 104.115 46.830 104.955 ;
        RECT 47.040 103.945 47.210 104.785 ;
        RECT 47.690 103.945 47.980 105.110 ;
        RECT 48.150 105.035 48.670 105.575 ;
        RECT 48.840 105.205 49.360 105.745 ;
        RECT 49.590 105.675 49.800 106.495 ;
        RECT 49.970 105.695 50.300 106.325 ;
        RECT 49.970 105.095 50.220 105.695 ;
        RECT 50.470 105.675 50.700 106.495 ;
        RECT 50.910 105.745 52.120 106.495 ;
        RECT 50.390 105.255 50.720 105.505 ;
        RECT 48.150 103.945 49.360 105.035 ;
        RECT 49.590 103.945 49.800 105.085 ;
        RECT 49.970 104.115 50.300 105.095 ;
        RECT 50.470 103.945 50.700 105.085 ;
        RECT 50.910 105.035 51.430 105.575 ;
        RECT 51.600 105.205 52.120 105.745 ;
        RECT 52.330 105.675 52.560 106.495 ;
        RECT 52.730 105.695 53.060 106.325 ;
        RECT 52.310 105.255 52.640 105.505 ;
        RECT 52.810 105.095 53.060 105.695 ;
        RECT 53.230 105.675 53.440 106.495 ;
        RECT 53.760 105.945 53.930 106.325 ;
        RECT 54.110 106.115 54.440 106.495 ;
        RECT 53.760 105.775 54.425 105.945 ;
        RECT 54.620 105.820 54.880 106.325 ;
        RECT 55.360 106.025 55.530 106.495 ;
        RECT 55.700 105.845 56.030 106.325 ;
        RECT 56.200 106.025 56.370 106.495 ;
        RECT 56.540 105.845 56.870 106.325 ;
        RECT 53.690 105.225 54.020 105.595 ;
        RECT 54.255 105.520 54.425 105.775 ;
        RECT 50.910 103.945 52.120 105.035 ;
        RECT 52.330 103.945 52.560 105.085 ;
        RECT 52.730 104.115 53.060 105.095 ;
        RECT 54.255 105.190 54.540 105.520 ;
        RECT 53.230 103.945 53.440 105.085 ;
        RECT 54.255 105.045 54.425 105.190 ;
        RECT 53.760 104.875 54.425 105.045 ;
        RECT 54.710 105.020 54.880 105.820 ;
        RECT 53.760 104.115 53.930 104.875 ;
        RECT 54.110 103.945 54.440 104.705 ;
        RECT 54.610 104.115 54.880 105.020 ;
        RECT 55.105 105.675 56.870 105.845 ;
        RECT 57.040 105.685 57.210 106.495 ;
        RECT 57.410 106.115 58.480 106.285 ;
        RECT 57.410 105.760 57.730 106.115 ;
        RECT 55.105 105.125 55.515 105.675 ;
        RECT 57.405 105.505 57.730 105.760 ;
        RECT 55.700 105.295 57.730 105.505 ;
        RECT 57.385 105.285 57.730 105.295 ;
        RECT 57.900 105.545 58.140 105.945 ;
        RECT 58.310 105.885 58.480 106.115 ;
        RECT 58.650 106.055 58.840 106.495 ;
        RECT 59.010 106.045 59.960 106.325 ;
        RECT 60.180 106.135 60.530 106.305 ;
        RECT 58.310 105.715 58.840 105.885 ;
        RECT 55.105 104.955 56.830 105.125 ;
        RECT 55.360 103.945 55.530 104.785 ;
        RECT 55.740 104.115 55.990 104.955 ;
        RECT 56.200 103.945 56.370 104.785 ;
        RECT 56.540 104.115 56.830 104.955 ;
        RECT 57.040 103.945 57.210 105.005 ;
        RECT 57.385 104.665 57.555 105.285 ;
        RECT 57.900 105.175 58.440 105.545 ;
        RECT 58.620 105.435 58.840 105.715 ;
        RECT 59.010 105.265 59.180 106.045 ;
        RECT 58.775 105.095 59.180 105.265 ;
        RECT 59.350 105.255 59.700 105.875 ;
        RECT 58.775 105.005 58.945 105.095 ;
        RECT 59.870 105.085 60.080 105.875 ;
        RECT 57.725 104.835 58.945 105.005 ;
        RECT 59.405 104.925 60.080 105.085 ;
        RECT 57.385 104.495 58.185 104.665 ;
        RECT 57.505 103.945 57.835 104.325 ;
        RECT 58.015 104.205 58.185 104.495 ;
        RECT 58.775 104.455 58.945 104.835 ;
        RECT 59.115 104.915 60.080 104.925 ;
        RECT 60.270 105.745 60.530 106.135 ;
        RECT 60.740 106.035 61.070 106.495 ;
        RECT 61.945 106.105 62.800 106.275 ;
        RECT 63.005 106.105 63.500 106.275 ;
        RECT 63.670 106.135 64.000 106.495 ;
        RECT 60.270 105.055 60.440 105.745 ;
        RECT 60.610 105.395 60.780 105.575 ;
        RECT 60.950 105.565 61.740 105.815 ;
        RECT 61.945 105.395 62.115 106.105 ;
        RECT 62.285 105.595 62.640 105.815 ;
        RECT 60.610 105.225 62.300 105.395 ;
        RECT 59.115 104.625 59.575 104.915 ;
        RECT 60.270 104.885 61.770 105.055 ;
        RECT 60.270 104.745 60.440 104.885 ;
        RECT 59.880 104.575 60.440 104.745 ;
        RECT 58.355 103.945 58.605 104.405 ;
        RECT 58.775 104.115 59.645 104.455 ;
        RECT 59.880 104.115 60.050 104.575 ;
        RECT 60.885 104.545 61.960 104.715 ;
        RECT 60.220 103.945 60.590 104.405 ;
        RECT 60.885 104.205 61.055 104.545 ;
        RECT 61.225 103.945 61.555 104.375 ;
        RECT 61.790 104.205 61.960 104.545 ;
        RECT 62.130 104.445 62.300 105.225 ;
        RECT 62.470 105.005 62.640 105.595 ;
        RECT 62.810 105.195 63.160 105.815 ;
        RECT 62.470 104.615 62.935 105.005 ;
        RECT 63.330 104.745 63.500 106.105 ;
        RECT 63.670 104.915 64.130 105.965 ;
        RECT 63.105 104.575 63.500 104.745 ;
        RECT 63.105 104.445 63.275 104.575 ;
        RECT 62.130 104.115 62.810 104.445 ;
        RECT 63.025 104.115 63.275 104.445 ;
        RECT 63.445 103.945 63.695 104.405 ;
        RECT 63.865 104.130 64.190 104.915 ;
        RECT 64.360 104.115 64.530 106.235 ;
        RECT 64.700 106.115 65.030 106.495 ;
        RECT 65.200 105.945 65.455 106.235 ;
        RECT 64.705 105.775 65.455 105.945 ;
        RECT 64.705 104.785 64.935 105.775 ;
        RECT 66.090 105.725 68.680 106.495 ;
        RECT 65.105 104.955 65.455 105.605 ;
        RECT 66.090 105.035 67.300 105.555 ;
        RECT 67.470 105.205 68.680 105.725 ;
        RECT 68.910 105.675 69.120 106.495 ;
        RECT 69.290 105.695 69.620 106.325 ;
        RECT 69.290 105.095 69.540 105.695 ;
        RECT 69.790 105.675 70.020 106.495 ;
        RECT 70.290 105.675 70.500 106.495 ;
        RECT 70.670 105.695 71.000 106.325 ;
        RECT 69.710 105.255 70.040 105.505 ;
        RECT 70.670 105.095 70.920 105.695 ;
        RECT 71.170 105.675 71.400 106.495 ;
        RECT 72.160 105.945 72.330 106.325 ;
        RECT 72.510 106.115 72.840 106.495 ;
        RECT 72.160 105.775 72.825 105.945 ;
        RECT 73.020 105.820 73.280 106.325 ;
        RECT 71.090 105.255 71.420 105.505 ;
        RECT 72.090 105.225 72.420 105.595 ;
        RECT 72.655 105.520 72.825 105.775 ;
        RECT 72.655 105.190 72.940 105.520 ;
        RECT 64.705 104.615 65.455 104.785 ;
        RECT 64.700 103.945 65.030 104.445 ;
        RECT 65.200 104.115 65.455 104.615 ;
        RECT 66.090 103.945 68.680 105.035 ;
        RECT 68.910 103.945 69.120 105.085 ;
        RECT 69.290 104.115 69.620 105.095 ;
        RECT 69.790 103.945 70.020 105.085 ;
        RECT 70.290 103.945 70.500 105.085 ;
        RECT 70.670 104.115 71.000 105.095 ;
        RECT 71.170 103.945 71.400 105.085 ;
        RECT 72.655 105.045 72.825 105.190 ;
        RECT 72.160 104.875 72.825 105.045 ;
        RECT 73.110 105.020 73.280 105.820 ;
        RECT 73.450 105.770 73.740 106.495 ;
        RECT 74.220 106.025 74.390 106.495 ;
        RECT 74.560 105.845 74.890 106.325 ;
        RECT 75.060 106.025 75.230 106.495 ;
        RECT 75.400 105.845 75.730 106.325 ;
        RECT 73.965 105.675 75.730 105.845 ;
        RECT 75.900 105.685 76.070 106.495 ;
        RECT 76.270 106.115 77.340 106.285 ;
        RECT 76.270 105.760 76.590 106.115 ;
        RECT 73.965 105.125 74.375 105.675 ;
        RECT 76.265 105.505 76.590 105.760 ;
        RECT 74.560 105.295 76.590 105.505 ;
        RECT 76.245 105.285 76.590 105.295 ;
        RECT 76.760 105.545 77.000 105.945 ;
        RECT 77.170 105.885 77.340 106.115 ;
        RECT 77.510 106.055 77.700 106.495 ;
        RECT 77.870 106.045 78.820 106.325 ;
        RECT 79.040 106.135 79.390 106.305 ;
        RECT 77.170 105.715 77.700 105.885 ;
        RECT 72.160 104.115 72.330 104.875 ;
        RECT 72.510 103.945 72.840 104.705 ;
        RECT 73.010 104.115 73.280 105.020 ;
        RECT 73.450 103.945 73.740 105.110 ;
        RECT 73.965 104.955 75.690 105.125 ;
        RECT 74.220 103.945 74.390 104.785 ;
        RECT 74.600 104.115 74.850 104.955 ;
        RECT 75.060 103.945 75.230 104.785 ;
        RECT 75.400 104.115 75.690 104.955 ;
        RECT 75.900 103.945 76.070 105.005 ;
        RECT 76.245 104.665 76.415 105.285 ;
        RECT 76.760 105.175 77.300 105.545 ;
        RECT 77.480 105.435 77.700 105.715 ;
        RECT 77.870 105.265 78.040 106.045 ;
        RECT 77.635 105.095 78.040 105.265 ;
        RECT 78.210 105.255 78.560 105.875 ;
        RECT 77.635 105.005 77.805 105.095 ;
        RECT 78.730 105.085 78.940 105.875 ;
        RECT 76.585 104.835 77.805 105.005 ;
        RECT 78.265 104.925 78.940 105.085 ;
        RECT 76.245 104.495 77.045 104.665 ;
        RECT 76.365 103.945 76.695 104.325 ;
        RECT 76.875 104.205 77.045 104.495 ;
        RECT 77.635 104.455 77.805 104.835 ;
        RECT 77.975 104.915 78.940 104.925 ;
        RECT 79.130 105.745 79.390 106.135 ;
        RECT 79.600 106.035 79.930 106.495 ;
        RECT 80.805 106.105 81.660 106.275 ;
        RECT 81.865 106.105 82.360 106.275 ;
        RECT 82.530 106.135 82.860 106.495 ;
        RECT 79.130 105.055 79.300 105.745 ;
        RECT 79.470 105.395 79.640 105.575 ;
        RECT 79.810 105.565 80.600 105.815 ;
        RECT 80.805 105.395 80.975 106.105 ;
        RECT 81.145 105.595 81.500 105.815 ;
        RECT 79.470 105.225 81.160 105.395 ;
        RECT 77.975 104.625 78.435 104.915 ;
        RECT 79.130 104.885 80.630 105.055 ;
        RECT 79.130 104.745 79.300 104.885 ;
        RECT 78.740 104.575 79.300 104.745 ;
        RECT 77.215 103.945 77.465 104.405 ;
        RECT 77.635 104.115 78.505 104.455 ;
        RECT 78.740 104.115 78.910 104.575 ;
        RECT 79.745 104.545 80.820 104.715 ;
        RECT 79.080 103.945 79.450 104.405 ;
        RECT 79.745 104.205 79.915 104.545 ;
        RECT 80.085 103.945 80.415 104.375 ;
        RECT 80.650 104.205 80.820 104.545 ;
        RECT 80.990 104.445 81.160 105.225 ;
        RECT 81.330 105.005 81.500 105.595 ;
        RECT 81.670 105.195 82.020 105.815 ;
        RECT 81.330 104.615 81.795 105.005 ;
        RECT 82.190 104.745 82.360 106.105 ;
        RECT 82.530 104.915 82.990 105.965 ;
        RECT 81.965 104.575 82.360 104.745 ;
        RECT 81.965 104.445 82.135 104.575 ;
        RECT 80.990 104.115 81.670 104.445 ;
        RECT 81.885 104.115 82.135 104.445 ;
        RECT 82.305 103.945 82.555 104.405 ;
        RECT 82.725 104.130 83.050 104.915 ;
        RECT 83.220 104.115 83.390 106.235 ;
        RECT 83.560 106.115 83.890 106.495 ;
        RECT 84.060 105.945 84.315 106.235 ;
        RECT 84.800 106.025 84.970 106.495 ;
        RECT 83.565 105.775 84.315 105.945 ;
        RECT 85.140 105.845 85.470 106.325 ;
        RECT 85.640 106.025 85.810 106.495 ;
        RECT 85.980 105.845 86.310 106.325 ;
        RECT 83.565 104.785 83.795 105.775 ;
        RECT 84.545 105.675 86.310 105.845 ;
        RECT 86.480 105.685 86.650 106.495 ;
        RECT 86.850 106.115 87.920 106.285 ;
        RECT 86.850 105.760 87.170 106.115 ;
        RECT 83.965 104.955 84.315 105.605 ;
        RECT 84.545 105.125 84.955 105.675 ;
        RECT 86.845 105.505 87.170 105.760 ;
        RECT 85.140 105.295 87.170 105.505 ;
        RECT 86.825 105.285 87.170 105.295 ;
        RECT 87.340 105.545 87.580 105.945 ;
        RECT 87.750 105.885 87.920 106.115 ;
        RECT 88.090 106.055 88.280 106.495 ;
        RECT 88.450 106.045 89.400 106.325 ;
        RECT 89.620 106.135 89.970 106.305 ;
        RECT 87.750 105.715 88.280 105.885 ;
        RECT 84.545 104.955 86.270 105.125 ;
        RECT 83.565 104.615 84.315 104.785 ;
        RECT 83.560 103.945 83.890 104.445 ;
        RECT 84.060 104.115 84.315 104.615 ;
        RECT 84.800 103.945 84.970 104.785 ;
        RECT 85.180 104.115 85.430 104.955 ;
        RECT 85.640 103.945 85.810 104.785 ;
        RECT 85.980 104.115 86.270 104.955 ;
        RECT 86.480 103.945 86.650 105.005 ;
        RECT 86.825 104.665 86.995 105.285 ;
        RECT 87.340 105.175 87.880 105.545 ;
        RECT 88.060 105.435 88.280 105.715 ;
        RECT 88.450 105.265 88.620 106.045 ;
        RECT 88.215 105.095 88.620 105.265 ;
        RECT 88.790 105.255 89.140 105.875 ;
        RECT 88.215 105.005 88.385 105.095 ;
        RECT 89.310 105.085 89.520 105.875 ;
        RECT 87.165 104.835 88.385 105.005 ;
        RECT 88.845 104.925 89.520 105.085 ;
        RECT 86.825 104.495 87.625 104.665 ;
        RECT 86.945 103.945 87.275 104.325 ;
        RECT 87.455 104.205 87.625 104.495 ;
        RECT 88.215 104.455 88.385 104.835 ;
        RECT 88.555 104.915 89.520 104.925 ;
        RECT 89.710 105.745 89.970 106.135 ;
        RECT 90.180 106.035 90.510 106.495 ;
        RECT 91.385 106.105 92.240 106.275 ;
        RECT 92.445 106.105 92.940 106.275 ;
        RECT 93.110 106.135 93.440 106.495 ;
        RECT 89.710 105.055 89.880 105.745 ;
        RECT 90.050 105.395 90.220 105.575 ;
        RECT 90.390 105.565 91.180 105.815 ;
        RECT 91.385 105.395 91.555 106.105 ;
        RECT 91.725 105.595 92.080 105.815 ;
        RECT 90.050 105.225 91.740 105.395 ;
        RECT 88.555 104.625 89.015 104.915 ;
        RECT 89.710 104.885 91.210 105.055 ;
        RECT 89.710 104.745 89.880 104.885 ;
        RECT 89.320 104.575 89.880 104.745 ;
        RECT 87.795 103.945 88.045 104.405 ;
        RECT 88.215 104.115 89.085 104.455 ;
        RECT 89.320 104.115 89.490 104.575 ;
        RECT 90.325 104.545 91.400 104.715 ;
        RECT 89.660 103.945 90.030 104.405 ;
        RECT 90.325 104.205 90.495 104.545 ;
        RECT 90.665 103.945 90.995 104.375 ;
        RECT 91.230 104.205 91.400 104.545 ;
        RECT 91.570 104.445 91.740 105.225 ;
        RECT 91.910 105.005 92.080 105.595 ;
        RECT 92.250 105.195 92.600 105.815 ;
        RECT 91.910 104.615 92.375 105.005 ;
        RECT 92.770 104.745 92.940 106.105 ;
        RECT 93.110 104.915 93.570 105.965 ;
        RECT 92.545 104.575 92.940 104.745 ;
        RECT 92.545 104.445 92.715 104.575 ;
        RECT 91.570 104.115 92.250 104.445 ;
        RECT 92.465 104.115 92.715 104.445 ;
        RECT 92.885 103.945 93.135 104.405 ;
        RECT 93.305 104.130 93.630 104.915 ;
        RECT 93.800 104.115 93.970 106.235 ;
        RECT 94.140 106.115 94.470 106.495 ;
        RECT 94.640 105.945 94.895 106.235 ;
        RECT 94.145 105.775 94.895 105.945 ;
        RECT 94.145 104.785 94.375 105.775 ;
        RECT 95.070 105.725 97.660 106.495 ;
        RECT 94.545 104.955 94.895 105.605 ;
        RECT 95.070 105.035 96.280 105.555 ;
        RECT 96.450 105.205 97.660 105.725 ;
        RECT 97.870 105.675 98.100 106.495 ;
        RECT 98.270 105.695 98.600 106.325 ;
        RECT 97.850 105.255 98.180 105.505 ;
        RECT 98.350 105.095 98.600 105.695 ;
        RECT 98.770 105.675 98.980 106.495 ;
        RECT 99.210 105.770 99.500 106.495 ;
        RECT 99.980 106.025 100.150 106.495 ;
        RECT 100.320 105.845 100.650 106.325 ;
        RECT 100.820 106.025 100.990 106.495 ;
        RECT 101.160 105.845 101.490 106.325 ;
        RECT 99.725 105.675 101.490 105.845 ;
        RECT 101.660 105.685 101.830 106.495 ;
        RECT 102.030 106.115 103.100 106.285 ;
        RECT 102.030 105.760 102.350 106.115 ;
        RECT 99.725 105.125 100.135 105.675 ;
        RECT 102.025 105.505 102.350 105.760 ;
        RECT 100.320 105.295 102.350 105.505 ;
        RECT 102.005 105.285 102.350 105.295 ;
        RECT 102.520 105.545 102.760 105.945 ;
        RECT 102.930 105.885 103.100 106.115 ;
        RECT 103.270 106.055 103.460 106.495 ;
        RECT 103.630 106.045 104.580 106.325 ;
        RECT 104.800 106.135 105.150 106.305 ;
        RECT 102.930 105.715 103.460 105.885 ;
        RECT 94.145 104.615 94.895 104.785 ;
        RECT 94.140 103.945 94.470 104.445 ;
        RECT 94.640 104.115 94.895 104.615 ;
        RECT 95.070 103.945 97.660 105.035 ;
        RECT 97.870 103.945 98.100 105.085 ;
        RECT 98.270 104.115 98.600 105.095 ;
        RECT 98.770 103.945 98.980 105.085 ;
        RECT 99.210 103.945 99.500 105.110 ;
        RECT 99.725 104.955 101.450 105.125 ;
        RECT 99.980 103.945 100.150 104.785 ;
        RECT 100.360 104.115 100.610 104.955 ;
        RECT 100.820 103.945 100.990 104.785 ;
        RECT 101.160 104.115 101.450 104.955 ;
        RECT 101.660 103.945 101.830 105.005 ;
        RECT 102.005 104.665 102.175 105.285 ;
        RECT 102.520 105.175 103.060 105.545 ;
        RECT 103.240 105.435 103.460 105.715 ;
        RECT 103.630 105.265 103.800 106.045 ;
        RECT 103.395 105.095 103.800 105.265 ;
        RECT 103.970 105.255 104.320 105.875 ;
        RECT 103.395 105.005 103.565 105.095 ;
        RECT 104.490 105.085 104.700 105.875 ;
        RECT 102.345 104.835 103.565 105.005 ;
        RECT 104.025 104.925 104.700 105.085 ;
        RECT 102.005 104.495 102.805 104.665 ;
        RECT 102.125 103.945 102.455 104.325 ;
        RECT 102.635 104.205 102.805 104.495 ;
        RECT 103.395 104.455 103.565 104.835 ;
        RECT 103.735 104.915 104.700 104.925 ;
        RECT 104.890 105.745 105.150 106.135 ;
        RECT 105.360 106.035 105.690 106.495 ;
        RECT 106.565 106.105 107.420 106.275 ;
        RECT 107.625 106.105 108.120 106.275 ;
        RECT 108.290 106.135 108.620 106.495 ;
        RECT 104.890 105.055 105.060 105.745 ;
        RECT 105.230 105.395 105.400 105.575 ;
        RECT 105.570 105.565 106.360 105.815 ;
        RECT 106.565 105.395 106.735 106.105 ;
        RECT 106.905 105.595 107.260 105.815 ;
        RECT 105.230 105.225 106.920 105.395 ;
        RECT 103.735 104.625 104.195 104.915 ;
        RECT 104.890 104.885 106.390 105.055 ;
        RECT 104.890 104.745 105.060 104.885 ;
        RECT 104.500 104.575 105.060 104.745 ;
        RECT 102.975 103.945 103.225 104.405 ;
        RECT 103.395 104.115 104.265 104.455 ;
        RECT 104.500 104.115 104.670 104.575 ;
        RECT 105.505 104.545 106.580 104.715 ;
        RECT 104.840 103.945 105.210 104.405 ;
        RECT 105.505 104.205 105.675 104.545 ;
        RECT 105.845 103.945 106.175 104.375 ;
        RECT 106.410 104.205 106.580 104.545 ;
        RECT 106.750 104.445 106.920 105.225 ;
        RECT 107.090 105.005 107.260 105.595 ;
        RECT 107.430 105.195 107.780 105.815 ;
        RECT 107.090 104.615 107.555 105.005 ;
        RECT 107.950 104.745 108.120 106.105 ;
        RECT 108.290 104.915 108.750 105.965 ;
        RECT 107.725 104.575 108.120 104.745 ;
        RECT 107.725 104.445 107.895 104.575 ;
        RECT 106.750 104.115 107.430 104.445 ;
        RECT 107.645 104.115 107.895 104.445 ;
        RECT 108.065 103.945 108.315 104.405 ;
        RECT 108.485 104.130 108.810 104.915 ;
        RECT 108.980 104.115 109.150 106.235 ;
        RECT 109.320 106.115 109.650 106.495 ;
        RECT 109.820 105.945 110.075 106.235 ;
        RECT 109.325 105.775 110.075 105.945 ;
        RECT 109.325 104.785 109.555 105.775 ;
        RECT 111.170 105.745 112.380 106.495 ;
        RECT 109.725 104.955 110.075 105.605 ;
        RECT 111.170 105.035 111.690 105.575 ;
        RECT 111.860 105.205 112.380 105.745 ;
        RECT 109.325 104.615 110.075 104.785 ;
        RECT 109.320 103.945 109.650 104.445 ;
        RECT 109.820 104.115 110.075 104.615 ;
        RECT 111.170 103.945 112.380 105.035 ;
        RECT 18.165 103.775 112.465 103.945 ;
        RECT 18.250 102.685 19.460 103.775 ;
        RECT 18.250 101.975 18.770 102.515 ;
        RECT 18.940 102.145 19.460 102.685 ;
        RECT 20.090 102.685 21.760 103.775 ;
        RECT 20.090 102.165 20.840 102.685 ;
        RECT 21.930 102.610 22.220 103.775 ;
        RECT 22.700 102.935 22.870 103.775 ;
        RECT 23.080 102.765 23.330 103.605 ;
        RECT 23.540 102.935 23.710 103.775 ;
        RECT 23.880 102.765 24.170 103.605 ;
        RECT 22.445 102.595 24.170 102.765 ;
        RECT 24.380 102.715 24.550 103.775 ;
        RECT 24.845 103.395 25.175 103.775 ;
        RECT 25.355 103.225 25.525 103.515 ;
        RECT 25.695 103.315 25.945 103.775 ;
        RECT 24.725 103.055 25.525 103.225 ;
        RECT 26.115 103.265 26.985 103.605 ;
        RECT 21.010 101.995 21.760 102.515 ;
        RECT 18.250 101.225 19.460 101.975 ;
        RECT 20.090 101.225 21.760 101.995 ;
        RECT 22.445 102.045 22.855 102.595 ;
        RECT 24.725 102.435 24.895 103.055 ;
        RECT 26.115 102.885 26.285 103.265 ;
        RECT 27.220 103.145 27.390 103.605 ;
        RECT 27.560 103.315 27.930 103.775 ;
        RECT 28.225 103.175 28.395 103.515 ;
        RECT 28.565 103.345 28.895 103.775 ;
        RECT 29.130 103.175 29.300 103.515 ;
        RECT 25.065 102.715 26.285 102.885 ;
        RECT 26.455 102.805 26.915 103.095 ;
        RECT 27.220 102.975 27.780 103.145 ;
        RECT 28.225 103.005 29.300 103.175 ;
        RECT 29.470 103.275 30.150 103.605 ;
        RECT 30.365 103.275 30.615 103.605 ;
        RECT 30.785 103.315 31.035 103.775 ;
        RECT 27.610 102.835 27.780 102.975 ;
        RECT 26.455 102.795 27.420 102.805 ;
        RECT 26.115 102.625 26.285 102.715 ;
        RECT 26.745 102.635 27.420 102.795 ;
        RECT 24.725 102.425 25.070 102.435 ;
        RECT 23.040 102.215 25.070 102.425 ;
        RECT 21.930 101.225 22.220 101.950 ;
        RECT 22.445 101.875 24.210 102.045 ;
        RECT 22.700 101.225 22.870 101.695 ;
        RECT 23.040 101.395 23.370 101.875 ;
        RECT 23.540 101.225 23.710 101.695 ;
        RECT 23.880 101.395 24.210 101.875 ;
        RECT 24.380 101.225 24.550 102.035 ;
        RECT 24.745 101.960 25.070 102.215 ;
        RECT 24.750 101.605 25.070 101.960 ;
        RECT 25.240 102.175 25.780 102.545 ;
        RECT 26.115 102.455 26.520 102.625 ;
        RECT 25.240 101.775 25.480 102.175 ;
        RECT 25.960 102.005 26.180 102.285 ;
        RECT 25.650 101.835 26.180 102.005 ;
        RECT 25.650 101.605 25.820 101.835 ;
        RECT 26.350 101.675 26.520 102.455 ;
        RECT 26.690 101.845 27.040 102.465 ;
        RECT 27.210 101.845 27.420 102.635 ;
        RECT 27.610 102.665 29.110 102.835 ;
        RECT 27.610 101.975 27.780 102.665 ;
        RECT 29.470 102.495 29.640 103.275 ;
        RECT 30.445 103.145 30.615 103.275 ;
        RECT 27.950 102.325 29.640 102.495 ;
        RECT 29.810 102.715 30.275 103.105 ;
        RECT 30.445 102.975 30.840 103.145 ;
        RECT 27.950 102.145 28.120 102.325 ;
        RECT 24.750 101.435 25.820 101.605 ;
        RECT 25.990 101.225 26.180 101.665 ;
        RECT 26.350 101.395 27.300 101.675 ;
        RECT 27.610 101.585 27.870 101.975 ;
        RECT 28.290 101.905 29.080 102.155 ;
        RECT 27.520 101.415 27.870 101.585 ;
        RECT 28.080 101.225 28.410 101.685 ;
        RECT 29.285 101.615 29.455 102.325 ;
        RECT 29.810 102.125 29.980 102.715 ;
        RECT 29.625 101.905 29.980 102.125 ;
        RECT 30.150 101.905 30.500 102.525 ;
        RECT 30.670 101.615 30.840 102.975 ;
        RECT 31.205 102.805 31.530 103.590 ;
        RECT 31.010 101.755 31.470 102.805 ;
        RECT 29.285 101.445 30.140 101.615 ;
        RECT 30.345 101.445 30.840 101.615 ;
        RECT 31.010 101.225 31.340 101.585 ;
        RECT 31.700 101.485 31.870 103.605 ;
        RECT 32.040 103.275 32.370 103.775 ;
        RECT 32.540 103.105 32.795 103.605 ;
        RECT 32.045 102.935 32.795 103.105 ;
        RECT 32.045 101.945 32.275 102.935 ;
        RECT 32.445 102.115 32.795 102.765 ;
        RECT 32.970 102.685 34.640 103.775 ;
        RECT 32.970 102.165 33.720 102.685 ;
        RECT 34.810 102.610 35.100 103.775 ;
        RECT 35.730 102.685 38.320 103.775 ;
        RECT 33.890 101.995 34.640 102.515 ;
        RECT 35.730 102.165 36.940 102.685 ;
        RECT 38.550 102.635 38.760 103.775 ;
        RECT 38.930 102.625 39.260 103.605 ;
        RECT 39.430 102.635 39.660 103.775 ;
        RECT 39.870 102.685 41.080 103.775 ;
        RECT 37.110 101.995 38.320 102.515 ;
        RECT 32.045 101.775 32.795 101.945 ;
        RECT 32.040 101.225 32.370 101.605 ;
        RECT 32.540 101.485 32.795 101.775 ;
        RECT 32.970 101.225 34.640 101.995 ;
        RECT 34.810 101.225 35.100 101.950 ;
        RECT 35.730 101.225 38.320 101.995 ;
        RECT 38.550 101.225 38.760 102.045 ;
        RECT 38.930 102.025 39.180 102.625 ;
        RECT 39.350 102.215 39.680 102.465 ;
        RECT 39.870 102.145 40.390 102.685 ;
        RECT 41.290 102.635 41.520 103.775 ;
        RECT 41.690 102.625 42.020 103.605 ;
        RECT 42.190 102.635 42.400 103.775 ;
        RECT 42.630 102.685 43.840 103.775 ;
        RECT 44.010 102.685 47.520 103.775 ;
        RECT 38.930 101.395 39.260 102.025 ;
        RECT 39.430 101.225 39.660 102.045 ;
        RECT 40.560 101.975 41.080 102.515 ;
        RECT 41.270 102.215 41.600 102.465 ;
        RECT 39.870 101.225 41.080 101.975 ;
        RECT 41.290 101.225 41.520 102.045 ;
        RECT 41.770 102.025 42.020 102.625 ;
        RECT 42.630 102.145 43.150 102.685 ;
        RECT 41.690 101.395 42.020 102.025 ;
        RECT 42.190 101.225 42.400 102.045 ;
        RECT 43.320 101.975 43.840 102.515 ;
        RECT 44.010 102.165 45.700 102.685 ;
        RECT 47.690 102.610 47.980 103.775 ;
        RECT 48.610 102.685 52.120 103.775 ;
        RECT 52.295 103.340 57.640 103.775 ;
        RECT 45.870 101.995 47.520 102.515 ;
        RECT 48.610 102.165 50.300 102.685 ;
        RECT 50.470 101.995 52.120 102.515 ;
        RECT 53.885 102.090 54.235 103.340 ;
        RECT 57.850 102.635 58.080 103.775 ;
        RECT 58.250 102.625 58.580 103.605 ;
        RECT 58.750 102.635 58.960 103.775 ;
        RECT 59.230 102.635 59.460 103.775 ;
        RECT 59.630 102.625 59.960 103.605 ;
        RECT 60.130 102.635 60.340 103.775 ;
        RECT 42.630 101.225 43.840 101.975 ;
        RECT 44.010 101.225 47.520 101.995 ;
        RECT 47.690 101.225 47.980 101.950 ;
        RECT 48.610 101.225 52.120 101.995 ;
        RECT 55.715 101.770 56.055 102.600 ;
        RECT 57.830 102.215 58.160 102.465 ;
        RECT 52.295 101.225 57.640 101.770 ;
        RECT 57.850 101.225 58.080 102.045 ;
        RECT 58.330 102.025 58.580 102.625 ;
        RECT 59.210 102.215 59.540 102.465 ;
        RECT 58.250 101.395 58.580 102.025 ;
        RECT 58.750 101.225 58.960 102.045 ;
        RECT 59.230 101.225 59.460 102.045 ;
        RECT 59.710 102.025 59.960 102.625 ;
        RECT 60.570 102.610 60.860 103.775 ;
        RECT 61.030 102.685 62.700 103.775 ;
        RECT 62.875 103.105 63.130 103.605 ;
        RECT 63.300 103.275 63.630 103.775 ;
        RECT 62.875 102.935 63.625 103.105 ;
        RECT 61.030 102.165 61.780 102.685 ;
        RECT 59.630 101.395 59.960 102.025 ;
        RECT 60.130 101.225 60.340 102.045 ;
        RECT 61.950 101.995 62.700 102.515 ;
        RECT 62.875 102.115 63.225 102.765 ;
        RECT 60.570 101.225 60.860 101.950 ;
        RECT 61.030 101.225 62.700 101.995 ;
        RECT 63.395 101.945 63.625 102.935 ;
        RECT 62.875 101.775 63.625 101.945 ;
        RECT 62.875 101.485 63.130 101.775 ;
        RECT 63.300 101.225 63.630 101.605 ;
        RECT 63.800 101.485 63.970 103.605 ;
        RECT 64.140 102.805 64.465 103.590 ;
        RECT 64.635 103.315 64.885 103.775 ;
        RECT 65.055 103.275 65.305 103.605 ;
        RECT 65.520 103.275 66.200 103.605 ;
        RECT 65.055 103.145 65.225 103.275 ;
        RECT 64.830 102.975 65.225 103.145 ;
        RECT 64.200 101.755 64.660 102.805 ;
        RECT 64.830 101.615 65.000 102.975 ;
        RECT 65.395 102.715 65.860 103.105 ;
        RECT 65.170 101.905 65.520 102.525 ;
        RECT 65.690 102.125 65.860 102.715 ;
        RECT 66.030 102.495 66.200 103.275 ;
        RECT 66.370 103.175 66.540 103.515 ;
        RECT 66.775 103.345 67.105 103.775 ;
        RECT 67.275 103.175 67.445 103.515 ;
        RECT 67.740 103.315 68.110 103.775 ;
        RECT 66.370 103.005 67.445 103.175 ;
        RECT 68.280 103.145 68.450 103.605 ;
        RECT 68.685 103.265 69.555 103.605 ;
        RECT 69.725 103.315 69.975 103.775 ;
        RECT 67.890 102.975 68.450 103.145 ;
        RECT 67.890 102.835 68.060 102.975 ;
        RECT 66.560 102.665 68.060 102.835 ;
        RECT 68.755 102.805 69.215 103.095 ;
        RECT 66.030 102.325 67.720 102.495 ;
        RECT 65.690 101.905 66.045 102.125 ;
        RECT 66.215 101.615 66.385 102.325 ;
        RECT 66.590 101.905 67.380 102.155 ;
        RECT 67.550 102.145 67.720 102.325 ;
        RECT 67.890 101.975 68.060 102.665 ;
        RECT 64.330 101.225 64.660 101.585 ;
        RECT 64.830 101.445 65.325 101.615 ;
        RECT 65.530 101.445 66.385 101.615 ;
        RECT 67.260 101.225 67.590 101.685 ;
        RECT 67.800 101.585 68.060 101.975 ;
        RECT 68.250 102.795 69.215 102.805 ;
        RECT 69.385 102.885 69.555 103.265 ;
        RECT 70.145 103.225 70.315 103.515 ;
        RECT 70.495 103.395 70.825 103.775 ;
        RECT 70.145 103.055 70.945 103.225 ;
        RECT 68.250 102.635 68.925 102.795 ;
        RECT 69.385 102.715 70.605 102.885 ;
        RECT 68.250 101.845 68.460 102.635 ;
        RECT 69.385 102.625 69.555 102.715 ;
        RECT 68.630 101.845 68.980 102.465 ;
        RECT 69.150 102.455 69.555 102.625 ;
        RECT 69.150 101.675 69.320 102.455 ;
        RECT 69.490 102.005 69.710 102.285 ;
        RECT 69.890 102.175 70.430 102.545 ;
        RECT 70.775 102.435 70.945 103.055 ;
        RECT 71.120 102.715 71.290 103.775 ;
        RECT 71.500 102.765 71.790 103.605 ;
        RECT 71.960 102.935 72.130 103.775 ;
        RECT 72.340 102.765 72.590 103.605 ;
        RECT 72.800 102.935 72.970 103.775 ;
        RECT 71.500 102.595 73.225 102.765 ;
        RECT 73.450 102.610 73.740 103.775 ;
        RECT 73.910 102.685 76.500 103.775 ;
        RECT 69.490 101.835 70.020 102.005 ;
        RECT 67.800 101.415 68.150 101.585 ;
        RECT 68.370 101.395 69.320 101.675 ;
        RECT 69.490 101.225 69.680 101.665 ;
        RECT 69.850 101.605 70.020 101.835 ;
        RECT 70.190 101.775 70.430 102.175 ;
        RECT 70.600 102.425 70.945 102.435 ;
        RECT 70.600 102.215 72.630 102.425 ;
        RECT 70.600 101.960 70.925 102.215 ;
        RECT 72.815 102.045 73.225 102.595 ;
        RECT 73.910 102.165 75.120 102.685 ;
        RECT 76.710 102.635 76.940 103.775 ;
        RECT 77.110 102.625 77.440 103.605 ;
        RECT 77.610 102.635 77.820 103.775 ;
        RECT 78.050 102.685 81.560 103.775 ;
        RECT 70.600 101.605 70.920 101.960 ;
        RECT 69.850 101.435 70.920 101.605 ;
        RECT 71.120 101.225 71.290 102.035 ;
        RECT 71.460 101.875 73.225 102.045 ;
        RECT 75.290 101.995 76.500 102.515 ;
        RECT 76.690 102.215 77.020 102.465 ;
        RECT 71.460 101.395 71.790 101.875 ;
        RECT 71.960 101.225 72.130 101.695 ;
        RECT 72.300 101.395 72.630 101.875 ;
        RECT 72.800 101.225 72.970 101.695 ;
        RECT 73.450 101.225 73.740 101.950 ;
        RECT 73.910 101.225 76.500 101.995 ;
        RECT 76.710 101.225 76.940 102.045 ;
        RECT 77.190 102.025 77.440 102.625 ;
        RECT 78.050 102.165 79.740 102.685 ;
        RECT 81.790 102.635 82.000 103.775 ;
        RECT 82.170 102.625 82.500 103.605 ;
        RECT 82.670 102.635 82.900 103.775 ;
        RECT 83.570 102.685 86.160 103.775 ;
        RECT 77.110 101.395 77.440 102.025 ;
        RECT 77.610 101.225 77.820 102.045 ;
        RECT 79.910 101.995 81.560 102.515 ;
        RECT 78.050 101.225 81.560 101.995 ;
        RECT 81.790 101.225 82.000 102.045 ;
        RECT 82.170 102.025 82.420 102.625 ;
        RECT 82.590 102.215 82.920 102.465 ;
        RECT 83.570 102.165 84.780 102.685 ;
        RECT 86.330 102.610 86.620 103.775 ;
        RECT 86.790 102.685 88.460 103.775 ;
        RECT 88.940 102.935 89.110 103.775 ;
        RECT 89.320 102.765 89.570 103.605 ;
        RECT 89.780 102.935 89.950 103.775 ;
        RECT 90.120 102.765 90.410 103.605 ;
        RECT 82.170 101.395 82.500 102.025 ;
        RECT 82.670 101.225 82.900 102.045 ;
        RECT 84.950 101.995 86.160 102.515 ;
        RECT 86.790 102.165 87.540 102.685 ;
        RECT 88.685 102.595 90.410 102.765 ;
        RECT 90.620 102.715 90.790 103.775 ;
        RECT 91.085 103.395 91.415 103.775 ;
        RECT 91.595 103.225 91.765 103.515 ;
        RECT 91.935 103.315 92.185 103.775 ;
        RECT 90.965 103.055 91.765 103.225 ;
        RECT 92.355 103.265 93.225 103.605 ;
        RECT 87.710 101.995 88.460 102.515 ;
        RECT 83.570 101.225 86.160 101.995 ;
        RECT 86.330 101.225 86.620 101.950 ;
        RECT 86.790 101.225 88.460 101.995 ;
        RECT 88.685 102.045 89.095 102.595 ;
        RECT 90.965 102.435 91.135 103.055 ;
        RECT 92.355 102.885 92.525 103.265 ;
        RECT 93.460 103.145 93.630 103.605 ;
        RECT 93.800 103.315 94.170 103.775 ;
        RECT 94.465 103.175 94.635 103.515 ;
        RECT 94.805 103.345 95.135 103.775 ;
        RECT 95.370 103.175 95.540 103.515 ;
        RECT 91.305 102.715 92.525 102.885 ;
        RECT 92.695 102.805 93.155 103.095 ;
        RECT 93.460 102.975 94.020 103.145 ;
        RECT 94.465 103.005 95.540 103.175 ;
        RECT 95.710 103.275 96.390 103.605 ;
        RECT 96.605 103.275 96.855 103.605 ;
        RECT 97.025 103.315 97.275 103.775 ;
        RECT 93.850 102.835 94.020 102.975 ;
        RECT 92.695 102.795 93.660 102.805 ;
        RECT 92.355 102.625 92.525 102.715 ;
        RECT 92.985 102.635 93.660 102.795 ;
        RECT 90.965 102.425 91.310 102.435 ;
        RECT 89.280 102.215 91.310 102.425 ;
        RECT 88.685 101.875 90.450 102.045 ;
        RECT 88.940 101.225 89.110 101.695 ;
        RECT 89.280 101.395 89.610 101.875 ;
        RECT 89.780 101.225 89.950 101.695 ;
        RECT 90.120 101.395 90.450 101.875 ;
        RECT 90.620 101.225 90.790 102.035 ;
        RECT 90.985 101.960 91.310 102.215 ;
        RECT 90.990 101.605 91.310 101.960 ;
        RECT 91.480 102.175 92.020 102.545 ;
        RECT 92.355 102.455 92.760 102.625 ;
        RECT 91.480 101.775 91.720 102.175 ;
        RECT 92.200 102.005 92.420 102.285 ;
        RECT 91.890 101.835 92.420 102.005 ;
        RECT 91.890 101.605 92.060 101.835 ;
        RECT 92.590 101.675 92.760 102.455 ;
        RECT 92.930 101.845 93.280 102.465 ;
        RECT 93.450 101.845 93.660 102.635 ;
        RECT 93.850 102.665 95.350 102.835 ;
        RECT 93.850 101.975 94.020 102.665 ;
        RECT 95.710 102.495 95.880 103.275 ;
        RECT 96.685 103.145 96.855 103.275 ;
        RECT 94.190 102.325 95.880 102.495 ;
        RECT 96.050 102.715 96.515 103.105 ;
        RECT 96.685 102.975 97.080 103.145 ;
        RECT 94.190 102.145 94.360 102.325 ;
        RECT 90.990 101.435 92.060 101.605 ;
        RECT 92.230 101.225 92.420 101.665 ;
        RECT 92.590 101.395 93.540 101.675 ;
        RECT 93.850 101.585 94.110 101.975 ;
        RECT 94.530 101.905 95.320 102.155 ;
        RECT 93.760 101.415 94.110 101.585 ;
        RECT 94.320 101.225 94.650 101.685 ;
        RECT 95.525 101.615 95.695 102.325 ;
        RECT 96.050 102.125 96.220 102.715 ;
        RECT 95.865 101.905 96.220 102.125 ;
        RECT 96.390 101.905 96.740 102.525 ;
        RECT 96.910 101.615 97.080 102.975 ;
        RECT 97.445 102.805 97.770 103.590 ;
        RECT 97.250 101.755 97.710 102.805 ;
        RECT 95.525 101.445 96.380 101.615 ;
        RECT 96.585 101.445 97.080 101.615 ;
        RECT 97.250 101.225 97.580 101.585 ;
        RECT 97.940 101.485 98.110 103.605 ;
        RECT 98.280 103.275 98.610 103.775 ;
        RECT 98.780 103.105 99.035 103.605 ;
        RECT 98.285 102.935 99.035 103.105 ;
        RECT 98.285 101.945 98.515 102.935 ;
        RECT 98.685 102.115 99.035 102.765 ;
        RECT 99.210 102.610 99.500 103.775 ;
        RECT 100.900 102.935 101.070 103.775 ;
        RECT 101.280 102.765 101.530 103.605 ;
        RECT 101.740 102.935 101.910 103.775 ;
        RECT 102.080 102.765 102.370 103.605 ;
        RECT 100.645 102.595 102.370 102.765 ;
        RECT 102.580 102.715 102.750 103.775 ;
        RECT 103.045 103.395 103.375 103.775 ;
        RECT 103.555 103.225 103.725 103.515 ;
        RECT 103.895 103.315 104.145 103.775 ;
        RECT 102.925 103.055 103.725 103.225 ;
        RECT 104.315 103.265 105.185 103.605 ;
        RECT 100.645 102.045 101.055 102.595 ;
        RECT 102.925 102.435 103.095 103.055 ;
        RECT 104.315 102.885 104.485 103.265 ;
        RECT 105.420 103.145 105.590 103.605 ;
        RECT 105.760 103.315 106.130 103.775 ;
        RECT 106.425 103.175 106.595 103.515 ;
        RECT 106.765 103.345 107.095 103.775 ;
        RECT 107.330 103.175 107.500 103.515 ;
        RECT 103.265 102.715 104.485 102.885 ;
        RECT 104.655 102.805 105.115 103.095 ;
        RECT 105.420 102.975 105.980 103.145 ;
        RECT 106.425 103.005 107.500 103.175 ;
        RECT 107.670 103.275 108.350 103.605 ;
        RECT 108.565 103.275 108.815 103.605 ;
        RECT 108.985 103.315 109.235 103.775 ;
        RECT 105.810 102.835 105.980 102.975 ;
        RECT 104.655 102.795 105.620 102.805 ;
        RECT 104.315 102.625 104.485 102.715 ;
        RECT 104.945 102.635 105.620 102.795 ;
        RECT 102.925 102.425 103.270 102.435 ;
        RECT 101.240 102.215 103.270 102.425 ;
        RECT 98.285 101.775 99.035 101.945 ;
        RECT 98.280 101.225 98.610 101.605 ;
        RECT 98.780 101.485 99.035 101.775 ;
        RECT 99.210 101.225 99.500 101.950 ;
        RECT 100.645 101.875 102.410 102.045 ;
        RECT 100.900 101.225 101.070 101.695 ;
        RECT 101.240 101.395 101.570 101.875 ;
        RECT 101.740 101.225 101.910 101.695 ;
        RECT 102.080 101.395 102.410 101.875 ;
        RECT 102.580 101.225 102.750 102.035 ;
        RECT 102.945 101.960 103.270 102.215 ;
        RECT 102.950 101.605 103.270 101.960 ;
        RECT 103.440 102.175 103.980 102.545 ;
        RECT 104.315 102.455 104.720 102.625 ;
        RECT 103.440 101.775 103.680 102.175 ;
        RECT 104.160 102.005 104.380 102.285 ;
        RECT 103.850 101.835 104.380 102.005 ;
        RECT 103.850 101.605 104.020 101.835 ;
        RECT 104.550 101.675 104.720 102.455 ;
        RECT 104.890 101.845 105.240 102.465 ;
        RECT 105.410 101.845 105.620 102.635 ;
        RECT 105.810 102.665 107.310 102.835 ;
        RECT 105.810 101.975 105.980 102.665 ;
        RECT 107.670 102.495 107.840 103.275 ;
        RECT 108.645 103.145 108.815 103.275 ;
        RECT 106.150 102.325 107.840 102.495 ;
        RECT 108.010 102.715 108.475 103.105 ;
        RECT 108.645 102.975 109.040 103.145 ;
        RECT 106.150 102.145 106.320 102.325 ;
        RECT 102.950 101.435 104.020 101.605 ;
        RECT 104.190 101.225 104.380 101.665 ;
        RECT 104.550 101.395 105.500 101.675 ;
        RECT 105.810 101.585 106.070 101.975 ;
        RECT 106.490 101.905 107.280 102.155 ;
        RECT 105.720 101.415 106.070 101.585 ;
        RECT 106.280 101.225 106.610 101.685 ;
        RECT 107.485 101.615 107.655 102.325 ;
        RECT 108.010 102.125 108.180 102.715 ;
        RECT 107.825 101.905 108.180 102.125 ;
        RECT 108.350 101.905 108.700 102.525 ;
        RECT 108.870 101.615 109.040 102.975 ;
        RECT 109.405 102.805 109.730 103.590 ;
        RECT 109.210 101.755 109.670 102.805 ;
        RECT 107.485 101.445 108.340 101.615 ;
        RECT 108.545 101.445 109.040 101.615 ;
        RECT 109.210 101.225 109.540 101.585 ;
        RECT 109.900 101.485 110.070 103.605 ;
        RECT 110.240 103.275 110.570 103.775 ;
        RECT 110.740 103.105 110.995 103.605 ;
        RECT 110.245 102.935 110.995 103.105 ;
        RECT 110.245 101.945 110.475 102.935 ;
        RECT 110.645 102.115 110.995 102.765 ;
        RECT 111.170 102.685 112.380 103.775 ;
        RECT 111.170 102.145 111.690 102.685 ;
        RECT 111.860 101.975 112.380 102.515 ;
        RECT 110.245 101.775 110.995 101.945 ;
        RECT 110.240 101.225 110.570 101.605 ;
        RECT 110.740 101.485 110.995 101.775 ;
        RECT 111.170 101.225 112.380 101.975 ;
        RECT 18.165 101.055 112.465 101.225 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 17.370 193.380 112.465 193.860 ;
        RECT 102.990 192.840 103.280 192.885 ;
        RECT 105.635 192.840 105.955 192.900 ;
        RECT 106.230 192.840 106.880 192.885 ;
        RECT 102.990 192.700 106.880 192.840 ;
        RECT 102.990 192.655 103.580 192.700 ;
        RECT 20.535 192.300 20.855 192.560 ;
        RECT 28.355 192.500 28.675 192.560 ;
        RECT 30.670 192.500 30.960 192.545 ;
        RECT 28.355 192.360 30.960 192.500 ;
        RECT 28.355 192.300 28.675 192.360 ;
        RECT 30.670 192.315 30.960 192.360 ;
        RECT 43.995 192.300 44.315 192.560 ;
        RECT 44.915 192.500 45.235 192.560 ;
        RECT 46.770 192.500 47.060 192.545 ;
        RECT 44.915 192.360 47.060 192.500 ;
        RECT 44.915 192.300 45.235 192.360 ;
        RECT 46.770 192.315 47.060 192.360 ;
        RECT 51.355 192.500 51.675 192.560 ;
        RECT 52.750 192.500 53.040 192.545 ;
        RECT 64.710 192.500 65.000 192.545 ;
        RECT 66.550 192.500 66.840 192.545 ;
        RECT 70.215 192.500 70.535 192.560 ;
        RECT 51.355 192.360 70.535 192.500 ;
        RECT 51.355 192.300 51.675 192.360 ;
        RECT 52.750 192.315 53.040 192.360 ;
        RECT 64.710 192.315 65.000 192.360 ;
        RECT 66.550 192.315 66.840 192.360 ;
        RECT 70.215 192.300 70.535 192.360 ;
        RECT 75.275 192.500 75.595 192.560 ;
        RECT 78.050 192.500 78.340 192.545 ;
        RECT 75.275 192.360 78.340 192.500 ;
        RECT 75.275 192.300 75.595 192.360 ;
        RECT 78.050 192.315 78.340 192.360 ;
        RECT 87.695 192.500 88.015 192.560 ;
        RECT 89.550 192.500 89.840 192.545 ;
        RECT 87.695 192.360 89.840 192.500 ;
        RECT 87.695 192.300 88.015 192.360 ;
        RECT 89.550 192.315 89.840 192.360 ;
        RECT 94.595 192.500 94.915 192.560 ;
        RECT 96.450 192.500 96.740 192.545 ;
        RECT 94.595 192.360 96.740 192.500 ;
        RECT 94.595 192.300 94.915 192.360 ;
        RECT 96.450 192.315 96.740 192.360 ;
        RECT 98.735 192.500 99.055 192.560 ;
        RECT 99.670 192.500 99.960 192.545 ;
        RECT 98.735 192.360 99.960 192.500 ;
        RECT 98.735 192.300 99.055 192.360 ;
        RECT 99.670 192.315 99.960 192.360 ;
        RECT 103.290 192.340 103.580 192.655 ;
        RECT 105.635 192.640 105.955 192.700 ;
        RECT 106.230 192.655 106.880 192.700 ;
        RECT 108.855 192.640 109.175 192.900 ;
        RECT 104.370 192.500 104.660 192.545 ;
        RECT 107.950 192.500 108.240 192.545 ;
        RECT 109.785 192.500 110.075 192.545 ;
        RECT 104.370 192.360 110.075 192.500 ;
        RECT 104.370 192.315 104.660 192.360 ;
        RECT 107.950 192.315 108.240 192.360 ;
        RECT 109.785 192.315 110.075 192.360 ;
        RECT 75.735 192.160 76.055 192.220 ;
        RECT 76.670 192.160 76.960 192.205 ;
        RECT 75.735 192.020 76.960 192.160 ;
        RECT 75.735 191.960 76.055 192.020 ;
        RECT 76.670 191.975 76.960 192.020 ;
        RECT 77.590 192.160 77.880 192.205 ;
        RECT 78.495 192.160 78.815 192.220 ;
        RECT 77.590 192.020 78.815 192.160 ;
        RECT 77.590 191.975 77.880 192.020 ;
        RECT 78.495 191.960 78.815 192.020 ;
        RECT 108.395 192.160 108.715 192.220 ;
        RECT 110.250 192.160 110.540 192.205 ;
        RECT 108.395 192.020 110.540 192.160 ;
        RECT 108.395 191.960 108.715 192.020 ;
        RECT 110.250 191.975 110.540 192.020 ;
        RECT 101.510 191.820 101.800 191.865 ;
        RECT 101.955 191.820 102.275 191.880 ;
        RECT 101.510 191.680 102.275 191.820 ;
        RECT 101.510 191.635 101.800 191.680 ;
        RECT 101.955 191.620 102.275 191.680 ;
        RECT 104.370 191.820 104.660 191.865 ;
        RECT 107.490 191.820 107.780 191.865 ;
        RECT 109.380 191.820 109.670 191.865 ;
        RECT 104.370 191.680 109.670 191.820 ;
        RECT 104.370 191.635 104.660 191.680 ;
        RECT 107.490 191.635 107.780 191.680 ;
        RECT 109.380 191.635 109.670 191.680 ;
        RECT 20.995 191.280 21.315 191.540 ;
        RECT 31.575 191.280 31.895 191.540 ;
        RECT 43.535 191.280 43.855 191.540 ;
        RECT 44.455 191.480 44.775 191.540 ;
        RECT 45.850 191.480 46.140 191.525 ;
        RECT 44.455 191.340 46.140 191.480 ;
        RECT 44.455 191.280 44.775 191.340 ;
        RECT 45.850 191.295 46.140 191.340 ;
        RECT 52.275 191.280 52.595 191.540 ;
        RECT 64.250 191.480 64.540 191.525 ;
        RECT 64.695 191.480 65.015 191.540 ;
        RECT 64.250 191.340 65.015 191.480 ;
        RECT 64.250 191.295 64.540 191.340 ;
        RECT 64.695 191.280 65.015 191.340 ;
        RECT 66.090 191.480 66.380 191.525 ;
        RECT 66.535 191.480 66.855 191.540 ;
        RECT 66.090 191.340 66.855 191.480 ;
        RECT 66.090 191.295 66.380 191.340 ;
        RECT 66.535 191.280 66.855 191.340 ;
        RECT 79.890 191.480 80.180 191.525 ;
        RECT 82.635 191.480 82.955 191.540 ;
        RECT 79.890 191.340 82.955 191.480 ;
        RECT 79.890 191.295 80.180 191.340 ;
        RECT 82.635 191.280 82.955 191.340 ;
        RECT 88.615 191.280 88.935 191.540 ;
        RECT 96.910 191.480 97.200 191.525 ;
        RECT 97.815 191.480 98.135 191.540 ;
        RECT 96.910 191.340 98.135 191.480 ;
        RECT 96.910 191.295 97.200 191.340 ;
        RECT 97.815 191.280 98.135 191.340 ;
        RECT 100.590 191.480 100.880 191.525 ;
        RECT 103.335 191.480 103.655 191.540 ;
        RECT 100.590 191.340 103.655 191.480 ;
        RECT 100.590 191.295 100.880 191.340 ;
        RECT 103.335 191.280 103.655 191.340 ;
        RECT 18.165 190.660 112.465 191.140 ;
        RECT 27.090 190.120 27.380 190.165 ;
        RECT 30.210 190.120 30.500 190.165 ;
        RECT 32.100 190.120 32.390 190.165 ;
        RECT 27.090 189.980 32.390 190.120 ;
        RECT 27.090 189.935 27.380 189.980 ;
        RECT 30.210 189.935 30.500 189.980 ;
        RECT 32.100 189.935 32.390 189.980 ;
        RECT 40.285 190.120 40.575 190.165 ;
        RECT 43.065 190.120 43.355 190.165 ;
        RECT 44.925 190.120 45.215 190.165 ;
        RECT 40.285 189.980 45.215 190.120 ;
        RECT 40.285 189.935 40.575 189.980 ;
        RECT 43.065 189.935 43.355 189.980 ;
        RECT 44.925 189.935 45.215 189.980 ;
        RECT 48.560 190.120 48.850 190.165 ;
        RECT 50.450 190.120 50.740 190.165 ;
        RECT 53.570 190.120 53.860 190.165 ;
        RECT 48.560 189.980 53.860 190.120 ;
        RECT 48.560 189.935 48.850 189.980 ;
        RECT 50.450 189.935 50.740 189.980 ;
        RECT 53.570 189.935 53.860 189.980 ;
        RECT 63.890 190.120 64.180 190.165 ;
        RECT 67.010 190.120 67.300 190.165 ;
        RECT 68.900 190.120 69.190 190.165 ;
        RECT 63.890 189.980 69.190 190.120 ;
        RECT 63.890 189.935 64.180 189.980 ;
        RECT 67.010 189.935 67.300 189.980 ;
        RECT 68.900 189.935 69.190 189.980 ;
        RECT 78.005 190.120 78.295 190.165 ;
        RECT 80.785 190.120 81.075 190.165 ;
        RECT 82.645 190.120 82.935 190.165 ;
        RECT 78.005 189.980 82.935 190.120 ;
        RECT 78.005 189.935 78.295 189.980 ;
        RECT 80.785 189.935 81.075 189.980 ;
        RECT 82.645 189.935 82.935 189.980 ;
        RECT 87.660 190.120 87.950 190.165 ;
        RECT 89.550 190.120 89.840 190.165 ;
        RECT 92.670 190.120 92.960 190.165 ;
        RECT 87.660 189.980 92.960 190.120 ;
        RECT 87.660 189.935 87.950 189.980 ;
        RECT 89.550 189.935 89.840 189.980 ;
        RECT 92.670 189.935 92.960 189.980 ;
        RECT 95.530 189.935 95.820 190.165 ;
        RECT 98.850 190.120 99.140 190.165 ;
        RECT 101.970 190.120 102.260 190.165 ;
        RECT 103.860 190.120 104.150 190.165 ;
        RECT 98.850 189.980 104.150 190.120 ;
        RECT 98.850 189.935 99.140 189.980 ;
        RECT 101.970 189.935 102.260 189.980 ;
        RECT 103.860 189.935 104.150 189.980 ;
        RECT 21.010 189.780 21.300 189.825 ;
        RECT 23.755 189.780 24.075 189.840 ;
        RECT 21.010 189.640 24.075 189.780 ;
        RECT 21.010 189.595 21.300 189.640 ;
        RECT 23.755 189.580 24.075 189.640 ;
        RECT 24.230 189.595 24.520 189.825 ;
        RECT 24.305 189.440 24.445 189.595 ;
        RECT 31.575 189.580 31.895 189.840 ;
        RECT 32.955 189.580 33.275 189.840 ;
        RECT 43.550 189.780 43.840 189.825 ;
        RECT 44.455 189.780 44.775 189.840 ;
        RECT 43.550 189.640 44.775 189.780 ;
        RECT 43.550 189.595 43.840 189.640 ;
        RECT 44.455 189.580 44.775 189.640 ;
        RECT 45.390 189.780 45.680 189.825 ;
        RECT 45.835 189.780 46.155 189.840 ;
        RECT 47.690 189.780 47.980 189.825 ;
        RECT 45.390 189.640 47.980 189.780 ;
        RECT 45.390 189.595 45.680 189.640 ;
        RECT 45.835 189.580 46.155 189.640 ;
        RECT 47.690 189.595 47.980 189.640 ;
        RECT 62.395 189.780 62.715 189.840 ;
        RECT 68.390 189.780 68.680 189.825 ;
        RECT 83.110 189.780 83.400 189.825 ;
        RECT 83.555 189.780 83.875 189.840 ;
        RECT 86.790 189.780 87.080 189.825 ;
        RECT 62.395 189.640 68.680 189.780 ;
        RECT 62.395 189.580 62.715 189.640 ;
        RECT 68.390 189.595 68.680 189.640 ;
        RECT 77.665 189.640 82.405 189.780 ;
        RECT 25.135 189.440 25.455 189.500 ;
        RECT 24.305 189.300 25.455 189.440 ;
        RECT 25.135 189.240 25.455 189.300 ;
        RECT 20.995 189.100 21.315 189.160 ;
        RECT 26.010 189.145 26.300 189.460 ;
        RECT 27.090 189.440 27.380 189.485 ;
        RECT 30.670 189.440 30.960 189.485 ;
        RECT 32.505 189.440 32.795 189.485 ;
        RECT 27.090 189.300 32.795 189.440 ;
        RECT 27.090 189.255 27.380 189.300 ;
        RECT 30.670 189.255 30.960 189.300 ;
        RECT 32.505 189.255 32.795 189.300 ;
        RECT 40.285 189.440 40.575 189.485 ;
        RECT 40.285 189.300 42.820 189.440 ;
        RECT 40.285 189.255 40.575 189.300 ;
        RECT 38.475 189.145 38.795 189.160 ;
        RECT 42.605 189.145 42.820 189.300 ;
        RECT 47.215 189.240 47.535 189.500 ;
        RECT 48.155 189.440 48.445 189.485 ;
        RECT 49.990 189.440 50.280 189.485 ;
        RECT 53.570 189.440 53.860 189.485 ;
        RECT 48.155 189.300 53.860 189.440 ;
        RECT 48.155 189.255 48.445 189.300 ;
        RECT 49.990 189.255 50.280 189.300 ;
        RECT 53.570 189.255 53.860 189.300 ;
        RECT 25.710 189.100 26.300 189.145 ;
        RECT 28.950 189.100 29.600 189.145 ;
        RECT 20.995 188.960 29.600 189.100 ;
        RECT 20.995 188.900 21.315 188.960 ;
        RECT 25.710 188.915 26.000 188.960 ;
        RECT 28.950 188.915 29.600 188.960 ;
        RECT 38.425 189.100 38.795 189.145 ;
        RECT 41.685 189.100 41.975 189.145 ;
        RECT 38.425 188.960 41.975 189.100 ;
        RECT 38.425 188.915 38.795 188.960 ;
        RECT 41.685 188.915 41.975 188.960 ;
        RECT 42.605 189.100 42.895 189.145 ;
        RECT 44.465 189.100 44.755 189.145 ;
        RECT 42.605 188.960 44.755 189.100 ;
        RECT 42.605 188.915 42.895 188.960 ;
        RECT 44.465 188.915 44.755 188.960 ;
        RECT 49.070 189.100 49.360 189.145 ;
        RECT 49.515 189.100 49.835 189.160 ;
        RECT 49.070 188.960 49.835 189.100 ;
        RECT 49.070 188.915 49.360 188.960 ;
        RECT 38.475 188.900 38.795 188.915 ;
        RECT 49.515 188.900 49.835 188.960 ;
        RECT 51.350 189.100 52.000 189.145 ;
        RECT 52.275 189.100 52.595 189.160 ;
        RECT 54.650 189.145 54.940 189.460 ;
        RECT 62.810 189.145 63.100 189.460 ;
        RECT 63.890 189.440 64.180 189.485 ;
        RECT 67.470 189.440 67.760 189.485 ;
        RECT 69.305 189.440 69.595 189.485 ;
        RECT 63.890 189.300 69.595 189.440 ;
        RECT 63.890 189.255 64.180 189.300 ;
        RECT 67.470 189.255 67.760 189.300 ;
        RECT 69.305 189.255 69.595 189.300 ;
        RECT 69.755 189.240 70.075 189.500 ;
        RECT 70.215 189.440 70.535 189.500 ;
        RECT 77.665 189.440 77.805 189.640 ;
        RECT 70.215 189.300 77.805 189.440 ;
        RECT 78.005 189.440 78.295 189.485 ;
        RECT 81.270 189.440 81.560 189.485 ;
        RECT 81.715 189.440 82.035 189.500 ;
        RECT 78.005 189.300 80.540 189.440 ;
        RECT 70.215 189.240 70.535 189.300 ;
        RECT 78.005 189.255 78.295 189.300 ;
        RECT 54.650 189.100 55.240 189.145 ;
        RECT 51.350 188.960 55.240 189.100 ;
        RECT 51.350 188.915 52.000 188.960 ;
        RECT 52.275 188.900 52.595 188.960 ;
        RECT 54.950 188.915 55.240 188.960 ;
        RECT 62.510 189.100 63.100 189.145 ;
        RECT 64.695 189.100 65.015 189.160 ;
        RECT 65.750 189.100 66.400 189.145 ;
        RECT 62.510 188.960 66.400 189.100 ;
        RECT 62.510 188.915 62.800 188.960 ;
        RECT 64.695 188.900 65.015 188.960 ;
        RECT 65.750 188.915 66.400 188.960 ;
        RECT 74.815 189.100 75.135 189.160 ;
        RECT 80.325 189.145 80.540 189.300 ;
        RECT 81.270 189.300 82.035 189.440 ;
        RECT 82.265 189.440 82.405 189.640 ;
        RECT 83.110 189.640 87.080 189.780 ;
        RECT 83.110 189.595 83.400 189.640 ;
        RECT 83.555 189.580 83.875 189.640 ;
        RECT 86.790 189.595 87.080 189.640 ;
        RECT 88.170 189.780 88.460 189.825 ;
        RECT 88.615 189.780 88.935 189.840 ;
        RECT 88.170 189.640 88.935 189.780 ;
        RECT 88.170 189.595 88.460 189.640 ;
        RECT 88.615 189.580 88.935 189.640 ;
        RECT 95.605 189.500 95.745 189.935 ;
        RECT 103.335 189.580 103.655 189.840 ;
        RECT 104.730 189.780 105.020 189.825 ;
        RECT 108.395 189.780 108.715 189.840 ;
        RECT 104.730 189.640 108.715 189.780 ;
        RECT 104.730 189.595 105.020 189.640 ;
        RECT 108.395 189.580 108.715 189.640 ;
        RECT 84.950 189.440 85.240 189.485 ;
        RECT 82.265 189.300 85.240 189.440 ;
        RECT 81.270 189.255 81.560 189.300 ;
        RECT 81.715 189.240 82.035 189.300 ;
        RECT 84.950 189.255 85.240 189.300 ;
        RECT 87.255 189.440 87.545 189.485 ;
        RECT 89.090 189.440 89.380 189.485 ;
        RECT 92.670 189.440 92.960 189.485 ;
        RECT 87.255 189.300 92.960 189.440 ;
        RECT 87.255 189.255 87.545 189.300 ;
        RECT 89.090 189.255 89.380 189.300 ;
        RECT 92.670 189.255 92.960 189.300 ;
        RECT 76.145 189.100 76.435 189.145 ;
        RECT 79.405 189.100 79.695 189.145 ;
        RECT 74.815 188.960 79.695 189.100 ;
        RECT 74.815 188.900 75.135 188.960 ;
        RECT 76.145 188.915 76.435 188.960 ;
        RECT 79.405 188.915 79.695 188.960 ;
        RECT 80.325 189.100 80.615 189.145 ;
        RECT 82.185 189.100 82.475 189.145 ;
        RECT 80.325 188.960 82.475 189.100 ;
        RECT 80.325 188.915 80.615 188.960 ;
        RECT 82.185 188.915 82.475 188.960 ;
        RECT 23.770 188.760 24.060 188.805 ;
        RECT 26.515 188.760 26.835 188.820 ;
        RECT 23.770 188.620 26.835 188.760 ;
        RECT 23.770 188.575 24.060 188.620 ;
        RECT 26.515 188.560 26.835 188.620 ;
        RECT 36.420 188.760 36.710 188.805 ;
        RECT 40.315 188.760 40.635 188.820 ;
        RECT 36.420 188.620 40.635 188.760 ;
        RECT 36.420 188.575 36.710 188.620 ;
        RECT 40.315 188.560 40.635 188.620 ;
        RECT 45.375 188.760 45.695 188.820 ;
        RECT 46.310 188.760 46.600 188.805 ;
        RECT 45.375 188.620 46.600 188.760 ;
        RECT 45.375 188.560 45.695 188.620 ;
        RECT 46.310 188.575 46.600 188.620 ;
        RECT 56.415 188.560 56.735 188.820 ;
        RECT 61.030 188.760 61.320 188.805 ;
        RECT 61.475 188.760 61.795 188.820 ;
        RECT 61.030 188.620 61.795 188.760 ;
        RECT 61.030 188.575 61.320 188.620 ;
        RECT 61.475 188.560 61.795 188.620 ;
        RECT 74.140 188.760 74.430 188.805 ;
        RECT 78.495 188.760 78.815 188.820 ;
        RECT 74.140 188.620 78.815 188.760 ;
        RECT 85.025 188.760 85.165 189.255 ;
        RECT 93.750 189.145 94.040 189.460 ;
        RECT 94.595 189.440 94.915 189.500 ;
        RECT 94.595 189.300 95.285 189.440 ;
        RECT 94.595 189.240 94.915 189.300 ;
        RECT 85.410 189.100 85.700 189.145 ;
        RECT 90.450 189.100 91.100 189.145 ;
        RECT 93.750 189.100 94.340 189.145 ;
        RECT 85.410 188.960 94.340 189.100 ;
        RECT 95.145 189.100 95.285 189.300 ;
        RECT 95.515 189.240 95.835 189.500 ;
        RECT 95.975 189.240 96.295 189.500 ;
        RECT 97.815 189.460 98.135 189.500 ;
        RECT 97.770 189.240 98.135 189.460 ;
        RECT 98.850 189.440 99.140 189.485 ;
        RECT 102.430 189.440 102.720 189.485 ;
        RECT 104.265 189.440 104.555 189.485 ;
        RECT 98.850 189.300 104.555 189.440 ;
        RECT 98.850 189.255 99.140 189.300 ;
        RECT 102.430 189.255 102.720 189.300 ;
        RECT 104.265 189.255 104.555 189.300 ;
        RECT 105.190 189.255 105.480 189.485 ;
        RECT 96.065 189.100 96.205 189.240 ;
        RECT 97.770 189.145 98.060 189.240 ;
        RECT 97.470 189.100 98.060 189.145 ;
        RECT 100.710 189.100 101.360 189.145 ;
        RECT 95.145 188.960 97.125 189.100 ;
        RECT 85.410 188.915 85.700 188.960 ;
        RECT 90.450 188.915 91.100 188.960 ;
        RECT 94.050 188.915 94.340 188.960 ;
        RECT 93.215 188.760 93.535 188.820 ;
        RECT 85.025 188.620 93.535 188.760 ;
        RECT 74.140 188.575 74.430 188.620 ;
        RECT 78.495 188.560 78.815 188.620 ;
        RECT 93.215 188.560 93.535 188.620 ;
        RECT 95.055 188.760 95.375 188.820 ;
        RECT 95.990 188.760 96.280 188.805 ;
        RECT 95.055 188.620 96.280 188.760 ;
        RECT 96.985 188.760 97.125 188.960 ;
        RECT 97.470 188.960 101.360 189.100 ;
        RECT 97.470 188.915 97.760 188.960 ;
        RECT 100.710 188.915 101.360 188.960 ;
        RECT 105.265 188.820 105.405 189.255 ;
        RECT 105.635 189.240 105.955 189.500 ;
        RECT 105.175 188.760 105.495 188.820 ;
        RECT 96.985 188.620 105.495 188.760 ;
        RECT 95.055 188.560 95.375 188.620 ;
        RECT 95.990 188.575 96.280 188.620 ;
        RECT 105.175 188.560 105.495 188.620 ;
        RECT 17.370 187.940 112.465 188.420 ;
        RECT 26.515 187.540 26.835 187.800 ;
        RECT 28.355 187.540 28.675 187.800 ;
        RECT 28.830 187.555 29.120 187.785 ;
        RECT 49.515 187.740 49.835 187.800 ;
        RECT 49.990 187.740 50.280 187.785 ;
        RECT 49.515 187.600 50.280 187.740 ;
        RECT 20.535 187.060 20.855 187.120 ;
        RECT 23.310 187.060 23.600 187.105 ;
        RECT 20.535 186.920 23.600 187.060 ;
        RECT 20.535 186.860 20.855 186.920 ;
        RECT 23.310 186.875 23.600 186.920 ;
        RECT 24.215 187.060 24.535 187.120 ;
        RECT 28.905 187.060 29.045 187.555 ;
        RECT 49.515 187.540 49.835 187.600 ;
        RECT 49.990 187.555 50.280 187.600 ;
        RECT 62.395 187.540 62.715 187.800 ;
        RECT 78.495 187.740 78.815 187.800 ;
        RECT 78.495 187.600 83.325 187.740 ;
        RECT 78.495 187.540 78.815 187.600 ;
        RECT 30.310 187.400 30.600 187.445 ;
        RECT 33.550 187.400 34.200 187.445 ;
        RECT 30.310 187.260 34.200 187.400 ;
        RECT 30.310 187.215 30.900 187.260 ;
        RECT 33.550 187.215 34.200 187.260 ;
        RECT 24.215 186.920 29.045 187.060 ;
        RECT 24.215 186.860 24.535 186.920 ;
        RECT 30.610 186.900 30.900 187.215 ;
        RECT 36.175 187.200 36.495 187.460 ;
        RECT 43.535 187.445 43.855 187.460 ;
        RECT 40.265 187.400 40.555 187.445 ;
        RECT 43.525 187.400 43.855 187.445 ;
        RECT 40.265 187.260 43.855 187.400 ;
        RECT 40.265 187.215 40.555 187.260 ;
        RECT 43.525 187.215 43.855 187.260 ;
        RECT 43.535 187.200 43.855 187.215 ;
        RECT 44.445 187.400 44.735 187.445 ;
        RECT 46.305 187.400 46.595 187.445 ;
        RECT 44.445 187.260 46.595 187.400 ;
        RECT 44.445 187.215 44.735 187.260 ;
        RECT 46.305 187.215 46.595 187.260 ;
        RECT 64.350 187.400 64.640 187.445 ;
        RECT 66.535 187.400 66.855 187.460 ;
        RECT 67.590 187.400 68.240 187.445 ;
        RECT 64.350 187.260 68.240 187.400 ;
        RECT 64.350 187.215 64.940 187.260 ;
        RECT 31.690 187.060 31.980 187.105 ;
        RECT 35.270 187.060 35.560 187.105 ;
        RECT 37.105 187.060 37.395 187.105 ;
        RECT 31.690 186.920 37.395 187.060 ;
        RECT 25.595 186.520 25.915 186.780 ;
        RECT 26.055 186.720 26.375 186.780 ;
        RECT 27.435 186.720 27.755 186.780 ;
        RECT 26.055 186.580 27.755 186.720 ;
        RECT 26.055 186.520 26.375 186.580 ;
        RECT 27.435 186.520 27.755 186.580 ;
        RECT 23.770 186.380 24.060 186.425 ;
        RECT 30.745 186.380 30.885 186.900 ;
        RECT 31.690 186.875 31.980 186.920 ;
        RECT 35.270 186.875 35.560 186.920 ;
        RECT 37.105 186.875 37.395 186.920 ;
        RECT 42.125 187.060 42.415 187.105 ;
        RECT 44.445 187.060 44.660 187.215 ;
        RECT 42.125 186.920 44.660 187.060 ;
        RECT 42.125 186.875 42.415 186.920 ;
        RECT 45.375 186.860 45.695 187.120 ;
        RECT 49.530 187.060 49.820 187.105 ;
        RECT 51.355 187.060 51.675 187.120 ;
        RECT 49.530 186.920 51.675 187.060 ;
        RECT 49.530 186.875 49.820 186.920 ;
        RECT 51.355 186.860 51.675 186.920 ;
        RECT 51.830 187.060 52.120 187.105 ;
        RECT 53.210 187.060 53.500 187.105 ;
        RECT 51.830 186.920 53.500 187.060 ;
        RECT 51.830 186.875 52.120 186.920 ;
        RECT 53.210 186.875 53.500 186.920 ;
        RECT 58.270 187.060 58.560 187.105 ;
        RECT 59.175 187.060 59.495 187.120 ;
        RECT 58.270 186.920 59.495 187.060 ;
        RECT 58.270 186.875 58.560 186.920 ;
        RECT 59.175 186.860 59.495 186.920 ;
        RECT 61.490 187.060 61.780 187.105 ;
        RECT 61.935 187.060 62.255 187.120 ;
        RECT 61.490 186.920 62.255 187.060 ;
        RECT 61.490 186.875 61.780 186.920 ;
        RECT 61.935 186.860 62.255 186.920 ;
        RECT 64.650 186.900 64.940 187.215 ;
        RECT 66.535 187.200 66.855 187.260 ;
        RECT 67.590 187.215 68.240 187.260 ;
        RECT 72.530 187.400 72.820 187.445 ;
        RECT 76.605 187.400 76.895 187.445 ;
        RECT 79.865 187.400 80.155 187.445 ;
        RECT 72.530 187.260 80.155 187.400 ;
        RECT 72.530 187.215 72.820 187.260 ;
        RECT 76.605 187.215 76.895 187.260 ;
        RECT 79.865 187.215 80.155 187.260 ;
        RECT 80.785 187.400 81.075 187.445 ;
        RECT 82.645 187.400 82.935 187.445 ;
        RECT 80.785 187.260 82.935 187.400 ;
        RECT 83.185 187.400 83.325 187.600 ;
        RECT 87.695 187.540 88.015 187.800 ;
        RECT 98.735 187.540 99.055 187.800 ;
        RECT 107.030 187.740 107.320 187.785 ;
        RECT 108.855 187.740 109.175 187.800 ;
        RECT 107.030 187.600 109.175 187.740 ;
        RECT 107.030 187.555 107.320 187.600 ;
        RECT 108.855 187.540 109.175 187.600 ;
        RECT 85.870 187.400 86.160 187.445 ;
        RECT 95.515 187.400 95.835 187.460 ;
        RECT 96.910 187.400 97.200 187.445 ;
        RECT 83.185 187.260 86.160 187.400 ;
        RECT 80.785 187.215 81.075 187.260 ;
        RECT 82.645 187.215 82.935 187.260 ;
        RECT 85.870 187.215 86.160 187.260 ;
        RECT 89.625 187.260 97.200 187.400 ;
        RECT 65.730 187.060 66.020 187.105 ;
        RECT 69.310 187.060 69.600 187.105 ;
        RECT 71.145 187.060 71.435 187.105 ;
        RECT 65.730 186.920 71.435 187.060 ;
        RECT 65.730 186.875 66.020 186.920 ;
        RECT 69.310 186.875 69.600 186.920 ;
        RECT 71.145 186.875 71.435 186.920 ;
        RECT 72.990 187.060 73.280 187.105 ;
        RECT 74.355 187.060 74.675 187.120 ;
        RECT 72.990 186.920 74.675 187.060 ;
        RECT 72.990 186.875 73.280 186.920 ;
        RECT 74.355 186.860 74.675 186.920 ;
        RECT 78.465 187.060 78.755 187.105 ;
        RECT 80.785 187.060 81.000 187.215 ;
        RECT 78.465 186.920 81.000 187.060 ;
        RECT 81.255 187.060 81.575 187.120 ;
        RECT 81.730 187.060 82.020 187.105 ;
        RECT 81.255 186.920 82.020 187.060 ;
        RECT 78.465 186.875 78.755 186.920 ;
        RECT 81.255 186.860 81.575 186.920 ;
        RECT 81.730 186.875 82.020 186.920 ;
        RECT 85.410 187.060 85.700 187.105 ;
        RECT 89.625 187.060 89.765 187.260 ;
        RECT 95.515 187.200 95.835 187.260 ;
        RECT 96.910 187.215 97.200 187.260 ;
        RECT 85.410 186.920 89.765 187.060 ;
        RECT 89.995 187.060 90.315 187.120 ;
        RECT 90.470 187.060 90.760 187.105 ;
        RECT 89.995 186.920 90.760 187.060 ;
        RECT 85.410 186.875 85.700 186.920 ;
        RECT 89.995 186.860 90.315 186.920 ;
        RECT 90.470 186.875 90.760 186.920 ;
        RECT 93.215 186.860 93.535 187.120 ;
        RECT 94.595 187.060 94.915 187.120 ;
        RECT 96.450 187.060 96.740 187.105 ;
        RECT 101.510 187.060 101.800 187.105 ;
        RECT 106.110 187.060 106.400 187.105 ;
        RECT 94.595 186.920 101.800 187.060 ;
        RECT 94.595 186.860 94.915 186.920 ;
        RECT 96.450 186.875 96.740 186.920 ;
        RECT 101.510 186.875 101.800 186.920 ;
        RECT 103.425 186.920 106.400 187.060 ;
        RECT 31.115 186.720 31.435 186.780 ;
        RECT 37.570 186.720 37.860 186.765 ;
        RECT 45.835 186.720 46.155 186.780 ;
        RECT 47.230 186.720 47.520 186.765 ;
        RECT 31.115 186.580 47.520 186.720 ;
        RECT 31.115 186.520 31.435 186.580 ;
        RECT 37.570 186.535 37.860 186.580 ;
        RECT 45.835 186.520 46.155 186.580 ;
        RECT 47.230 186.535 47.520 186.580 ;
        RECT 52.290 186.720 52.580 186.765 ;
        RECT 55.955 186.720 56.275 186.780 ;
        RECT 52.290 186.580 56.275 186.720 ;
        RECT 52.290 186.535 52.580 186.580 ;
        RECT 23.770 186.240 30.885 186.380 ;
        RECT 31.690 186.380 31.980 186.425 ;
        RECT 34.810 186.380 35.100 186.425 ;
        RECT 36.700 186.380 36.990 186.425 ;
        RECT 31.690 186.240 36.990 186.380 ;
        RECT 23.770 186.195 24.060 186.240 ;
        RECT 31.690 186.195 31.980 186.240 ;
        RECT 34.810 186.195 35.100 186.240 ;
        RECT 36.700 186.195 36.990 186.240 ;
        RECT 42.125 186.380 42.415 186.425 ;
        RECT 44.905 186.380 45.195 186.425 ;
        RECT 46.765 186.380 47.055 186.425 ;
        RECT 42.125 186.240 47.055 186.380 ;
        RECT 47.305 186.380 47.445 186.535 ;
        RECT 55.955 186.520 56.275 186.580 ;
        RECT 56.415 186.520 56.735 186.780 ;
        RECT 59.650 186.720 59.940 186.765 ;
        RECT 60.095 186.720 60.415 186.780 ;
        RECT 64.235 186.720 64.555 186.780 ;
        RECT 59.650 186.580 64.555 186.720 ;
        RECT 59.650 186.535 59.940 186.580 ;
        RECT 60.095 186.520 60.415 186.580 ;
        RECT 64.235 186.520 64.555 186.580 ;
        RECT 69.755 186.720 70.075 186.780 ;
        RECT 71.610 186.720 71.900 186.765 ;
        RECT 83.555 186.720 83.875 186.780 ;
        RECT 84.490 186.720 84.780 186.765 ;
        RECT 93.675 186.720 93.995 186.780 ;
        RECT 95.530 186.720 95.820 186.765 ;
        RECT 100.130 186.720 100.420 186.765 ;
        RECT 69.755 186.580 83.875 186.720 ;
        RECT 69.755 186.520 70.075 186.580 ;
        RECT 71.610 186.535 71.900 186.580 ;
        RECT 83.555 186.520 83.875 186.580 ;
        RECT 84.105 186.580 100.420 186.720 ;
        RECT 54.575 186.380 54.895 186.440 ;
        RECT 47.305 186.240 54.895 186.380 ;
        RECT 56.505 186.380 56.645 186.520 ;
        RECT 63.775 186.380 64.095 186.440 ;
        RECT 56.505 186.240 64.095 186.380 ;
        RECT 42.125 186.195 42.415 186.240 ;
        RECT 44.905 186.195 45.195 186.240 ;
        RECT 46.765 186.195 47.055 186.240 ;
        RECT 54.575 186.180 54.895 186.240 ;
        RECT 21.010 186.040 21.300 186.085 ;
        RECT 24.675 186.040 24.995 186.100 ;
        RECT 21.010 185.900 24.995 186.040 ;
        RECT 21.010 185.855 21.300 185.900 ;
        RECT 24.675 185.840 24.995 185.900 ;
        RECT 38.260 186.040 38.550 186.085 ;
        RECT 40.775 186.040 41.095 186.100 ;
        RECT 38.260 185.900 41.095 186.040 ;
        RECT 38.260 185.855 38.550 185.900 ;
        RECT 40.775 185.840 41.095 185.900 ;
        RECT 49.055 185.840 49.375 186.100 ;
        RECT 59.725 186.085 59.865 186.240 ;
        RECT 63.775 186.180 64.095 186.240 ;
        RECT 65.730 186.380 66.020 186.425 ;
        RECT 68.850 186.380 69.140 186.425 ;
        RECT 70.740 186.380 71.030 186.425 ;
        RECT 65.730 186.240 71.030 186.380 ;
        RECT 65.730 186.195 66.020 186.240 ;
        RECT 68.850 186.195 69.140 186.240 ;
        RECT 70.740 186.195 71.030 186.240 ;
        RECT 78.465 186.380 78.755 186.425 ;
        RECT 81.245 186.380 81.535 186.425 ;
        RECT 83.105 186.380 83.395 186.425 ;
        RECT 78.465 186.240 83.395 186.380 ;
        RECT 78.465 186.195 78.755 186.240 ;
        RECT 81.245 186.195 81.535 186.240 ;
        RECT 83.105 186.195 83.395 186.240 ;
        RECT 59.650 185.855 59.940 186.085 ;
        RECT 61.015 185.840 61.335 186.100 ;
        RECT 62.395 186.040 62.715 186.100 ;
        RECT 62.870 186.040 63.160 186.085 ;
        RECT 62.395 185.900 63.160 186.040 ;
        RECT 62.395 185.840 62.715 185.900 ;
        RECT 62.870 185.855 63.160 185.900 ;
        RECT 70.325 186.040 70.615 186.085 ;
        RECT 71.135 186.040 71.455 186.100 ;
        RECT 70.325 185.900 71.455 186.040 ;
        RECT 70.325 185.855 70.615 185.900 ;
        RECT 71.135 185.840 71.455 185.900 ;
        RECT 74.600 186.040 74.890 186.085 ;
        RECT 75.275 186.040 75.595 186.100 ;
        RECT 74.600 185.900 75.595 186.040 ;
        RECT 74.600 185.855 74.890 185.900 ;
        RECT 75.275 185.840 75.595 185.900 ;
        RECT 75.735 186.040 76.055 186.100 ;
        RECT 84.105 186.040 84.245 186.580 ;
        RECT 84.490 186.535 84.780 186.580 ;
        RECT 93.675 186.520 93.995 186.580 ;
        RECT 95.530 186.535 95.820 186.580 ;
        RECT 100.130 186.535 100.420 186.580 ;
        RECT 101.050 186.720 101.340 186.765 ;
        RECT 101.955 186.720 102.275 186.780 ;
        RECT 101.050 186.580 102.275 186.720 ;
        RECT 101.050 186.535 101.340 186.580 ;
        RECT 101.955 186.520 102.275 186.580 ;
        RECT 103.425 186.425 103.565 186.920 ;
        RECT 106.110 186.875 106.400 186.920 ;
        RECT 103.350 186.195 103.640 186.425 ;
        RECT 75.735 185.900 84.245 186.040 ;
        RECT 90.010 186.040 90.300 186.085 ;
        RECT 90.455 186.040 90.775 186.100 ;
        RECT 90.010 185.900 90.775 186.040 ;
        RECT 75.735 185.840 76.055 185.900 ;
        RECT 90.010 185.855 90.300 185.900 ;
        RECT 90.455 185.840 90.775 185.900 ;
        RECT 94.135 185.840 94.455 186.100 ;
        RECT 18.165 185.220 112.465 185.700 ;
        RECT 25.595 185.020 25.915 185.080 ;
        RECT 28.815 185.020 29.135 185.080 ;
        RECT 31.115 185.020 31.435 185.080 ;
        RECT 36.175 185.020 36.495 185.080 ;
        RECT 36.650 185.020 36.940 185.065 ;
        RECT 25.595 184.880 28.585 185.020 ;
        RECT 25.595 184.820 25.915 184.880 ;
        RECT 21.880 184.680 22.170 184.725 ;
        RECT 23.770 184.680 24.060 184.725 ;
        RECT 26.890 184.680 27.180 184.725 ;
        RECT 21.880 184.540 27.180 184.680 ;
        RECT 28.445 184.680 28.585 184.880 ;
        RECT 28.815 184.880 31.435 185.020 ;
        RECT 28.815 184.820 29.135 184.880 ;
        RECT 31.115 184.820 31.435 184.880 ;
        RECT 33.965 184.880 35.945 185.020 ;
        RECT 33.965 184.680 34.105 184.880 ;
        RECT 28.445 184.540 34.105 184.680 ;
        RECT 21.880 184.495 22.170 184.540 ;
        RECT 23.770 184.495 24.060 184.540 ;
        RECT 26.890 184.495 27.180 184.540 ;
        RECT 24.215 184.340 24.535 184.400 ;
        RECT 24.215 184.200 29.045 184.340 ;
        RECT 24.215 184.140 24.535 184.200 ;
        RECT 20.535 183.800 20.855 184.060 ;
        RECT 21.010 183.815 21.300 184.045 ;
        RECT 21.475 184.000 21.765 184.045 ;
        RECT 23.310 184.000 23.600 184.045 ;
        RECT 26.890 184.000 27.180 184.045 ;
        RECT 21.475 183.860 27.180 184.000 ;
        RECT 21.475 183.815 21.765 183.860 ;
        RECT 23.310 183.815 23.600 183.860 ;
        RECT 26.890 183.815 27.180 183.860 ;
        RECT 20.075 183.120 20.395 183.380 ;
        RECT 21.085 183.320 21.225 183.815 ;
        RECT 22.375 183.460 22.695 183.720 ;
        RECT 24.675 183.705 24.995 183.720 ;
        RECT 27.970 183.705 28.260 184.020 ;
        RECT 28.905 184.000 29.045 184.200 ;
        RECT 29.735 184.140 30.055 184.400 ;
        RECT 31.205 184.385 31.345 184.540 ;
        RECT 34.350 184.495 34.640 184.725 ;
        RECT 31.130 184.155 31.420 184.385 ;
        RECT 32.050 184.000 32.340 184.045 ;
        RECT 33.875 184.000 34.195 184.060 ;
        RECT 28.905 183.860 34.195 184.000 ;
        RECT 34.425 184.000 34.565 184.495 ;
        RECT 35.805 184.340 35.945 184.880 ;
        RECT 36.175 184.880 36.940 185.020 ;
        RECT 36.175 184.820 36.495 184.880 ;
        RECT 36.650 184.835 36.940 184.880 ;
        RECT 38.030 185.020 38.320 185.065 ;
        RECT 38.475 185.020 38.795 185.080 ;
        RECT 38.030 184.880 38.795 185.020 ;
        RECT 38.030 184.835 38.320 184.880 ;
        RECT 38.475 184.820 38.795 184.880 ;
        RECT 42.630 185.020 42.920 185.065 ;
        RECT 44.915 185.020 45.235 185.080 ;
        RECT 42.630 184.880 45.235 185.020 ;
        RECT 42.630 184.835 42.920 184.880 ;
        RECT 44.915 184.820 45.235 184.880 ;
        RECT 46.770 185.020 47.060 185.065 ;
        RECT 47.215 185.020 47.535 185.080 ;
        RECT 46.770 184.880 47.535 185.020 ;
        RECT 46.770 184.835 47.060 184.880 ;
        RECT 47.215 184.820 47.535 184.880 ;
        RECT 55.955 185.020 56.275 185.080 ;
        RECT 63.315 185.020 63.635 185.080 ;
        RECT 65.615 185.020 65.935 185.080 ;
        RECT 55.955 184.880 59.405 185.020 ;
        RECT 55.955 184.820 56.275 184.880 ;
        RECT 52.390 184.680 52.680 184.725 ;
        RECT 55.510 184.680 55.800 184.725 ;
        RECT 57.400 184.680 57.690 184.725 ;
        RECT 39.485 184.540 44.225 184.680 ;
        RECT 38.935 184.340 39.255 184.400 ;
        RECT 39.485 184.385 39.625 184.540 ;
        RECT 39.410 184.340 39.700 184.385 ;
        RECT 43.535 184.340 43.855 184.400 ;
        RECT 44.085 184.385 44.225 184.540 ;
        RECT 52.390 184.540 57.690 184.680 ;
        RECT 52.390 184.495 52.680 184.540 ;
        RECT 55.510 184.495 55.800 184.540 ;
        RECT 57.400 184.495 57.690 184.540 ;
        RECT 58.730 184.495 59.020 184.725 ;
        RECT 59.265 184.680 59.405 184.880 ;
        RECT 63.315 184.880 65.935 185.020 ;
        RECT 63.315 184.820 63.635 184.880 ;
        RECT 65.615 184.820 65.935 184.880 ;
        RECT 71.135 184.820 71.455 185.080 ;
        RECT 71.595 185.020 71.915 185.080 ;
        RECT 72.530 185.020 72.820 185.065 ;
        RECT 71.595 184.880 72.820 185.020 ;
        RECT 71.595 184.820 71.915 184.880 ;
        RECT 72.530 184.835 72.820 184.880 ;
        RECT 74.815 184.820 75.135 185.080 ;
        RECT 81.255 184.820 81.575 185.080 ;
        RECT 81.715 184.820 82.035 185.080 ;
        RECT 93.675 185.020 93.995 185.080 ;
        RECT 93.675 184.880 95.285 185.020 ;
        RECT 93.675 184.820 93.995 184.880 ;
        RECT 64.710 184.680 65.000 184.725 ;
        RECT 89.650 184.680 89.940 184.725 ;
        RECT 92.770 184.680 93.060 184.725 ;
        RECT 94.660 184.680 94.950 184.725 ;
        RECT 59.265 184.540 65.000 184.680 ;
        RECT 64.710 184.495 65.000 184.540 ;
        RECT 67.545 184.540 72.745 184.680 ;
        RECT 35.805 184.200 39.700 184.340 ;
        RECT 38.935 184.140 39.255 184.200 ;
        RECT 39.410 184.155 39.700 184.200 ;
        RECT 40.405 184.200 43.855 184.340 ;
        RECT 35.730 184.000 36.020 184.045 ;
        RECT 34.425 183.860 36.020 184.000 ;
        RECT 32.050 183.815 32.340 183.860 ;
        RECT 33.875 183.800 34.195 183.860 ;
        RECT 35.730 183.815 36.020 183.860 ;
        RECT 37.570 184.000 37.860 184.045 ;
        RECT 40.405 184.000 40.545 184.200 ;
        RECT 43.535 184.140 43.855 184.200 ;
        RECT 44.010 184.155 44.300 184.385 ;
        RECT 56.890 184.340 57.180 184.385 ;
        RECT 58.805 184.340 58.945 184.495 ;
        RECT 56.890 184.200 58.945 184.340 ;
        RECT 61.015 184.340 61.335 184.400 ;
        RECT 62.410 184.340 62.700 184.385 ;
        RECT 61.015 184.200 62.700 184.340 ;
        RECT 56.890 184.155 57.180 184.200 ;
        RECT 61.015 184.140 61.335 184.200 ;
        RECT 62.410 184.155 62.700 184.200 ;
        RECT 64.235 184.340 64.555 184.400 ;
        RECT 67.545 184.340 67.685 184.540 ;
        RECT 64.235 184.200 67.685 184.340 ;
        RECT 64.235 184.140 64.555 184.200 ;
        RECT 37.570 183.860 40.545 184.000 ;
        RECT 40.775 184.000 41.095 184.060 ;
        RECT 42.615 184.000 42.935 184.060 ;
        RECT 44.470 184.000 44.760 184.045 ;
        RECT 40.775 183.860 44.760 184.000 ;
        RECT 37.570 183.815 37.860 183.860 ;
        RECT 40.775 183.800 41.095 183.860 ;
        RECT 42.615 183.800 42.935 183.860 ;
        RECT 44.470 183.815 44.760 183.860 ;
        RECT 48.150 184.000 48.440 184.045 ;
        RECT 50.435 184.000 50.755 184.060 ;
        RECT 48.150 183.860 50.755 184.000 ;
        RECT 48.150 183.815 48.440 183.860 ;
        RECT 50.435 183.800 50.755 183.860 ;
        RECT 24.670 183.660 25.320 183.705 ;
        RECT 27.970 183.660 28.560 183.705 ;
        RECT 24.670 183.520 28.560 183.660 ;
        RECT 24.670 183.475 25.320 183.520 ;
        RECT 28.270 183.475 28.560 183.520 ;
        RECT 32.510 183.660 32.800 183.705 ;
        RECT 49.055 183.660 49.375 183.720 ;
        RECT 51.310 183.705 51.600 184.020 ;
        RECT 52.390 184.000 52.680 184.045 ;
        RECT 55.970 184.000 56.260 184.045 ;
        RECT 57.805 184.000 58.095 184.045 ;
        RECT 52.390 183.860 58.095 184.000 ;
        RECT 52.390 183.815 52.680 183.860 ;
        RECT 55.970 183.815 56.260 183.860 ;
        RECT 57.805 183.815 58.095 183.860 ;
        RECT 58.270 183.815 58.560 184.045 ;
        RECT 59.650 184.000 59.940 184.045 ;
        RECT 58.805 183.860 59.940 184.000 ;
        RECT 51.010 183.660 51.600 183.705 ;
        RECT 54.250 183.660 54.900 183.705 ;
        RECT 58.345 183.660 58.485 183.815 ;
        RECT 32.510 183.520 40.545 183.660 ;
        RECT 32.510 183.475 32.800 183.520 ;
        RECT 24.675 183.460 24.995 183.475 ;
        RECT 40.405 183.380 40.545 183.520 ;
        RECT 49.055 183.520 54.900 183.660 ;
        RECT 49.055 183.460 49.375 183.520 ;
        RECT 51.010 183.475 51.300 183.520 ;
        RECT 54.250 183.475 54.900 183.520 ;
        RECT 55.125 183.520 58.485 183.660 ;
        RECT 55.125 183.380 55.265 183.520 ;
        RECT 32.955 183.320 33.275 183.380 ;
        RECT 21.085 183.180 33.275 183.320 ;
        RECT 32.955 183.120 33.275 183.180 ;
        RECT 40.315 183.120 40.635 183.380 ;
        RECT 44.930 183.320 45.220 183.365 ;
        RECT 48.135 183.320 48.455 183.380 ;
        RECT 44.930 183.180 48.455 183.320 ;
        RECT 44.930 183.135 45.220 183.180 ;
        RECT 48.135 183.120 48.455 183.180 ;
        RECT 55.035 183.120 55.355 183.380 ;
        RECT 57.335 183.320 57.655 183.380 ;
        RECT 58.805 183.320 58.945 183.860 ;
        RECT 59.650 183.815 59.940 183.860 ;
        RECT 62.855 184.000 63.175 184.060 ;
        RECT 63.790 184.000 64.080 184.045 ;
        RECT 66.090 184.000 66.380 184.045 ;
        RECT 62.855 183.860 66.380 184.000 ;
        RECT 62.855 183.800 63.175 183.860 ;
        RECT 63.790 183.815 64.080 183.860 ;
        RECT 66.090 183.815 66.380 183.860 ;
        RECT 66.535 183.800 66.855 184.060 ;
        RECT 67.545 184.045 67.685 184.200 ;
        RECT 69.295 184.340 69.615 184.400 ;
        RECT 71.595 184.340 71.915 184.400 ;
        RECT 69.295 184.200 71.915 184.340 ;
        RECT 69.295 184.140 69.615 184.200 ;
        RECT 71.595 184.140 71.915 184.200 ;
        RECT 67.470 183.815 67.760 184.045 ;
        RECT 68.375 183.800 68.695 184.060 ;
        RECT 69.770 183.980 70.060 184.045 ;
        RECT 69.385 183.840 70.060 183.980 ;
        RECT 59.175 183.660 59.495 183.720 ;
        RECT 65.615 183.660 65.935 183.720 ;
        RECT 69.385 183.660 69.525 183.840 ;
        RECT 69.770 183.815 70.060 183.840 ;
        RECT 72.070 184.000 72.360 184.045 ;
        RECT 72.605 184.000 72.745 184.540 ;
        RECT 89.650 184.540 94.950 184.680 ;
        RECT 89.650 184.495 89.940 184.540 ;
        RECT 92.770 184.495 93.060 184.540 ;
        RECT 94.660 184.495 94.950 184.540 ;
        RECT 75.735 184.340 76.055 184.400 ;
        RECT 76.210 184.340 76.500 184.385 ;
        RECT 75.735 184.200 76.500 184.340 ;
        RECT 75.735 184.140 76.055 184.200 ;
        RECT 76.210 184.155 76.500 184.200 ;
        RECT 94.135 184.140 94.455 184.400 ;
        RECT 95.145 184.340 95.285 184.880 ;
        RECT 96.525 184.540 100.805 184.680 ;
        RECT 96.525 184.385 96.665 184.540 ;
        RECT 100.665 184.385 100.805 184.540 ;
        RECT 103.810 184.495 104.100 184.725 ;
        RECT 96.450 184.340 96.740 184.385 ;
        RECT 95.145 184.200 96.740 184.340 ;
        RECT 96.450 184.155 96.740 184.200 ;
        RECT 100.590 184.155 100.880 184.385 ;
        RECT 103.885 184.340 104.025 184.495 ;
        RECT 103.885 184.200 106.325 184.340 ;
        RECT 72.070 183.860 72.745 184.000 ;
        RECT 72.070 183.815 72.360 183.860 ;
        RECT 72.990 183.815 73.280 184.045 ;
        RECT 73.065 183.660 73.205 183.815 ;
        RECT 74.355 183.800 74.675 184.060 ;
        RECT 80.350 184.000 80.640 184.045 ;
        RECT 79.505 183.860 80.640 184.000 ;
        RECT 59.175 183.520 65.385 183.660 ;
        RECT 59.175 183.460 59.495 183.520 ;
        RECT 57.335 183.180 58.945 183.320 ;
        RECT 57.335 183.120 57.655 183.180 ;
        RECT 61.015 183.120 61.335 183.380 ;
        RECT 65.245 183.365 65.385 183.520 ;
        RECT 65.615 183.520 69.525 183.660 ;
        RECT 71.225 183.520 73.205 183.660 ;
        RECT 65.615 183.460 65.935 183.520 ;
        RECT 65.170 183.320 65.460 183.365 ;
        RECT 68.375 183.320 68.695 183.380 ;
        RECT 71.225 183.320 71.365 183.520 ;
        RECT 65.170 183.180 71.365 183.320 ;
        RECT 71.595 183.320 71.915 183.380 ;
        RECT 75.275 183.320 75.595 183.380 ;
        RECT 77.130 183.320 77.420 183.365 ;
        RECT 71.595 183.180 77.420 183.320 ;
        RECT 65.170 183.135 65.460 183.180 ;
        RECT 68.375 183.120 68.695 183.180 ;
        RECT 71.595 183.120 71.915 183.180 ;
        RECT 75.275 183.120 75.595 183.180 ;
        RECT 77.130 183.135 77.420 183.180 ;
        RECT 77.575 183.120 77.895 183.380 ;
        RECT 79.505 183.365 79.645 183.860 ;
        RECT 80.350 183.815 80.640 183.860 ;
        RECT 82.635 183.800 82.955 184.060 ;
        RECT 88.570 183.705 88.860 184.020 ;
        RECT 89.650 184.000 89.940 184.045 ;
        RECT 93.230 184.000 93.520 184.045 ;
        RECT 95.065 184.000 95.355 184.045 ;
        RECT 89.650 183.860 95.355 184.000 ;
        RECT 89.650 183.815 89.940 183.860 ;
        RECT 93.230 183.815 93.520 183.860 ;
        RECT 95.065 183.815 95.355 183.860 ;
        RECT 95.530 184.000 95.820 184.045 ;
        RECT 96.895 184.000 97.215 184.060 ;
        RECT 95.530 183.860 97.215 184.000 ;
        RECT 95.530 183.815 95.820 183.860 ;
        RECT 96.895 183.800 97.215 183.860 ;
        RECT 98.275 184.000 98.595 184.060 ;
        RECT 101.955 184.000 102.275 184.060 ;
        RECT 98.275 183.860 102.275 184.000 ;
        RECT 98.275 183.800 98.595 183.860 ;
        RECT 101.955 183.800 102.275 183.860 ;
        RECT 105.175 183.800 105.495 184.060 ;
        RECT 106.185 184.045 106.325 184.200 ;
        RECT 106.110 183.815 106.400 184.045 ;
        RECT 88.270 183.660 88.860 183.705 ;
        RECT 90.455 183.660 90.775 183.720 ;
        RECT 91.510 183.660 92.160 183.705 ;
        RECT 88.270 183.520 92.160 183.660 ;
        RECT 88.270 183.475 88.560 183.520 ;
        RECT 90.455 183.460 90.775 183.520 ;
        RECT 91.510 183.475 92.160 183.520 ;
        RECT 97.830 183.660 98.120 183.705 ;
        RECT 97.830 183.520 101.265 183.660 ;
        RECT 97.830 183.475 98.120 183.520 ;
        RECT 101.125 183.380 101.265 183.520 ;
        RECT 79.430 183.135 79.720 183.365 ;
        RECT 85.855 183.320 86.175 183.380 ;
        RECT 86.790 183.320 87.080 183.365 ;
        RECT 85.855 183.180 87.080 183.320 ;
        RECT 85.855 183.120 86.175 183.180 ;
        RECT 86.790 183.135 87.080 183.180 ;
        RECT 92.295 183.320 92.615 183.380 ;
        RECT 97.370 183.320 97.660 183.365 ;
        RECT 92.295 183.180 97.660 183.320 ;
        RECT 92.295 183.120 92.615 183.180 ;
        RECT 97.370 183.135 97.660 183.180 ;
        RECT 99.670 183.320 99.960 183.365 ;
        RECT 100.575 183.320 100.895 183.380 ;
        RECT 99.670 183.180 100.895 183.320 ;
        RECT 99.670 183.135 99.960 183.180 ;
        RECT 100.575 183.120 100.895 183.180 ;
        RECT 101.035 183.320 101.355 183.380 ;
        RECT 101.510 183.320 101.800 183.365 ;
        RECT 101.035 183.180 101.800 183.320 ;
        RECT 101.035 183.120 101.355 183.180 ;
        RECT 101.510 183.135 101.800 183.180 ;
        RECT 104.715 183.120 105.035 183.380 ;
        RECT 107.030 183.320 107.320 183.365 ;
        RECT 108.395 183.320 108.715 183.380 ;
        RECT 107.030 183.180 108.715 183.320 ;
        RECT 107.030 183.135 107.320 183.180 ;
        RECT 108.395 183.120 108.715 183.180 ;
        RECT 17.370 182.500 112.465 182.980 ;
        RECT 21.470 182.300 21.760 182.345 ;
        RECT 22.375 182.300 22.695 182.360 ;
        RECT 21.470 182.160 22.695 182.300 ;
        RECT 21.470 182.115 21.760 182.160 ;
        RECT 22.375 182.100 22.695 182.160 ;
        RECT 26.990 182.115 27.280 182.345 ;
        RECT 33.415 182.300 33.735 182.360 ;
        RECT 33.415 182.160 39.165 182.300 ;
        RECT 27.065 181.960 27.205 182.115 ;
        RECT 33.415 182.100 33.735 182.160 ;
        RECT 39.025 182.020 39.165 182.160 ;
        RECT 57.335 182.100 57.655 182.360 ;
        RECT 57.810 182.115 58.100 182.345 ;
        RECT 61.935 182.300 62.255 182.360 ;
        RECT 66.090 182.300 66.380 182.345 ;
        RECT 61.935 182.160 66.380 182.300 ;
        RECT 35.715 182.005 36.035 182.020 ;
        RECT 20.625 181.820 27.205 181.960 ;
        RECT 32.610 181.960 32.900 182.005 ;
        RECT 35.715 181.960 36.500 182.005 ;
        RECT 32.610 181.820 36.500 181.960 ;
        RECT 20.625 181.665 20.765 181.820 ;
        RECT 32.610 181.775 33.200 181.820 ;
        RECT 20.550 181.435 20.840 181.665 ;
        RECT 27.435 181.620 27.755 181.680 ;
        RECT 28.830 181.620 29.120 181.665 ;
        RECT 31.115 181.620 31.435 181.680 ;
        RECT 27.435 181.480 31.435 181.620 ;
        RECT 27.435 181.420 27.755 181.480 ;
        RECT 28.830 181.435 29.120 181.480 ;
        RECT 31.115 181.420 31.435 181.480 ;
        RECT 32.910 181.460 33.200 181.775 ;
        RECT 35.715 181.775 36.500 181.820 ;
        RECT 38.935 181.960 39.255 182.020 ;
        RECT 38.935 181.820 40.085 181.960 ;
        RECT 35.715 181.760 36.035 181.775 ;
        RECT 38.935 181.760 39.255 181.820 ;
        RECT 39.945 181.665 40.085 181.820 ;
        RECT 55.510 181.775 55.800 182.005 ;
        RECT 56.590 181.960 56.880 182.005 ;
        RECT 57.885 181.960 58.025 182.115 ;
        RECT 61.935 182.100 62.255 182.160 ;
        RECT 66.090 182.115 66.380 182.160 ;
        RECT 99.670 182.115 99.960 182.345 ;
        RECT 61.015 181.960 61.335 182.020 ;
        RECT 66.850 181.960 67.140 182.005 ;
        RECT 56.590 181.820 58.025 181.960 ;
        RECT 58.345 181.820 67.140 181.960 ;
        RECT 56.590 181.775 56.880 181.820 ;
        RECT 33.990 181.620 34.280 181.665 ;
        RECT 37.570 181.620 37.860 181.665 ;
        RECT 39.405 181.620 39.695 181.665 ;
        RECT 33.990 181.480 39.695 181.620 ;
        RECT 33.990 181.435 34.280 181.480 ;
        RECT 37.570 181.435 37.860 181.480 ;
        RECT 39.405 181.435 39.695 181.480 ;
        RECT 39.870 181.435 40.160 181.665 ;
        RECT 55.585 181.620 55.725 181.775 ;
        RECT 58.345 181.620 58.485 181.820 ;
        RECT 61.015 181.760 61.335 181.820 ;
        RECT 66.850 181.775 67.140 181.820 ;
        RECT 67.930 181.960 68.220 182.005 ;
        RECT 69.295 181.960 69.615 182.020 ;
        RECT 95.055 182.005 95.375 182.020 ;
        RECT 67.930 181.820 69.615 181.960 ;
        RECT 67.930 181.775 68.220 181.820 ;
        RECT 69.295 181.760 69.615 181.820 ;
        RECT 91.490 181.960 91.780 182.005 ;
        RECT 94.730 181.960 95.380 182.005 ;
        RECT 91.490 181.820 95.380 181.960 ;
        RECT 91.490 181.775 92.080 181.820 ;
        RECT 94.730 181.775 95.380 181.820 ;
        RECT 97.370 181.960 97.660 182.005 ;
        RECT 99.745 181.960 99.885 182.115 ;
        RECT 97.370 181.820 99.885 181.960 ;
        RECT 102.530 181.960 102.820 182.005 ;
        RECT 104.715 181.960 105.035 182.020 ;
        RECT 105.770 181.960 106.420 182.005 ;
        RECT 102.530 181.820 106.420 181.960 ;
        RECT 97.370 181.775 97.660 181.820 ;
        RECT 102.530 181.775 103.120 181.820 ;
        RECT 55.585 181.480 58.485 181.620 ;
        RECT 58.715 181.420 59.035 181.680 ;
        RECT 59.635 181.420 59.955 181.680 ;
        RECT 62.395 181.420 62.715 181.680 ;
        RECT 74.815 181.620 75.135 181.680 ;
        RECT 77.575 181.620 77.895 181.680 ;
        RECT 74.815 181.480 77.895 181.620 ;
        RECT 74.815 181.420 75.135 181.480 ;
        RECT 77.575 181.420 77.895 181.480 ;
        RECT 78.050 181.620 78.340 181.665 ;
        RECT 81.715 181.620 82.035 181.680 ;
        RECT 78.050 181.480 82.035 181.620 ;
        RECT 78.050 181.435 78.340 181.480 ;
        RECT 81.715 181.420 82.035 181.480 ;
        RECT 91.790 181.460 92.080 181.775 ;
        RECT 95.055 181.760 95.375 181.775 ;
        RECT 92.870 181.620 93.160 181.665 ;
        RECT 96.450 181.620 96.740 181.665 ;
        RECT 98.285 181.620 98.575 181.665 ;
        RECT 92.870 181.480 98.575 181.620 ;
        RECT 92.870 181.435 93.160 181.480 ;
        RECT 96.450 181.435 96.740 181.480 ;
        RECT 98.285 181.435 98.575 181.480 ;
        RECT 100.575 181.420 100.895 181.680 ;
        RECT 102.830 181.460 103.120 181.775 ;
        RECT 104.715 181.760 105.035 181.820 ;
        RECT 105.770 181.775 106.420 181.820 ;
        RECT 108.395 181.760 108.715 182.020 ;
        RECT 108.855 181.960 109.175 182.020 ;
        RECT 108.855 181.820 110.005 181.960 ;
        RECT 108.855 181.760 109.175 181.820 ;
        RECT 109.865 181.665 110.005 181.820 ;
        RECT 103.910 181.620 104.200 181.665 ;
        RECT 107.490 181.620 107.780 181.665 ;
        RECT 109.325 181.620 109.615 181.665 ;
        RECT 103.910 181.480 109.615 181.620 ;
        RECT 103.910 181.435 104.200 181.480 ;
        RECT 107.490 181.435 107.780 181.480 ;
        RECT 109.325 181.435 109.615 181.480 ;
        RECT 109.790 181.435 110.080 181.665 ;
        RECT 22.850 181.280 23.140 181.325 ;
        RECT 29.290 181.280 29.580 181.325 ;
        RECT 22.850 181.140 29.580 181.280 ;
        RECT 22.850 181.095 23.140 181.140 ;
        RECT 29.290 181.095 29.580 181.140 ;
        RECT 30.210 181.280 30.500 181.325 ;
        RECT 32.495 181.280 32.815 181.340 ;
        RECT 34.795 181.280 35.115 181.340 ;
        RECT 30.210 181.140 32.815 181.280 ;
        RECT 30.210 181.095 30.500 181.140 ;
        RECT 29.365 180.940 29.505 181.095 ;
        RECT 32.495 181.080 32.815 181.140 ;
        RECT 33.045 181.140 35.115 181.280 ;
        RECT 29.735 180.940 30.055 181.000 ;
        RECT 33.045 180.940 33.185 181.140 ;
        RECT 34.795 181.080 35.115 181.140 ;
        RECT 38.015 181.280 38.335 181.340 ;
        RECT 38.490 181.280 38.780 181.325 ;
        RECT 38.015 181.140 38.780 181.280 ;
        RECT 38.015 181.080 38.335 181.140 ;
        RECT 38.490 181.095 38.780 181.140 ;
        RECT 57.795 181.280 58.115 181.340 ;
        RECT 59.175 181.280 59.495 181.340 ;
        RECT 57.795 181.140 59.495 181.280 ;
        RECT 57.795 181.080 58.115 181.140 ;
        RECT 59.175 181.080 59.495 181.140 ;
        RECT 60.110 181.280 60.400 181.325 ;
        RECT 62.855 181.280 63.175 181.340 ;
        RECT 60.110 181.140 63.175 181.280 ;
        RECT 60.110 181.095 60.400 181.140 ;
        RECT 29.365 180.800 33.185 180.940 ;
        RECT 33.990 180.940 34.280 180.985 ;
        RECT 37.110 180.940 37.400 180.985 ;
        RECT 39.000 180.940 39.290 180.985 ;
        RECT 33.990 180.800 39.290 180.940 ;
        RECT 29.735 180.740 30.055 180.800 ;
        RECT 33.990 180.755 34.280 180.800 ;
        RECT 37.110 180.755 37.400 180.800 ;
        RECT 39.000 180.755 39.290 180.800 ;
        RECT 56.875 180.940 57.195 181.000 ;
        RECT 60.185 180.940 60.325 181.095 ;
        RECT 62.855 181.080 63.175 181.140 ;
        RECT 73.895 181.280 74.215 181.340 ;
        RECT 75.735 181.280 76.055 181.340 ;
        RECT 76.670 181.280 76.960 181.325 ;
        RECT 73.895 181.140 76.960 181.280 ;
        RECT 73.895 181.080 74.215 181.140 ;
        RECT 75.735 181.080 76.055 181.140 ;
        RECT 76.670 181.095 76.960 181.140 ;
        RECT 96.895 181.280 97.215 181.340 ;
        RECT 98.750 181.280 99.040 181.325 ;
        RECT 96.895 181.140 99.040 181.280 ;
        RECT 96.895 181.080 97.215 181.140 ;
        RECT 98.750 181.095 99.040 181.140 ;
        RECT 56.875 180.800 60.325 180.940 ;
        RECT 92.870 180.940 93.160 180.985 ;
        RECT 95.990 180.940 96.280 180.985 ;
        RECT 97.880 180.940 98.170 180.985 ;
        RECT 92.870 180.800 98.170 180.940 ;
        RECT 56.875 180.740 57.195 180.800 ;
        RECT 92.870 180.755 93.160 180.800 ;
        RECT 95.990 180.755 96.280 180.800 ;
        RECT 97.880 180.755 98.170 180.800 ;
        RECT 103.910 180.940 104.200 180.985 ;
        RECT 107.030 180.940 107.320 180.985 ;
        RECT 108.920 180.940 109.210 180.985 ;
        RECT 103.910 180.800 109.210 180.940 ;
        RECT 103.910 180.755 104.200 180.800 ;
        RECT 107.030 180.755 107.320 180.800 ;
        RECT 108.920 180.755 109.210 180.800 ;
        RECT 25.610 180.600 25.900 180.645 ;
        RECT 26.055 180.600 26.375 180.660 ;
        RECT 25.610 180.460 26.375 180.600 ;
        RECT 25.610 180.415 25.900 180.460 ;
        RECT 26.055 180.400 26.375 180.460 ;
        RECT 31.130 180.600 31.420 180.645 ;
        RECT 33.415 180.600 33.735 180.660 ;
        RECT 31.130 180.460 33.735 180.600 ;
        RECT 31.130 180.415 31.420 180.460 ;
        RECT 33.415 180.400 33.735 180.460 ;
        RECT 55.955 180.600 56.275 180.660 ;
        RECT 56.430 180.600 56.720 180.645 ;
        RECT 55.955 180.460 56.720 180.600 ;
        RECT 55.955 180.400 56.275 180.460 ;
        RECT 56.430 180.415 56.720 180.460 ;
        RECT 58.715 180.600 59.035 180.660 ;
        RECT 61.015 180.600 61.335 180.660 ;
        RECT 61.490 180.600 61.780 180.645 ;
        RECT 63.315 180.600 63.635 180.660 ;
        RECT 58.715 180.460 63.635 180.600 ;
        RECT 58.715 180.400 59.035 180.460 ;
        RECT 61.015 180.400 61.335 180.460 ;
        RECT 61.490 180.415 61.780 180.460 ;
        RECT 63.315 180.400 63.635 180.460 ;
        RECT 66.535 180.600 66.855 180.660 ;
        RECT 67.010 180.600 67.300 180.645 ;
        RECT 66.535 180.460 67.300 180.600 ;
        RECT 66.535 180.400 66.855 180.460 ;
        RECT 67.010 180.415 67.300 180.460 ;
        RECT 79.875 180.400 80.195 180.660 ;
        RECT 90.010 180.600 90.300 180.645 ;
        RECT 92.295 180.600 92.615 180.660 ;
        RECT 90.010 180.460 92.615 180.600 ;
        RECT 90.010 180.415 90.300 180.460 ;
        RECT 92.295 180.400 92.615 180.460 ;
        RECT 99.195 180.600 99.515 180.660 ;
        RECT 101.035 180.600 101.355 180.660 ;
        RECT 99.195 180.460 101.355 180.600 ;
        RECT 99.195 180.400 99.515 180.460 ;
        RECT 101.035 180.400 101.355 180.460 ;
        RECT 18.165 179.780 112.465 180.260 ;
        RECT 35.715 179.380 36.035 179.640 ;
        RECT 38.015 179.380 38.335 179.640 ;
        RECT 60.095 179.580 60.415 179.640 ;
        RECT 61.935 179.580 62.255 179.640 ;
        RECT 60.095 179.440 62.255 179.580 ;
        RECT 60.095 179.380 60.415 179.440 ;
        RECT 61.935 179.380 62.255 179.440 ;
        RECT 93.215 179.580 93.535 179.640 ;
        RECT 94.150 179.580 94.440 179.625 ;
        RECT 93.215 179.440 94.440 179.580 ;
        RECT 93.215 179.380 93.535 179.440 ;
        RECT 94.150 179.395 94.440 179.440 ;
        RECT 95.055 179.580 95.375 179.640 ;
        RECT 95.530 179.580 95.820 179.625 ;
        RECT 95.055 179.440 95.820 179.580 ;
        RECT 95.055 179.380 95.375 179.440 ;
        RECT 95.530 179.395 95.820 179.440 ;
        RECT 22.950 179.240 23.240 179.285 ;
        RECT 26.070 179.240 26.360 179.285 ;
        RECT 27.960 179.240 28.250 179.285 ;
        RECT 22.950 179.100 28.250 179.240 ;
        RECT 22.950 179.055 23.240 179.100 ;
        RECT 26.070 179.055 26.360 179.100 ;
        RECT 27.960 179.055 28.250 179.100 ;
        RECT 29.290 179.055 29.580 179.285 ;
        RECT 34.350 179.055 34.640 179.285 ;
        RECT 49.025 179.240 49.315 179.285 ;
        RECT 51.805 179.240 52.095 179.285 ;
        RECT 53.665 179.240 53.955 179.285 ;
        RECT 49.025 179.100 53.955 179.240 ;
        RECT 49.025 179.055 49.315 179.100 ;
        RECT 51.805 179.055 52.095 179.100 ;
        RECT 53.665 179.055 53.955 179.100 ;
        RECT 76.770 179.240 77.060 179.285 ;
        RECT 79.890 179.240 80.180 179.285 ;
        RECT 81.780 179.240 82.070 179.285 ;
        RECT 93.675 179.240 93.995 179.300 ;
        RECT 76.770 179.100 82.070 179.240 ;
        RECT 76.770 179.055 77.060 179.100 ;
        RECT 79.890 179.055 80.180 179.100 ;
        RECT 81.780 179.055 82.070 179.100 ;
        RECT 91.465 179.100 93.995 179.240 ;
        RECT 20.090 178.900 20.380 178.945 ;
        RECT 24.675 178.900 24.995 178.960 ;
        RECT 20.090 178.760 24.995 178.900 ;
        RECT 20.090 178.715 20.380 178.760 ;
        RECT 24.675 178.700 24.995 178.760 ;
        RECT 27.450 178.900 27.740 178.945 ;
        RECT 29.365 178.900 29.505 179.055 ;
        RECT 27.450 178.760 29.505 178.900 ;
        RECT 31.590 178.900 31.880 178.945 ;
        RECT 32.495 178.900 32.815 178.960 ;
        RECT 34.425 178.900 34.565 179.055 ;
        RECT 50.435 178.900 50.755 178.960 ;
        RECT 56.875 178.900 57.195 178.960 ;
        RECT 31.590 178.760 34.105 178.900 ;
        RECT 34.425 178.760 37.325 178.900 ;
        RECT 27.450 178.715 27.740 178.760 ;
        RECT 31.590 178.715 31.880 178.760 ;
        RECT 32.495 178.700 32.815 178.760 ;
        RECT 20.075 178.220 20.395 178.280 ;
        RECT 21.870 178.265 22.160 178.580 ;
        RECT 22.950 178.560 23.240 178.605 ;
        RECT 26.530 178.560 26.820 178.605 ;
        RECT 28.365 178.560 28.655 178.605 ;
        RECT 22.950 178.420 28.655 178.560 ;
        RECT 22.950 178.375 23.240 178.420 ;
        RECT 26.530 178.375 26.820 178.420 ;
        RECT 28.365 178.375 28.655 178.420 ;
        RECT 28.815 178.360 29.135 178.620 ;
        RECT 30.210 178.375 30.500 178.605 ;
        RECT 21.570 178.220 22.160 178.265 ;
        RECT 24.810 178.220 25.460 178.265 ;
        RECT 20.075 178.080 25.460 178.220 ;
        RECT 20.075 178.020 20.395 178.080 ;
        RECT 21.570 178.035 21.860 178.080 ;
        RECT 24.810 178.035 25.460 178.080 ;
        RECT 27.895 178.220 28.215 178.280 ;
        RECT 30.285 178.220 30.425 178.375 ;
        RECT 27.895 178.080 30.425 178.220 ;
        RECT 32.050 178.220 32.340 178.265 ;
        RECT 33.415 178.220 33.735 178.280 ;
        RECT 32.050 178.080 33.735 178.220 ;
        RECT 33.965 178.220 34.105 178.760 ;
        RECT 35.255 178.560 35.575 178.620 ;
        RECT 37.185 178.605 37.325 178.760 ;
        RECT 50.435 178.760 57.195 178.900 ;
        RECT 50.435 178.700 50.755 178.760 ;
        RECT 56.875 178.700 57.195 178.760 ;
        RECT 58.270 178.900 58.560 178.945 ;
        RECT 62.395 178.900 62.715 178.960 ;
        RECT 70.215 178.900 70.535 178.960 ;
        RECT 70.690 178.900 70.980 178.945 ;
        RECT 89.995 178.900 90.315 178.960 ;
        RECT 91.465 178.945 91.605 179.100 ;
        RECT 93.675 179.040 93.995 179.100 ;
        RECT 58.270 178.760 62.715 178.900 ;
        RECT 58.270 178.715 58.560 178.760 ;
        RECT 62.395 178.700 62.715 178.760 ;
        RECT 68.005 178.760 70.980 178.900 ;
        RECT 36.190 178.560 36.480 178.605 ;
        RECT 35.255 178.420 36.480 178.560 ;
        RECT 35.255 178.360 35.575 178.420 ;
        RECT 36.190 178.375 36.480 178.420 ;
        RECT 37.110 178.375 37.400 178.605 ;
        RECT 38.015 178.560 38.335 178.620 ;
        RECT 39.410 178.560 39.700 178.605 ;
        RECT 38.015 178.420 39.700 178.560 ;
        RECT 38.015 178.360 38.335 178.420 ;
        RECT 39.410 178.375 39.700 178.420 ;
        RECT 43.995 178.560 44.315 178.620 ;
        RECT 44.470 178.560 44.760 178.605 ;
        RECT 44.915 178.560 45.235 178.620 ;
        RECT 43.995 178.420 45.235 178.560 ;
        RECT 43.995 178.360 44.315 178.420 ;
        RECT 44.470 178.375 44.760 178.420 ;
        RECT 44.915 178.360 45.235 178.420 ;
        RECT 49.025 178.560 49.315 178.605 ;
        RECT 49.025 178.420 51.560 178.560 ;
        RECT 49.025 178.375 49.315 178.420 ;
        RECT 37.555 178.220 37.875 178.280 ;
        RECT 50.435 178.265 50.755 178.280 ;
        RECT 33.965 178.080 37.875 178.220 ;
        RECT 27.895 178.020 28.215 178.080 ;
        RECT 32.050 178.035 32.340 178.080 ;
        RECT 33.415 178.020 33.735 178.080 ;
        RECT 37.555 178.020 37.875 178.080 ;
        RECT 47.165 178.220 47.455 178.265 ;
        RECT 50.425 178.220 50.755 178.265 ;
        RECT 47.165 178.080 50.755 178.220 ;
        RECT 47.165 178.035 47.455 178.080 ;
        RECT 50.425 178.035 50.755 178.080 ;
        RECT 51.345 178.265 51.560 178.420 ;
        RECT 52.275 178.360 52.595 178.620 ;
        RECT 54.130 178.560 54.420 178.605 ;
        RECT 54.575 178.560 54.895 178.620 ;
        RECT 54.130 178.420 54.895 178.560 ;
        RECT 54.130 178.375 54.420 178.420 ;
        RECT 54.575 178.360 54.895 178.420 ;
        RECT 59.315 178.560 59.605 178.605 ;
        RECT 61.475 178.560 61.795 178.620 ;
        RECT 68.005 178.605 68.145 178.760 ;
        RECT 70.215 178.700 70.535 178.760 ;
        RECT 70.690 178.715 70.980 178.760 ;
        RECT 74.445 178.760 85.625 178.900 ;
        RECT 74.445 178.620 74.585 178.760 ;
        RECT 59.315 178.420 61.795 178.560 ;
        RECT 59.315 178.375 59.605 178.420 ;
        RECT 61.475 178.360 61.795 178.420 ;
        RECT 67.930 178.375 68.220 178.605 ;
        RECT 68.375 178.360 68.695 178.620 ;
        RECT 69.770 178.560 70.060 178.605 ;
        RECT 72.515 178.560 72.835 178.620 ;
        RECT 69.770 178.420 72.835 178.560 ;
        RECT 69.770 178.375 70.060 178.420 ;
        RECT 72.515 178.360 72.835 178.420 ;
        RECT 73.450 178.560 73.740 178.605 ;
        RECT 74.355 178.560 74.675 178.620 ;
        RECT 73.450 178.420 74.675 178.560 ;
        RECT 73.450 178.375 73.740 178.420 ;
        RECT 74.355 178.360 74.675 178.420 ;
        RECT 75.690 178.265 75.980 178.580 ;
        RECT 76.770 178.560 77.060 178.605 ;
        RECT 80.350 178.560 80.640 178.605 ;
        RECT 82.185 178.560 82.475 178.605 ;
        RECT 76.770 178.420 82.475 178.560 ;
        RECT 76.770 178.375 77.060 178.420 ;
        RECT 80.350 178.375 80.640 178.420 ;
        RECT 82.185 178.375 82.475 178.420 ;
        RECT 82.635 178.360 82.955 178.620 ;
        RECT 85.485 178.605 85.625 178.760 ;
        RECT 86.865 178.760 90.315 178.900 ;
        RECT 86.865 178.605 87.005 178.760 ;
        RECT 89.995 178.700 90.315 178.760 ;
        RECT 91.390 178.715 91.680 178.945 ;
        RECT 85.410 178.560 85.700 178.605 ;
        RECT 86.790 178.560 87.080 178.605 ;
        RECT 85.410 178.420 87.080 178.560 ;
        RECT 85.410 178.375 85.700 178.420 ;
        RECT 86.790 178.375 87.080 178.420 ;
        RECT 87.235 178.560 87.555 178.620 ;
        RECT 88.170 178.560 88.460 178.605 ;
        RECT 87.235 178.420 88.460 178.560 ;
        RECT 87.235 178.360 87.555 178.420 ;
        RECT 88.170 178.375 88.460 178.420 ;
        RECT 95.975 178.360 96.295 178.620 ;
        RECT 96.435 178.560 96.755 178.620 ;
        RECT 102.430 178.560 102.720 178.605 ;
        RECT 96.435 178.420 102.720 178.560 ;
        RECT 96.435 178.360 96.755 178.420 ;
        RECT 102.430 178.375 102.720 178.420 ;
        RECT 105.635 178.360 105.955 178.620 ;
        RECT 51.345 178.220 51.635 178.265 ;
        RECT 53.205 178.220 53.495 178.265 ;
        RECT 51.345 178.080 53.495 178.220 ;
        RECT 51.345 178.035 51.635 178.080 ;
        RECT 53.205 178.035 53.495 178.080 ;
        RECT 72.990 178.220 73.280 178.265 ;
        RECT 75.390 178.220 75.980 178.265 ;
        RECT 78.630 178.220 79.280 178.265 ;
        RECT 72.990 178.080 79.280 178.220 ;
        RECT 72.990 178.035 73.280 178.080 ;
        RECT 75.390 178.035 75.680 178.080 ;
        RECT 78.630 178.035 79.280 178.080 ;
        RECT 50.435 178.020 50.755 178.035 ;
        RECT 81.255 178.020 81.575 178.280 ;
        RECT 85.855 178.220 86.175 178.280 ;
        RECT 91.850 178.220 92.140 178.265 ;
        RECT 85.855 178.080 92.140 178.220 ;
        RECT 85.855 178.020 86.175 178.080 ;
        RECT 91.850 178.035 92.140 178.080 ;
        RECT 31.575 177.880 31.895 177.940 ;
        RECT 32.510 177.880 32.800 177.925 ;
        RECT 31.575 177.740 32.800 177.880 ;
        RECT 31.575 177.680 31.895 177.740 ;
        RECT 32.510 177.695 32.800 177.740 ;
        RECT 38.475 177.680 38.795 177.940 ;
        RECT 43.995 177.680 44.315 177.940 ;
        RECT 45.160 177.880 45.450 177.925 ;
        RECT 49.515 177.880 49.835 177.940 ;
        RECT 45.160 177.740 49.835 177.880 ;
        RECT 45.160 177.695 45.450 177.740 ;
        RECT 49.515 177.680 49.835 177.740 ;
        RECT 58.715 177.680 59.035 177.940 ;
        RECT 60.095 177.680 60.415 177.940 ;
        RECT 67.455 177.680 67.775 177.940 ;
        RECT 68.850 177.880 69.140 177.925 ;
        RECT 71.135 177.880 71.455 177.940 ;
        RECT 68.850 177.740 71.455 177.880 ;
        RECT 68.850 177.695 69.140 177.740 ;
        RECT 71.135 177.680 71.455 177.740 ;
        RECT 73.910 177.880 74.200 177.925 ;
        RECT 74.815 177.880 75.135 177.940 ;
        RECT 73.910 177.740 75.135 177.880 ;
        RECT 73.910 177.695 74.200 177.740 ;
        RECT 74.815 177.680 75.135 177.740 ;
        RECT 84.950 177.880 85.240 177.925 ;
        RECT 85.395 177.880 85.715 177.940 ;
        RECT 84.950 177.740 85.715 177.880 ;
        RECT 84.950 177.695 85.240 177.740 ;
        RECT 85.395 177.680 85.715 177.740 ;
        RECT 87.250 177.880 87.540 177.925 ;
        RECT 87.695 177.880 88.015 177.940 ;
        RECT 87.250 177.740 88.015 177.880 ;
        RECT 87.250 177.695 87.540 177.740 ;
        RECT 87.695 177.680 88.015 177.740 ;
        RECT 89.090 177.880 89.380 177.925 ;
        RECT 89.995 177.880 90.315 177.940 ;
        RECT 89.090 177.740 90.315 177.880 ;
        RECT 89.090 177.695 89.380 177.740 ;
        RECT 89.995 177.680 90.315 177.740 ;
        RECT 92.295 177.880 92.615 177.940 ;
        RECT 93.675 177.880 93.995 177.940 ;
        RECT 92.295 177.740 93.995 177.880 ;
        RECT 92.295 177.680 92.615 177.740 ;
        RECT 93.675 177.680 93.995 177.740 ;
        RECT 102.415 177.880 102.735 177.940 ;
        RECT 102.890 177.880 103.180 177.925 ;
        RECT 102.415 177.740 103.180 177.880 ;
        RECT 102.415 177.680 102.735 177.740 ;
        RECT 102.890 177.695 103.180 177.740 ;
        RECT 106.570 177.880 106.860 177.925 ;
        RECT 107.015 177.880 107.335 177.940 ;
        RECT 106.570 177.740 107.335 177.880 ;
        RECT 106.570 177.695 106.860 177.740 ;
        RECT 107.015 177.680 107.335 177.740 ;
        RECT 17.370 177.060 112.465 177.540 ;
        RECT 26.055 176.660 26.375 176.920 ;
        RECT 27.895 176.660 28.215 176.920 ;
        RECT 28.600 176.860 28.890 176.905 ;
        RECT 37.095 176.860 37.415 176.920 ;
        RECT 47.000 176.860 47.290 176.905 ;
        RECT 48.135 176.860 48.455 176.920 ;
        RECT 28.600 176.720 45.605 176.860 ;
        RECT 28.600 176.675 28.890 176.720 ;
        RECT 37.095 176.660 37.415 176.720 ;
        RECT 30.605 176.520 30.895 176.565 ;
        RECT 32.035 176.520 32.355 176.580 ;
        RECT 33.865 176.520 34.155 176.565 ;
        RECT 30.605 176.380 34.155 176.520 ;
        RECT 30.605 176.335 30.895 176.380 ;
        RECT 32.035 176.320 32.355 176.380 ;
        RECT 33.865 176.335 34.155 176.380 ;
        RECT 34.785 176.520 35.075 176.565 ;
        RECT 36.645 176.520 36.935 176.565 ;
        RECT 34.785 176.380 36.935 176.520 ;
        RECT 34.785 176.335 35.075 176.380 ;
        RECT 36.645 176.335 36.935 176.380 ;
        RECT 38.955 176.520 39.245 176.565 ;
        RECT 40.815 176.520 41.105 176.565 ;
        RECT 38.955 176.380 41.105 176.520 ;
        RECT 38.955 176.335 39.245 176.380 ;
        RECT 40.815 176.335 41.105 176.380 ;
        RECT 41.735 176.520 42.025 176.565 ;
        RECT 43.995 176.520 44.315 176.580 ;
        RECT 44.995 176.520 45.285 176.565 ;
        RECT 41.735 176.380 45.285 176.520 ;
        RECT 45.465 176.520 45.605 176.720 ;
        RECT 47.000 176.720 48.455 176.860 ;
        RECT 47.000 176.675 47.290 176.720 ;
        RECT 48.135 176.660 48.455 176.720 ;
        RECT 49.515 176.660 49.835 176.920 ;
        RECT 51.830 176.675 52.120 176.905 ;
        RECT 52.275 176.860 52.595 176.920 ;
        RECT 53.210 176.860 53.500 176.905 ;
        RECT 52.275 176.720 53.500 176.860 ;
        RECT 49.990 176.520 50.280 176.565 ;
        RECT 45.465 176.380 50.280 176.520 ;
        RECT 41.735 176.335 42.025 176.380 ;
        RECT 24.675 176.180 24.995 176.240 ;
        RECT 25.610 176.180 25.900 176.225 ;
        RECT 24.675 176.040 25.900 176.180 ;
        RECT 24.675 175.980 24.995 176.040 ;
        RECT 25.610 175.995 25.900 176.040 ;
        RECT 32.465 176.180 32.755 176.225 ;
        RECT 34.785 176.180 35.000 176.335 ;
        RECT 32.465 176.040 35.000 176.180 ;
        RECT 35.730 176.180 36.020 176.225 ;
        RECT 38.475 176.180 38.795 176.240 ;
        RECT 35.730 176.040 38.795 176.180 ;
        RECT 40.890 176.180 41.105 176.335 ;
        RECT 43.995 176.320 44.315 176.380 ;
        RECT 44.995 176.335 45.285 176.380 ;
        RECT 49.990 176.335 50.280 176.380 ;
        RECT 43.135 176.180 43.425 176.225 ;
        RECT 40.890 176.040 43.425 176.180 ;
        RECT 51.905 176.180 52.045 176.675 ;
        RECT 52.275 176.660 52.595 176.720 ;
        RECT 53.210 176.675 53.500 176.720 ;
        RECT 57.795 176.660 58.115 176.920 ;
        RECT 61.475 176.860 61.795 176.920 ;
        RECT 61.950 176.860 62.240 176.905 ;
        RECT 61.475 176.720 62.240 176.860 ;
        RECT 61.475 176.660 61.795 176.720 ;
        RECT 61.950 176.675 62.240 176.720 ;
        RECT 80.810 176.860 81.100 176.905 ;
        RECT 81.255 176.860 81.575 176.920 ;
        RECT 89.995 176.860 90.315 176.920 ;
        RECT 80.810 176.720 81.575 176.860 ;
        RECT 80.810 176.675 81.100 176.720 ;
        RECT 81.255 176.660 81.575 176.720 ;
        RECT 89.165 176.720 90.315 176.860 ;
        RECT 56.875 176.520 57.195 176.580 ;
        RECT 59.635 176.520 59.955 176.580 ;
        RECT 56.875 176.380 59.955 176.520 ;
        RECT 56.875 176.320 57.195 176.380 ;
        RECT 59.635 176.320 59.955 176.380 ;
        RECT 65.270 176.520 65.560 176.565 ;
        RECT 67.455 176.520 67.775 176.580 ;
        RECT 68.510 176.520 69.160 176.565 ;
        RECT 65.270 176.380 69.160 176.520 ;
        RECT 65.270 176.335 65.860 176.380 ;
        RECT 52.290 176.180 52.580 176.225 ;
        RECT 51.905 176.040 52.580 176.180 ;
        RECT 32.465 175.995 32.755 176.040 ;
        RECT 35.730 175.995 36.020 176.040 ;
        RECT 38.475 175.980 38.795 176.040 ;
        RECT 43.135 175.995 43.425 176.040 ;
        RECT 52.290 175.995 52.580 176.040 ;
        RECT 58.715 175.980 59.035 176.240 ;
        RECT 65.570 176.020 65.860 176.335 ;
        RECT 67.455 176.320 67.775 176.380 ;
        RECT 68.510 176.335 69.160 176.380 ;
        RECT 71.135 176.320 71.455 176.580 ;
        RECT 83.210 176.520 83.500 176.565 ;
        RECT 85.395 176.520 85.715 176.580 ;
        RECT 89.165 176.565 89.305 176.720 ;
        RECT 89.995 176.660 90.315 176.720 ;
        RECT 86.450 176.520 87.100 176.565 ;
        RECT 83.210 176.380 87.100 176.520 ;
        RECT 83.210 176.335 83.800 176.380 ;
        RECT 66.650 176.180 66.940 176.225 ;
        RECT 70.230 176.180 70.520 176.225 ;
        RECT 72.065 176.180 72.355 176.225 ;
        RECT 66.650 176.040 72.355 176.180 ;
        RECT 66.650 175.995 66.940 176.040 ;
        RECT 70.230 175.995 70.520 176.040 ;
        RECT 72.065 175.995 72.355 176.040 ;
        RECT 79.875 175.980 80.195 176.240 ;
        RECT 83.510 176.020 83.800 176.335 ;
        RECT 85.395 176.320 85.715 176.380 ;
        RECT 86.450 176.335 87.100 176.380 ;
        RECT 89.090 176.335 89.380 176.565 ;
        RECT 90.455 176.320 90.775 176.580 ;
        RECT 101.610 176.520 101.900 176.565 ;
        RECT 102.415 176.520 102.735 176.580 ;
        RECT 104.850 176.520 105.500 176.565 ;
        RECT 101.610 176.380 105.500 176.520 ;
        RECT 101.610 176.335 102.200 176.380 ;
        RECT 84.590 176.180 84.880 176.225 ;
        RECT 88.170 176.180 88.460 176.225 ;
        RECT 90.005 176.180 90.295 176.225 ;
        RECT 84.590 176.040 90.295 176.180 ;
        RECT 90.545 176.180 90.685 176.320 ;
        RECT 96.435 176.180 96.755 176.240 ;
        RECT 97.830 176.180 98.120 176.225 ;
        RECT 90.545 176.040 98.120 176.180 ;
        RECT 84.590 175.995 84.880 176.040 ;
        RECT 88.170 175.995 88.460 176.040 ;
        RECT 90.005 175.995 90.295 176.040 ;
        RECT 96.435 175.980 96.755 176.040 ;
        RECT 97.830 175.995 98.120 176.040 ;
        RECT 101.910 176.020 102.200 176.335 ;
        RECT 102.415 176.320 102.735 176.380 ;
        RECT 104.850 176.335 105.500 176.380 ;
        RECT 102.990 176.180 103.280 176.225 ;
        RECT 106.570 176.180 106.860 176.225 ;
        RECT 108.405 176.180 108.695 176.225 ;
        RECT 102.990 176.040 108.695 176.180 ;
        RECT 102.990 175.995 103.280 176.040 ;
        RECT 106.570 175.995 106.860 176.040 ;
        RECT 108.405 175.995 108.695 176.040 ;
        RECT 25.150 175.840 25.440 175.885 ;
        RECT 32.955 175.840 33.275 175.900 ;
        RECT 25.150 175.700 33.275 175.840 ;
        RECT 25.150 175.655 25.440 175.700 ;
        RECT 32.955 175.640 33.275 175.700 ;
        RECT 37.570 175.840 37.860 175.885 ;
        RECT 38.030 175.840 38.320 175.885 ;
        RECT 38.935 175.840 39.255 175.900 ;
        RECT 37.570 175.700 39.255 175.840 ;
        RECT 37.570 175.655 37.860 175.700 ;
        RECT 38.030 175.655 38.320 175.700 ;
        RECT 38.935 175.640 39.255 175.700 ;
        RECT 39.870 175.840 40.160 175.885 ;
        RECT 44.455 175.840 44.775 175.900 ;
        RECT 39.870 175.700 44.775 175.840 ;
        RECT 39.870 175.655 40.160 175.700 ;
        RECT 44.455 175.640 44.775 175.700 ;
        RECT 48.610 175.655 48.900 175.885 ;
        RECT 58.805 175.840 58.945 175.980 ;
        RECT 62.410 175.840 62.700 175.885 ;
        RECT 63.790 175.840 64.080 175.885 ;
        RECT 58.805 175.700 64.080 175.840 ;
        RECT 62.410 175.655 62.700 175.700 ;
        RECT 63.790 175.655 64.080 175.700 ;
        RECT 72.530 175.840 72.820 175.885 ;
        RECT 90.455 175.840 90.775 175.900 ;
        RECT 96.895 175.840 97.215 175.900 ;
        RECT 72.530 175.700 74.125 175.840 ;
        RECT 72.530 175.655 72.820 175.700 ;
        RECT 32.465 175.500 32.755 175.545 ;
        RECT 35.245 175.500 35.535 175.545 ;
        RECT 37.105 175.500 37.395 175.545 ;
        RECT 32.465 175.360 37.395 175.500 ;
        RECT 32.465 175.315 32.755 175.360 ;
        RECT 35.245 175.315 35.535 175.360 ;
        RECT 37.105 175.315 37.395 175.360 ;
        RECT 38.495 175.500 38.785 175.545 ;
        RECT 40.355 175.500 40.645 175.545 ;
        RECT 43.135 175.500 43.425 175.545 ;
        RECT 38.495 175.360 43.425 175.500 ;
        RECT 38.495 175.315 38.785 175.360 ;
        RECT 40.355 175.315 40.645 175.360 ;
        RECT 43.135 175.315 43.425 175.360 ;
        RECT 48.685 175.500 48.825 175.655 ;
        RECT 49.055 175.500 49.375 175.560 ;
        RECT 48.685 175.360 49.375 175.500 ;
        RECT 37.555 175.160 37.875 175.220 ;
        RECT 48.685 175.160 48.825 175.360 ;
        RECT 49.055 175.300 49.375 175.360 ;
        RECT 59.650 175.500 59.940 175.545 ;
        RECT 61.475 175.500 61.795 175.560 ;
        RECT 59.650 175.360 61.795 175.500 ;
        RECT 59.650 175.315 59.940 175.360 ;
        RECT 61.475 175.300 61.795 175.360 ;
        RECT 66.650 175.500 66.940 175.545 ;
        RECT 69.770 175.500 70.060 175.545 ;
        RECT 71.660 175.500 71.950 175.545 ;
        RECT 66.650 175.360 71.950 175.500 ;
        RECT 73.985 175.500 74.125 175.700 ;
        RECT 90.455 175.700 97.215 175.840 ;
        RECT 90.455 175.640 90.775 175.700 ;
        RECT 96.895 175.640 97.215 175.700 ;
        RECT 98.275 175.640 98.595 175.900 ;
        RECT 108.855 175.640 109.175 175.900 ;
        RECT 82.635 175.500 82.955 175.560 ;
        RECT 73.985 175.360 82.955 175.500 ;
        RECT 66.650 175.315 66.940 175.360 ;
        RECT 69.770 175.315 70.060 175.360 ;
        RECT 71.660 175.315 71.950 175.360 ;
        RECT 82.635 175.300 82.955 175.360 ;
        RECT 84.590 175.500 84.880 175.545 ;
        RECT 87.710 175.500 88.000 175.545 ;
        RECT 89.600 175.500 89.890 175.545 ;
        RECT 84.590 175.360 89.890 175.500 ;
        RECT 84.590 175.315 84.880 175.360 ;
        RECT 87.710 175.315 88.000 175.360 ;
        RECT 89.600 175.315 89.890 175.360 ;
        RECT 102.990 175.500 103.280 175.545 ;
        RECT 106.110 175.500 106.400 175.545 ;
        RECT 108.000 175.500 108.290 175.545 ;
        RECT 102.990 175.360 108.290 175.500 ;
        RECT 102.990 175.315 103.280 175.360 ;
        RECT 106.110 175.315 106.400 175.360 ;
        RECT 108.000 175.315 108.290 175.360 ;
        RECT 37.555 175.020 48.825 175.160 ;
        RECT 62.395 175.160 62.715 175.220 ;
        RECT 63.330 175.160 63.620 175.205 ;
        RECT 62.395 175.020 63.620 175.160 ;
        RECT 37.555 174.960 37.875 175.020 ;
        RECT 62.395 174.960 62.715 175.020 ;
        RECT 63.330 174.975 63.620 175.020 ;
        RECT 81.715 174.960 82.035 175.220 ;
        RECT 100.130 175.160 100.420 175.205 ;
        RECT 101.955 175.160 102.275 175.220 ;
        RECT 100.130 175.020 102.275 175.160 ;
        RECT 100.130 174.975 100.420 175.020 ;
        RECT 101.955 174.960 102.275 175.020 ;
        RECT 107.585 175.160 107.875 175.205 ;
        RECT 108.395 175.160 108.715 175.220 ;
        RECT 107.585 175.020 108.715 175.160 ;
        RECT 107.585 174.975 107.875 175.020 ;
        RECT 108.395 174.960 108.715 175.020 ;
        RECT 18.165 174.340 112.465 174.820 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 26.070 174.140 26.360 174.185 ;
        RECT 31.575 174.140 31.895 174.200 ;
        RECT 26.070 174.000 31.895 174.140 ;
        RECT 26.070 173.955 26.360 174.000 ;
        RECT 31.575 173.940 31.895 174.000 ;
        RECT 32.035 173.940 32.355 174.200 ;
        RECT 34.350 174.140 34.640 174.185 ;
        RECT 38.015 174.140 38.335 174.200 ;
        RECT 34.350 174.000 38.335 174.140 ;
        RECT 34.350 173.955 34.640 174.000 ;
        RECT 38.015 173.940 38.335 174.000 ;
        RECT 44.455 173.940 44.775 174.200 ;
        RECT 50.435 173.940 50.755 174.200 ;
        RECT 88.170 174.140 88.460 174.185 ;
        RECT 94.595 174.140 94.915 174.200 ;
        RECT 88.170 174.000 94.915 174.140 ;
        RECT 88.170 173.955 88.460 174.000 ;
        RECT 94.595 173.940 94.915 174.000 ;
        RECT 96.895 174.140 97.215 174.200 ;
        RECT 108.395 174.140 108.715 174.200 ;
        RECT 108.870 174.140 109.160 174.185 ;
        RECT 96.895 174.000 108.165 174.140 ;
        RECT 96.895 173.940 97.215 174.000 ;
        RECT 32.125 173.800 32.265 173.940 ;
        RECT 38.950 173.800 39.240 173.845 ;
        RECT 32.125 173.660 39.240 173.800 ;
        RECT 38.950 173.615 39.240 173.660 ;
        RECT 59.635 173.800 59.955 173.860 ;
        RECT 79.990 173.800 80.280 173.845 ;
        RECT 83.110 173.800 83.400 173.845 ;
        RECT 85.000 173.800 85.290 173.845 ;
        RECT 59.635 173.660 62.625 173.800 ;
        RECT 59.635 173.600 59.955 173.660 ;
        RECT 31.590 173.275 31.880 173.505 ;
        RECT 32.050 173.460 32.340 173.505 ;
        RECT 37.095 173.460 37.415 173.520 ;
        RECT 44.915 173.460 45.235 173.520 ;
        RECT 32.050 173.320 37.415 173.460 ;
        RECT 32.050 173.275 32.340 173.320 ;
        RECT 23.310 172.935 23.600 173.165 ;
        RECT 31.665 173.120 31.805 173.275 ;
        RECT 37.095 173.260 37.415 173.320 ;
        RECT 39.485 173.320 46.525 173.460 ;
        RECT 37.555 173.120 37.875 173.180 ;
        RECT 39.485 173.165 39.625 173.320 ;
        RECT 44.915 173.260 45.235 173.320 ;
        RECT 31.665 172.980 37.875 173.120 ;
        RECT 23.385 172.780 23.525 172.935 ;
        RECT 37.555 172.920 37.875 172.980 ;
        RECT 39.410 172.935 39.700 173.165 ;
        RECT 45.390 173.120 45.680 173.165 ;
        RECT 45.390 172.980 46.065 173.120 ;
        RECT 45.390 172.935 45.680 172.980 ;
        RECT 24.675 172.780 24.995 172.840 ;
        RECT 32.035 172.780 32.355 172.840 ;
        RECT 23.385 172.640 32.355 172.780 ;
        RECT 24.675 172.580 24.995 172.640 ;
        RECT 32.035 172.580 32.355 172.640 ;
        RECT 32.510 172.440 32.800 172.485 ;
        RECT 33.415 172.440 33.735 172.500 ;
        RECT 32.510 172.300 33.735 172.440 ;
        RECT 32.510 172.255 32.800 172.300 ;
        RECT 33.415 172.240 33.735 172.300 ;
        RECT 34.795 172.440 35.115 172.500 ;
        RECT 37.555 172.440 37.875 172.500 ;
        RECT 45.925 172.485 46.065 172.980 ;
        RECT 46.385 172.840 46.525 173.320 ;
        RECT 48.135 173.260 48.455 173.520 ;
        RECT 49.055 173.460 49.375 173.520 ;
        RECT 54.115 173.460 54.435 173.520 ;
        RECT 49.055 173.320 54.435 173.460 ;
        RECT 49.055 173.260 49.375 173.320 ;
        RECT 54.115 173.260 54.435 173.320 ;
        RECT 61.475 173.260 61.795 173.520 ;
        RECT 61.935 173.260 62.255 173.520 ;
        RECT 62.485 173.505 62.625 173.660 ;
        RECT 79.990 173.660 85.290 173.800 ;
        RECT 79.990 173.615 80.280 173.660 ;
        RECT 83.110 173.615 83.400 173.660 ;
        RECT 85.000 173.615 85.290 173.660 ;
        RECT 91.030 173.800 91.320 173.845 ;
        RECT 94.150 173.800 94.440 173.845 ;
        RECT 96.040 173.800 96.330 173.845 ;
        RECT 91.030 173.660 96.330 173.800 ;
        RECT 91.030 173.615 91.320 173.660 ;
        RECT 94.150 173.615 94.440 173.660 ;
        RECT 96.040 173.615 96.330 173.660 ;
        RECT 98.290 173.800 98.580 173.845 ;
        RECT 98.735 173.800 99.055 173.860 ;
        RECT 98.290 173.660 99.055 173.800 ;
        RECT 98.290 173.615 98.580 173.660 ;
        RECT 98.735 173.600 99.055 173.660 ;
        RECT 102.530 173.800 102.820 173.845 ;
        RECT 105.650 173.800 105.940 173.845 ;
        RECT 107.540 173.800 107.830 173.845 ;
        RECT 102.530 173.660 107.830 173.800 ;
        RECT 102.530 173.615 102.820 173.660 ;
        RECT 105.650 173.615 105.940 173.660 ;
        RECT 107.540 173.615 107.830 173.660 ;
        RECT 62.410 173.275 62.700 173.505 ;
        RECT 62.870 173.460 63.160 173.505 ;
        RECT 63.775 173.460 64.095 173.520 ;
        RECT 62.870 173.320 64.095 173.460 ;
        RECT 62.870 173.275 63.160 173.320 ;
        RECT 63.775 173.260 64.095 173.320 ;
        RECT 74.355 173.460 74.675 173.520 ;
        RECT 84.490 173.460 84.780 173.505 ;
        RECT 95.515 173.460 95.835 173.520 ;
        RECT 74.355 173.320 75.965 173.460 ;
        RECT 74.355 173.260 74.675 173.320 ;
        RECT 46.755 173.120 47.075 173.180 ;
        RECT 47.690 173.120 47.980 173.165 ;
        RECT 49.515 173.120 49.835 173.180 ;
        RECT 46.755 172.980 49.835 173.120 ;
        RECT 46.755 172.920 47.075 172.980 ;
        RECT 47.690 172.935 47.980 172.980 ;
        RECT 49.515 172.920 49.835 172.980 ;
        RECT 50.910 172.935 51.200 173.165 ;
        RECT 59.635 173.120 59.955 173.180 ;
        RECT 70.230 173.120 70.520 173.165 ;
        RECT 59.635 172.980 70.520 173.120 ;
        RECT 46.295 172.780 46.615 172.840 ;
        RECT 50.985 172.780 51.125 172.935 ;
        RECT 59.635 172.920 59.955 172.980 ;
        RECT 70.230 172.935 70.520 172.980 ;
        RECT 72.515 173.120 72.835 173.180 ;
        RECT 75.825 173.165 75.965 173.320 ;
        RECT 84.490 173.320 95.835 173.460 ;
        RECT 84.490 173.275 84.780 173.320 ;
        RECT 95.515 173.260 95.835 173.320 ;
        RECT 96.895 173.260 97.215 173.520 ;
        RECT 107.015 173.260 107.335 173.520 ;
        RECT 108.025 173.460 108.165 174.000 ;
        RECT 108.395 174.000 109.160 174.140 ;
        RECT 108.395 173.940 108.715 174.000 ;
        RECT 108.870 173.955 109.160 174.000 ;
        RECT 108.410 173.460 108.700 173.505 ;
        RECT 108.855 173.460 109.175 173.520 ;
        RECT 108.025 173.320 109.175 173.460 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 108.410 173.275 108.700 173.320 ;
        RECT 108.855 173.260 109.175 173.320 ;
        RECT 72.990 173.120 73.280 173.165 ;
        RECT 72.515 172.980 73.280 173.120 ;
        RECT 72.515 172.920 72.835 172.980 ;
        RECT 72.990 172.935 73.280 172.980 ;
        RECT 75.750 172.935 76.040 173.165 ;
        RECT 46.295 172.640 51.125 172.780 ;
        RECT 63.315 172.780 63.635 172.840 ;
        RECT 63.790 172.780 64.080 172.825 ;
        RECT 63.315 172.640 64.080 172.780 ;
        RECT 46.295 172.580 46.615 172.640 ;
        RECT 63.315 172.580 63.635 172.640 ;
        RECT 63.790 172.595 64.080 172.640 ;
        RECT 66.535 172.780 66.855 172.840 ;
        RECT 67.470 172.780 67.760 172.825 ;
        RECT 66.535 172.640 67.760 172.780 ;
        RECT 66.535 172.580 66.855 172.640 ;
        RECT 67.470 172.595 67.760 172.640 ;
        RECT 69.310 172.780 69.600 172.825 ;
        RECT 73.895 172.780 74.215 172.840 ;
        RECT 78.910 172.825 79.200 173.140 ;
        RECT 79.990 173.120 80.280 173.165 ;
        RECT 83.570 173.120 83.860 173.165 ;
        RECT 85.405 173.120 85.695 173.165 ;
        RECT 79.990 172.980 85.695 173.120 ;
        RECT 79.990 172.935 80.280 172.980 ;
        RECT 83.570 172.935 83.860 172.980 ;
        RECT 85.405 172.935 85.695 172.980 ;
        RECT 85.870 172.935 86.160 173.165 ;
        RECT 69.310 172.640 74.215 172.780 ;
        RECT 69.310 172.595 69.600 172.640 ;
        RECT 73.895 172.580 74.215 172.640 ;
        RECT 76.210 172.780 76.500 172.825 ;
        RECT 78.610 172.780 79.200 172.825 ;
        RECT 81.850 172.780 82.500 172.825 ;
        RECT 85.945 172.780 86.085 172.935 ;
        RECT 87.695 172.920 88.015 173.180 ;
        RECT 76.210 172.640 82.500 172.780 ;
        RECT 76.210 172.595 76.500 172.640 ;
        RECT 78.610 172.595 78.900 172.640 ;
        RECT 81.850 172.595 82.500 172.640 ;
        RECT 82.725 172.640 86.085 172.780 ;
        RECT 88.155 172.780 88.475 172.840 ;
        RECT 89.950 172.825 90.240 173.140 ;
        RECT 91.030 173.120 91.320 173.165 ;
        RECT 94.610 173.120 94.900 173.165 ;
        RECT 96.445 173.120 96.735 173.165 ;
        RECT 97.830 173.120 98.120 173.165 ;
        RECT 91.030 172.980 96.735 173.120 ;
        RECT 91.030 172.935 91.320 172.980 ;
        RECT 94.610 172.935 94.900 172.980 ;
        RECT 96.445 172.935 96.735 172.980 ;
        RECT 97.445 172.980 98.120 173.120 ;
        RECT 89.650 172.780 90.240 172.825 ;
        RECT 92.890 172.780 93.540 172.825 ;
        RECT 88.155 172.640 93.540 172.780 ;
        RECT 82.725 172.500 82.865 172.640 ;
        RECT 88.155 172.580 88.475 172.640 ;
        RECT 89.650 172.595 89.940 172.640 ;
        RECT 92.890 172.595 93.540 172.640 ;
        RECT 95.530 172.780 95.820 172.825 ;
        RECT 96.895 172.780 97.215 172.840 ;
        RECT 95.530 172.640 97.215 172.780 ;
        RECT 95.530 172.595 95.820 172.640 ;
        RECT 96.895 172.580 97.215 172.640 ;
        RECT 34.795 172.300 37.875 172.440 ;
        RECT 34.795 172.240 35.115 172.300 ;
        RECT 37.555 172.240 37.875 172.300 ;
        RECT 45.850 172.255 46.140 172.485 ;
        RECT 70.215 172.440 70.535 172.500 ;
        RECT 70.690 172.440 70.980 172.485 ;
        RECT 70.215 172.300 70.980 172.440 ;
        RECT 70.215 172.240 70.535 172.300 ;
        RECT 70.690 172.255 70.980 172.300 ;
        RECT 77.130 172.440 77.420 172.485 ;
        RECT 81.255 172.440 81.575 172.500 ;
        RECT 77.130 172.300 81.575 172.440 ;
        RECT 77.130 172.255 77.420 172.300 ;
        RECT 81.255 172.240 81.575 172.300 ;
        RECT 82.635 172.240 82.955 172.500 ;
        RECT 86.775 172.440 87.095 172.500 ;
        RECT 87.250 172.440 87.540 172.485 ;
        RECT 86.775 172.300 87.540 172.440 ;
        RECT 86.775 172.240 87.095 172.300 ;
        RECT 87.250 172.255 87.540 172.300 ;
        RECT 96.435 172.440 96.755 172.500 ;
        RECT 97.445 172.440 97.585 172.980 ;
        RECT 97.830 172.935 98.120 172.980 ;
        RECT 98.275 172.780 98.595 172.840 ;
        RECT 101.450 172.825 101.740 173.140 ;
        RECT 102.530 173.120 102.820 173.165 ;
        RECT 106.110 173.120 106.400 173.165 ;
        RECT 107.945 173.120 108.235 173.165 ;
        RECT 102.530 172.980 108.235 173.120 ;
        RECT 102.530 172.935 102.820 172.980 ;
        RECT 106.110 172.935 106.400 172.980 ;
        RECT 107.945 172.935 108.235 172.980 ;
        RECT 109.790 172.935 110.080 173.165 ;
        RECT 101.150 172.780 101.740 172.825 ;
        RECT 104.390 172.780 105.040 172.825 ;
        RECT 98.275 172.640 105.040 172.780 ;
        RECT 98.275 172.580 98.595 172.640 ;
        RECT 101.150 172.595 101.440 172.640 ;
        RECT 104.390 172.595 105.040 172.640 ;
        RECT 96.435 172.300 97.585 172.440 ;
        RECT 99.670 172.440 99.960 172.485 ;
        RECT 102.875 172.440 103.195 172.500 ;
        RECT 99.670 172.300 103.195 172.440 ;
        RECT 96.435 172.240 96.755 172.300 ;
        RECT 99.670 172.255 99.960 172.300 ;
        RECT 102.875 172.240 103.195 172.300 ;
        RECT 103.795 172.440 104.115 172.500 ;
        RECT 109.865 172.440 110.005 172.935 ;
        RECT 103.795 172.300 110.005 172.440 ;
        RECT 103.795 172.240 104.115 172.300 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 17.370 171.620 112.465 172.100 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 21.010 171.420 21.300 171.465 ;
        RECT 31.130 171.420 31.420 171.465 ;
        RECT 32.035 171.420 32.355 171.480 ;
        RECT 49.055 171.420 49.375 171.480 ;
        RECT 21.010 171.280 25.825 171.420 ;
        RECT 21.010 171.235 21.300 171.280 ;
        RECT 23.755 170.880 24.075 171.140 ;
        RECT 25.685 171.080 25.825 171.280 ;
        RECT 31.130 171.280 32.355 171.420 ;
        RECT 31.130 171.235 31.420 171.280 ;
        RECT 32.035 171.220 32.355 171.280 ;
        RECT 43.625 171.280 47.905 171.420 ;
        RECT 26.050 171.080 26.700 171.125 ;
        RECT 29.650 171.080 29.940 171.125 ;
        RECT 38.015 171.080 38.335 171.140 ;
        RECT 25.685 170.940 29.940 171.080 ;
        RECT 26.050 170.895 26.700 170.940 ;
        RECT 29.350 170.895 29.940 170.940 ;
        RECT 33.045 170.940 38.335 171.080 ;
        RECT 20.535 170.740 20.855 170.800 ;
        RECT 21.915 170.740 22.235 170.800 ;
        RECT 20.535 170.600 22.235 170.740 ;
        RECT 20.535 170.540 20.855 170.600 ;
        RECT 21.915 170.540 22.235 170.600 ;
        RECT 22.855 170.740 23.145 170.785 ;
        RECT 24.690 170.740 24.980 170.785 ;
        RECT 28.270 170.740 28.560 170.785 ;
        RECT 22.855 170.600 28.560 170.740 ;
        RECT 22.855 170.555 23.145 170.600 ;
        RECT 24.690 170.555 24.980 170.600 ;
        RECT 28.270 170.555 28.560 170.600 ;
        RECT 29.350 170.580 29.640 170.895 ;
        RECT 33.045 170.800 33.185 170.940 ;
        RECT 31.590 170.555 31.880 170.785 ;
        RECT 22.390 170.400 22.680 170.445 ;
        RECT 28.815 170.400 29.135 170.460 ;
        RECT 22.390 170.260 29.135 170.400 ;
        RECT 22.390 170.215 22.680 170.260 ;
        RECT 28.815 170.200 29.135 170.260 ;
        RECT 31.115 170.400 31.435 170.460 ;
        RECT 31.665 170.400 31.805 170.555 ;
        RECT 32.495 170.540 32.815 170.800 ;
        RECT 32.955 170.540 33.275 170.800 ;
        RECT 33.430 170.740 33.720 170.785 ;
        RECT 34.335 170.740 34.655 170.800 ;
        RECT 36.635 170.740 36.955 170.800 ;
        RECT 37.185 170.785 37.325 170.940 ;
        RECT 38.015 170.880 38.335 170.940 ;
        RECT 40.315 171.080 40.635 171.140 ;
        RECT 43.625 171.080 43.765 171.280 ;
        RECT 46.755 171.080 47.075 171.140 ;
        RECT 40.315 170.940 43.765 171.080 ;
        RECT 45.465 170.940 47.075 171.080 ;
        RECT 47.765 171.080 47.905 171.280 ;
        RECT 49.055 171.280 51.125 171.420 ;
        RECT 49.055 171.220 49.375 171.280 ;
        RECT 47.765 170.940 50.665 171.080 ;
        RECT 40.315 170.880 40.635 170.940 ;
        RECT 33.430 170.600 36.955 170.740 ;
        RECT 33.430 170.555 33.720 170.600 ;
        RECT 34.335 170.540 34.655 170.600 ;
        RECT 36.635 170.540 36.955 170.600 ;
        RECT 37.110 170.555 37.400 170.785 ;
        RECT 37.555 170.540 37.875 170.800 ;
        RECT 38.490 170.555 38.780 170.785 ;
        RECT 42.155 170.740 42.475 170.800 ;
        RECT 44.470 170.740 44.760 170.785 ;
        RECT 42.155 170.600 44.760 170.740 ;
        RECT 38.565 170.400 38.705 170.555 ;
        RECT 42.155 170.540 42.475 170.600 ;
        RECT 44.470 170.555 44.760 170.600 ;
        RECT 40.315 170.400 40.635 170.460 ;
        RECT 31.115 170.260 40.635 170.400 ;
        RECT 31.115 170.200 31.435 170.260 ;
        RECT 40.315 170.200 40.635 170.260 ;
        RECT 23.260 170.060 23.550 170.105 ;
        RECT 25.150 170.060 25.440 170.105 ;
        RECT 28.270 170.060 28.560 170.105 ;
        RECT 23.260 169.920 28.560 170.060 ;
        RECT 23.260 169.875 23.550 169.920 ;
        RECT 25.150 169.875 25.440 169.920 ;
        RECT 28.270 169.875 28.560 169.920 ;
        RECT 34.810 170.060 35.100 170.105 ;
        RECT 36.635 170.060 36.955 170.120 ;
        RECT 34.810 169.920 36.955 170.060 ;
        RECT 44.545 170.060 44.685 170.555 ;
        RECT 44.915 170.540 45.235 170.800 ;
        RECT 45.465 170.785 45.605 170.940 ;
        RECT 46.755 170.880 47.075 170.940 ;
        RECT 45.390 170.555 45.680 170.785 ;
        RECT 46.310 170.740 46.600 170.785 ;
        RECT 47.675 170.740 47.995 170.800 ;
        RECT 49.055 170.740 49.375 170.800 ;
        RECT 46.310 170.600 49.375 170.740 ;
        RECT 46.310 170.555 46.600 170.600 ;
        RECT 47.675 170.540 47.995 170.600 ;
        RECT 49.055 170.540 49.375 170.600 ;
        RECT 49.530 170.555 49.820 170.785 ;
        RECT 49.605 170.120 49.745 170.555 ;
        RECT 49.975 170.540 50.295 170.800 ;
        RECT 50.525 170.785 50.665 170.940 ;
        RECT 50.450 170.555 50.740 170.785 ;
        RECT 50.985 170.740 51.125 171.280 ;
        RECT 54.115 171.220 54.435 171.480 ;
        RECT 61.475 171.420 61.795 171.480 ;
        RECT 66.550 171.420 66.840 171.465 ;
        RECT 60.645 171.280 70.445 171.420 ;
        RECT 55.510 171.080 55.800 171.125 ;
        RECT 59.635 171.080 59.955 171.140 ;
        RECT 55.510 170.940 59.955 171.080 ;
        RECT 55.510 170.895 55.800 170.940 ;
        RECT 59.635 170.880 59.955 170.940 ;
        RECT 51.340 170.740 51.630 170.785 ;
        RECT 50.985 170.600 51.630 170.740 ;
        RECT 51.340 170.555 51.630 170.600 ;
        RECT 57.335 170.540 57.655 170.800 ;
        RECT 59.175 170.740 59.495 170.800 ;
        RECT 60.645 170.785 60.785 171.280 ;
        RECT 61.475 171.220 61.795 171.280 ;
        RECT 66.550 171.235 66.840 171.280 ;
        RECT 61.935 171.080 62.255 171.140 ;
        RECT 62.855 171.080 63.175 171.140 ;
        RECT 61.565 170.940 63.175 171.080 ;
        RECT 61.565 170.785 61.705 170.940 ;
        RECT 61.935 170.880 62.255 170.940 ;
        RECT 62.855 170.880 63.175 170.940 ;
        RECT 64.235 170.880 64.555 171.140 ;
        RECT 66.625 170.940 69.525 171.080 ;
        RECT 60.110 170.740 60.400 170.785 ;
        RECT 59.175 170.600 60.400 170.740 ;
        RECT 59.175 170.540 59.495 170.600 ;
        RECT 60.110 170.555 60.400 170.600 ;
        RECT 60.570 170.555 60.860 170.785 ;
        RECT 61.490 170.555 61.780 170.785 ;
        RECT 62.945 170.740 63.085 170.880 ;
        RECT 66.625 170.760 66.765 170.940 ;
        RECT 67.010 170.760 67.300 170.785 ;
        RECT 66.625 170.740 67.300 170.760 ;
        RECT 62.945 170.620 67.300 170.740 ;
        RECT 62.945 170.600 66.765 170.620 ;
        RECT 67.010 170.555 67.300 170.620 ;
        RECT 67.455 170.740 67.775 170.800 ;
        RECT 69.385 170.785 69.525 170.940 ;
        RECT 70.305 170.785 70.445 171.280 ;
        RECT 72.990 171.235 73.280 171.465 ;
        RECT 73.895 171.420 74.215 171.480 ;
        RECT 84.015 171.420 84.335 171.480 ;
        RECT 73.895 171.280 84.335 171.420 ;
        RECT 68.850 170.740 69.140 170.785 ;
        RECT 67.455 170.600 69.140 170.740 ;
        RECT 67.455 170.540 67.775 170.600 ;
        RECT 68.850 170.555 69.140 170.600 ;
        RECT 69.310 170.555 69.600 170.785 ;
        RECT 70.230 170.555 70.520 170.785 ;
        RECT 72.055 170.540 72.375 170.800 ;
        RECT 73.065 170.740 73.205 171.235 ;
        RECT 73.895 171.220 74.215 171.280 ;
        RECT 84.015 171.220 84.335 171.280 ;
        RECT 87.235 171.220 87.555 171.480 ;
        RECT 92.770 171.420 93.060 171.465 ;
        RECT 94.595 171.420 94.915 171.480 ;
        RECT 92.770 171.280 94.915 171.420 ;
        RECT 92.770 171.235 93.060 171.280 ;
        RECT 94.595 171.220 94.915 171.280 ;
        RECT 95.070 171.235 95.360 171.465 ;
        RECT 74.835 171.080 75.125 171.125 ;
        RECT 76.695 171.080 76.985 171.125 ;
        RECT 74.835 170.940 76.985 171.080 ;
        RECT 74.835 170.895 75.125 170.940 ;
        RECT 76.695 170.895 76.985 170.940 ;
        RECT 77.615 171.080 77.905 171.125 ;
        RECT 80.875 171.080 81.165 171.125 ;
        RECT 86.775 171.080 87.095 171.140 ;
        RECT 77.615 170.940 87.095 171.080 ;
        RECT 77.615 170.895 77.905 170.940 ;
        RECT 80.875 170.895 81.165 170.940 ;
        RECT 75.750 170.740 76.040 170.785 ;
        RECT 73.065 170.600 76.040 170.740 ;
        RECT 76.770 170.740 76.985 170.895 ;
        RECT 86.775 170.880 87.095 170.940 ;
        RECT 90.930 171.080 91.220 171.125 ;
        RECT 93.230 171.080 93.520 171.125 ;
        RECT 90.930 170.940 93.520 171.080 ;
        RECT 95.145 171.080 95.285 171.235 ;
        RECT 95.515 171.220 95.835 171.480 ;
        RECT 96.895 171.220 97.215 171.480 ;
        RECT 103.795 171.420 104.115 171.480 ;
        RECT 104.270 171.420 104.560 171.465 ;
        RECT 103.795 171.280 104.560 171.420 ;
        RECT 103.795 171.220 104.115 171.280 ;
        RECT 104.270 171.235 104.560 171.280 ;
        RECT 104.730 171.420 105.020 171.465 ;
        RECT 105.635 171.420 105.955 171.480 ;
        RECT 104.730 171.280 105.955 171.420 ;
        RECT 104.730 171.235 105.020 171.280 ;
        RECT 105.635 171.220 105.955 171.280 ;
        RECT 101.495 171.080 101.815 171.140 ;
        RECT 101.970 171.080 102.260 171.125 ;
        RECT 106.570 171.080 106.860 171.125 ;
        RECT 95.145 170.940 98.045 171.080 ;
        RECT 90.930 170.895 91.220 170.940 ;
        RECT 93.230 170.895 93.520 170.940 ;
        RECT 79.015 170.740 79.305 170.785 ;
        RECT 76.770 170.600 79.305 170.740 ;
        RECT 75.750 170.555 76.040 170.600 ;
        RECT 79.015 170.555 79.305 170.600 ;
        RECT 81.715 170.740 82.035 170.800 ;
        RECT 84.950 170.740 85.240 170.785 ;
        RECT 81.715 170.600 85.240 170.740 ;
        RECT 81.715 170.540 82.035 170.600 ;
        RECT 84.950 170.555 85.240 170.600 ;
        RECT 85.395 170.540 85.715 170.800 ;
        RECT 89.535 170.740 89.855 170.800 ;
        RECT 97.905 170.785 98.045 170.940 ;
        RECT 101.495 170.940 106.860 171.080 ;
        RECT 101.495 170.880 101.815 170.940 ;
        RECT 101.970 170.895 102.260 170.940 ;
        RECT 106.570 170.895 106.860 170.940 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 96.450 170.740 96.740 170.785 ;
        RECT 89.535 170.600 96.740 170.740 ;
        RECT 89.535 170.540 89.855 170.600 ;
        RECT 96.450 170.555 96.740 170.600 ;
        RECT 97.830 170.555 98.120 170.785 ;
        RECT 102.430 170.740 102.720 170.785 ;
        RECT 98.365 170.600 102.720 170.740 ;
        RECT 61.030 170.400 61.320 170.445 ;
        RECT 61.935 170.400 62.255 170.460 ;
        RECT 68.375 170.400 68.695 170.460 ;
        RECT 69.770 170.400 70.060 170.445 ;
        RECT 61.030 170.260 70.060 170.400 ;
        RECT 61.030 170.215 61.320 170.260 ;
        RECT 61.935 170.200 62.255 170.260 ;
        RECT 49.515 170.060 49.835 170.120 ;
        RECT 58.255 170.060 58.575 170.120 ;
        RECT 64.325 170.105 64.465 170.260 ;
        RECT 68.375 170.200 68.695 170.260 ;
        RECT 69.770 170.215 70.060 170.260 ;
        RECT 73.910 170.400 74.200 170.445 ;
        RECT 82.635 170.400 82.955 170.460 ;
        RECT 73.910 170.260 82.955 170.400 ;
        RECT 73.910 170.215 74.200 170.260 ;
        RECT 82.635 170.200 82.955 170.260 ;
        RECT 84.015 170.200 84.335 170.460 ;
        RECT 87.710 170.215 88.000 170.445 ;
        RECT 89.995 170.400 90.315 170.460 ;
        RECT 91.850 170.400 92.140 170.445 ;
        RECT 89.995 170.260 92.140 170.400 ;
        RECT 44.545 169.920 58.575 170.060 ;
        RECT 34.810 169.875 35.100 169.920 ;
        RECT 36.635 169.860 36.955 169.920 ;
        RECT 49.515 169.860 49.835 169.920 ;
        RECT 58.255 169.860 58.575 169.920 ;
        RECT 64.250 169.875 64.540 170.105 ;
        RECT 64.695 170.060 65.015 170.120 ;
        RECT 67.455 170.060 67.775 170.120 ;
        RECT 64.695 169.920 67.775 170.060 ;
        RECT 64.695 169.860 65.015 169.920 ;
        RECT 67.455 169.860 67.775 169.920 ;
        RECT 67.915 169.860 68.235 170.120 ;
        RECT 74.375 170.060 74.665 170.105 ;
        RECT 76.235 170.060 76.525 170.105 ;
        RECT 79.015 170.060 79.305 170.105 ;
        RECT 74.375 169.920 79.305 170.060 ;
        RECT 74.375 169.875 74.665 169.920 ;
        RECT 76.235 169.875 76.525 169.920 ;
        RECT 79.015 169.875 79.305 169.920 ;
        RECT 81.255 170.060 81.575 170.120 ;
        RECT 87.785 170.060 87.925 170.215 ;
        RECT 89.995 170.200 90.315 170.260 ;
        RECT 91.850 170.215 92.140 170.260 ;
        RECT 94.595 170.400 94.915 170.460 ;
        RECT 98.365 170.400 98.505 170.600 ;
        RECT 102.430 170.555 102.720 170.600 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 94.595 170.260 98.505 170.400 ;
        RECT 91.375 170.060 91.695 170.120 ;
        RECT 81.255 169.920 91.695 170.060 ;
        RECT 91.925 170.060 92.065 170.215 ;
        RECT 94.595 170.200 94.915 170.260 ;
        RECT 101.050 170.215 101.340 170.445 ;
        RECT 102.875 170.400 103.195 170.460 ;
        RECT 107.030 170.400 107.320 170.445 ;
        RECT 102.875 170.260 107.320 170.400 ;
        RECT 101.125 170.060 101.265 170.215 ;
        RECT 102.875 170.200 103.195 170.260 ;
        RECT 107.030 170.215 107.320 170.260 ;
        RECT 107.490 170.215 107.780 170.445 ;
        RECT 101.955 170.060 102.275 170.120 ;
        RECT 107.565 170.060 107.705 170.215 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 91.925 169.920 107.705 170.060 ;
        RECT 81.255 169.860 81.575 169.920 ;
        RECT 91.375 169.860 91.695 169.920 ;
        RECT 101.955 169.860 102.275 169.920 ;
        RECT 35.270 169.720 35.560 169.765 ;
        RECT 36.175 169.720 36.495 169.780 ;
        RECT 35.270 169.580 36.495 169.720 ;
        RECT 35.270 169.535 35.560 169.580 ;
        RECT 36.175 169.520 36.495 169.580 ;
        RECT 43.090 169.720 43.380 169.765 ;
        RECT 44.455 169.720 44.775 169.780 ;
        RECT 43.090 169.580 44.775 169.720 ;
        RECT 43.090 169.535 43.380 169.580 ;
        RECT 44.455 169.520 44.775 169.580 ;
        RECT 45.835 169.720 46.155 169.780 ;
        RECT 48.150 169.720 48.440 169.765 ;
        RECT 45.835 169.580 48.440 169.720 ;
        RECT 45.835 169.520 46.155 169.580 ;
        RECT 48.150 169.535 48.440 169.580 ;
        RECT 57.795 169.720 58.115 169.780 ;
        RECT 59.190 169.720 59.480 169.765 ;
        RECT 57.795 169.580 59.480 169.720 ;
        RECT 57.795 169.520 58.115 169.580 ;
        RECT 59.190 169.535 59.480 169.580 ;
        RECT 66.995 169.720 67.315 169.780 ;
        RECT 71.150 169.720 71.440 169.765 ;
        RECT 66.995 169.580 71.440 169.720 ;
        RECT 66.995 169.520 67.315 169.580 ;
        RECT 71.150 169.535 71.440 169.580 ;
        RECT 82.175 169.720 82.495 169.780 ;
        RECT 82.880 169.720 83.170 169.765 ;
        RECT 82.175 169.580 83.170 169.720 ;
        RECT 82.175 169.520 82.495 169.580 ;
        RECT 82.880 169.535 83.170 169.580 ;
        RECT 87.235 169.720 87.555 169.780 ;
        RECT 101.495 169.720 101.815 169.780 ;
        RECT 87.235 169.580 101.815 169.720 ;
        RECT 87.235 169.520 87.555 169.580 ;
        RECT 101.495 169.520 101.815 169.580 ;
        RECT 18.165 168.900 112.465 169.380 ;
        RECT 23.310 168.700 23.600 168.745 ;
        RECT 23.755 168.700 24.075 168.760 ;
        RECT 23.310 168.560 24.075 168.700 ;
        RECT 23.310 168.515 23.600 168.560 ;
        RECT 23.755 168.500 24.075 168.560 ;
        RECT 32.035 168.700 32.355 168.760 ;
        RECT 48.595 168.700 48.915 168.760 ;
        RECT 32.035 168.560 48.915 168.700 ;
        RECT 32.035 168.500 32.355 168.560 ;
        RECT 48.595 168.500 48.915 168.560 ;
        RECT 58.270 168.700 58.560 168.745 ;
        RECT 59.175 168.700 59.495 168.760 ;
        RECT 58.270 168.560 59.495 168.700 ;
        RECT 58.270 168.515 58.560 168.560 ;
        RECT 32.125 168.360 32.265 168.500 ;
        RECT 34.335 168.360 34.655 168.420 ;
        RECT 27.065 168.220 32.265 168.360 ;
        RECT 33.045 168.220 34.655 168.360 ;
        RECT 27.065 168.065 27.205 168.220 ;
        RECT 26.990 167.835 27.280 168.065 ;
        RECT 27.435 167.820 27.755 168.080 ;
        RECT 27.895 168.020 28.215 168.080 ;
        RECT 33.045 168.020 33.185 168.220 ;
        RECT 34.335 168.160 34.655 168.220 ;
        RECT 37.095 168.360 37.415 168.420 ;
        RECT 37.095 168.220 41.005 168.360 ;
        RECT 37.095 168.160 37.415 168.220 ;
        RECT 27.895 167.880 33.185 168.020 ;
        RECT 27.895 167.820 28.215 167.880 ;
        RECT 21.915 167.480 22.235 167.740 ;
        RECT 24.230 167.680 24.520 167.725 ;
        RECT 24.230 167.540 24.905 167.680 ;
        RECT 24.230 167.495 24.520 167.540 ;
        RECT 22.390 167.000 22.680 167.045 ;
        RECT 22.835 167.000 23.155 167.060 ;
        RECT 24.765 167.045 24.905 167.540 ;
        RECT 28.815 167.480 29.135 167.740 ;
        RECT 31.115 167.480 31.435 167.740 ;
        RECT 31.575 167.680 31.895 167.740 ;
        RECT 32.050 167.680 32.340 167.725 ;
        RECT 31.575 167.540 32.340 167.680 ;
        RECT 31.575 167.480 31.895 167.540 ;
        RECT 32.050 167.495 32.340 167.540 ;
        RECT 32.495 167.480 32.815 167.740 ;
        RECT 33.045 167.725 33.185 167.880 ;
        RECT 33.875 168.020 34.195 168.080 ;
        RECT 33.875 167.880 37.785 168.020 ;
        RECT 33.875 167.820 34.195 167.880 ;
        RECT 32.970 167.680 33.260 167.725 ;
        RECT 36.550 167.680 36.840 167.725 ;
        RECT 32.970 167.660 35.945 167.680 ;
        RECT 36.495 167.660 36.840 167.680 ;
        RECT 32.970 167.540 36.840 167.660 ;
        RECT 32.970 167.495 33.260 167.540 ;
        RECT 35.805 167.520 36.840 167.540 ;
        RECT 36.550 167.495 36.840 167.520 ;
        RECT 37.095 167.480 37.415 167.740 ;
        RECT 37.645 167.725 37.785 167.880 ;
        RECT 38.335 167.880 40.545 168.020 ;
        RECT 38.335 167.725 38.475 167.880 ;
        RECT 40.405 167.740 40.545 167.880 ;
        RECT 37.570 167.495 37.860 167.725 ;
        RECT 38.335 167.540 38.660 167.725 ;
        RECT 38.370 167.495 38.660 167.540 ;
        RECT 38.950 167.495 39.240 167.725 ;
        RECT 25.595 167.340 25.915 167.400 ;
        RECT 31.205 167.340 31.345 167.480 ;
        RECT 25.595 167.200 31.345 167.340 ;
        RECT 34.350 167.340 34.640 167.385 ;
        RECT 34.795 167.340 35.115 167.400 ;
        RECT 34.350 167.200 35.115 167.340 ;
        RECT 25.595 167.140 25.915 167.200 ;
        RECT 34.350 167.155 34.640 167.200 ;
        RECT 34.795 167.140 35.115 167.200 ;
        RECT 39.025 167.340 39.165 167.495 ;
        RECT 40.315 167.480 40.635 167.740 ;
        RECT 40.865 167.680 41.005 168.220 ;
        RECT 45.005 168.220 49.285 168.360 ;
        RECT 45.005 168.080 45.145 168.220 ;
        RECT 44.915 168.020 45.235 168.080 ;
        RECT 41.785 167.880 45.235 168.020 ;
        RECT 41.785 167.725 41.925 167.880 ;
        RECT 44.915 167.820 45.235 167.880 ;
        RECT 49.145 168.020 49.285 168.220 ;
        RECT 56.430 168.175 56.720 168.405 ;
        RECT 49.975 168.020 50.295 168.080 ;
        RECT 56.505 168.020 56.645 168.175 ;
        RECT 58.345 168.020 58.485 168.515 ;
        RECT 59.175 168.500 59.495 168.560 ;
        RECT 59.635 168.500 59.955 168.760 ;
        RECT 65.630 168.700 65.920 168.745 ;
        RECT 66.995 168.700 67.315 168.760 ;
        RECT 84.950 168.700 85.240 168.745 ;
        RECT 89.535 168.700 89.855 168.760 ;
        RECT 63.405 168.560 65.385 168.700 ;
        RECT 61.475 168.360 61.795 168.420 ;
        RECT 63.405 168.360 63.545 168.560 ;
        RECT 64.695 168.360 65.015 168.420 ;
        RECT 59.725 168.220 63.545 168.360 ;
        RECT 63.865 168.220 65.015 168.360 ;
        RECT 65.245 168.360 65.385 168.560 ;
        RECT 65.630 168.560 67.315 168.700 ;
        RECT 65.630 168.515 65.920 168.560 ;
        RECT 66.995 168.500 67.315 168.560 ;
        RECT 79.965 168.560 84.705 168.700 ;
        RECT 65.245 168.220 67.225 168.360 ;
        RECT 59.725 168.065 59.865 168.220 ;
        RECT 61.475 168.160 61.795 168.220 ;
        RECT 49.145 167.880 56.645 168.020 ;
        RECT 41.250 167.680 41.540 167.725 ;
        RECT 40.865 167.540 41.540 167.680 ;
        RECT 41.250 167.495 41.540 167.540 ;
        RECT 41.710 167.495 42.000 167.725 ;
        RECT 42.155 167.480 42.475 167.740 ;
        RECT 47.230 167.495 47.520 167.725 ;
        RECT 46.755 167.340 47.075 167.400 ;
        RECT 39.025 167.200 47.075 167.340 ;
        RECT 22.390 166.860 23.155 167.000 ;
        RECT 22.390 166.815 22.680 166.860 ;
        RECT 22.835 166.800 23.155 166.860 ;
        RECT 24.690 166.815 24.980 167.045 ;
        RECT 26.530 167.000 26.820 167.045 ;
        RECT 27.435 167.000 27.755 167.060 ;
        RECT 26.530 166.860 27.755 167.000 ;
        RECT 26.530 166.815 26.820 166.860 ;
        RECT 27.435 166.800 27.755 166.860 ;
        RECT 29.735 166.800 30.055 167.060 ;
        RECT 32.955 167.000 33.275 167.060 ;
        RECT 35.270 167.000 35.560 167.045 ;
        RECT 32.955 166.860 35.560 167.000 ;
        RECT 32.955 166.800 33.275 166.860 ;
        RECT 35.270 166.815 35.560 166.860 ;
        RECT 35.715 167.000 36.035 167.060 ;
        RECT 39.025 167.000 39.165 167.200 ;
        RECT 46.755 167.140 47.075 167.200 ;
        RECT 35.715 166.860 39.165 167.000 ;
        RECT 35.715 166.800 36.035 166.860 ;
        RECT 39.395 166.800 39.715 167.060 ;
        RECT 43.535 166.800 43.855 167.060 ;
        RECT 44.010 167.000 44.300 167.045 ;
        RECT 45.375 167.000 45.695 167.060 ;
        RECT 44.010 166.860 45.695 167.000 ;
        RECT 47.305 167.000 47.445 167.495 ;
        RECT 47.675 167.480 47.995 167.740 ;
        RECT 48.135 167.680 48.455 167.740 ;
        RECT 49.145 167.725 49.285 167.880 ;
        RECT 49.975 167.820 50.295 167.880 ;
        RECT 48.610 167.680 48.900 167.725 ;
        RECT 48.135 167.540 48.900 167.680 ;
        RECT 48.135 167.480 48.455 167.540 ;
        RECT 48.610 167.495 48.900 167.540 ;
        RECT 49.070 167.495 49.360 167.725 ;
        RECT 49.515 167.480 49.835 167.740 ;
        RECT 56.505 167.680 56.645 167.880 ;
        RECT 57.425 167.880 58.485 168.020 ;
        RECT 57.425 167.725 57.565 167.880 ;
        RECT 59.650 167.835 59.940 168.065 ;
        RECT 61.935 168.020 62.255 168.080 ;
        RECT 62.410 168.020 62.700 168.065 ;
        RECT 61.935 167.880 62.700 168.020 ;
        RECT 61.935 167.820 62.255 167.880 ;
        RECT 62.410 167.835 62.700 167.880 ;
        RECT 62.855 167.820 63.175 168.080 ;
        RECT 63.865 168.065 64.005 168.220 ;
        RECT 64.695 168.160 65.015 168.220 ;
        RECT 63.790 167.835 64.080 168.065 ;
        RECT 64.235 168.020 64.555 168.080 ;
        RECT 66.075 168.020 66.395 168.080 ;
        RECT 67.085 168.065 67.225 168.220 ;
        RECT 66.550 168.020 66.840 168.065 ;
        RECT 64.235 167.880 65.845 168.020 ;
        RECT 64.235 167.820 64.555 167.880 ;
        RECT 56.505 167.540 57.105 167.680 ;
        RECT 50.435 167.000 50.755 167.060 ;
        RECT 47.305 166.860 50.755 167.000 ;
        RECT 44.010 166.815 44.300 166.860 ;
        RECT 45.375 166.800 45.695 166.860 ;
        RECT 50.435 166.800 50.755 166.860 ;
        RECT 50.910 167.000 51.200 167.045 ;
        RECT 51.815 167.000 52.135 167.060 ;
        RECT 50.910 166.860 52.135 167.000 ;
        RECT 56.965 167.000 57.105 167.540 ;
        RECT 57.350 167.495 57.640 167.725 ;
        RECT 57.795 167.480 58.115 167.740 ;
        RECT 59.175 167.480 59.495 167.740 ;
        RECT 61.015 167.680 61.335 167.740 ;
        RECT 63.330 167.680 63.620 167.725 ;
        RECT 61.015 167.540 63.620 167.680 ;
        RECT 61.015 167.480 61.335 167.540 ;
        RECT 63.330 167.495 63.620 167.540 ;
        RECT 64.695 167.680 65.015 167.740 ;
        RECT 65.170 167.680 65.460 167.725 ;
        RECT 64.695 167.540 65.460 167.680 ;
        RECT 65.705 167.680 65.845 167.880 ;
        RECT 66.075 167.880 66.840 168.020 ;
        RECT 66.075 167.820 66.395 167.880 ;
        RECT 66.550 167.835 66.840 167.880 ;
        RECT 67.010 168.020 67.300 168.065 ;
        RECT 68.390 168.020 68.680 168.065 ;
        RECT 67.010 167.880 68.680 168.020 ;
        RECT 67.010 167.835 67.300 167.880 ;
        RECT 68.390 167.835 68.680 167.880 ;
        RECT 67.930 167.680 68.220 167.725 ;
        RECT 65.705 167.540 68.220 167.680 ;
        RECT 64.695 167.480 65.015 167.540 ;
        RECT 65.170 167.495 65.460 167.540 ;
        RECT 67.930 167.495 68.220 167.540 ;
        RECT 79.965 167.340 80.105 168.560 ;
        RECT 81.255 168.360 81.575 168.420 ;
        RECT 84.565 168.360 84.705 168.560 ;
        RECT 84.950 168.560 89.855 168.700 ;
        RECT 84.950 168.515 85.240 168.560 ;
        RECT 89.535 168.500 89.855 168.560 ;
        RECT 89.075 168.360 89.395 168.420 ;
        RECT 81.255 168.220 82.865 168.360 ;
        RECT 84.565 168.220 89.395 168.360 ;
        RECT 81.255 168.160 81.575 168.220 ;
        RECT 80.795 168.020 81.115 168.080 ;
        RECT 82.725 168.065 82.865 168.220 ;
        RECT 81.730 168.020 82.020 168.065 ;
        RECT 80.795 167.880 82.020 168.020 ;
        RECT 80.795 167.820 81.115 167.880 ;
        RECT 81.730 167.835 82.020 167.880 ;
        RECT 82.650 167.835 82.940 168.065 ;
        RECT 80.350 167.495 80.640 167.725 ;
        RECT 62.485 167.200 80.105 167.340 ;
        RECT 80.425 167.340 80.565 167.495 ;
        RECT 86.775 167.480 87.095 167.740 ;
        RECT 87.235 167.680 87.555 167.740 ;
        RECT 88.245 167.725 88.385 168.220 ;
        RECT 89.075 168.160 89.395 168.220 ;
        RECT 101.955 167.820 102.275 168.080 ;
        RECT 87.710 167.680 88.000 167.725 ;
        RECT 87.235 167.540 88.000 167.680 ;
        RECT 87.235 167.480 87.555 167.540 ;
        RECT 87.710 167.495 88.000 167.540 ;
        RECT 88.185 167.495 88.475 167.725 ;
        RECT 88.630 167.570 88.920 167.725 ;
        RECT 90.470 167.680 90.760 167.725 ;
        RECT 90.915 167.680 91.235 167.740 ;
        RECT 88.630 167.495 89.305 167.570 ;
        RECT 90.470 167.540 91.235 167.680 ;
        RECT 90.470 167.495 90.760 167.540 ;
        RECT 88.705 167.430 89.305 167.495 ;
        RECT 90.915 167.480 91.235 167.540 ;
        RECT 91.375 167.480 91.695 167.740 ;
        RECT 91.850 167.495 92.140 167.725 ;
        RECT 82.635 167.340 82.955 167.400 ;
        RECT 80.425 167.200 82.955 167.340 ;
        RECT 62.485 167.000 62.625 167.200 ;
        RECT 82.635 167.140 82.955 167.200 ;
        RECT 56.965 166.860 62.625 167.000 ;
        RECT 62.855 167.000 63.175 167.060 ;
        RECT 66.535 167.000 66.855 167.060 ;
        RECT 67.010 167.000 67.300 167.045 ;
        RECT 62.855 166.860 67.300 167.000 ;
        RECT 50.910 166.815 51.200 166.860 ;
        RECT 51.815 166.800 52.135 166.860 ;
        RECT 62.855 166.800 63.175 166.860 ;
        RECT 66.535 166.800 66.855 166.860 ;
        RECT 67.010 166.815 67.300 166.860 ;
        RECT 82.175 167.000 82.495 167.060 ;
        RECT 83.110 167.000 83.400 167.045 ;
        RECT 82.175 166.860 83.400 167.000 ;
        RECT 82.175 166.800 82.495 166.860 ;
        RECT 83.110 166.815 83.400 166.860 ;
        RECT 87.235 167.000 87.555 167.060 ;
        RECT 89.165 167.000 89.305 167.430 ;
        RECT 89.535 167.340 89.855 167.400 ;
        RECT 91.925 167.340 92.065 167.495 ;
        RECT 92.295 167.480 92.615 167.740 ;
        RECT 92.755 167.680 93.075 167.740 ;
        RECT 94.150 167.680 94.440 167.725 ;
        RECT 92.755 167.540 94.440 167.680 ;
        RECT 92.755 167.480 93.075 167.540 ;
        RECT 94.150 167.495 94.440 167.540 ;
        RECT 94.595 167.680 94.915 167.740 ;
        RECT 95.070 167.680 95.360 167.725 ;
        RECT 94.595 167.540 95.360 167.680 ;
        RECT 94.595 167.480 94.915 167.540 ;
        RECT 95.070 167.495 95.360 167.540 ;
        RECT 95.530 167.495 95.820 167.725 ;
        RECT 95.990 167.495 96.280 167.725 ;
        RECT 105.650 167.680 105.940 167.725 ;
        RECT 104.805 167.540 105.940 167.680 ;
        RECT 95.605 167.340 95.745 167.495 ;
        RECT 89.535 167.200 95.745 167.340 ;
        RECT 89.535 167.140 89.855 167.200 ;
        RECT 95.145 167.060 95.285 167.200 ;
        RECT 87.235 166.860 89.305 167.000 ;
        RECT 90.010 167.000 90.300 167.045 ;
        RECT 92.295 167.000 92.615 167.060 ;
        RECT 90.010 166.860 92.615 167.000 ;
        RECT 87.235 166.800 87.555 166.860 ;
        RECT 90.010 166.815 90.300 166.860 ;
        RECT 92.295 166.800 92.615 166.860 ;
        RECT 92.755 167.000 93.075 167.060 ;
        RECT 93.690 167.000 93.980 167.045 ;
        RECT 92.755 166.860 93.980 167.000 ;
        RECT 92.755 166.800 93.075 166.860 ;
        RECT 93.690 166.815 93.980 166.860 ;
        RECT 95.055 166.800 95.375 167.060 ;
        RECT 95.515 167.000 95.835 167.060 ;
        RECT 96.065 167.000 96.205 167.495 ;
        RECT 95.515 166.860 96.205 167.000 ;
        RECT 96.895 167.000 97.215 167.060 ;
        RECT 97.370 167.000 97.660 167.045 ;
        RECT 96.895 166.860 97.660 167.000 ;
        RECT 95.515 166.800 95.835 166.860 ;
        RECT 96.895 166.800 97.215 166.860 ;
        RECT 97.370 166.815 97.660 166.860 ;
        RECT 101.955 167.000 102.275 167.060 ;
        RECT 102.430 167.000 102.720 167.045 ;
        RECT 101.955 166.860 102.720 167.000 ;
        RECT 101.955 166.800 102.275 166.860 ;
        RECT 102.430 166.815 102.720 166.860 ;
        RECT 102.875 166.800 103.195 167.060 ;
        RECT 104.805 167.045 104.945 167.540 ;
        RECT 105.650 167.495 105.940 167.540 ;
        RECT 104.730 166.815 105.020 167.045 ;
        RECT 106.570 167.000 106.860 167.045 ;
        RECT 107.475 167.000 107.795 167.060 ;
        RECT 106.570 166.860 107.795 167.000 ;
        RECT 106.570 166.815 106.860 166.860 ;
        RECT 107.475 166.800 107.795 166.860 ;
        RECT 17.370 166.180 112.465 166.660 ;
        RECT 24.675 165.980 24.995 166.040 ;
        RECT 32.495 165.980 32.815 166.040 ;
        RECT 24.675 165.840 32.815 165.980 ;
        RECT 24.675 165.780 24.995 165.840 ;
        RECT 32.495 165.780 32.815 165.840 ;
        RECT 34.350 165.980 34.640 166.025 ;
        RECT 35.255 165.980 35.575 166.040 ;
        RECT 48.150 165.980 48.440 166.025 ;
        RECT 34.350 165.840 35.575 165.980 ;
        RECT 34.350 165.795 34.640 165.840 ;
        RECT 35.255 165.780 35.575 165.840 ;
        RECT 46.385 165.840 48.440 165.980 ;
        RECT 22.835 165.640 23.155 165.700 ;
        RECT 23.870 165.640 24.160 165.685 ;
        RECT 27.110 165.640 27.760 165.685 ;
        RECT 22.835 165.500 27.760 165.640 ;
        RECT 22.835 165.440 23.155 165.500 ;
        RECT 23.870 165.455 24.460 165.500 ;
        RECT 27.110 165.455 27.760 165.500 ;
        RECT 24.170 165.140 24.460 165.455 ;
        RECT 29.735 165.440 30.055 165.700 ;
        RECT 39.395 165.685 39.715 165.700 ;
        RECT 34.810 165.455 35.100 165.685 ;
        RECT 39.345 165.640 39.715 165.685 ;
        RECT 42.605 165.640 42.895 165.685 ;
        RECT 39.345 165.500 42.895 165.640 ;
        RECT 39.345 165.455 39.715 165.500 ;
        RECT 42.605 165.455 42.895 165.500 ;
        RECT 43.525 165.640 43.815 165.685 ;
        RECT 45.385 165.640 45.675 165.685 ;
        RECT 43.525 165.500 45.675 165.640 ;
        RECT 43.525 165.455 43.815 165.500 ;
        RECT 45.385 165.455 45.675 165.500 ;
        RECT 25.250 165.300 25.540 165.345 ;
        RECT 28.830 165.300 29.120 165.345 ;
        RECT 30.665 165.300 30.955 165.345 ;
        RECT 25.250 165.160 30.955 165.300 ;
        RECT 25.250 165.115 25.540 165.160 ;
        RECT 28.830 165.115 29.120 165.160 ;
        RECT 30.665 165.115 30.955 165.160 ;
        RECT 31.130 165.300 31.420 165.345 ;
        RECT 32.495 165.300 32.815 165.360 ;
        RECT 31.130 165.160 32.815 165.300 ;
        RECT 31.130 165.115 31.420 165.160 ;
        RECT 32.495 165.100 32.815 165.160 ;
        RECT 32.035 164.960 32.355 165.020 ;
        RECT 33.430 164.960 33.720 165.005 ;
        RECT 32.035 164.820 33.720 164.960 ;
        RECT 32.035 164.760 32.355 164.820 ;
        RECT 33.430 164.775 33.720 164.820 ;
        RECT 25.250 164.620 25.540 164.665 ;
        RECT 28.370 164.620 28.660 164.665 ;
        RECT 30.260 164.620 30.550 164.665 ;
        RECT 25.250 164.480 30.550 164.620 ;
        RECT 34.885 164.620 35.025 165.455 ;
        RECT 39.395 165.440 39.715 165.455 ;
        RECT 41.205 165.300 41.495 165.345 ;
        RECT 43.525 165.300 43.740 165.455 ;
        RECT 41.205 165.160 43.740 165.300 ;
        RECT 44.470 165.300 44.760 165.345 ;
        RECT 46.385 165.300 46.525 165.840 ;
        RECT 48.150 165.795 48.440 165.840 ;
        RECT 48.595 165.980 48.915 166.040 ;
        RECT 50.435 165.980 50.755 166.040 ;
        RECT 52.750 165.980 53.040 166.025 ;
        RECT 48.595 165.840 53.040 165.980 ;
        RECT 48.595 165.780 48.915 165.840 ;
        RECT 50.435 165.780 50.755 165.840 ;
        RECT 52.750 165.795 53.040 165.840 ;
        RECT 56.890 165.980 57.180 166.025 ;
        RECT 57.335 165.980 57.655 166.040 ;
        RECT 56.890 165.840 57.655 165.980 ;
        RECT 56.890 165.795 57.180 165.840 ;
        RECT 57.335 165.780 57.655 165.840 ;
        RECT 58.255 165.980 58.575 166.040 ;
        RECT 71.595 165.980 71.915 166.040 ;
        RECT 58.255 165.840 71.915 165.980 ;
        RECT 58.255 165.780 58.575 165.840 ;
        RECT 71.595 165.780 71.915 165.840 ;
        RECT 72.055 165.980 72.375 166.040 ;
        RECT 72.990 165.980 73.280 166.025 ;
        RECT 102.875 165.980 103.195 166.040 ;
        RECT 72.055 165.840 73.280 165.980 ;
        RECT 72.055 165.780 72.375 165.840 ;
        RECT 72.990 165.795 73.280 165.840 ;
        RECT 96.985 165.840 103.195 165.980 ;
        RECT 46.755 165.640 47.075 165.700 ;
        RECT 56.415 165.640 56.735 165.700 ;
        RECT 46.755 165.500 56.735 165.640 ;
        RECT 46.755 165.440 47.075 165.500 ;
        RECT 44.470 165.160 46.525 165.300 ;
        RECT 41.205 165.115 41.495 165.160 ;
        RECT 44.470 165.115 44.760 165.160 ;
        RECT 49.055 165.100 49.375 165.360 ;
        RECT 49.605 165.345 49.745 165.500 ;
        RECT 56.415 165.440 56.735 165.500 ;
        RECT 49.530 165.115 49.820 165.345 ;
        RECT 50.895 165.300 51.215 165.360 ;
        RECT 52.290 165.300 52.580 165.345 ;
        RECT 50.895 165.160 52.580 165.300 ;
        RECT 50.895 165.100 51.215 165.160 ;
        RECT 52.290 165.115 52.580 165.160 ;
        RECT 55.970 165.300 56.260 165.345 ;
        RECT 56.875 165.300 57.195 165.360 ;
        RECT 57.425 165.345 57.565 165.780 ;
        RECT 62.855 165.440 63.175 165.700 ;
        RECT 70.690 165.640 70.980 165.685 ;
        RECT 66.625 165.500 70.980 165.640 ;
        RECT 55.970 165.160 57.195 165.300 ;
        RECT 55.970 165.115 56.260 165.160 ;
        RECT 56.875 165.100 57.195 165.160 ;
        RECT 57.350 165.115 57.640 165.345 ;
        RECT 59.190 165.300 59.480 165.345 ;
        RECT 60.095 165.300 60.415 165.360 ;
        RECT 59.190 165.160 60.415 165.300 ;
        RECT 59.190 165.115 59.480 165.160 ;
        RECT 60.095 165.100 60.415 165.160 ;
        RECT 63.775 165.300 64.095 165.360 ;
        RECT 64.710 165.300 65.000 165.345 ;
        RECT 63.775 165.160 65.000 165.300 ;
        RECT 63.775 165.100 64.095 165.160 ;
        RECT 64.710 165.115 65.000 165.160 ;
        RECT 65.615 165.100 65.935 165.360 ;
        RECT 66.625 165.345 66.765 165.500 ;
        RECT 70.690 165.455 70.980 165.500 ;
        RECT 71.150 165.640 71.440 165.685 ;
        RECT 74.355 165.640 74.675 165.700 ;
        RECT 85.855 165.685 86.175 165.700 ;
        RECT 71.150 165.500 74.675 165.640 ;
        RECT 71.150 165.455 71.440 165.500 ;
        RECT 66.550 165.115 66.840 165.345 ;
        RECT 67.010 165.115 67.300 165.345 ;
        RECT 67.470 165.115 67.760 165.345 ;
        RECT 38.935 164.960 39.255 165.020 ;
        RECT 46.310 164.960 46.600 165.005 ;
        RECT 38.935 164.820 46.600 164.960 ;
        RECT 38.935 164.760 39.255 164.820 ;
        RECT 46.310 164.775 46.600 164.820 ;
        RECT 51.830 164.960 52.120 165.005 ;
        RECT 61.490 164.960 61.780 165.005 ;
        RECT 51.830 164.820 61.780 164.960 ;
        RECT 51.830 164.775 52.120 164.820 ;
        RECT 61.490 164.775 61.780 164.820 ;
        RECT 66.075 164.960 66.395 165.020 ;
        RECT 67.085 164.960 67.225 165.115 ;
        RECT 66.075 164.820 67.225 164.960 ;
        RECT 67.545 164.960 67.685 165.115 ;
        RECT 69.755 164.960 70.075 165.020 ;
        RECT 67.545 164.820 70.075 164.960 ;
        RECT 37.340 164.620 37.630 164.665 ;
        RECT 41.205 164.620 41.495 164.665 ;
        RECT 43.985 164.620 44.275 164.665 ;
        RECT 45.845 164.620 46.135 164.665 ;
        RECT 34.885 164.480 41.005 164.620 ;
        RECT 25.250 164.435 25.540 164.480 ;
        RECT 28.370 164.435 28.660 164.480 ;
        RECT 30.260 164.435 30.550 164.480 ;
        RECT 37.340 164.435 37.630 164.480 ;
        RECT 22.390 164.280 22.680 164.325 ;
        RECT 27.435 164.280 27.755 164.340 ;
        RECT 22.390 164.140 27.755 164.280 ;
        RECT 22.390 164.095 22.680 164.140 ;
        RECT 27.435 164.080 27.755 164.140 ;
        RECT 36.650 164.280 36.940 164.325 ;
        RECT 39.395 164.280 39.715 164.340 ;
        RECT 36.650 164.140 39.715 164.280 ;
        RECT 40.865 164.280 41.005 164.480 ;
        RECT 41.205 164.480 46.135 164.620 ;
        RECT 41.205 164.435 41.495 164.480 ;
        RECT 43.985 164.435 44.275 164.480 ;
        RECT 45.845 164.435 46.135 164.480 ;
        RECT 47.215 164.620 47.535 164.680 ;
        RECT 51.905 164.620 52.045 164.775 ;
        RECT 66.075 164.760 66.395 164.820 ;
        RECT 47.215 164.480 52.045 164.620 ;
        RECT 52.275 164.620 52.595 164.680 ;
        RECT 58.270 164.620 58.560 164.665 ;
        RECT 67.545 164.620 67.685 164.820 ;
        RECT 69.755 164.760 70.075 164.820 ;
        RECT 70.215 164.760 70.535 165.020 ;
        RECT 70.765 164.960 70.905 165.455 ;
        RECT 74.355 165.440 74.675 165.500 ;
        RECT 85.805 165.640 86.175 165.685 ;
        RECT 89.065 165.640 89.355 165.685 ;
        RECT 85.805 165.500 89.355 165.640 ;
        RECT 85.805 165.455 86.175 165.500 ;
        RECT 89.065 165.455 89.355 165.500 ;
        RECT 89.985 165.640 90.275 165.685 ;
        RECT 91.845 165.640 92.135 165.685 ;
        RECT 89.985 165.500 92.135 165.640 ;
        RECT 89.985 165.455 90.275 165.500 ;
        RECT 91.845 165.455 92.135 165.500 ;
        RECT 95.055 165.640 95.375 165.700 ;
        RECT 95.055 165.500 96.665 165.640 ;
        RECT 85.855 165.440 86.175 165.455 ;
        RECT 73.895 165.100 74.215 165.360 ;
        RECT 87.665 165.300 87.955 165.345 ;
        RECT 89.985 165.300 90.200 165.455 ;
        RECT 95.055 165.440 95.375 165.500 ;
        RECT 96.525 165.360 96.665 165.500 ;
        RECT 87.665 165.160 90.200 165.300 ;
        RECT 87.665 165.115 87.955 165.160 ;
        RECT 90.915 165.100 91.235 165.360 ;
        RECT 91.375 165.300 91.695 165.360 ;
        RECT 95.515 165.300 95.835 165.360 ;
        RECT 95.990 165.300 96.280 165.345 ;
        RECT 91.375 165.160 96.280 165.300 ;
        RECT 91.375 165.100 91.695 165.160 ;
        RECT 95.515 165.100 95.835 165.160 ;
        RECT 95.990 165.115 96.280 165.160 ;
        RECT 96.435 165.100 96.755 165.360 ;
        RECT 96.985 165.345 97.125 165.840 ;
        RECT 102.875 165.780 103.195 165.840 ;
        RECT 98.735 165.640 99.055 165.700 ;
        RECT 101.610 165.640 101.900 165.685 ;
        RECT 104.850 165.640 105.500 165.685 ;
        RECT 98.735 165.500 105.500 165.640 ;
        RECT 98.735 165.440 99.055 165.500 ;
        RECT 101.610 165.455 102.200 165.500 ;
        RECT 104.850 165.455 105.500 165.500 ;
        RECT 96.910 165.115 97.200 165.345 ;
        RECT 97.355 165.300 97.675 165.360 ;
        RECT 97.830 165.300 98.120 165.345 ;
        RECT 97.355 165.160 98.120 165.300 ;
        RECT 97.355 165.100 97.675 165.160 ;
        RECT 97.830 165.115 98.120 165.160 ;
        RECT 101.910 165.140 102.200 165.455 ;
        RECT 107.475 165.440 107.795 165.700 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 102.990 165.300 103.280 165.345 ;
        RECT 106.570 165.300 106.860 165.345 ;
        RECT 108.405 165.300 108.695 165.345 ;
        RECT 102.990 165.160 108.695 165.300 ;
        RECT 102.990 165.115 103.280 165.160 ;
        RECT 106.570 165.115 106.860 165.160 ;
        RECT 108.405 165.115 108.695 165.160 ;
        RECT 108.855 165.100 109.175 165.360 ;
        RECT 82.175 164.960 82.495 165.020 ;
        RECT 70.765 164.820 82.495 164.960 ;
        RECT 82.175 164.760 82.495 164.820 ;
        RECT 82.635 164.960 82.955 165.020 ;
        RECT 92.770 164.960 93.060 165.005 ;
        RECT 82.635 164.820 93.060 164.960 ;
        RECT 82.635 164.760 82.955 164.820 ;
        RECT 92.770 164.775 93.060 164.820 ;
        RECT 52.275 164.480 67.685 164.620 ;
        RECT 71.595 164.620 71.915 164.680 ;
        RECT 87.665 164.620 87.955 164.665 ;
        RECT 90.445 164.620 90.735 164.665 ;
        RECT 92.305 164.620 92.595 164.665 ;
        RECT 71.595 164.480 87.465 164.620 ;
        RECT 47.215 164.420 47.535 164.480 ;
        RECT 52.275 164.420 52.595 164.480 ;
        RECT 58.270 164.435 58.560 164.480 ;
        RECT 71.595 164.420 71.915 164.480 ;
        RECT 87.325 164.340 87.465 164.480 ;
        RECT 87.665 164.480 92.595 164.620 ;
        RECT 87.665 164.435 87.955 164.480 ;
        RECT 90.445 164.435 90.735 164.480 ;
        RECT 92.305 164.435 92.595 164.480 ;
        RECT 102.990 164.620 103.280 164.665 ;
        RECT 106.110 164.620 106.400 164.665 ;
        RECT 108.000 164.620 108.290 164.665 ;
        RECT 102.990 164.480 108.290 164.620 ;
        RECT 102.990 164.435 103.280 164.480 ;
        RECT 106.110 164.435 106.400 164.480 ;
        RECT 108.000 164.435 108.290 164.480 ;
        RECT 44.915 164.280 45.235 164.340 ;
        RECT 40.865 164.140 45.235 164.280 ;
        RECT 36.650 164.095 36.940 164.140 ;
        RECT 39.395 164.080 39.715 164.140 ;
        RECT 44.915 164.080 45.235 164.140 ;
        RECT 49.975 164.080 50.295 164.340 ;
        RECT 54.590 164.280 54.880 164.325 ;
        RECT 59.175 164.280 59.495 164.340 ;
        RECT 54.590 164.140 59.495 164.280 ;
        RECT 54.590 164.095 54.880 164.140 ;
        RECT 59.175 164.080 59.495 164.140 ;
        RECT 60.095 164.080 60.415 164.340 ;
        RECT 63.775 164.080 64.095 164.340 ;
        RECT 64.235 164.280 64.555 164.340 ;
        RECT 68.375 164.280 68.695 164.340 ;
        RECT 64.235 164.140 68.695 164.280 ;
        RECT 64.235 164.080 64.555 164.140 ;
        RECT 68.375 164.080 68.695 164.140 ;
        RECT 68.835 164.080 69.155 164.340 ;
        RECT 80.335 164.280 80.655 164.340 ;
        RECT 83.800 164.280 84.090 164.325 ;
        RECT 80.335 164.140 84.090 164.280 ;
        RECT 80.335 164.080 80.655 164.140 ;
        RECT 83.800 164.095 84.090 164.140 ;
        RECT 87.235 164.280 87.555 164.340 ;
        RECT 88.155 164.280 88.475 164.340 ;
        RECT 91.375 164.280 91.695 164.340 ;
        RECT 87.235 164.140 91.695 164.280 ;
        RECT 87.235 164.080 87.555 164.140 ;
        RECT 88.155 164.080 88.475 164.140 ;
        RECT 91.375 164.080 91.695 164.140 ;
        RECT 91.835 164.280 92.155 164.340 ;
        RECT 94.610 164.280 94.900 164.325 ;
        RECT 91.835 164.140 94.900 164.280 ;
        RECT 91.835 164.080 92.155 164.140 ;
        RECT 94.610 164.095 94.900 164.140 ;
        RECT 100.130 164.280 100.420 164.325 ;
        RECT 101.955 164.280 102.275 164.340 ;
        RECT 100.130 164.140 102.275 164.280 ;
        RECT 100.130 164.095 100.420 164.140 ;
        RECT 101.955 164.080 102.275 164.140 ;
        RECT 18.165 163.460 112.465 163.940 ;
        RECT 26.975 163.260 27.295 163.320 ;
        RECT 32.035 163.260 32.355 163.320 ;
        RECT 40.315 163.260 40.635 163.320 ;
        RECT 63.790 163.260 64.080 163.305 ;
        RECT 65.615 163.260 65.935 163.320 ;
        RECT 70.215 163.260 70.535 163.320 ;
        RECT 80.335 163.260 80.655 163.320 ;
        RECT 84.030 163.260 84.320 163.305 ;
        RECT 85.855 163.260 86.175 163.320 ;
        RECT 26.975 163.120 40.085 163.260 ;
        RECT 26.975 163.060 27.295 163.120 ;
        RECT 32.035 163.060 32.355 163.120 ;
        RECT 21.930 162.735 22.220 162.965 ;
        RECT 25.250 162.920 25.540 162.965 ;
        RECT 28.370 162.920 28.660 162.965 ;
        RECT 30.260 162.920 30.550 162.965 ;
        RECT 25.250 162.780 30.550 162.920 ;
        RECT 25.250 162.735 25.540 162.780 ;
        RECT 28.370 162.735 28.660 162.780 ;
        RECT 30.260 162.735 30.550 162.780 ;
        RECT 39.410 162.735 39.700 162.965 ;
        RECT 39.945 162.920 40.085 163.120 ;
        RECT 40.315 163.120 66.995 163.260 ;
        RECT 40.315 163.060 40.635 163.120 ;
        RECT 63.790 163.075 64.080 163.120 ;
        RECT 65.615 163.060 65.935 163.120 ;
        RECT 43.535 162.920 43.855 162.980 ;
        RECT 47.215 162.920 47.535 162.980 ;
        RECT 39.945 162.780 47.535 162.920 ;
        RECT 20.090 162.580 20.380 162.625 ;
        RECT 22.005 162.580 22.145 162.735 ;
        RECT 29.750 162.580 30.040 162.625 ;
        RECT 20.090 162.440 21.685 162.580 ;
        RECT 22.005 162.440 30.040 162.580 ;
        RECT 20.090 162.395 20.380 162.440 ;
        RECT 20.550 162.055 20.840 162.285 ;
        RECT 20.625 161.900 20.765 162.055 ;
        RECT 20.995 162.040 21.315 162.300 ;
        RECT 21.545 162.240 21.685 162.440 ;
        RECT 29.750 162.395 30.040 162.440 ;
        RECT 31.130 162.580 31.420 162.625 ;
        RECT 32.495 162.580 32.815 162.640 ;
        RECT 38.935 162.580 39.255 162.640 ;
        RECT 31.130 162.440 39.255 162.580 ;
        RECT 39.485 162.580 39.625 162.735 ;
        RECT 43.535 162.720 43.855 162.780 ;
        RECT 47.215 162.720 47.535 162.780 ;
        RECT 49.530 162.920 49.820 162.965 ;
        RECT 50.895 162.920 51.215 162.980 ;
        RECT 49.530 162.780 51.215 162.920 ;
        RECT 49.530 162.735 49.820 162.780 ;
        RECT 50.895 162.720 51.215 162.780 ;
        RECT 52.390 162.920 52.680 162.965 ;
        RECT 55.510 162.920 55.800 162.965 ;
        RECT 57.400 162.920 57.690 162.965 ;
        RECT 52.390 162.780 57.690 162.920 ;
        RECT 52.390 162.735 52.680 162.780 ;
        RECT 55.510 162.735 55.800 162.780 ;
        RECT 57.400 162.735 57.690 162.780 ;
        RECT 61.935 162.920 62.255 162.980 ;
        RECT 64.235 162.920 64.555 162.980 ;
        RECT 61.935 162.780 64.555 162.920 ;
        RECT 66.855 162.920 66.995 163.120 ;
        RECT 70.215 163.120 77.115 163.260 ;
        RECT 70.215 163.060 70.535 163.120 ;
        RECT 72.975 162.920 73.295 162.980 ;
        RECT 76.975 162.920 77.115 163.120 ;
        RECT 80.335 163.120 83.785 163.260 ;
        RECT 80.335 163.060 80.655 163.120 ;
        RECT 66.855 162.780 74.125 162.920 ;
        RECT 76.975 162.780 77.345 162.920 ;
        RECT 61.935 162.720 62.255 162.780 ;
        RECT 64.235 162.720 64.555 162.780 ;
        RECT 72.975 162.720 73.295 162.780 ;
        RECT 43.995 162.580 44.315 162.640 ;
        RECT 54.575 162.580 54.895 162.640 ;
        RECT 58.270 162.580 58.560 162.625 ;
        RECT 39.485 162.440 58.560 162.580 ;
        RECT 31.130 162.395 31.420 162.440 ;
        RECT 32.495 162.380 32.815 162.440 ;
        RECT 38.935 162.380 39.255 162.440 ;
        RECT 43.995 162.380 44.315 162.440 ;
        RECT 24.170 162.240 24.460 162.260 ;
        RECT 21.545 162.100 24.460 162.240 ;
        RECT 21.915 161.900 22.235 161.960 ;
        RECT 24.170 161.945 24.460 162.100 ;
        RECT 25.250 162.240 25.540 162.285 ;
        RECT 28.830 162.240 29.120 162.285 ;
        RECT 30.665 162.240 30.955 162.285 ;
        RECT 25.250 162.100 30.955 162.240 ;
        RECT 25.250 162.055 25.540 162.100 ;
        RECT 28.830 162.055 29.120 162.100 ;
        RECT 30.665 162.055 30.955 162.100 ;
        RECT 42.615 162.240 42.935 162.300 ;
        RECT 46.845 162.285 46.985 162.440 ;
        RECT 54.575 162.380 54.895 162.440 ;
        RECT 58.270 162.395 58.560 162.440 ;
        RECT 69.295 162.580 69.615 162.640 ;
        RECT 70.690 162.580 70.980 162.625 ;
        RECT 69.295 162.440 70.980 162.580 ;
        RECT 69.295 162.380 69.615 162.440 ;
        RECT 70.690 162.395 70.980 162.440 ;
        RECT 45.850 162.240 46.140 162.285 ;
        RECT 42.615 162.100 46.140 162.240 ;
        RECT 42.615 162.040 42.935 162.100 ;
        RECT 45.850 162.055 46.140 162.100 ;
        RECT 46.770 162.055 47.060 162.285 ;
        RECT 49.975 162.240 50.295 162.300 ;
        RECT 51.310 162.240 51.600 162.260 ;
        RECT 49.975 162.100 51.600 162.240 ;
        RECT 49.975 162.040 50.295 162.100 ;
        RECT 51.310 161.945 51.600 162.100 ;
        RECT 52.390 162.240 52.680 162.285 ;
        RECT 55.970 162.240 56.260 162.285 ;
        RECT 57.805 162.240 58.095 162.285 ;
        RECT 52.390 162.100 58.095 162.240 ;
        RECT 52.390 162.055 52.680 162.100 ;
        RECT 55.970 162.055 56.260 162.100 ;
        RECT 57.805 162.055 58.095 162.100 ;
        RECT 61.475 162.240 61.795 162.300 ;
        RECT 64.710 162.240 65.000 162.285 ;
        RECT 66.535 162.240 66.855 162.300 ;
        RECT 61.475 162.100 66.855 162.240 ;
        RECT 61.475 162.040 61.795 162.100 ;
        RECT 64.710 162.055 65.000 162.100 ;
        RECT 66.535 162.040 66.855 162.100 ;
        RECT 66.995 162.240 67.315 162.300 ;
        RECT 68.850 162.240 69.140 162.285 ;
        RECT 66.995 162.100 69.140 162.240 ;
        RECT 66.995 162.040 67.315 162.100 ;
        RECT 68.850 162.055 69.140 162.100 ;
        RECT 69.755 162.240 70.075 162.300 ;
        RECT 73.985 162.285 74.125 162.780 ;
        RECT 74.355 162.580 74.675 162.640 ;
        RECT 77.205 162.625 77.345 162.780 ;
        RECT 82.190 162.735 82.480 162.965 ;
        RECT 83.645 162.920 83.785 163.120 ;
        RECT 84.030 163.120 86.175 163.260 ;
        RECT 84.030 163.075 84.320 163.120 ;
        RECT 85.855 163.060 86.175 163.120 ;
        RECT 87.695 163.260 88.015 163.320 ;
        RECT 90.915 163.260 91.235 163.320 ;
        RECT 91.850 163.260 92.140 163.305 ;
        RECT 87.695 163.120 89.765 163.260 ;
        RECT 87.695 163.060 88.015 163.120 ;
        RECT 83.645 162.780 89.305 162.920 ;
        RECT 76.670 162.580 76.960 162.625 ;
        RECT 74.355 162.440 76.960 162.580 ;
        RECT 74.355 162.380 74.675 162.440 ;
        RECT 76.670 162.395 76.960 162.440 ;
        RECT 77.130 162.580 77.420 162.625 ;
        RECT 79.430 162.580 79.720 162.625 ;
        RECT 80.795 162.580 81.115 162.640 ;
        RECT 77.130 162.440 81.115 162.580 ;
        RECT 82.265 162.580 82.405 162.735 ;
        RECT 87.235 162.580 87.555 162.640 ;
        RECT 89.165 162.625 89.305 162.780 ;
        RECT 88.170 162.580 88.460 162.625 ;
        RECT 82.265 162.440 86.085 162.580 ;
        RECT 77.130 162.395 77.420 162.440 ;
        RECT 79.430 162.395 79.720 162.440 ;
        RECT 80.795 162.380 81.115 162.440 ;
        RECT 72.070 162.240 72.360 162.285 ;
        RECT 69.755 162.100 72.360 162.240 ;
        RECT 69.755 162.040 70.075 162.100 ;
        RECT 72.070 162.055 72.360 162.100 ;
        RECT 72.530 162.055 72.820 162.285 ;
        RECT 72.990 162.240 73.280 162.285 ;
        RECT 72.990 162.100 73.665 162.240 ;
        RECT 72.990 162.055 73.280 162.100 ;
        RECT 20.625 161.760 22.235 161.900 ;
        RECT 21.915 161.700 22.235 161.760 ;
        RECT 23.870 161.900 24.460 161.945 ;
        RECT 27.110 161.900 27.760 161.945 ;
        RECT 23.870 161.760 27.760 161.900 ;
        RECT 23.870 161.715 24.160 161.760 ;
        RECT 27.110 161.715 27.760 161.760 ;
        RECT 51.010 161.900 51.600 161.945 ;
        RECT 54.250 161.900 54.900 161.945 ;
        RECT 51.010 161.760 54.900 161.900 ;
        RECT 51.010 161.715 51.300 161.760 ;
        RECT 54.250 161.715 54.900 161.760 ;
        RECT 56.890 161.900 57.180 161.945 ;
        RECT 58.255 161.900 58.575 161.960 ;
        RECT 71.595 161.900 71.915 161.960 ;
        RECT 72.605 161.900 72.745 162.055 ;
        RECT 56.890 161.760 58.575 161.900 ;
        RECT 56.890 161.715 57.180 161.760 ;
        RECT 58.255 161.700 58.575 161.760 ;
        RECT 66.855 161.760 72.745 161.900 ;
        RECT 73.525 161.900 73.665 162.100 ;
        RECT 73.910 162.055 74.200 162.285 ;
        RECT 78.955 162.240 79.275 162.300 ;
        RECT 85.945 162.285 86.085 162.440 ;
        RECT 87.235 162.440 88.460 162.580 ;
        RECT 87.235 162.380 87.555 162.440 ;
        RECT 88.170 162.395 88.460 162.440 ;
        RECT 89.090 162.395 89.380 162.625 ;
        RECT 89.625 162.580 89.765 163.120 ;
        RECT 90.915 163.120 92.140 163.260 ;
        RECT 90.915 163.060 91.235 163.120 ;
        RECT 91.850 163.075 92.140 163.120 ;
        RECT 103.795 162.920 104.115 162.980 ;
        RECT 91.925 162.780 104.115 162.920 ;
        RECT 91.925 162.580 92.065 162.780 ;
        RECT 103.795 162.720 104.115 162.780 ;
        RECT 104.270 162.920 104.560 162.965 ;
        RECT 104.270 162.780 109.085 162.920 ;
        RECT 104.270 162.735 104.560 162.780 ;
        RECT 89.625 162.440 92.065 162.580 ;
        RECT 83.570 162.240 83.860 162.285 ;
        RECT 78.955 162.100 85.625 162.240 ;
        RECT 78.955 162.040 79.275 162.100 ;
        RECT 83.570 162.055 83.860 162.100 ;
        RECT 76.210 161.900 76.500 161.945 ;
        RECT 77.115 161.900 77.435 161.960 ;
        RECT 79.890 161.900 80.180 161.945 ;
        RECT 73.525 161.760 80.180 161.900 ;
        RECT 85.485 161.900 85.625 162.100 ;
        RECT 85.870 162.055 86.160 162.285 ;
        RECT 87.695 162.240 88.015 162.300 ;
        RECT 86.405 162.100 88.015 162.240 ;
        RECT 88.245 162.240 88.385 162.395 ;
        RECT 94.595 162.380 94.915 162.640 ;
        RECT 101.510 162.580 101.800 162.625 ;
        RECT 102.875 162.580 103.195 162.640 ;
        RECT 95.145 162.440 96.665 162.580 ;
        RECT 89.995 162.240 90.315 162.300 ;
        RECT 92.770 162.240 93.060 162.285 ;
        RECT 88.245 162.100 90.315 162.240 ;
        RECT 86.405 161.900 86.545 162.100 ;
        RECT 87.695 162.040 88.015 162.100 ;
        RECT 89.995 162.040 90.315 162.100 ;
        RECT 90.545 162.100 93.060 162.240 ;
        RECT 85.485 161.760 86.545 161.900 ;
        RECT 22.390 161.560 22.680 161.605 ;
        RECT 26.055 161.560 26.375 161.620 ;
        RECT 22.390 161.420 26.375 161.560 ;
        RECT 22.390 161.375 22.680 161.420 ;
        RECT 26.055 161.360 26.375 161.420 ;
        RECT 38.015 161.560 38.335 161.620 ;
        RECT 49.975 161.560 50.295 161.620 ;
        RECT 60.095 161.560 60.415 161.620 ;
        RECT 66.075 161.560 66.395 161.620 ;
        RECT 66.855 161.560 66.995 161.760 ;
        RECT 71.595 161.700 71.915 161.760 ;
        RECT 76.210 161.715 76.500 161.760 ;
        RECT 77.115 161.700 77.435 161.760 ;
        RECT 79.890 161.715 80.180 161.760 ;
        RECT 38.015 161.420 66.995 161.560 ;
        RECT 38.015 161.360 38.335 161.420 ;
        RECT 49.975 161.360 50.295 161.420 ;
        RECT 60.095 161.360 60.415 161.420 ;
        RECT 66.075 161.360 66.395 161.420 ;
        RECT 67.915 161.360 68.235 161.620 ;
        RECT 74.370 161.560 74.660 161.605 ;
        RECT 75.275 161.560 75.595 161.620 ;
        RECT 74.370 161.420 75.595 161.560 ;
        RECT 74.370 161.375 74.660 161.420 ;
        RECT 75.275 161.360 75.595 161.420 ;
        RECT 75.735 161.560 76.055 161.620 ;
        RECT 80.335 161.560 80.655 161.620 ;
        RECT 75.735 161.420 80.655 161.560 ;
        RECT 75.735 161.360 76.055 161.420 ;
        RECT 80.335 161.360 80.655 161.420 ;
        RECT 84.015 161.560 84.335 161.620 ;
        RECT 84.950 161.560 85.240 161.605 ;
        RECT 84.015 161.420 85.240 161.560 ;
        RECT 84.015 161.360 84.335 161.420 ;
        RECT 84.950 161.375 85.240 161.420 ;
        RECT 89.550 161.560 89.840 161.605 ;
        RECT 89.995 161.560 90.315 161.620 ;
        RECT 89.550 161.420 90.315 161.560 ;
        RECT 90.545 161.560 90.685 162.100 ;
        RECT 92.770 162.055 93.060 162.100 ;
        RECT 90.915 161.900 91.235 161.960 ;
        RECT 95.145 161.900 95.285 162.440 ;
        RECT 96.525 162.300 96.665 162.440 ;
        RECT 96.985 162.440 99.425 162.580 ;
        RECT 95.990 162.055 96.280 162.285 ;
        RECT 90.915 161.760 95.285 161.900 ;
        RECT 95.515 161.900 95.835 161.960 ;
        RECT 96.065 161.900 96.205 162.055 ;
        RECT 96.435 162.040 96.755 162.300 ;
        RECT 96.985 162.285 97.125 162.440 ;
        RECT 96.910 162.055 97.200 162.285 ;
        RECT 97.355 162.240 97.675 162.300 ;
        RECT 97.830 162.240 98.120 162.285 ;
        RECT 97.355 162.100 98.120 162.240 ;
        RECT 99.285 162.240 99.425 162.440 ;
        RECT 101.510 162.440 103.195 162.580 ;
        RECT 101.510 162.395 101.800 162.440 ;
        RECT 102.875 162.380 103.195 162.440 ;
        RECT 101.955 162.240 102.275 162.300 ;
        RECT 102.430 162.240 102.720 162.285 ;
        RECT 99.285 162.100 102.720 162.240 ;
        RECT 97.355 162.040 97.675 162.100 ;
        RECT 97.830 162.055 98.120 162.100 ;
        RECT 101.955 162.040 102.275 162.100 ;
        RECT 102.430 162.055 102.720 162.100 ;
        RECT 103.795 162.240 104.115 162.300 ;
        RECT 104.730 162.240 105.020 162.285 ;
        RECT 103.795 162.100 105.020 162.240 ;
        RECT 103.795 162.040 104.115 162.100 ;
        RECT 104.730 162.055 105.020 162.100 ;
        RECT 105.175 162.040 105.495 162.300 ;
        RECT 107.935 162.040 108.255 162.300 ;
        RECT 108.945 162.285 109.085 162.780 ;
        RECT 108.870 162.055 109.160 162.285 ;
        RECT 95.515 161.760 96.205 161.900 ;
        RECT 90.915 161.700 91.235 161.760 ;
        RECT 95.515 161.700 95.835 161.760 ;
        RECT 91.390 161.560 91.680 161.605 ;
        RECT 90.545 161.420 91.680 161.560 ;
        RECT 89.550 161.375 89.840 161.420 ;
        RECT 89.995 161.360 90.315 161.420 ;
        RECT 91.390 161.375 91.680 161.420 ;
        RECT 96.435 161.560 96.755 161.620 ;
        RECT 97.445 161.560 97.585 162.040 ;
        RECT 96.435 161.420 97.585 161.560 ;
        RECT 96.435 161.360 96.755 161.420 ;
        RECT 101.955 161.360 102.275 161.620 ;
        RECT 102.415 161.560 102.735 161.620 ;
        RECT 107.490 161.560 107.780 161.605 ;
        RECT 102.415 161.420 107.780 161.560 ;
        RECT 102.415 161.360 102.735 161.420 ;
        RECT 107.490 161.375 107.780 161.420 ;
        RECT 109.775 161.360 110.095 161.620 ;
        RECT 17.370 160.740 112.465 161.220 ;
        RECT 27.895 160.540 28.215 160.600 ;
        RECT 24.305 160.400 28.215 160.540 ;
        RECT 24.305 160.200 24.445 160.400 ;
        RECT 27.895 160.340 28.215 160.400 ;
        RECT 28.815 160.540 29.135 160.600 ;
        RECT 29.750 160.540 30.040 160.585 ;
        RECT 28.815 160.400 30.040 160.540 ;
        RECT 28.815 160.340 29.135 160.400 ;
        RECT 29.750 160.355 30.040 160.400 ;
        RECT 45.375 160.340 45.695 160.600 ;
        RECT 47.230 160.540 47.520 160.585 ;
        RECT 49.055 160.540 49.375 160.600 ;
        RECT 47.230 160.400 49.375 160.540 ;
        RECT 47.230 160.355 47.520 160.400 ;
        RECT 49.055 160.340 49.375 160.400 ;
        RECT 49.515 160.540 49.835 160.600 ;
        RECT 52.275 160.540 52.595 160.600 ;
        RECT 49.515 160.400 52.595 160.540 ;
        RECT 49.515 160.340 49.835 160.400 ;
        RECT 52.275 160.340 52.595 160.400 ;
        RECT 58.255 160.340 58.575 160.600 ;
        RECT 61.935 160.540 62.255 160.600 ;
        RECT 65.630 160.540 65.920 160.585 ;
        RECT 89.995 160.540 90.315 160.600 ;
        RECT 91.375 160.540 91.695 160.600 ;
        RECT 101.955 160.585 102.275 160.600 ;
        RECT 101.740 160.540 102.275 160.585 ;
        RECT 61.935 160.400 65.920 160.540 ;
        RECT 61.935 160.340 62.255 160.400 ;
        RECT 65.630 160.355 65.920 160.400 ;
        RECT 69.385 160.400 89.765 160.540 ;
        RECT 33.415 160.200 33.735 160.260 ;
        RECT 23.845 160.060 24.445 160.200 ;
        RECT 24.765 160.060 33.735 160.200 ;
        RECT 23.845 159.905 23.985 160.060 ;
        RECT 23.770 159.675 24.060 159.905 ;
        RECT 24.215 159.660 24.535 159.920 ;
        RECT 24.765 159.905 24.905 160.060 ;
        RECT 33.415 160.000 33.735 160.060 ;
        RECT 43.075 160.200 43.395 160.260 ;
        RECT 43.075 160.060 50.665 160.200 ;
        RECT 43.075 160.000 43.395 160.060 ;
        RECT 24.690 159.675 24.980 159.905 ;
        RECT 25.595 159.660 25.915 159.920 ;
        RECT 26.055 159.860 26.375 159.920 ;
        RECT 27.910 159.860 28.200 159.905 ;
        RECT 31.575 159.860 31.895 159.920 ;
        RECT 26.055 159.720 31.895 159.860 ;
        RECT 26.055 159.660 26.375 159.720 ;
        RECT 27.910 159.675 28.200 159.720 ;
        RECT 31.575 159.660 31.895 159.720 ;
        RECT 38.935 159.860 39.255 159.920 ;
        RECT 39.870 159.860 40.160 159.905 ;
        RECT 38.935 159.720 40.160 159.860 ;
        RECT 38.935 159.660 39.255 159.720 ;
        RECT 39.870 159.675 40.160 159.720 ;
        RECT 49.515 159.660 49.835 159.920 ;
        RECT 49.975 159.660 50.295 159.920 ;
        RECT 50.525 159.905 50.665 160.060 ;
        RECT 50.985 160.060 54.805 160.200 ;
        RECT 50.450 159.675 50.740 159.905 ;
        RECT 26.975 159.320 27.295 159.580 ;
        RECT 27.435 159.320 27.755 159.580 ;
        RECT 43.535 159.520 43.855 159.580 ;
        RECT 44.010 159.520 44.300 159.565 ;
        RECT 43.535 159.380 44.300 159.520 ;
        RECT 43.535 159.320 43.855 159.380 ;
        RECT 44.010 159.335 44.300 159.380 ;
        RECT 44.915 159.320 45.235 159.580 ;
        RECT 50.985 159.520 51.125 160.060 ;
        RECT 51.370 159.675 51.660 159.905 ;
        RECT 53.210 159.675 53.500 159.905 ;
        RECT 45.465 159.380 51.125 159.520 ;
        RECT 27.525 159.180 27.665 159.320 ;
        RECT 45.465 159.180 45.605 159.380 ;
        RECT 27.525 159.040 45.605 159.180 ;
        RECT 49.055 159.180 49.375 159.240 ;
        RECT 51.445 159.180 51.585 159.675 ;
        RECT 53.285 159.520 53.425 159.675 ;
        RECT 53.655 159.660 53.975 159.920 ;
        RECT 54.130 159.875 54.420 159.905 ;
        RECT 54.665 159.875 54.805 160.060 ;
        RECT 56.415 160.000 56.735 160.260 ;
        RECT 67.915 160.200 68.235 160.260 ;
        RECT 64.785 160.060 68.235 160.200 ;
        RECT 54.130 159.735 54.805 159.875 ;
        RECT 55.050 159.860 55.340 159.905 ;
        RECT 54.130 159.675 54.420 159.735 ;
        RECT 55.050 159.720 57.105 159.860 ;
        RECT 55.050 159.675 55.340 159.720 ;
        RECT 54.575 159.520 54.895 159.580 ;
        RECT 53.285 159.380 54.895 159.520 ;
        RECT 54.575 159.320 54.895 159.380 ;
        RECT 56.965 159.520 57.105 159.720 ;
        RECT 57.795 159.660 58.115 159.920 ;
        RECT 59.175 159.660 59.495 159.920 ;
        RECT 61.030 159.860 61.320 159.905 ;
        RECT 61.475 159.860 61.795 159.920 ;
        RECT 61.030 159.720 61.795 159.860 ;
        RECT 61.030 159.675 61.320 159.720 ;
        RECT 61.475 159.660 61.795 159.720 ;
        RECT 62.870 159.860 63.160 159.905 ;
        RECT 63.775 159.860 64.095 159.920 ;
        RECT 64.785 159.905 64.925 160.060 ;
        RECT 67.915 160.000 68.235 160.060 ;
        RECT 62.870 159.720 64.095 159.860 ;
        RECT 62.870 159.675 63.160 159.720 ;
        RECT 63.775 159.660 64.095 159.720 ;
        RECT 64.710 159.675 65.000 159.905 ;
        RECT 66.535 159.660 66.855 159.920 ;
        RECT 69.385 159.520 69.525 160.400 ;
        RECT 74.370 160.200 74.660 160.245 ;
        RECT 78.905 160.200 79.195 160.245 ;
        RECT 82.165 160.200 82.455 160.245 ;
        RECT 74.370 160.060 82.455 160.200 ;
        RECT 74.370 160.015 74.660 160.060 ;
        RECT 78.905 160.015 79.195 160.060 ;
        RECT 82.165 160.015 82.455 160.060 ;
        RECT 83.085 160.200 83.375 160.245 ;
        RECT 84.945 160.200 85.235 160.245 ;
        RECT 83.085 160.060 85.235 160.200 ;
        RECT 89.625 160.200 89.765 160.400 ;
        RECT 89.995 160.400 102.275 160.540 ;
        RECT 89.995 160.340 90.315 160.400 ;
        RECT 91.375 160.340 91.695 160.400 ;
        RECT 101.740 160.355 102.275 160.400 ;
        RECT 101.955 160.340 102.275 160.355 ;
        RECT 93.215 160.200 93.535 160.260 ;
        RECT 103.745 160.200 104.035 160.245 ;
        RECT 105.175 160.200 105.495 160.260 ;
        RECT 107.005 160.200 107.295 160.245 ;
        RECT 89.625 160.060 98.965 160.200 ;
        RECT 83.085 160.015 83.375 160.060 ;
        RECT 84.945 160.015 85.235 160.060 ;
        RECT 69.755 159.860 70.075 159.920 ;
        RECT 71.150 159.860 71.440 159.905 ;
        RECT 69.755 159.720 71.440 159.860 ;
        RECT 69.755 159.660 70.075 159.720 ;
        RECT 71.150 159.675 71.440 159.720 ;
        RECT 71.595 159.660 71.915 159.920 ;
        RECT 72.070 159.675 72.360 159.905 ;
        RECT 56.965 159.380 69.525 159.520 ;
        RECT 72.145 159.520 72.285 159.675 ;
        RECT 72.975 159.660 73.295 159.920 ;
        RECT 74.830 159.675 75.120 159.905 ;
        RECT 74.355 159.520 74.675 159.580 ;
        RECT 72.145 159.380 74.675 159.520 ;
        RECT 74.905 159.520 75.045 159.675 ;
        RECT 75.275 159.660 75.595 159.920 ;
        RECT 77.115 159.905 77.435 159.920 ;
        RECT 76.900 159.675 77.435 159.905 ;
        RECT 80.765 159.860 81.055 159.905 ;
        RECT 83.085 159.860 83.300 160.015 ;
        RECT 93.215 160.000 93.535 160.060 ;
        RECT 98.825 159.920 98.965 160.060 ;
        RECT 103.745 160.060 107.295 160.200 ;
        RECT 103.745 160.015 104.035 160.060 ;
        RECT 105.175 160.000 105.495 160.060 ;
        RECT 107.005 160.015 107.295 160.060 ;
        RECT 107.925 160.200 108.215 160.245 ;
        RECT 109.785 160.200 110.075 160.245 ;
        RECT 107.925 160.060 110.075 160.200 ;
        RECT 107.925 160.015 108.215 160.060 ;
        RECT 109.785 160.015 110.075 160.060 ;
        RECT 80.765 159.720 83.300 159.860 ;
        RECT 80.765 159.675 81.055 159.720 ;
        RECT 77.115 159.660 77.435 159.675 ;
        RECT 84.015 159.660 84.335 159.920 ;
        RECT 95.055 159.660 95.375 159.920 ;
        RECT 95.515 159.860 95.835 159.920 ;
        RECT 96.910 159.860 97.200 159.905 ;
        RECT 95.515 159.720 97.200 159.860 ;
        RECT 95.515 159.660 95.835 159.720 ;
        RECT 96.910 159.675 97.200 159.720 ;
        RECT 97.355 159.660 97.675 159.920 ;
        RECT 97.815 159.660 98.135 159.920 ;
        RECT 98.735 159.660 99.055 159.920 ;
        RECT 105.605 159.860 105.895 159.905 ;
        RECT 107.925 159.860 108.140 160.015 ;
        RECT 105.605 159.720 108.140 159.860 ;
        RECT 109.315 159.860 109.635 159.920 ;
        RECT 110.710 159.860 111.000 159.905 ;
        RECT 109.315 159.720 111.000 159.860 ;
        RECT 105.605 159.675 105.895 159.720 ;
        RECT 109.315 159.660 109.635 159.720 ;
        RECT 110.710 159.675 111.000 159.720 ;
        RECT 78.955 159.520 79.275 159.580 ;
        RECT 74.905 159.380 79.275 159.520 ;
        RECT 56.965 159.180 57.105 159.380 ;
        RECT 60.185 159.225 60.325 159.380 ;
        RECT 74.355 159.320 74.675 159.380 ;
        RECT 78.955 159.320 79.275 159.380 ;
        RECT 82.635 159.520 82.955 159.580 ;
        RECT 85.870 159.520 86.160 159.565 ;
        RECT 82.635 159.380 86.160 159.520 ;
        RECT 82.635 159.320 82.955 159.380 ;
        RECT 85.870 159.335 86.160 159.380 ;
        RECT 108.870 159.520 109.160 159.565 ;
        RECT 109.775 159.520 110.095 159.580 ;
        RECT 108.870 159.380 110.095 159.520 ;
        RECT 108.870 159.335 109.160 159.380 ;
        RECT 109.775 159.320 110.095 159.380 ;
        RECT 49.055 159.040 57.105 159.180 ;
        RECT 49.055 158.980 49.375 159.040 ;
        RECT 60.110 158.995 60.400 159.225 ;
        RECT 61.950 159.180 62.240 159.225 ;
        RECT 80.765 159.180 81.055 159.225 ;
        RECT 83.545 159.180 83.835 159.225 ;
        RECT 85.405 159.180 85.695 159.225 ;
        RECT 60.645 159.040 80.565 159.180 ;
        RECT 22.390 158.840 22.680 158.885 ;
        RECT 23.295 158.840 23.615 158.900 ;
        RECT 22.390 158.700 23.615 158.840 ;
        RECT 22.390 158.655 22.680 158.700 ;
        RECT 23.295 158.640 23.615 158.700 ;
        RECT 47.675 158.840 47.995 158.900 ;
        RECT 48.150 158.840 48.440 158.885 ;
        RECT 47.675 158.700 48.440 158.840 ;
        RECT 47.675 158.640 47.995 158.700 ;
        RECT 48.150 158.655 48.440 158.700 ;
        RECT 51.355 158.840 51.675 158.900 ;
        RECT 51.830 158.840 52.120 158.885 ;
        RECT 51.355 158.700 52.120 158.840 ;
        RECT 51.355 158.640 51.675 158.700 ;
        RECT 51.830 158.655 52.120 158.700 ;
        RECT 54.575 158.840 54.895 158.900 ;
        RECT 60.645 158.840 60.785 159.040 ;
        RECT 61.950 158.995 62.240 159.040 ;
        RECT 54.575 158.700 60.785 158.840 ;
        RECT 61.475 158.840 61.795 158.900 ;
        RECT 63.790 158.840 64.080 158.885 ;
        RECT 61.475 158.700 64.080 158.840 ;
        RECT 54.575 158.640 54.895 158.700 ;
        RECT 61.475 158.640 61.795 158.700 ;
        RECT 63.790 158.655 64.080 158.700 ;
        RECT 69.770 158.840 70.060 158.885 ;
        RECT 71.135 158.840 71.455 158.900 ;
        RECT 69.770 158.700 71.455 158.840 ;
        RECT 69.770 158.655 70.060 158.700 ;
        RECT 71.135 158.640 71.455 158.700 ;
        RECT 76.210 158.840 76.500 158.885 ;
        RECT 78.035 158.840 78.355 158.900 ;
        RECT 76.210 158.700 78.355 158.840 ;
        RECT 80.425 158.840 80.565 159.040 ;
        RECT 80.765 159.040 85.695 159.180 ;
        RECT 80.765 158.995 81.055 159.040 ;
        RECT 83.545 158.995 83.835 159.040 ;
        RECT 85.405 158.995 85.695 159.040 ;
        RECT 86.315 159.180 86.635 159.240 ;
        RECT 102.415 159.180 102.735 159.240 ;
        RECT 86.315 159.040 102.735 159.180 ;
        RECT 86.315 158.980 86.635 159.040 ;
        RECT 102.415 158.980 102.735 159.040 ;
        RECT 105.605 159.180 105.895 159.225 ;
        RECT 108.385 159.180 108.675 159.225 ;
        RECT 110.245 159.180 110.535 159.225 ;
        RECT 105.605 159.040 110.535 159.180 ;
        RECT 105.605 158.995 105.895 159.040 ;
        RECT 108.385 158.995 108.675 159.040 ;
        RECT 110.245 158.995 110.535 159.040 ;
        RECT 87.695 158.840 88.015 158.900 ;
        RECT 80.425 158.700 88.015 158.840 ;
        RECT 76.210 158.655 76.500 158.700 ;
        RECT 78.035 158.640 78.355 158.700 ;
        RECT 87.695 158.640 88.015 158.700 ;
        RECT 88.630 158.840 88.920 158.885 ;
        RECT 89.995 158.840 90.315 158.900 ;
        RECT 88.630 158.700 90.315 158.840 ;
        RECT 88.630 158.655 88.920 158.700 ;
        RECT 89.995 158.640 90.315 158.700 ;
        RECT 94.595 158.840 94.915 158.900 ;
        RECT 95.530 158.840 95.820 158.885 ;
        RECT 94.595 158.700 95.820 158.840 ;
        RECT 94.595 158.640 94.915 158.700 ;
        RECT 95.530 158.655 95.820 158.700 ;
        RECT 18.165 158.020 112.465 158.500 ;
        RECT 20.995 157.820 21.315 157.880 ;
        RECT 21.470 157.820 21.760 157.865 ;
        RECT 20.995 157.680 21.760 157.820 ;
        RECT 20.995 157.620 21.315 157.680 ;
        RECT 21.470 157.635 21.760 157.680 ;
        RECT 22.835 157.820 23.155 157.880 ;
        RECT 49.515 157.820 49.835 157.880 ;
        RECT 57.335 157.820 57.655 157.880 ;
        RECT 61.015 157.820 61.335 157.880 ;
        RECT 62.410 157.820 62.700 157.865 ;
        RECT 72.055 157.820 72.375 157.880 ;
        RECT 22.835 157.680 53.195 157.820 ;
        RECT 22.835 157.620 23.155 157.680 ;
        RECT 49.515 157.620 49.835 157.680 ;
        RECT 26.975 157.480 27.295 157.540 ;
        RECT 24.765 157.340 27.295 157.480 ;
        RECT 24.765 157.185 24.905 157.340 ;
        RECT 26.975 157.280 27.295 157.340 ;
        RECT 28.470 157.480 28.760 157.525 ;
        RECT 31.590 157.480 31.880 157.525 ;
        RECT 33.480 157.480 33.770 157.525 ;
        RECT 28.470 157.340 33.770 157.480 ;
        RECT 28.470 157.295 28.760 157.340 ;
        RECT 31.590 157.295 31.880 157.340 ;
        RECT 33.480 157.295 33.770 157.340 ;
        RECT 38.130 157.480 38.420 157.525 ;
        RECT 41.250 157.480 41.540 157.525 ;
        RECT 43.140 157.480 43.430 157.525 ;
        RECT 38.130 157.340 43.430 157.480 ;
        RECT 38.130 157.295 38.420 157.340 ;
        RECT 41.250 157.295 41.540 157.340 ;
        RECT 43.140 157.295 43.430 157.340 ;
        RECT 47.215 157.480 47.535 157.540 ;
        RECT 53.055 157.480 53.195 157.680 ;
        RECT 57.335 157.680 72.375 157.820 ;
        RECT 57.335 157.620 57.655 157.680 ;
        RECT 61.015 157.620 61.335 157.680 ;
        RECT 62.410 157.635 62.700 157.680 ;
        RECT 72.055 157.620 72.375 157.680 ;
        RECT 73.680 157.820 73.970 157.865 ;
        RECT 74.355 157.820 74.675 157.880 ;
        RECT 86.315 157.820 86.635 157.880 ;
        RECT 73.680 157.680 74.675 157.820 ;
        RECT 73.680 157.635 73.970 157.680 ;
        RECT 74.355 157.620 74.675 157.680 ;
        RECT 74.905 157.680 86.635 157.820 ;
        RECT 74.905 157.480 75.045 157.680 ;
        RECT 86.315 157.620 86.635 157.680 ;
        RECT 47.215 157.340 50.665 157.480 ;
        RECT 53.055 157.340 66.305 157.480 ;
        RECT 47.215 157.280 47.535 157.340 ;
        RECT 24.690 156.955 24.980 157.185 ;
        RECT 25.610 157.140 25.900 157.185 ;
        RECT 29.275 157.140 29.595 157.200 ;
        RECT 25.610 157.000 29.595 157.140 ;
        RECT 25.610 156.955 25.900 157.000 ;
        RECT 29.275 156.940 29.595 157.000 ;
        RECT 31.115 157.140 31.435 157.200 ;
        RECT 32.970 157.140 33.260 157.185 ;
        RECT 31.115 157.000 33.260 157.140 ;
        RECT 31.115 156.940 31.435 157.000 ;
        RECT 32.970 156.955 33.260 157.000 ;
        RECT 34.335 157.140 34.655 157.200 ;
        RECT 38.935 157.140 39.255 157.200 ;
        RECT 34.335 157.000 39.255 157.140 ;
        RECT 34.335 156.940 34.655 157.000 ;
        RECT 38.935 156.940 39.255 157.000 ;
        RECT 43.995 156.940 44.315 157.200 ;
        RECT 44.915 157.140 45.235 157.200 ;
        RECT 50.525 157.140 50.665 157.340 ;
        RECT 52.275 157.140 52.595 157.200 ;
        RECT 44.915 157.000 47.905 157.140 ;
        RECT 44.915 156.940 45.235 157.000 ;
        RECT 21.010 156.800 21.300 156.845 ;
        RECT 22.835 156.800 23.155 156.860 ;
        RECT 21.010 156.660 23.155 156.800 ;
        RECT 21.010 156.615 21.300 156.660 ;
        RECT 22.835 156.600 23.155 156.660 ;
        RECT 23.770 156.800 24.060 156.845 ;
        RECT 26.055 156.800 26.375 156.860 ;
        RECT 23.770 156.660 26.375 156.800 ;
        RECT 23.770 156.615 24.060 156.660 ;
        RECT 26.055 156.600 26.375 156.660 ;
        RECT 21.915 156.460 22.235 156.520 ;
        RECT 27.390 156.505 27.680 156.820 ;
        RECT 28.470 156.800 28.760 156.845 ;
        RECT 32.050 156.800 32.340 156.845 ;
        RECT 33.885 156.800 34.175 156.845 ;
        RECT 28.470 156.660 34.175 156.800 ;
        RECT 28.470 156.615 28.760 156.660 ;
        RECT 32.050 156.615 32.340 156.660 ;
        RECT 33.885 156.615 34.175 156.660 ;
        RECT 37.050 156.505 37.340 156.820 ;
        RECT 38.130 156.800 38.420 156.845 ;
        RECT 41.710 156.800 42.000 156.845 ;
        RECT 43.545 156.800 43.835 156.845 ;
        RECT 46.755 156.800 47.075 156.860 ;
        RECT 38.130 156.660 43.835 156.800 ;
        RECT 38.130 156.615 38.420 156.660 ;
        RECT 41.710 156.615 42.000 156.660 ;
        RECT 43.545 156.615 43.835 156.660 ;
        RECT 46.385 156.660 47.075 156.800 ;
        RECT 27.090 156.460 27.680 156.505 ;
        RECT 30.330 156.460 30.980 156.505 ;
        RECT 36.750 156.460 37.340 156.505 ;
        RECT 39.990 156.460 40.640 156.505 ;
        RECT 21.915 156.320 30.980 156.460 ;
        RECT 21.915 156.260 22.235 156.320 ;
        RECT 27.090 156.275 27.380 156.320 ;
        RECT 30.330 156.275 30.980 156.320 ;
        RECT 31.205 156.320 40.640 156.460 ;
        RECT 20.535 155.920 20.855 156.180 ;
        RECT 23.310 156.120 23.600 156.165 ;
        RECT 23.755 156.120 24.075 156.180 ;
        RECT 23.310 155.980 24.075 156.120 ;
        RECT 23.310 155.935 23.600 155.980 ;
        RECT 23.755 155.920 24.075 155.980 ;
        RECT 25.595 156.120 25.915 156.180 ;
        RECT 31.205 156.120 31.345 156.320 ;
        RECT 36.750 156.275 37.040 156.320 ;
        RECT 39.990 156.275 40.640 156.320 ;
        RECT 42.630 156.460 42.920 156.505 ;
        RECT 43.075 156.460 43.395 156.520 ;
        RECT 42.630 156.320 43.395 156.460 ;
        RECT 46.385 156.460 46.525 156.660 ;
        RECT 46.755 156.600 47.075 156.660 ;
        RECT 47.215 156.600 47.535 156.860 ;
        RECT 47.765 156.845 47.905 157.000 ;
        RECT 50.525 157.000 52.595 157.140 ;
        RECT 47.690 156.615 47.980 156.845 ;
        RECT 48.610 156.800 48.900 156.845 ;
        RECT 49.055 156.800 49.375 156.860 ;
        RECT 48.610 156.660 49.375 156.800 ;
        RECT 48.610 156.615 48.900 156.660 ;
        RECT 49.055 156.600 49.375 156.660 ;
        RECT 49.975 156.600 50.295 156.860 ;
        RECT 50.525 156.845 50.665 157.000 ;
        RECT 52.275 156.940 52.595 157.000 ;
        RECT 53.195 157.140 53.515 157.200 ;
        RECT 53.670 157.140 53.960 157.185 ;
        RECT 57.795 157.140 58.115 157.200 ;
        RECT 63.775 157.140 64.095 157.200 ;
        RECT 66.165 157.185 66.305 157.340 ;
        RECT 67.545 157.340 75.045 157.480 ;
        RECT 77.545 157.480 77.835 157.525 ;
        RECT 80.325 157.480 80.615 157.525 ;
        RECT 82.185 157.480 82.475 157.525 ;
        RECT 96.435 157.480 96.755 157.540 ;
        RECT 77.545 157.340 82.475 157.480 ;
        RECT 53.195 157.000 53.960 157.140 ;
        RECT 53.195 156.940 53.515 157.000 ;
        RECT 53.670 156.955 53.960 157.000 ;
        RECT 55.125 157.000 58.115 157.140 ;
        RECT 50.450 156.615 50.740 156.845 ;
        RECT 50.910 156.800 51.200 156.845 ;
        RECT 54.575 156.800 54.895 156.860 ;
        RECT 55.125 156.845 55.265 157.000 ;
        RECT 57.795 156.940 58.115 157.000 ;
        RECT 60.185 157.000 64.095 157.140 ;
        RECT 50.910 156.660 54.895 156.800 ;
        RECT 50.910 156.615 51.200 156.660 ;
        RECT 50.985 156.460 51.125 156.615 ;
        RECT 54.575 156.600 54.895 156.660 ;
        RECT 55.050 156.615 55.340 156.845 ;
        RECT 57.335 156.600 57.655 156.860 ;
        RECT 46.385 156.320 51.125 156.460 ;
        RECT 57.885 156.460 58.025 156.940 ;
        RECT 60.185 156.845 60.325 157.000 ;
        RECT 63.775 156.940 64.095 157.000 ;
        RECT 66.090 156.955 66.380 157.185 ;
        RECT 60.110 156.615 60.400 156.845 ;
        RECT 65.170 156.800 65.460 156.845 ;
        RECT 67.545 156.800 67.685 157.340 ;
        RECT 77.545 157.295 77.835 157.340 ;
        RECT 80.325 157.295 80.615 157.340 ;
        RECT 82.185 157.295 82.475 157.340 ;
        RECT 92.845 157.340 96.755 157.480 ;
        RECT 75.735 157.140 76.055 157.200 ;
        RECT 72.145 157.000 76.055 157.140 ;
        RECT 65.170 156.660 67.685 156.800 ;
        RECT 65.170 156.615 65.460 156.660 ;
        RECT 62.870 156.460 63.160 156.505 ;
        RECT 65.245 156.460 65.385 156.615 ;
        RECT 67.915 156.600 68.235 156.860 ;
        RECT 69.755 156.800 70.075 156.860 ;
        RECT 71.150 156.800 71.440 156.845 ;
        RECT 69.755 156.660 71.440 156.800 ;
        RECT 69.755 156.600 70.075 156.660 ;
        RECT 71.150 156.615 71.440 156.660 ;
        RECT 71.595 156.600 71.915 156.860 ;
        RECT 72.145 156.845 72.285 157.000 ;
        RECT 75.735 156.940 76.055 157.000 ;
        RECT 78.035 157.140 78.355 157.200 ;
        RECT 80.810 157.140 81.100 157.185 ;
        RECT 78.035 157.000 81.100 157.140 ;
        RECT 78.035 156.940 78.355 157.000 ;
        RECT 80.810 156.955 81.100 157.000 ;
        RECT 88.155 157.140 88.475 157.200 ;
        RECT 88.155 157.000 90.685 157.140 ;
        RECT 88.155 156.940 88.475 157.000 ;
        RECT 72.070 156.615 72.360 156.845 ;
        RECT 72.975 156.600 73.295 156.860 ;
        RECT 77.545 156.800 77.835 156.845 ;
        RECT 77.545 156.660 80.080 156.800 ;
        RECT 77.545 156.615 77.835 156.660 ;
        RECT 75.685 156.460 75.975 156.505 ;
        RECT 78.035 156.460 78.355 156.520 ;
        RECT 79.865 156.505 80.080 156.660 ;
        RECT 82.635 156.600 82.955 156.860 ;
        RECT 88.630 156.800 88.920 156.845 ;
        RECT 89.995 156.800 90.315 156.860 ;
        RECT 90.545 156.845 90.685 157.000 ;
        RECT 88.630 156.660 90.315 156.800 ;
        RECT 88.630 156.615 88.920 156.660 ;
        RECT 89.995 156.600 90.315 156.660 ;
        RECT 90.470 156.615 90.760 156.845 ;
        RECT 90.915 156.600 91.235 156.860 ;
        RECT 91.375 156.600 91.695 156.860 ;
        RECT 92.310 156.800 92.600 156.845 ;
        RECT 92.845 156.800 92.985 157.340 ;
        RECT 96.435 157.280 96.755 157.340 ;
        RECT 98.735 157.480 99.055 157.540 ;
        RECT 98.735 157.340 99.885 157.480 ;
        RECT 98.735 157.280 99.055 157.340 ;
        RECT 95.515 157.140 95.835 157.200 ;
        RECT 97.355 157.140 97.675 157.200 ;
        RECT 94.685 157.000 98.965 157.140 ;
        RECT 92.310 156.660 92.985 156.800 ;
        RECT 92.310 156.615 92.600 156.660 ;
        RECT 93.215 156.600 93.535 156.860 ;
        RECT 93.675 156.800 93.995 156.860 ;
        RECT 94.685 156.845 94.825 157.000 ;
        RECT 95.515 156.940 95.835 157.000 ;
        RECT 97.355 156.940 97.675 157.000 ;
        RECT 94.150 156.800 94.440 156.845 ;
        RECT 93.675 156.660 94.440 156.800 ;
        RECT 93.675 156.600 93.995 156.660 ;
        RECT 94.150 156.615 94.440 156.660 ;
        RECT 94.610 156.615 94.900 156.845 ;
        RECT 95.055 156.800 95.375 156.860 ;
        RECT 98.825 156.845 98.965 157.000 ;
        RECT 98.290 156.800 98.580 156.845 ;
        RECT 95.055 156.660 98.580 156.800 ;
        RECT 95.055 156.600 95.375 156.660 ;
        RECT 98.290 156.615 98.580 156.660 ;
        RECT 98.750 156.615 99.040 156.845 ;
        RECT 99.195 156.600 99.515 156.860 ;
        RECT 99.745 156.800 99.885 157.340 ;
        RECT 103.795 156.940 104.115 157.200 ;
        RECT 100.130 156.800 100.420 156.845 ;
        RECT 99.745 156.660 100.420 156.800 ;
        RECT 100.130 156.615 100.420 156.660 ;
        RECT 102.415 156.800 102.735 156.860 ;
        RECT 105.190 156.800 105.480 156.845 ;
        RECT 102.415 156.660 105.480 156.800 ;
        RECT 102.415 156.600 102.735 156.660 ;
        RECT 105.190 156.615 105.480 156.660 ;
        RECT 78.945 156.460 79.235 156.505 ;
        RECT 57.885 156.320 65.385 156.460 ;
        RECT 68.925 156.320 75.505 156.460 ;
        RECT 42.630 156.275 42.920 156.320 ;
        RECT 43.075 156.260 43.395 156.320 ;
        RECT 62.870 156.275 63.160 156.320 ;
        RECT 25.595 155.980 31.345 156.120 ;
        RECT 25.595 155.920 25.915 155.980 ;
        RECT 35.255 155.920 35.575 156.180 ;
        RECT 44.915 156.120 45.235 156.180 ;
        RECT 45.390 156.120 45.680 156.165 ;
        RECT 44.915 155.980 45.680 156.120 ;
        RECT 44.915 155.920 45.235 155.980 ;
        RECT 45.390 155.935 45.680 155.980 ;
        RECT 52.275 155.920 52.595 156.180 ;
        RECT 57.795 155.920 58.115 156.180 ;
        RECT 59.175 155.920 59.495 156.180 ;
        RECT 60.095 156.120 60.415 156.180 ;
        RECT 68.925 156.165 69.065 156.320 ;
        RECT 68.850 156.120 69.140 156.165 ;
        RECT 60.095 155.980 69.140 156.120 ;
        RECT 60.095 155.920 60.415 155.980 ;
        RECT 68.850 155.935 69.140 155.980 ;
        RECT 69.755 155.920 70.075 156.180 ;
        RECT 75.365 156.120 75.505 156.320 ;
        RECT 75.685 156.320 79.235 156.460 ;
        RECT 75.685 156.275 75.975 156.320 ;
        RECT 78.035 156.260 78.355 156.320 ;
        RECT 78.945 156.275 79.235 156.320 ;
        RECT 79.865 156.460 80.155 156.505 ;
        RECT 81.725 156.460 82.015 156.505 ;
        RECT 96.910 156.460 97.200 156.505 ;
        RECT 79.865 156.320 82.015 156.460 ;
        RECT 79.865 156.275 80.155 156.320 ;
        RECT 81.725 156.275 82.015 156.320 ;
        RECT 91.465 156.320 97.200 156.460 ;
        RECT 91.465 156.180 91.605 156.320 ;
        RECT 96.910 156.275 97.200 156.320 ;
        RECT 84.475 156.120 84.795 156.180 ;
        RECT 75.365 155.980 84.795 156.120 ;
        RECT 84.475 155.920 84.795 155.980 ;
        RECT 84.935 156.120 85.255 156.180 ;
        RECT 89.090 156.120 89.380 156.165 ;
        RECT 84.935 155.980 89.380 156.120 ;
        RECT 84.935 155.920 85.255 155.980 ;
        RECT 89.090 155.935 89.380 155.980 ;
        RECT 91.375 155.920 91.695 156.180 ;
        RECT 93.215 156.120 93.535 156.180 ;
        RECT 95.515 156.120 95.835 156.180 ;
        RECT 93.215 155.980 95.835 156.120 ;
        RECT 93.215 155.920 93.535 155.980 ;
        RECT 95.515 155.920 95.835 155.980 ;
        RECT 96.450 156.120 96.740 156.165 ;
        RECT 97.355 156.120 97.675 156.180 ;
        RECT 96.450 155.980 97.675 156.120 ;
        RECT 96.450 155.935 96.740 155.980 ;
        RECT 97.355 155.920 97.675 155.980 ;
        RECT 17.370 155.300 112.465 155.780 ;
        RECT 27.895 155.100 28.215 155.160 ;
        RECT 29.275 155.100 29.595 155.160 ;
        RECT 27.895 154.960 29.595 155.100 ;
        RECT 27.895 154.900 28.215 154.960 ;
        RECT 29.275 154.900 29.595 154.960 ;
        RECT 34.335 154.900 34.655 155.160 ;
        RECT 42.170 155.100 42.460 155.145 ;
        RECT 43.075 155.100 43.395 155.160 ;
        RECT 42.170 154.960 43.395 155.100 ;
        RECT 42.170 154.915 42.460 154.960 ;
        RECT 43.075 154.900 43.395 154.960 ;
        RECT 66.535 155.100 66.855 155.160 ;
        RECT 87.235 155.100 87.555 155.160 ;
        RECT 95.055 155.100 95.375 155.160 ;
        RECT 66.535 154.960 69.065 155.100 ;
        RECT 66.535 154.900 66.855 154.960 ;
        RECT 21.010 154.760 21.300 154.805 ;
        RECT 21.915 154.760 22.235 154.820 ;
        RECT 21.010 154.620 22.235 154.760 ;
        RECT 21.010 154.575 21.300 154.620 ;
        RECT 21.915 154.560 22.235 154.620 ;
        RECT 23.310 154.760 23.600 154.805 ;
        RECT 25.595 154.760 25.915 154.820 ;
        RECT 23.310 154.620 25.915 154.760 ;
        RECT 23.310 154.575 23.600 154.620 ;
        RECT 25.595 154.560 25.915 154.620 ;
        RECT 27.450 154.760 27.740 154.805 ;
        RECT 29.750 154.760 30.040 154.805 ;
        RECT 27.450 154.620 30.040 154.760 ;
        RECT 27.450 154.575 27.740 154.620 ;
        RECT 29.750 154.575 30.040 154.620 ;
        RECT 40.790 154.760 41.080 154.805 ;
        RECT 42.615 154.760 42.935 154.820 ;
        RECT 47.215 154.760 47.535 154.820 ;
        RECT 57.795 154.805 58.115 154.820 ;
        RECT 40.790 154.620 42.935 154.760 ;
        RECT 40.790 154.575 41.080 154.620 ;
        RECT 42.615 154.560 42.935 154.620 ;
        RECT 45.465 154.620 47.535 154.760 ;
        RECT 21.470 154.420 21.760 154.465 ;
        RECT 22.835 154.420 23.155 154.480 ;
        RECT 21.470 154.280 23.155 154.420 ;
        RECT 21.470 154.235 21.760 154.280 ;
        RECT 20.995 154.080 21.315 154.140 ;
        RECT 21.545 154.080 21.685 154.235 ;
        RECT 22.835 154.220 23.155 154.280 ;
        RECT 24.690 154.420 24.980 154.465 ;
        RECT 35.255 154.420 35.575 154.480 ;
        RECT 24.690 154.280 35.575 154.420 ;
        RECT 24.690 154.235 24.980 154.280 ;
        RECT 35.255 154.220 35.575 154.280 ;
        RECT 39.395 154.420 39.715 154.480 ;
        RECT 41.250 154.420 41.540 154.465 ;
        RECT 39.395 154.280 41.540 154.420 ;
        RECT 39.395 154.220 39.715 154.280 ;
        RECT 41.250 154.235 41.540 154.280 ;
        RECT 43.995 154.220 44.315 154.480 ;
        RECT 45.465 154.465 45.605 154.620 ;
        RECT 47.215 154.560 47.535 154.620 ;
        RECT 57.745 154.760 58.115 154.805 ;
        RECT 61.005 154.760 61.295 154.805 ;
        RECT 57.745 154.620 61.295 154.760 ;
        RECT 57.745 154.575 58.115 154.620 ;
        RECT 61.005 154.575 61.295 154.620 ;
        RECT 61.925 154.760 62.215 154.805 ;
        RECT 63.785 154.760 64.075 154.805 ;
        RECT 68.375 154.760 68.695 154.820 ;
        RECT 61.925 154.620 64.075 154.760 ;
        RECT 61.925 154.575 62.215 154.620 ;
        RECT 63.785 154.575 64.075 154.620 ;
        RECT 66.660 154.620 68.695 154.760 ;
        RECT 57.795 154.560 58.115 154.575 ;
        RECT 44.930 154.235 45.220 154.465 ;
        RECT 45.390 154.235 45.680 154.465 ;
        RECT 45.850 154.420 46.140 154.465 ;
        RECT 46.755 154.420 47.075 154.480 ;
        RECT 52.735 154.420 53.055 154.480 ;
        RECT 45.850 154.280 47.075 154.420 ;
        RECT 45.850 154.235 46.140 154.280 ;
        RECT 20.995 153.940 21.685 154.080 ;
        RECT 26.975 154.080 27.295 154.140 ;
        RECT 28.370 154.080 28.660 154.125 ;
        RECT 26.975 153.940 28.660 154.080 ;
        RECT 20.995 153.880 21.315 153.940 ;
        RECT 26.975 153.880 27.295 153.940 ;
        RECT 28.370 153.895 28.660 153.940 ;
        RECT 31.575 154.080 31.895 154.140 ;
        RECT 45.005 154.080 45.145 154.235 ;
        RECT 46.755 154.220 47.075 154.280 ;
        RECT 47.305 154.280 53.055 154.420 ;
        RECT 47.305 154.140 47.445 154.280 ;
        RECT 52.735 154.220 53.055 154.280 ;
        RECT 59.605 154.420 59.895 154.465 ;
        RECT 61.925 154.420 62.140 154.575 ;
        RECT 66.030 154.530 66.320 154.575 ;
        RECT 59.605 154.280 62.140 154.420 ;
        RECT 62.395 154.420 62.715 154.480 ;
        RECT 65.705 154.420 66.320 154.530 ;
        RECT 66.660 154.465 66.800 154.620 ;
        RECT 68.375 154.560 68.695 154.620 ;
        RECT 62.395 154.390 66.320 154.420 ;
        RECT 62.395 154.280 65.845 154.390 ;
        RECT 66.030 154.345 66.320 154.390 ;
        RECT 59.605 154.235 59.895 154.280 ;
        RECT 62.395 154.220 62.715 154.280 ;
        RECT 66.550 154.235 66.840 154.465 ;
        RECT 67.455 154.220 67.775 154.480 ;
        RECT 68.925 154.465 69.065 154.960 ;
        RECT 87.235 154.960 95.375 155.100 ;
        RECT 87.235 154.900 87.555 154.960 ;
        RECT 78.035 154.760 78.355 154.820 ;
        RECT 78.510 154.760 78.800 154.805 ;
        RECT 74.445 154.620 77.805 154.760 ;
        RECT 67.930 154.420 68.220 154.465 ;
        RECT 68.850 154.420 69.140 154.465 ;
        RECT 67.930 154.280 69.140 154.420 ;
        RECT 67.930 154.235 68.220 154.280 ;
        RECT 68.850 154.235 69.140 154.280 ;
        RECT 31.575 153.940 45.145 154.080 ;
        RECT 46.295 154.080 46.615 154.140 ;
        RECT 47.215 154.080 47.535 154.140 ;
        RECT 46.295 153.940 47.535 154.080 ;
        RECT 31.575 153.880 31.895 153.940 ;
        RECT 46.295 153.880 46.615 153.940 ;
        RECT 47.215 153.880 47.535 153.940 ;
        RECT 62.855 153.880 63.175 154.140 ;
        RECT 64.695 153.880 65.015 154.140 ;
        RECT 66.075 154.080 66.395 154.140 ;
        RECT 74.445 154.080 74.585 154.620 ;
        RECT 74.830 154.420 75.120 154.465 ;
        RECT 75.275 154.420 75.595 154.480 ;
        RECT 74.830 154.280 75.595 154.420 ;
        RECT 74.830 154.235 75.120 154.280 ;
        RECT 75.275 154.220 75.595 154.280 ;
        RECT 66.075 153.940 74.585 154.080 ;
        RECT 77.665 154.080 77.805 154.620 ;
        RECT 78.035 154.620 78.800 154.760 ;
        RECT 78.035 154.560 78.355 154.620 ;
        RECT 78.510 154.575 78.800 154.620 ;
        RECT 85.395 154.760 85.715 154.820 ;
        RECT 93.215 154.760 93.535 154.820 ;
        RECT 85.395 154.620 90.685 154.760 ;
        RECT 85.395 154.560 85.715 154.620 ;
        RECT 78.955 154.220 79.275 154.480 ;
        RECT 87.235 154.420 87.555 154.480 ;
        RECT 90.545 154.465 90.685 154.620 ;
        RECT 91.465 154.620 93.535 154.760 ;
        RECT 91.465 154.465 91.605 154.620 ;
        RECT 93.215 154.560 93.535 154.620 ;
        RECT 93.765 154.465 93.905 154.960 ;
        RECT 95.055 154.900 95.375 154.960 ;
        RECT 95.975 154.760 96.295 154.820 ;
        RECT 103.810 154.760 104.100 154.805 ;
        RECT 94.685 154.620 96.295 154.760 ;
        RECT 94.685 154.465 94.825 154.620 ;
        RECT 95.975 154.560 96.295 154.620 ;
        RECT 101.355 154.620 104.100 154.760 ;
        RECT 89.550 154.420 89.840 154.465 ;
        RECT 87.235 154.280 89.840 154.420 ;
        RECT 87.235 154.220 87.555 154.280 ;
        RECT 89.550 154.235 89.840 154.280 ;
        RECT 90.010 154.235 90.300 154.465 ;
        RECT 90.470 154.235 90.760 154.465 ;
        RECT 91.390 154.235 91.680 154.465 ;
        RECT 93.690 154.235 93.980 154.465 ;
        RECT 94.150 154.235 94.440 154.465 ;
        RECT 94.610 154.235 94.900 154.465 ;
        RECT 82.635 154.080 82.955 154.140 ;
        RECT 77.665 153.940 82.955 154.080 ;
        RECT 66.075 153.880 66.395 153.940 ;
        RECT 82.635 153.880 82.955 153.940 ;
        RECT 84.475 154.080 84.795 154.140 ;
        RECT 90.085 154.080 90.225 154.235 ;
        RECT 93.215 154.080 93.535 154.140 ;
        RECT 94.225 154.080 94.365 154.235 ;
        RECT 95.515 154.220 95.835 154.480 ;
        RECT 101.355 154.420 101.495 154.620 ;
        RECT 103.810 154.575 104.100 154.620 ;
        RECT 96.065 154.280 101.495 154.420 ;
        RECT 84.475 153.940 94.365 154.080 ;
        RECT 84.475 153.880 84.795 153.940 ;
        RECT 93.215 153.880 93.535 153.940 ;
        RECT 38.475 153.740 38.795 153.800 ;
        RECT 43.995 153.740 44.315 153.800 ;
        RECT 59.605 153.740 59.895 153.785 ;
        RECT 62.385 153.740 62.675 153.785 ;
        RECT 64.245 153.740 64.535 153.785 ;
        RECT 90.455 153.740 90.775 153.800 ;
        RECT 96.065 153.740 96.205 154.280 ;
        RECT 102.415 154.220 102.735 154.480 ;
        RECT 105.650 154.235 105.940 154.465 ;
        RECT 98.735 154.080 99.055 154.140 ;
        RECT 105.725 154.080 105.865 154.235 ;
        RECT 98.735 153.940 105.865 154.080 ;
        RECT 98.735 153.880 99.055 153.940 ;
        RECT 38.475 153.600 56.645 153.740 ;
        RECT 38.475 153.540 38.795 153.600 ;
        RECT 43.995 153.540 44.315 153.600 ;
        RECT 31.575 153.200 31.895 153.460 ;
        RECT 47.230 153.400 47.520 153.445 ;
        RECT 48.595 153.400 48.915 153.460 ;
        RECT 47.230 153.260 48.915 153.400 ;
        RECT 47.230 153.215 47.520 153.260 ;
        RECT 48.595 153.200 48.915 153.260 ;
        RECT 55.035 153.400 55.355 153.460 ;
        RECT 55.740 153.400 56.030 153.445 ;
        RECT 55.035 153.260 56.030 153.400 ;
        RECT 56.505 153.400 56.645 153.600 ;
        RECT 59.605 153.600 64.535 153.740 ;
        RECT 59.605 153.555 59.895 153.600 ;
        RECT 62.385 153.555 62.675 153.600 ;
        RECT 64.245 153.555 64.535 153.600 ;
        RECT 64.785 153.600 69.985 153.740 ;
        RECT 64.785 153.400 64.925 153.600 ;
        RECT 56.505 153.260 64.925 153.400 ;
        RECT 66.075 153.400 66.395 153.460 ;
        RECT 67.915 153.400 68.235 153.460 ;
        RECT 69.845 153.445 69.985 153.600 ;
        RECT 90.455 153.600 96.205 153.740 ;
        RECT 90.455 153.540 90.775 153.600 ;
        RECT 66.075 153.260 68.235 153.400 ;
        RECT 55.035 153.200 55.355 153.260 ;
        RECT 55.740 153.215 56.030 153.260 ;
        RECT 66.075 153.200 66.395 153.260 ;
        RECT 67.915 153.200 68.235 153.260 ;
        RECT 69.770 153.400 70.060 153.445 ;
        RECT 70.215 153.400 70.535 153.460 ;
        RECT 69.770 153.260 70.535 153.400 ;
        RECT 69.770 153.215 70.060 153.260 ;
        RECT 70.215 153.200 70.535 153.260 ;
        RECT 76.210 153.400 76.500 153.445 ;
        RECT 82.635 153.400 82.955 153.460 ;
        RECT 76.210 153.260 82.955 153.400 ;
        RECT 76.210 153.215 76.500 153.260 ;
        RECT 82.635 153.200 82.955 153.260 ;
        RECT 88.170 153.400 88.460 153.445 ;
        RECT 90.915 153.400 91.235 153.460 ;
        RECT 88.170 153.260 91.235 153.400 ;
        RECT 88.170 153.215 88.460 153.260 ;
        RECT 90.915 153.200 91.235 153.260 ;
        RECT 92.310 153.400 92.600 153.445 ;
        RECT 93.215 153.400 93.535 153.460 ;
        RECT 92.310 153.260 93.535 153.400 ;
        RECT 92.310 153.215 92.600 153.260 ;
        RECT 93.215 153.200 93.535 153.260 ;
        RECT 106.555 153.200 106.875 153.460 ;
        RECT 18.165 152.580 112.465 153.060 ;
        RECT 26.515 152.380 26.835 152.440 ;
        RECT 31.115 152.380 31.435 152.440 ;
        RECT 31.590 152.380 31.880 152.425 ;
        RECT 26.515 152.240 30.885 152.380 ;
        RECT 26.515 152.180 26.835 152.240 ;
        RECT 22.950 152.040 23.240 152.085 ;
        RECT 26.070 152.040 26.360 152.085 ;
        RECT 27.960 152.040 28.250 152.085 ;
        RECT 22.950 151.900 28.250 152.040 ;
        RECT 30.745 152.040 30.885 152.240 ;
        RECT 31.115 152.240 31.880 152.380 ;
        RECT 31.115 152.180 31.435 152.240 ;
        RECT 31.590 152.195 31.880 152.240 ;
        RECT 34.350 152.380 34.640 152.425 ;
        RECT 35.255 152.380 35.575 152.440 ;
        RECT 34.350 152.240 35.575 152.380 ;
        RECT 34.350 152.195 34.640 152.240 ;
        RECT 35.255 152.180 35.575 152.240 ;
        RECT 43.995 152.180 44.315 152.440 ;
        RECT 45.375 152.380 45.695 152.440 ;
        RECT 45.850 152.380 46.140 152.425 ;
        RECT 45.375 152.240 46.140 152.380 ;
        RECT 45.375 152.180 45.695 152.240 ;
        RECT 45.850 152.195 46.140 152.240 ;
        RECT 48.135 152.180 48.455 152.440 ;
        RECT 57.335 152.380 57.655 152.440 ;
        RECT 62.870 152.380 63.160 152.425 ;
        RECT 57.335 152.240 97.125 152.380 ;
        RECT 57.335 152.180 57.655 152.240 ;
        RECT 62.870 152.195 63.160 152.240 ;
        RECT 43.090 152.040 43.380 152.085 ;
        RECT 49.975 152.040 50.295 152.100 ;
        RECT 63.775 152.040 64.095 152.100 ;
        RECT 74.355 152.040 74.675 152.100 ;
        RECT 95.515 152.040 95.835 152.100 ;
        RECT 30.745 151.900 43.380 152.040 ;
        RECT 22.950 151.855 23.240 151.900 ;
        RECT 26.070 151.855 26.360 151.900 ;
        RECT 27.960 151.855 28.250 151.900 ;
        RECT 43.090 151.855 43.380 151.900 ;
        RECT 43.625 151.900 50.295 152.040 ;
        RECT 28.815 151.700 29.135 151.760 ;
        RECT 33.415 151.700 33.735 151.760 ;
        RECT 28.815 151.560 33.735 151.700 ;
        RECT 28.815 151.500 29.135 151.560 ;
        RECT 33.415 151.500 33.735 151.560 ;
        RECT 33.890 151.700 34.180 151.745 ;
        RECT 35.270 151.700 35.560 151.745 ;
        RECT 33.890 151.560 35.560 151.700 ;
        RECT 33.890 151.515 34.180 151.560 ;
        RECT 35.270 151.515 35.560 151.560 ;
        RECT 35.715 151.700 36.035 151.760 ;
        RECT 35.715 151.560 37.785 151.700 ;
        RECT 35.715 151.500 36.035 151.560 ;
        RECT 20.535 151.020 20.855 151.080 ;
        RECT 21.870 151.065 22.160 151.380 ;
        RECT 22.950 151.360 23.240 151.405 ;
        RECT 26.530 151.360 26.820 151.405 ;
        RECT 28.365 151.360 28.655 151.405 ;
        RECT 22.950 151.220 28.655 151.360 ;
        RECT 22.950 151.175 23.240 151.220 ;
        RECT 26.530 151.175 26.820 151.220 ;
        RECT 28.365 151.175 28.655 151.220 ;
        RECT 30.195 151.160 30.515 151.420 ;
        RECT 30.670 151.360 30.960 151.405 ;
        RECT 31.575 151.360 31.895 151.420 ;
        RECT 30.670 151.220 31.895 151.360 ;
        RECT 30.670 151.175 30.960 151.220 ;
        RECT 31.575 151.160 31.895 151.220 ;
        RECT 32.955 151.160 33.275 151.420 ;
        RECT 36.650 151.175 36.940 151.405 ;
        RECT 21.570 151.020 22.160 151.065 ;
        RECT 24.810 151.020 25.460 151.065 ;
        RECT 20.535 150.880 25.460 151.020 ;
        RECT 20.535 150.820 20.855 150.880 ;
        RECT 21.570 150.835 21.860 150.880 ;
        RECT 24.810 150.835 25.460 150.880 ;
        RECT 27.450 150.835 27.740 151.065 ;
        RECT 20.075 150.480 20.395 150.740 ;
        RECT 27.525 150.680 27.665 150.835 ;
        RECT 34.335 150.820 34.655 151.080 ;
        RECT 36.725 151.020 36.865 151.175 ;
        RECT 37.095 151.160 37.415 151.420 ;
        RECT 37.645 151.405 37.785 151.560 ;
        RECT 37.570 151.175 37.860 151.405 ;
        RECT 38.475 151.160 38.795 151.420 ;
        RECT 38.015 151.020 38.335 151.080 ;
        RECT 43.625 151.020 43.765 151.900 ;
        RECT 49.975 151.840 50.295 151.900 ;
        RECT 50.985 151.900 57.565 152.040 ;
        RECT 44.915 151.500 45.235 151.760 ;
        RECT 45.835 151.500 46.155 151.760 ;
        RECT 47.675 151.500 47.995 151.760 ;
        RECT 48.610 151.700 48.900 151.745 ;
        RECT 50.985 151.700 51.125 151.900 ;
        RECT 48.225 151.560 48.900 151.700 ;
        RECT 44.010 151.360 44.300 151.405 ;
        RECT 45.925 151.360 46.065 151.500 ;
        RECT 44.010 151.220 46.065 151.360 ;
        RECT 44.010 151.175 44.300 151.220 ;
        RECT 46.755 151.160 47.075 151.420 ;
        RECT 36.725 150.880 43.765 151.020 ;
        RECT 45.390 151.020 45.680 151.065 ;
        RECT 45.835 151.020 46.155 151.080 ;
        RECT 48.225 151.065 48.365 151.560 ;
        RECT 48.610 151.515 48.900 151.560 ;
        RECT 50.525 151.560 51.125 151.700 ;
        RECT 52.735 151.700 53.055 151.760 ;
        RECT 53.210 151.700 53.500 151.745 ;
        RECT 55.495 151.700 55.815 151.760 ;
        RECT 52.735 151.560 55.815 151.700 ;
        RECT 49.975 151.160 50.295 151.420 ;
        RECT 50.525 151.405 50.665 151.560 ;
        RECT 52.735 151.500 53.055 151.560 ;
        RECT 53.210 151.515 53.500 151.560 ;
        RECT 55.495 151.500 55.815 151.560 ;
        RECT 50.450 151.175 50.740 151.405 ;
        RECT 45.390 150.880 46.155 151.020 ;
        RECT 29.290 150.680 29.580 150.725 ;
        RECT 27.525 150.540 29.580 150.680 ;
        RECT 29.290 150.495 29.580 150.540 ;
        RECT 32.035 150.480 32.355 150.740 ;
        RECT 32.495 150.680 32.815 150.740 ;
        RECT 36.725 150.680 36.865 150.880 ;
        RECT 38.015 150.820 38.335 150.880 ;
        RECT 45.390 150.835 45.680 150.880 ;
        RECT 45.835 150.820 46.155 150.880 ;
        RECT 48.150 150.835 48.440 151.065 ;
        RECT 50.525 151.020 50.665 151.175 ;
        RECT 50.895 151.160 51.215 151.420 ;
        RECT 51.830 151.360 52.120 151.405 ;
        RECT 54.575 151.360 54.895 151.420 ;
        RECT 56.890 151.360 57.180 151.405 ;
        RECT 51.830 151.220 54.895 151.360 ;
        RECT 51.830 151.175 52.120 151.220 ;
        RECT 54.575 151.160 54.895 151.220 ;
        RECT 55.125 151.220 57.180 151.360 ;
        RECT 57.425 151.360 57.565 151.900 ;
        RECT 63.775 151.900 69.065 152.040 ;
        RECT 63.775 151.840 64.095 151.900 ;
        RECT 66.995 151.700 67.315 151.760 ;
        RECT 62.945 151.560 67.315 151.700 ;
        RECT 61.950 151.360 62.240 151.405 ;
        RECT 62.395 151.360 62.715 151.420 ;
        RECT 57.425 151.220 61.705 151.360 ;
        RECT 48.685 150.880 50.665 151.020 ;
        RECT 32.495 150.540 36.865 150.680 ;
        RECT 37.095 150.680 37.415 150.740 ;
        RECT 48.685 150.680 48.825 150.880 ;
        RECT 55.125 150.740 55.265 151.220 ;
        RECT 56.890 151.175 57.180 151.220 ;
        RECT 61.565 151.080 61.705 151.220 ;
        RECT 61.950 151.220 62.715 151.360 ;
        RECT 61.950 151.175 62.240 151.220 ;
        RECT 62.395 151.160 62.715 151.220 ;
        RECT 61.475 151.020 61.795 151.080 ;
        RECT 62.945 151.020 63.085 151.560 ;
        RECT 66.995 151.500 67.315 151.560 ;
        RECT 63.775 151.160 64.095 151.420 ;
        RECT 65.615 151.160 65.935 151.420 ;
        RECT 66.535 151.405 66.855 151.420 ;
        RECT 66.535 151.360 66.875 151.405 ;
        RECT 66.375 151.220 66.875 151.360 ;
        RECT 66.535 151.175 66.875 151.220 ;
        RECT 66.535 151.160 66.855 151.175 ;
        RECT 68.375 151.160 68.695 151.420 ;
        RECT 68.925 151.360 69.065 151.900 ;
        RECT 74.355 151.900 78.265 152.040 ;
        RECT 74.355 151.840 74.675 151.900 ;
        RECT 73.985 151.560 77.805 151.700 ;
        RECT 72.055 151.360 72.375 151.420 ;
        RECT 73.985 151.405 74.125 151.560 ;
        RECT 73.910 151.360 74.200 151.405 ;
        RECT 68.925 151.220 74.200 151.360 ;
        RECT 72.055 151.160 72.375 151.220 ;
        RECT 73.910 151.175 74.200 151.220 ;
        RECT 74.355 151.160 74.675 151.420 ;
        RECT 74.815 151.160 75.135 151.420 ;
        RECT 77.665 151.405 77.805 151.560 ;
        RECT 78.125 151.405 78.265 151.900 ;
        RECT 92.385 151.900 95.835 152.040 ;
        RECT 81.715 151.700 82.035 151.760 ;
        RECT 78.585 151.560 82.035 151.700 ;
        RECT 78.585 151.405 78.725 151.560 ;
        RECT 81.715 151.500 82.035 151.560 ;
        RECT 82.635 151.500 82.955 151.760 ;
        RECT 75.750 151.175 76.040 151.405 ;
        RECT 77.590 151.175 77.880 151.405 ;
        RECT 78.050 151.175 78.340 151.405 ;
        RECT 78.510 151.175 78.800 151.405 ;
        RECT 79.430 151.175 79.720 151.405 ;
        RECT 79.875 151.360 80.195 151.420 ;
        RECT 80.810 151.360 81.100 151.405 ;
        RECT 87.710 151.360 88.000 151.405 ;
        RECT 79.875 151.220 81.100 151.360 ;
        RECT 61.475 150.880 63.085 151.020 ;
        RECT 70.215 151.020 70.535 151.080 ;
        RECT 75.825 151.020 75.965 151.175 ;
        RECT 77.115 151.020 77.435 151.080 ;
        RECT 79.505 151.020 79.645 151.175 ;
        RECT 79.875 151.160 80.195 151.220 ;
        RECT 80.810 151.175 81.100 151.220 ;
        RECT 85.945 151.220 88.000 151.360 ;
        RECT 70.215 150.880 79.645 151.020 ;
        RECT 81.715 151.020 82.035 151.080 ;
        RECT 84.030 151.020 84.320 151.065 ;
        RECT 81.715 150.880 84.320 151.020 ;
        RECT 61.475 150.820 61.795 150.880 ;
        RECT 70.215 150.820 70.535 150.880 ;
        RECT 77.115 150.820 77.435 150.880 ;
        RECT 81.715 150.820 82.035 150.880 ;
        RECT 84.030 150.835 84.320 150.880 ;
        RECT 37.095 150.540 48.825 150.680 ;
        RECT 49.055 150.680 49.375 150.740 ;
        RECT 53.670 150.680 53.960 150.725 ;
        RECT 49.055 150.540 53.960 150.680 ;
        RECT 32.495 150.480 32.815 150.540 ;
        RECT 37.095 150.480 37.415 150.540 ;
        RECT 49.055 150.480 49.375 150.540 ;
        RECT 53.670 150.495 53.960 150.540 ;
        RECT 54.130 150.680 54.420 150.725 ;
        RECT 55.035 150.680 55.355 150.740 ;
        RECT 54.130 150.540 55.355 150.680 ;
        RECT 54.130 150.495 54.420 150.540 ;
        RECT 55.035 150.480 55.355 150.540 ;
        RECT 55.970 150.680 56.260 150.725 ;
        RECT 58.715 150.680 59.035 150.740 ;
        RECT 55.970 150.540 59.035 150.680 ;
        RECT 55.970 150.495 56.260 150.540 ;
        RECT 58.715 150.480 59.035 150.540 ;
        RECT 60.110 150.680 60.400 150.725 ;
        RECT 63.775 150.680 64.095 150.740 ;
        RECT 60.110 150.540 64.095 150.680 ;
        RECT 60.110 150.495 60.400 150.540 ;
        RECT 63.775 150.480 64.095 150.540 ;
        RECT 67.470 150.680 67.760 150.725 ;
        RECT 67.915 150.680 68.235 150.740 ;
        RECT 67.470 150.540 68.235 150.680 ;
        RECT 67.470 150.495 67.760 150.540 ;
        RECT 67.915 150.480 68.235 150.540 ;
        RECT 68.375 150.680 68.695 150.740 ;
        RECT 69.310 150.680 69.600 150.725 ;
        RECT 68.375 150.540 69.600 150.680 ;
        RECT 68.375 150.480 68.695 150.540 ;
        RECT 69.310 150.495 69.600 150.540 ;
        RECT 72.515 150.480 72.835 150.740 ;
        RECT 72.975 150.680 73.295 150.740 ;
        RECT 76.210 150.680 76.500 150.725 ;
        RECT 72.975 150.540 76.500 150.680 ;
        RECT 72.975 150.480 73.295 150.540 ;
        RECT 76.210 150.495 76.500 150.540 ;
        RECT 81.255 150.480 81.575 150.740 ;
        RECT 83.555 150.480 83.875 150.740 ;
        RECT 85.945 150.725 86.085 151.220 ;
        RECT 87.710 151.175 88.000 151.220 ;
        RECT 91.850 151.360 92.140 151.405 ;
        RECT 92.385 151.360 92.525 151.900 ;
        RECT 95.515 151.840 95.835 151.900 ;
        RECT 94.135 151.700 94.455 151.760 ;
        RECT 92.845 151.560 94.455 151.700 ;
        RECT 92.845 151.405 92.985 151.560 ;
        RECT 94.135 151.500 94.455 151.560 ;
        RECT 91.850 151.220 92.525 151.360 ;
        RECT 91.850 151.175 92.140 151.220 ;
        RECT 92.770 151.175 93.060 151.405 ;
        RECT 93.230 151.175 93.520 151.405 ;
        RECT 93.690 151.360 93.980 151.405 ;
        RECT 95.055 151.360 95.375 151.420 ;
        RECT 93.690 151.220 95.375 151.360 ;
        RECT 93.690 151.175 93.980 151.220 ;
        RECT 93.305 151.020 93.445 151.175 ;
        RECT 95.055 151.160 95.375 151.220 ;
        RECT 96.435 151.360 96.755 151.420 ;
        RECT 96.985 151.405 97.125 152.240 ;
        RECT 103.910 152.040 104.200 152.085 ;
        RECT 107.030 152.040 107.320 152.085 ;
        RECT 108.920 152.040 109.210 152.085 ;
        RECT 103.910 151.900 109.210 152.040 ;
        RECT 103.910 151.855 104.200 151.900 ;
        RECT 107.030 151.855 107.320 151.900 ;
        RECT 108.920 151.855 109.210 151.900 ;
        RECT 103.335 151.700 103.655 151.760 ;
        RECT 101.355 151.560 103.655 151.700 ;
        RECT 96.910 151.360 97.200 151.405 ;
        RECT 96.435 151.220 97.200 151.360 ;
        RECT 96.435 151.160 96.755 151.220 ;
        RECT 96.910 151.175 97.200 151.220 ;
        RECT 97.370 151.175 97.660 151.405 ;
        RECT 97.830 151.175 98.120 151.405 ;
        RECT 98.275 151.360 98.595 151.420 ;
        RECT 98.750 151.360 99.040 151.405 ;
        RECT 98.275 151.220 99.040 151.360 ;
        RECT 94.135 151.020 94.455 151.080 ;
        RECT 96.525 151.020 96.665 151.160 ;
        RECT 93.305 150.880 93.905 151.020 ;
        RECT 93.765 150.740 93.905 150.880 ;
        RECT 94.135 150.880 96.665 151.020 ;
        RECT 94.135 150.820 94.455 150.880 ;
        RECT 85.870 150.495 86.160 150.725 ;
        RECT 87.695 150.680 88.015 150.740 ;
        RECT 88.630 150.680 88.920 150.725 ;
        RECT 87.695 150.540 88.920 150.680 ;
        RECT 87.695 150.480 88.015 150.540 ;
        RECT 88.630 150.495 88.920 150.540 ;
        RECT 93.675 150.480 93.995 150.740 ;
        RECT 95.055 150.480 95.375 150.740 ;
        RECT 95.515 150.480 95.835 150.740 ;
        RECT 97.445 150.680 97.585 151.175 ;
        RECT 97.905 151.020 98.045 151.175 ;
        RECT 98.275 151.160 98.595 151.220 ;
        RECT 98.750 151.175 99.040 151.220 ;
        RECT 99.670 151.360 99.960 151.405 ;
        RECT 101.355 151.360 101.495 151.560 ;
        RECT 103.335 151.500 103.655 151.560 ;
        RECT 106.555 151.700 106.875 151.760 ;
        RECT 108.410 151.700 108.700 151.745 ;
        RECT 106.555 151.560 108.700 151.700 ;
        RECT 106.555 151.500 106.875 151.560 ;
        RECT 108.410 151.515 108.700 151.560 ;
        RECT 99.670 151.220 101.495 151.360 ;
        RECT 99.670 151.175 99.960 151.220 ;
        RECT 102.830 151.065 103.120 151.380 ;
        RECT 103.910 151.360 104.200 151.405 ;
        RECT 107.490 151.360 107.780 151.405 ;
        RECT 109.325 151.360 109.615 151.405 ;
        RECT 103.910 151.220 109.615 151.360 ;
        RECT 103.910 151.175 104.200 151.220 ;
        RECT 107.490 151.175 107.780 151.220 ;
        RECT 109.325 151.175 109.615 151.220 ;
        RECT 109.790 151.175 110.080 151.405 ;
        RECT 100.130 151.020 100.420 151.065 ;
        RECT 102.530 151.020 103.120 151.065 ;
        RECT 105.770 151.020 106.420 151.065 ;
        RECT 97.905 150.880 99.425 151.020 ;
        RECT 99.285 150.740 99.425 150.880 ;
        RECT 100.130 150.880 106.420 151.020 ;
        RECT 100.130 150.835 100.420 150.880 ;
        RECT 102.530 150.835 102.820 150.880 ;
        RECT 105.770 150.835 106.420 150.880 ;
        RECT 108.855 151.020 109.175 151.080 ;
        RECT 109.865 151.020 110.005 151.175 ;
        RECT 110.695 151.020 111.015 151.080 ;
        RECT 108.855 150.880 111.015 151.020 ;
        RECT 108.855 150.820 109.175 150.880 ;
        RECT 110.695 150.820 111.015 150.880 ;
        RECT 97.815 150.680 98.135 150.740 ;
        RECT 97.445 150.540 98.135 150.680 ;
        RECT 97.815 150.480 98.135 150.540 ;
        RECT 99.195 150.680 99.515 150.740 ;
        RECT 101.050 150.680 101.340 150.725 ;
        RECT 99.195 150.540 101.340 150.680 ;
        RECT 99.195 150.480 99.515 150.540 ;
        RECT 101.050 150.495 101.340 150.540 ;
        RECT 17.370 149.860 112.465 150.340 ;
        RECT 27.450 149.660 27.740 149.705 ;
        RECT 30.195 149.660 30.515 149.720 ;
        RECT 27.450 149.520 30.515 149.660 ;
        RECT 27.450 149.475 27.740 149.520 ;
        RECT 30.195 149.460 30.515 149.520 ;
        RECT 34.335 149.660 34.655 149.720 ;
        RECT 36.190 149.660 36.480 149.705 ;
        RECT 34.335 149.520 36.480 149.660 ;
        RECT 34.335 149.460 34.655 149.520 ;
        RECT 36.190 149.475 36.480 149.520 ;
        RECT 38.475 149.460 38.795 149.720 ;
        RECT 40.315 149.660 40.635 149.720 ;
        RECT 48.610 149.660 48.900 149.705 ;
        RECT 49.055 149.660 49.375 149.720 ;
        RECT 40.315 149.520 49.375 149.660 ;
        RECT 40.315 149.460 40.635 149.520 ;
        RECT 48.610 149.475 48.900 149.520 ;
        RECT 49.055 149.460 49.375 149.520 ;
        RECT 49.605 149.520 55.725 149.660 ;
        RECT 20.075 149.320 20.395 149.380 ;
        RECT 23.755 149.320 24.075 149.380 ;
        RECT 25.150 149.320 25.440 149.365 ;
        RECT 38.565 149.320 38.705 149.460 ;
        RECT 20.075 149.180 34.105 149.320 ;
        RECT 20.075 149.120 20.395 149.180 ;
        RECT 23.755 149.120 24.075 149.180 ;
        RECT 25.150 149.135 25.440 149.180 ;
        RECT 25.595 148.780 25.915 149.040 ;
        RECT 31.115 148.780 31.435 149.040 ;
        RECT 32.495 148.980 32.815 149.040 ;
        RECT 33.965 149.025 34.105 149.180 ;
        RECT 34.885 149.180 38.705 149.320 ;
        RECT 38.935 149.320 39.255 149.380 ;
        RECT 46.755 149.320 47.075 149.380 ;
        RECT 49.605 149.320 49.745 149.520 ;
        RECT 38.935 149.180 46.065 149.320 ;
        RECT 34.885 149.025 35.025 149.180 ;
        RECT 38.935 149.120 39.255 149.180 ;
        RECT 32.970 148.980 33.260 149.025 ;
        RECT 32.495 148.840 33.260 148.980 ;
        RECT 32.495 148.780 32.815 148.840 ;
        RECT 32.970 148.795 33.260 148.840 ;
        RECT 33.430 148.795 33.720 149.025 ;
        RECT 33.890 148.795 34.180 149.025 ;
        RECT 34.810 148.795 35.100 149.025 ;
        RECT 24.690 148.640 24.980 148.685 ;
        RECT 26.975 148.640 27.295 148.700 ;
        RECT 33.505 148.640 33.645 148.795 ;
        RECT 37.555 148.780 37.875 149.040 ;
        RECT 38.030 148.795 38.320 149.025 ;
        RECT 38.490 148.795 38.780 149.025 ;
        RECT 39.410 148.980 39.700 149.025 ;
        RECT 39.855 148.980 40.175 149.040 ;
        RECT 39.410 148.840 40.175 148.980 ;
        RECT 39.410 148.795 39.700 148.840 ;
        RECT 37.095 148.640 37.415 148.700 ;
        RECT 24.690 148.500 27.295 148.640 ;
        RECT 24.690 148.455 24.980 148.500 ;
        RECT 26.975 148.440 27.295 148.500 ;
        RECT 32.585 148.500 37.415 148.640 ;
        RECT 32.585 148.360 32.725 148.500 ;
        RECT 37.095 148.440 37.415 148.500 ;
        RECT 31.590 148.300 31.880 148.345 ;
        RECT 32.035 148.300 32.355 148.360 ;
        RECT 31.590 148.160 32.355 148.300 ;
        RECT 31.590 148.115 31.880 148.160 ;
        RECT 32.035 148.100 32.355 148.160 ;
        RECT 32.495 148.100 32.815 148.360 ;
        RECT 38.105 148.300 38.245 148.795 ;
        RECT 38.565 148.640 38.705 148.795 ;
        RECT 39.855 148.780 40.175 148.840 ;
        RECT 40.315 148.780 40.635 149.040 ;
        RECT 43.090 148.980 43.380 149.025 ;
        RECT 45.390 148.980 45.680 149.025 ;
        RECT 43.090 148.840 45.680 148.980 ;
        RECT 43.090 148.795 43.380 148.840 ;
        RECT 45.390 148.795 45.680 148.840 ;
        RECT 40.405 148.640 40.545 148.780 ;
        RECT 38.565 148.500 40.545 148.640 ;
        RECT 44.470 148.455 44.760 148.685 ;
        RECT 39.395 148.300 39.715 148.360 ;
        RECT 38.105 148.160 39.715 148.300 ;
        RECT 39.395 148.100 39.715 148.160 ;
        RECT 30.670 147.960 30.960 148.005 ;
        RECT 38.935 147.960 39.255 148.020 ;
        RECT 30.670 147.820 39.255 147.960 ;
        RECT 44.545 147.960 44.685 148.455 ;
        RECT 44.915 148.440 45.235 148.700 ;
        RECT 45.925 148.640 46.065 149.180 ;
        RECT 46.755 149.180 49.745 149.320 ;
        RECT 50.090 149.320 50.380 149.365 ;
        RECT 50.895 149.320 51.215 149.380 ;
        RECT 53.330 149.320 53.980 149.365 ;
        RECT 50.090 149.180 53.980 149.320 ;
        RECT 55.585 149.320 55.725 149.520 ;
        RECT 62.855 149.460 63.175 149.720 ;
        RECT 63.775 149.660 64.095 149.720 ;
        RECT 74.355 149.660 74.675 149.720 ;
        RECT 87.695 149.660 88.015 149.720 ;
        RECT 93.675 149.660 93.995 149.720 ;
        RECT 96.910 149.660 97.200 149.705 ;
        RECT 63.775 149.520 65.385 149.660 ;
        RECT 63.775 149.460 64.095 149.520 ;
        RECT 59.190 149.320 59.480 149.365 ;
        RECT 55.585 149.180 64.005 149.320 ;
        RECT 46.755 149.120 47.075 149.180 ;
        RECT 50.090 149.135 50.680 149.180 ;
        RECT 50.390 148.820 50.680 149.135 ;
        RECT 50.895 149.120 51.215 149.180 ;
        RECT 53.330 149.135 53.980 149.180 ;
        RECT 59.190 149.135 59.480 149.180 ;
        RECT 51.470 148.980 51.760 149.025 ;
        RECT 55.050 148.980 55.340 149.025 ;
        RECT 56.885 148.980 57.175 149.025 ;
        RECT 51.470 148.840 57.175 148.980 ;
        RECT 51.470 148.795 51.760 148.840 ;
        RECT 55.050 148.795 55.340 148.840 ;
        RECT 56.885 148.795 57.175 148.840 ;
        RECT 58.715 148.780 59.035 149.040 ;
        RECT 60.570 148.995 60.860 149.025 ;
        RECT 60.185 148.855 60.860 148.995 ;
        RECT 57.350 148.640 57.640 148.685 ;
        RECT 45.925 148.500 57.640 148.640 ;
        RECT 57.350 148.455 57.640 148.500 ;
        RECT 57.795 148.640 58.115 148.700 ;
        RECT 60.185 148.640 60.325 148.855 ;
        RECT 60.570 148.795 60.860 148.855 ;
        RECT 61.030 148.795 61.320 149.025 ;
        RECT 57.795 148.500 60.325 148.640 ;
        RECT 57.795 148.440 58.115 148.500 ;
        RECT 51.470 148.300 51.760 148.345 ;
        RECT 54.590 148.300 54.880 148.345 ;
        RECT 56.480 148.300 56.770 148.345 ;
        RECT 46.845 148.160 51.125 148.300 ;
        RECT 44.915 147.960 45.235 148.020 ;
        RECT 46.845 147.960 46.985 148.160 ;
        RECT 44.545 147.820 46.985 147.960 ;
        RECT 47.230 147.960 47.520 148.005 ;
        RECT 49.975 147.960 50.295 148.020 ;
        RECT 47.230 147.820 50.295 147.960 ;
        RECT 50.985 147.960 51.125 148.160 ;
        RECT 51.470 148.160 56.770 148.300 ;
        RECT 51.470 148.115 51.760 148.160 ;
        RECT 54.590 148.115 54.880 148.160 ;
        RECT 56.480 148.115 56.770 148.160 ;
        RECT 58.255 148.300 58.575 148.360 ;
        RECT 61.105 148.300 61.245 148.795 ;
        RECT 61.475 148.780 61.795 149.040 ;
        RECT 61.935 148.980 62.255 149.040 ;
        RECT 63.865 149.025 64.005 149.180 ;
        RECT 64.695 149.120 65.015 149.380 ;
        RECT 62.410 148.980 62.700 149.025 ;
        RECT 61.935 148.840 62.700 148.980 ;
        RECT 61.935 148.780 62.255 148.840 ;
        RECT 62.410 148.795 62.700 148.840 ;
        RECT 63.790 148.795 64.080 149.025 ;
        RECT 64.250 148.795 64.540 149.025 ;
        RECT 65.245 148.980 65.385 149.520 ;
        RECT 71.225 149.520 75.965 149.660 ;
        RECT 66.995 149.320 67.315 149.380 ;
        RECT 71.225 149.320 71.365 149.520 ;
        RECT 74.355 149.460 74.675 149.520 ;
        RECT 66.995 149.180 71.365 149.320 ;
        RECT 66.995 149.120 67.315 149.180 ;
        RECT 65.630 148.980 65.920 149.025 ;
        RECT 65.245 148.840 65.920 148.980 ;
        RECT 65.630 148.795 65.920 148.840 ;
        RECT 66.090 148.980 66.380 149.025 ;
        RECT 66.535 148.980 66.855 149.040 ;
        RECT 66.090 148.840 66.855 148.980 ;
        RECT 66.090 148.795 66.380 148.840 ;
        RECT 64.325 148.640 64.465 148.795 ;
        RECT 66.535 148.780 66.855 148.840 ;
        RECT 67.455 148.980 67.775 149.040 ;
        RECT 67.930 148.980 68.220 149.025 ;
        RECT 67.455 148.840 68.220 148.980 ;
        RECT 67.455 148.780 67.775 148.840 ;
        RECT 67.930 148.795 68.220 148.840 ;
        RECT 69.770 148.980 70.060 149.025 ;
        RECT 70.215 148.980 70.535 149.040 ;
        RECT 69.770 148.840 70.535 148.980 ;
        RECT 69.770 148.795 70.060 148.840 ;
        RECT 70.215 148.780 70.535 148.840 ;
        RECT 70.675 148.780 70.995 149.040 ;
        RECT 71.225 149.025 71.365 149.180 ;
        RECT 72.145 149.180 75.505 149.320 ;
        RECT 72.145 149.040 72.285 149.180 ;
        RECT 71.150 148.795 71.440 149.025 ;
        RECT 71.610 148.980 71.900 149.025 ;
        RECT 72.055 148.980 72.375 149.040 ;
        RECT 73.895 148.980 74.215 149.040 ;
        RECT 75.365 149.025 75.505 149.180 ;
        RECT 75.825 149.025 75.965 149.520 ;
        RECT 87.695 149.520 89.765 149.660 ;
        RECT 87.695 149.460 88.015 149.520 ;
        RECT 78.495 149.320 78.815 149.380 ;
        RECT 76.285 149.180 78.815 149.320 ;
        RECT 76.285 149.025 76.425 149.180 ;
        RECT 78.495 149.120 78.815 149.180 ;
        RECT 81.255 149.320 81.575 149.380 ;
        RECT 89.625 149.365 89.765 149.520 ;
        RECT 92.385 149.520 97.200 149.660 ;
        RECT 83.670 149.320 83.960 149.365 ;
        RECT 86.910 149.320 87.560 149.365 ;
        RECT 81.255 149.180 87.560 149.320 ;
        RECT 81.255 149.120 81.575 149.180 ;
        RECT 83.670 149.135 84.260 149.180 ;
        RECT 86.910 149.135 87.560 149.180 ;
        RECT 89.550 149.135 89.840 149.365 ;
        RECT 89.995 149.320 90.315 149.380 ;
        RECT 89.995 149.180 91.145 149.320 ;
        RECT 71.610 148.840 72.375 148.980 ;
        RECT 71.610 148.795 71.900 148.840 ;
        RECT 72.055 148.780 72.375 148.840 ;
        RECT 72.605 148.840 74.215 148.980 ;
        RECT 72.605 148.640 72.745 148.840 ;
        RECT 73.895 148.780 74.215 148.840 ;
        RECT 75.290 148.795 75.580 149.025 ;
        RECT 75.750 148.795 76.040 149.025 ;
        RECT 76.210 148.795 76.500 149.025 ;
        RECT 77.115 148.780 77.435 149.040 ;
        RECT 83.970 148.820 84.260 149.135 ;
        RECT 89.995 149.120 90.315 149.180 ;
        RECT 91.005 149.025 91.145 149.180 ;
        RECT 92.385 149.025 92.525 149.520 ;
        RECT 93.675 149.460 93.995 149.520 ;
        RECT 96.910 149.475 97.200 149.520 ;
        RECT 98.735 149.460 99.055 149.720 ;
        RECT 96.450 149.320 96.740 149.365 ;
        RECT 99.195 149.320 99.515 149.380 ;
        RECT 96.450 149.180 99.515 149.320 ;
        RECT 96.450 149.135 96.740 149.180 ;
        RECT 99.195 149.120 99.515 149.180 ;
        RECT 103.745 149.320 104.035 149.365 ;
        RECT 105.175 149.320 105.495 149.380 ;
        RECT 107.005 149.320 107.295 149.365 ;
        RECT 103.745 149.180 107.295 149.320 ;
        RECT 103.745 149.135 104.035 149.180 ;
        RECT 105.175 149.120 105.495 149.180 ;
        RECT 107.005 149.135 107.295 149.180 ;
        RECT 107.925 149.320 108.215 149.365 ;
        RECT 109.785 149.320 110.075 149.365 ;
        RECT 107.925 149.180 110.075 149.320 ;
        RECT 107.925 149.135 108.215 149.180 ;
        RECT 109.785 149.135 110.075 149.180 ;
        RECT 85.050 148.980 85.340 149.025 ;
        RECT 88.630 148.980 88.920 149.025 ;
        RECT 90.465 148.980 90.755 149.025 ;
        RECT 85.050 148.840 90.755 148.980 ;
        RECT 85.050 148.795 85.340 148.840 ;
        RECT 88.630 148.795 88.920 148.840 ;
        RECT 90.465 148.795 90.755 148.840 ;
        RECT 90.930 148.795 91.220 149.025 ;
        RECT 91.390 148.795 91.680 149.025 ;
        RECT 92.310 148.795 92.600 149.025 ;
        RECT 92.770 148.795 93.060 149.025 ;
        RECT 93.230 148.995 93.520 149.025 ;
        RECT 94.135 149.010 94.455 149.040 ;
        RECT 93.765 148.995 94.455 149.010 ;
        RECT 93.230 148.870 94.455 148.995 ;
        RECT 97.815 148.980 98.135 149.040 ;
        RECT 93.230 148.855 93.905 148.870 ;
        RECT 93.230 148.795 93.520 148.855 ;
        RECT 64.325 148.500 66.765 148.640 ;
        RECT 66.625 148.360 66.765 148.500 ;
        RECT 67.085 148.500 72.745 148.640 ;
        RECT 72.990 148.640 73.280 148.685 ;
        RECT 73.435 148.640 73.755 148.700 ;
        RECT 72.990 148.500 73.755 148.640 ;
        RECT 58.255 148.160 61.705 148.300 ;
        RECT 58.255 148.100 58.575 148.160 ;
        RECT 52.735 147.960 53.055 148.020 ;
        RECT 50.985 147.820 53.055 147.960 ;
        RECT 30.670 147.775 30.960 147.820 ;
        RECT 38.935 147.760 39.255 147.820 ;
        RECT 44.915 147.760 45.235 147.820 ;
        RECT 47.230 147.775 47.520 147.820 ;
        RECT 49.975 147.760 50.295 147.820 ;
        RECT 52.735 147.760 53.055 147.820 ;
        RECT 56.065 147.960 56.355 148.005 ;
        RECT 57.810 147.960 58.100 148.005 ;
        RECT 56.065 147.820 58.100 147.960 ;
        RECT 61.565 147.960 61.705 148.160 ;
        RECT 66.535 148.100 66.855 148.360 ;
        RECT 67.085 148.345 67.225 148.500 ;
        RECT 72.990 148.455 73.280 148.500 ;
        RECT 73.435 148.440 73.755 148.500 ;
        RECT 82.190 148.640 82.480 148.685 ;
        RECT 83.555 148.640 83.875 148.700 ;
        RECT 91.465 148.640 91.605 148.795 ;
        RECT 82.190 148.500 83.875 148.640 ;
        RECT 82.190 148.455 82.480 148.500 ;
        RECT 83.555 148.440 83.875 148.500 ;
        RECT 91.060 148.500 91.605 148.640 ;
        RECT 92.845 148.640 92.985 148.795 ;
        RECT 94.135 148.780 94.455 148.870 ;
        RECT 94.685 148.840 98.135 148.980 ;
        RECT 94.685 148.640 94.825 148.840 ;
        RECT 97.815 148.780 98.135 148.840 ;
        RECT 105.605 148.980 105.895 149.025 ;
        RECT 107.925 148.980 108.140 149.135 ;
        RECT 105.605 148.840 108.140 148.980 ;
        RECT 105.605 148.795 105.895 148.840 ;
        RECT 110.695 148.780 111.015 149.040 ;
        RECT 92.845 148.500 94.825 148.640 ;
        RECT 95.990 148.640 96.280 148.685 ;
        RECT 95.990 148.500 101.495 148.640 ;
        RECT 67.010 148.115 67.300 148.345 ;
        RECT 67.455 148.100 67.775 148.360 ;
        RECT 72.055 148.300 72.375 148.360 ;
        RECT 73.910 148.300 74.200 148.345 ;
        RECT 72.055 148.160 74.200 148.300 ;
        RECT 72.055 148.100 72.375 148.160 ;
        RECT 73.910 148.115 74.200 148.160 ;
        RECT 85.050 148.300 85.340 148.345 ;
        RECT 88.170 148.300 88.460 148.345 ;
        RECT 90.060 148.300 90.350 148.345 ;
        RECT 91.060 148.300 91.200 148.500 ;
        RECT 95.990 148.455 96.280 148.500 ;
        RECT 94.135 148.300 94.455 148.360 ;
        RECT 94.610 148.300 94.900 148.345 ;
        RECT 85.050 148.160 90.350 148.300 ;
        RECT 85.050 148.115 85.340 148.160 ;
        RECT 88.170 148.115 88.460 148.160 ;
        RECT 90.060 148.115 90.350 148.160 ;
        RECT 90.545 148.160 93.905 148.300 ;
        RECT 67.545 147.960 67.685 148.100 ;
        RECT 61.565 147.820 67.685 147.960 ;
        RECT 68.850 147.960 69.140 148.005 ;
        RECT 74.815 147.960 75.135 148.020 ;
        RECT 68.850 147.820 75.135 147.960 ;
        RECT 56.065 147.775 56.355 147.820 ;
        RECT 57.810 147.775 58.100 147.820 ;
        RECT 68.850 147.775 69.140 147.820 ;
        RECT 74.815 147.760 75.135 147.820 ;
        RECT 86.775 147.960 87.095 148.020 ;
        RECT 90.545 147.960 90.685 148.160 ;
        RECT 86.775 147.820 90.685 147.960 ;
        RECT 93.765 147.960 93.905 148.160 ;
        RECT 94.135 148.160 94.900 148.300 ;
        RECT 101.355 148.300 101.495 148.500 ;
        RECT 108.855 148.440 109.175 148.700 ;
        RECT 105.605 148.300 105.895 148.345 ;
        RECT 108.385 148.300 108.675 148.345 ;
        RECT 110.245 148.300 110.535 148.345 ;
        RECT 101.355 148.160 102.645 148.300 ;
        RECT 94.135 148.100 94.455 148.160 ;
        RECT 94.610 148.115 94.900 148.160 ;
        RECT 102.505 148.020 102.645 148.160 ;
        RECT 105.605 148.160 110.535 148.300 ;
        RECT 105.605 148.115 105.895 148.160 ;
        RECT 108.385 148.115 108.675 148.160 ;
        RECT 110.245 148.115 110.535 148.160 ;
        RECT 98.275 147.960 98.595 148.020 ;
        RECT 101.955 148.005 102.275 148.020 ;
        RECT 93.765 147.820 98.595 147.960 ;
        RECT 86.775 147.760 87.095 147.820 ;
        RECT 98.275 147.760 98.595 147.820 ;
        RECT 101.740 147.775 102.275 148.005 ;
        RECT 101.955 147.760 102.275 147.775 ;
        RECT 102.415 147.760 102.735 148.020 ;
        RECT 18.165 147.140 112.465 147.620 ;
        RECT 19.630 146.940 19.920 146.985 ;
        RECT 25.135 146.940 25.455 147.000 ;
        RECT 31.575 146.940 31.895 147.000 ;
        RECT 38.475 146.940 38.795 147.000 ;
        RECT 19.630 146.800 31.895 146.940 ;
        RECT 19.630 146.755 19.920 146.800 ;
        RECT 25.135 146.740 25.455 146.800 ;
        RECT 31.575 146.740 31.895 146.800 ;
        RECT 32.125 146.800 38.795 146.940 ;
        RECT 22.490 146.600 22.780 146.645 ;
        RECT 25.610 146.600 25.900 146.645 ;
        RECT 27.500 146.600 27.790 146.645 ;
        RECT 22.490 146.460 27.790 146.600 ;
        RECT 22.490 146.415 22.780 146.460 ;
        RECT 25.610 146.415 25.900 146.460 ;
        RECT 27.500 146.415 27.790 146.460 ;
        RECT 28.815 146.400 29.135 146.660 ;
        RECT 28.370 146.260 28.660 146.305 ;
        RECT 28.905 146.260 29.045 146.400 ;
        RECT 32.125 146.260 32.265 146.800 ;
        RECT 38.475 146.740 38.795 146.800 ;
        RECT 45.835 146.940 46.155 147.000 ;
        RECT 50.895 146.940 51.215 147.000 ;
        RECT 51.370 146.940 51.660 146.985 ;
        RECT 45.835 146.800 49.745 146.940 ;
        RECT 45.835 146.740 46.155 146.800 ;
        RECT 34.335 146.600 34.655 146.660 ;
        RECT 38.015 146.600 38.335 146.660 ;
        RECT 33.505 146.460 38.335 146.600 ;
        RECT 33.505 146.260 33.645 146.460 ;
        RECT 34.335 146.400 34.655 146.460 ;
        RECT 28.370 146.120 29.045 146.260 ;
        RECT 31.205 146.120 32.265 146.260 ;
        RECT 33.045 146.120 33.645 146.260 ;
        RECT 28.370 146.075 28.660 146.120 ;
        RECT 31.205 145.980 31.345 146.120 ;
        RECT 20.535 145.580 20.855 145.640 ;
        RECT 21.410 145.625 21.700 145.940 ;
        RECT 22.490 145.920 22.780 145.965 ;
        RECT 26.070 145.920 26.360 145.965 ;
        RECT 27.905 145.920 28.195 145.965 ;
        RECT 28.830 145.920 29.120 145.965 ;
        RECT 22.490 145.780 28.195 145.920 ;
        RECT 22.490 145.735 22.780 145.780 ;
        RECT 26.070 145.735 26.360 145.780 ;
        RECT 27.905 145.735 28.195 145.780 ;
        RECT 28.445 145.780 29.120 145.920 ;
        RECT 28.445 145.640 28.585 145.780 ;
        RECT 28.830 145.735 29.120 145.780 ;
        RECT 31.115 145.720 31.435 145.980 ;
        RECT 31.575 145.920 31.895 145.980 ;
        RECT 32.050 145.920 32.340 145.965 ;
        RECT 31.575 145.780 32.340 145.920 ;
        RECT 31.575 145.720 31.895 145.780 ;
        RECT 32.050 145.735 32.340 145.780 ;
        RECT 32.495 145.720 32.815 145.980 ;
        RECT 33.045 145.965 33.185 146.120 ;
        RECT 36.725 145.965 36.865 146.460 ;
        RECT 38.015 146.400 38.335 146.460 ;
        RECT 43.505 146.600 43.795 146.645 ;
        RECT 46.285 146.600 46.575 146.645 ;
        RECT 48.145 146.600 48.435 146.645 ;
        RECT 43.505 146.460 48.435 146.600 ;
        RECT 43.505 146.415 43.795 146.460 ;
        RECT 46.285 146.415 46.575 146.460 ;
        RECT 48.145 146.415 48.435 146.460 ;
        RECT 49.070 146.415 49.360 146.645 ;
        RECT 49.605 146.600 49.745 146.800 ;
        RECT 50.895 146.800 51.660 146.940 ;
        RECT 50.895 146.740 51.215 146.800 ;
        RECT 51.370 146.755 51.660 146.800 ;
        RECT 54.575 146.940 54.895 147.000 ;
        RECT 55.955 146.940 56.275 147.000 ;
        RECT 67.915 146.940 68.235 147.000 ;
        RECT 54.575 146.800 68.235 146.940 ;
        RECT 54.575 146.740 54.895 146.800 ;
        RECT 55.955 146.740 56.275 146.800 ;
        RECT 67.915 146.740 68.235 146.800 ;
        RECT 70.675 146.940 70.995 147.000 ;
        RECT 71.150 146.940 71.440 146.985 ;
        RECT 76.900 146.940 77.190 146.985 ;
        RECT 81.715 146.940 82.035 147.000 ;
        RECT 70.675 146.800 71.440 146.940 ;
        RECT 70.675 146.740 70.995 146.800 ;
        RECT 71.150 146.755 71.440 146.800 ;
        RECT 75.365 146.800 82.035 146.940 ;
        RECT 52.750 146.600 53.040 146.645 ;
        RECT 58.255 146.600 58.575 146.660 ;
        RECT 49.605 146.460 53.040 146.600 ;
        RECT 52.750 146.415 53.040 146.460 ;
        RECT 54.665 146.460 58.575 146.600 ;
        RECT 39.640 146.260 39.930 146.305 ;
        RECT 45.375 146.260 45.695 146.320 ;
        RECT 39.640 146.120 45.695 146.260 ;
        RECT 39.640 146.075 39.930 146.120 ;
        RECT 45.375 146.060 45.695 146.120 ;
        RECT 46.770 146.260 47.060 146.305 ;
        RECT 49.145 146.260 49.285 146.415 ;
        RECT 46.770 146.120 49.285 146.260 ;
        RECT 46.770 146.075 47.060 146.120 ;
        RECT 32.970 145.735 33.260 145.965 ;
        RECT 33.505 145.780 35.945 145.920 ;
        RECT 21.110 145.580 21.700 145.625 ;
        RECT 24.350 145.580 25.000 145.625 ;
        RECT 20.535 145.440 25.000 145.580 ;
        RECT 20.535 145.380 20.855 145.440 ;
        RECT 21.110 145.395 21.400 145.440 ;
        RECT 24.350 145.395 25.000 145.440 ;
        RECT 26.990 145.395 27.280 145.625 ;
        RECT 21.915 145.240 22.235 145.300 ;
        RECT 27.065 145.240 27.205 145.395 ;
        RECT 28.355 145.380 28.675 145.640 ;
        RECT 33.505 145.580 33.645 145.780 ;
        RECT 29.365 145.440 33.645 145.580 ;
        RECT 34.350 145.580 34.640 145.625 ;
        RECT 34.795 145.580 35.115 145.640 ;
        RECT 34.350 145.440 35.115 145.580 ;
        RECT 21.915 145.100 27.205 145.240 ;
        RECT 27.895 145.240 28.215 145.300 ;
        RECT 29.365 145.240 29.505 145.440 ;
        RECT 34.350 145.395 34.640 145.440 ;
        RECT 34.795 145.380 35.115 145.440 ;
        RECT 27.895 145.100 29.505 145.240 ;
        RECT 21.915 145.040 22.235 145.100 ;
        RECT 27.895 145.040 28.215 145.100 ;
        RECT 29.735 145.040 30.055 145.300 ;
        RECT 33.875 145.240 34.195 145.300 ;
        RECT 35.270 145.240 35.560 145.285 ;
        RECT 33.875 145.100 35.560 145.240 ;
        RECT 35.805 145.240 35.945 145.780 ;
        RECT 36.650 145.735 36.940 145.965 ;
        RECT 37.095 145.720 37.415 145.980 ;
        RECT 37.570 145.735 37.860 145.965 ;
        RECT 37.645 145.240 37.785 145.735 ;
        RECT 38.475 145.720 38.795 145.980 ;
        RECT 43.505 145.920 43.795 145.965 ;
        RECT 46.295 145.920 46.615 145.980 ;
        RECT 48.610 145.920 48.900 145.965 ;
        RECT 43.505 145.780 46.040 145.920 ;
        RECT 43.505 145.735 43.795 145.780 ;
        RECT 38.935 145.580 39.255 145.640 ;
        RECT 45.825 145.625 46.040 145.780 ;
        RECT 46.295 145.780 48.900 145.920 ;
        RECT 46.295 145.720 46.615 145.780 ;
        RECT 48.610 145.735 48.900 145.780 ;
        RECT 49.975 145.720 50.295 145.980 ;
        RECT 54.665 145.965 54.805 146.460 ;
        RECT 58.255 146.400 58.575 146.460 ;
        RECT 60.110 146.415 60.400 146.645 ;
        RECT 64.250 146.600 64.540 146.645 ;
        RECT 64.250 146.460 74.585 146.600 ;
        RECT 64.250 146.415 64.540 146.460 ;
        RECT 55.495 146.260 55.815 146.320 ;
        RECT 56.890 146.260 57.180 146.305 ;
        RECT 55.495 146.120 57.180 146.260 ;
        RECT 60.185 146.260 60.325 146.415 ;
        RECT 60.185 146.120 66.765 146.260 ;
        RECT 55.495 146.060 55.815 146.120 ;
        RECT 56.890 146.075 57.180 146.120 ;
        RECT 50.910 145.735 51.200 145.965 ;
        RECT 54.130 145.735 54.420 145.965 ;
        RECT 54.590 145.735 54.880 145.965 ;
        RECT 41.645 145.580 41.935 145.625 ;
        RECT 44.905 145.580 45.195 145.625 ;
        RECT 38.935 145.440 45.195 145.580 ;
        RECT 38.935 145.380 39.255 145.440 ;
        RECT 41.645 145.395 41.935 145.440 ;
        RECT 44.905 145.395 45.195 145.440 ;
        RECT 45.825 145.580 46.115 145.625 ;
        RECT 47.685 145.580 47.975 145.625 ;
        RECT 45.825 145.440 47.975 145.580 ;
        RECT 45.825 145.395 46.115 145.440 ;
        RECT 47.685 145.395 47.975 145.440 ;
        RECT 49.515 145.580 49.835 145.640 ;
        RECT 50.985 145.580 51.125 145.735 ;
        RECT 49.515 145.440 51.125 145.580 ;
        RECT 54.205 145.580 54.345 145.735 ;
        RECT 55.035 145.720 55.355 145.980 ;
        RECT 55.955 145.720 56.275 145.980 ;
        RECT 61.015 145.920 61.335 145.980 ;
        RECT 62.395 145.920 62.715 145.980 ;
        RECT 66.625 145.965 66.765 146.120 ;
        RECT 72.055 146.060 72.375 146.320 ;
        RECT 74.445 145.980 74.585 146.460 ;
        RECT 63.330 145.920 63.620 145.965 ;
        RECT 61.015 145.780 62.165 145.920 ;
        RECT 61.015 145.720 61.335 145.780 ;
        RECT 57.335 145.580 57.655 145.640 ;
        RECT 54.205 145.440 57.655 145.580 ;
        RECT 49.515 145.380 49.835 145.440 ;
        RECT 57.335 145.380 57.655 145.440 ;
        RECT 57.810 145.580 58.100 145.625 ;
        RECT 61.475 145.580 61.795 145.640 ;
        RECT 57.810 145.440 61.795 145.580 ;
        RECT 62.025 145.580 62.165 145.780 ;
        RECT 62.395 145.780 63.620 145.920 ;
        RECT 62.395 145.720 62.715 145.780 ;
        RECT 63.330 145.735 63.620 145.780 ;
        RECT 66.090 145.735 66.380 145.965 ;
        RECT 66.550 145.735 66.840 145.965 ;
        RECT 68.835 145.920 69.155 145.980 ;
        RECT 71.150 145.920 71.440 145.965 ;
        RECT 68.835 145.780 71.440 145.920 ;
        RECT 66.165 145.580 66.305 145.735 ;
        RECT 68.835 145.720 69.155 145.780 ;
        RECT 71.150 145.735 71.440 145.780 ;
        RECT 74.355 145.720 74.675 145.980 ;
        RECT 74.815 145.720 75.135 145.980 ;
        RECT 75.365 145.965 75.505 146.800 ;
        RECT 76.900 146.755 77.190 146.800 ;
        RECT 81.715 146.740 82.035 146.800 ;
        RECT 93.675 146.740 93.995 147.000 ;
        RECT 95.975 146.740 96.295 147.000 ;
        RECT 105.175 146.740 105.495 147.000 ;
        RECT 107.490 146.940 107.780 146.985 ;
        RECT 108.855 146.940 109.175 147.000 ;
        RECT 107.490 146.800 109.175 146.940 ;
        RECT 107.490 146.755 107.780 146.800 ;
        RECT 108.855 146.740 109.175 146.800 ;
        RECT 80.765 146.600 81.055 146.645 ;
        RECT 83.545 146.600 83.835 146.645 ;
        RECT 85.405 146.600 85.695 146.645 ;
        RECT 102.415 146.600 102.735 146.660 ;
        RECT 80.765 146.460 85.695 146.600 ;
        RECT 80.765 146.415 81.055 146.460 ;
        RECT 83.545 146.415 83.835 146.460 ;
        RECT 85.405 146.415 85.695 146.460 ;
        RECT 101.585 146.460 102.735 146.600 ;
        RECT 93.215 146.060 93.535 146.320 ;
        RECT 95.055 146.060 95.375 146.320 ;
        RECT 101.585 146.305 101.725 146.460 ;
        RECT 102.415 146.400 102.735 146.460 ;
        RECT 104.270 146.415 104.560 146.645 ;
        RECT 101.510 146.075 101.800 146.305 ;
        RECT 101.955 146.060 102.275 146.320 ;
        RECT 104.345 146.260 104.485 146.415 ;
        RECT 104.345 146.120 106.785 146.260 ;
        RECT 75.290 145.735 75.580 145.965 ;
        RECT 76.210 145.735 76.500 145.965 ;
        RECT 80.765 145.920 81.055 145.965 ;
        RECT 80.765 145.780 83.300 145.920 ;
        RECT 80.765 145.735 81.055 145.780 ;
        RECT 62.025 145.440 66.305 145.580 ;
        RECT 57.810 145.395 58.100 145.440 ;
        RECT 61.475 145.380 61.795 145.440 ;
        RECT 35.805 145.100 37.785 145.240 ;
        RECT 58.270 145.240 58.560 145.285 ;
        RECT 58.715 145.240 59.035 145.300 ;
        RECT 58.270 145.100 59.035 145.240 ;
        RECT 33.875 145.040 34.195 145.100 ;
        RECT 35.270 145.055 35.560 145.100 ;
        RECT 58.270 145.055 58.560 145.100 ;
        RECT 58.715 145.040 59.035 145.100 ;
        RECT 63.775 145.240 64.095 145.300 ;
        RECT 65.630 145.240 65.920 145.285 ;
        RECT 63.775 145.100 65.920 145.240 ;
        RECT 66.165 145.240 66.305 145.440 ;
        RECT 72.530 145.580 72.820 145.625 ;
        RECT 72.990 145.580 73.280 145.625 ;
        RECT 72.530 145.440 73.280 145.580 ;
        RECT 72.530 145.395 72.820 145.440 ;
        RECT 72.990 145.395 73.280 145.440 ;
        RECT 73.895 145.580 74.215 145.640 ;
        RECT 75.735 145.580 76.055 145.640 ;
        RECT 76.285 145.580 76.425 145.735 ;
        RECT 83.085 145.625 83.300 145.780 ;
        RECT 84.015 145.720 84.335 145.980 ;
        RECT 85.855 145.720 86.175 145.980 ;
        RECT 87.695 145.920 88.015 145.980 ;
        RECT 90.455 145.920 90.775 145.980 ;
        RECT 87.695 145.780 90.775 145.920 ;
        RECT 87.695 145.720 88.015 145.780 ;
        RECT 90.455 145.720 90.775 145.780 ;
        RECT 92.755 145.720 93.075 145.980 ;
        RECT 94.135 145.720 94.455 145.980 ;
        RECT 94.610 145.920 94.900 145.965 ;
        RECT 95.515 145.920 95.835 145.980 ;
        RECT 94.610 145.780 95.835 145.920 ;
        RECT 94.610 145.735 94.900 145.780 ;
        RECT 95.515 145.720 95.835 145.780 ;
        RECT 95.990 145.920 96.280 145.965 ;
        RECT 96.895 145.920 97.215 145.980 ;
        RECT 95.990 145.780 97.215 145.920 ;
        RECT 95.990 145.735 96.280 145.780 ;
        RECT 96.895 145.720 97.215 145.780 ;
        RECT 99.195 145.920 99.515 145.980 ;
        RECT 102.430 145.920 102.720 145.965 ;
        RECT 99.195 145.780 102.720 145.920 ;
        RECT 99.195 145.720 99.515 145.780 ;
        RECT 102.430 145.735 102.720 145.780 ;
        RECT 103.795 145.920 104.115 145.980 ;
        RECT 106.645 145.965 106.785 146.120 ;
        RECT 104.730 145.920 105.020 145.965 ;
        RECT 103.795 145.780 105.020 145.920 ;
        RECT 103.795 145.720 104.115 145.780 ;
        RECT 104.730 145.735 105.020 145.780 ;
        RECT 106.570 145.735 106.860 145.965 ;
        RECT 73.895 145.440 76.425 145.580 ;
        RECT 78.905 145.580 79.195 145.625 ;
        RECT 82.165 145.580 82.455 145.625 ;
        RECT 83.085 145.580 83.375 145.625 ;
        RECT 84.945 145.580 85.235 145.625 ;
        RECT 107.475 145.580 107.795 145.640 ;
        RECT 78.905 145.440 82.865 145.580 ;
        RECT 73.895 145.380 74.215 145.440 ;
        RECT 75.735 145.380 76.055 145.440 ;
        RECT 78.905 145.395 79.195 145.440 ;
        RECT 82.165 145.395 82.455 145.440 ;
        RECT 66.535 145.240 66.855 145.300 ;
        RECT 66.165 145.100 66.855 145.240 ;
        RECT 63.775 145.040 64.095 145.100 ;
        RECT 65.630 145.055 65.920 145.100 ;
        RECT 66.535 145.040 66.855 145.100 ;
        RECT 67.470 145.240 67.760 145.285 ;
        RECT 68.835 145.240 69.155 145.300 ;
        RECT 67.470 145.100 69.155 145.240 ;
        RECT 67.470 145.055 67.760 145.100 ;
        RECT 68.835 145.040 69.155 145.100 ;
        RECT 70.215 145.040 70.535 145.300 ;
        RECT 82.725 145.240 82.865 145.440 ;
        RECT 83.085 145.440 85.235 145.580 ;
        RECT 83.085 145.395 83.375 145.440 ;
        RECT 84.945 145.395 85.235 145.440 ;
        RECT 91.925 145.440 107.795 145.580 ;
        RECT 91.925 145.285 92.065 145.440 ;
        RECT 107.475 145.380 107.795 145.440 ;
        RECT 87.250 145.240 87.540 145.285 ;
        RECT 82.725 145.100 87.540 145.240 ;
        RECT 87.250 145.055 87.540 145.100 ;
        RECT 91.850 145.055 92.140 145.285 ;
        RECT 96.910 145.240 97.200 145.285 ;
        RECT 105.635 145.240 105.955 145.300 ;
        RECT 96.910 145.100 105.955 145.240 ;
        RECT 96.910 145.055 97.200 145.100 ;
        RECT 105.635 145.040 105.955 145.100 ;
        RECT 17.370 144.420 112.465 144.900 ;
        RECT 21.455 144.020 21.775 144.280 ;
        RECT 32.495 144.020 32.815 144.280 ;
        RECT 45.375 144.020 45.695 144.280 ;
        RECT 61.475 144.265 61.795 144.280 ;
        RECT 61.475 144.035 62.010 144.265 ;
        RECT 80.810 144.220 81.100 144.265 ;
        RECT 81.715 144.220 82.035 144.280 ;
        RECT 80.810 144.080 82.035 144.220 ;
        RECT 80.810 144.035 81.100 144.080 ;
        RECT 61.475 144.020 61.795 144.035 ;
        RECT 81.715 144.020 82.035 144.080 ;
        RECT 84.015 144.220 84.335 144.280 ;
        RECT 84.490 144.220 84.780 144.265 ;
        RECT 97.815 144.220 98.135 144.280 ;
        RECT 84.015 144.080 84.780 144.220 ;
        RECT 84.015 144.020 84.335 144.080 ;
        RECT 84.490 144.035 84.780 144.080 ;
        RECT 97.445 144.080 98.135 144.220 ;
        RECT 21.915 143.880 22.235 143.940 ;
        RECT 23.870 143.880 24.160 143.925 ;
        RECT 27.110 143.880 27.760 143.925 ;
        RECT 21.915 143.740 27.760 143.880 ;
        RECT 21.915 143.680 22.235 143.740 ;
        RECT 23.870 143.695 24.460 143.740 ;
        RECT 27.110 143.695 27.760 143.740 ;
        RECT 20.550 143.540 20.840 143.585 ;
        RECT 22.835 143.540 23.155 143.600 ;
        RECT 20.550 143.400 23.155 143.540 ;
        RECT 20.550 143.355 20.840 143.400 ;
        RECT 22.835 143.340 23.155 143.400 ;
        RECT 24.170 143.380 24.460 143.695 ;
        RECT 29.735 143.680 30.055 143.940 ;
        RECT 31.115 143.680 31.435 143.940 ;
        RECT 32.585 143.880 32.725 144.020 ;
        RECT 45.465 143.880 45.605 144.020 ;
        RECT 63.775 143.925 64.095 143.940 ;
        RECT 32.585 143.740 34.105 143.880 ;
        RECT 25.250 143.540 25.540 143.585 ;
        RECT 28.830 143.540 29.120 143.585 ;
        RECT 30.665 143.540 30.955 143.585 ;
        RECT 25.250 143.400 30.955 143.540 ;
        RECT 31.205 143.540 31.345 143.680 ;
        RECT 33.965 143.585 34.105 143.740 ;
        RECT 39.945 143.740 45.605 143.880 ;
        RECT 63.725 143.880 64.095 143.925 ;
        RECT 66.985 143.880 67.275 143.925 ;
        RECT 63.725 143.740 67.275 143.880 ;
        RECT 32.510 143.540 32.800 143.585 ;
        RECT 31.205 143.400 32.800 143.540 ;
        RECT 25.250 143.355 25.540 143.400 ;
        RECT 28.830 143.355 29.120 143.400 ;
        RECT 30.665 143.355 30.955 143.400 ;
        RECT 32.510 143.355 32.800 143.400 ;
        RECT 33.430 143.355 33.720 143.585 ;
        RECT 33.890 143.355 34.180 143.585 ;
        RECT 29.275 143.200 29.595 143.260 ;
        RECT 31.130 143.200 31.420 143.245 ;
        RECT 29.275 143.060 31.420 143.200 ;
        RECT 29.275 143.000 29.595 143.060 ;
        RECT 31.130 143.015 31.420 143.060 ;
        RECT 31.575 143.200 31.895 143.260 ;
        RECT 33.505 143.200 33.645 143.355 ;
        RECT 34.335 143.340 34.655 143.600 ;
        RECT 37.555 143.540 37.875 143.600 ;
        RECT 38.935 143.540 39.255 143.600 ;
        RECT 37.555 143.400 39.255 143.540 ;
        RECT 37.555 143.340 37.875 143.400 ;
        RECT 38.935 143.340 39.255 143.400 ;
        RECT 39.395 143.340 39.715 143.600 ;
        RECT 39.945 143.585 40.085 143.740 ;
        RECT 63.725 143.695 64.095 143.740 ;
        RECT 66.985 143.695 67.275 143.740 ;
        RECT 67.905 143.880 68.195 143.925 ;
        RECT 69.765 143.880 70.055 143.925 ;
        RECT 67.905 143.740 70.055 143.880 ;
        RECT 67.905 143.695 68.195 143.740 ;
        RECT 69.765 143.695 70.055 143.740 ;
        RECT 95.070 143.880 95.360 143.925 ;
        RECT 95.530 143.880 95.820 143.925 ;
        RECT 95.070 143.740 95.820 143.880 ;
        RECT 95.070 143.695 95.360 143.740 ;
        RECT 95.530 143.695 95.820 143.740 ;
        RECT 63.775 143.680 64.095 143.695 ;
        RECT 39.870 143.355 40.160 143.585 ;
        RECT 40.315 143.540 40.635 143.600 ;
        RECT 40.790 143.540 41.080 143.585 ;
        RECT 40.315 143.400 41.080 143.540 ;
        RECT 40.315 143.340 40.635 143.400 ;
        RECT 40.790 143.355 41.080 143.400 ;
        RECT 61.015 143.340 61.335 143.600 ;
        RECT 65.585 143.540 65.875 143.585 ;
        RECT 67.905 143.540 68.120 143.695 ;
        RECT 65.585 143.400 68.120 143.540 ;
        RECT 65.585 143.355 65.875 143.400 ;
        RECT 68.835 143.340 69.155 143.600 ;
        RECT 79.875 143.540 80.195 143.600 ;
        RECT 81.270 143.540 81.560 143.585 ;
        RECT 85.410 143.540 85.700 143.585 ;
        RECT 79.875 143.400 81.560 143.540 ;
        RECT 79.875 143.340 80.195 143.400 ;
        RECT 81.270 143.355 81.560 143.400 ;
        RECT 83.185 143.400 85.700 143.540 ;
        RECT 31.575 143.060 33.645 143.200 ;
        RECT 43.075 143.200 43.395 143.260 ;
        RECT 45.850 143.200 46.140 143.245 ;
        RECT 43.075 143.060 46.140 143.200 ;
        RECT 31.575 143.000 31.895 143.060 ;
        RECT 43.075 143.000 43.395 143.060 ;
        RECT 45.850 143.015 46.140 143.060 ;
        RECT 46.310 143.015 46.600 143.245 ;
        RECT 70.690 143.200 70.980 143.245 ;
        RECT 71.135 143.200 71.455 143.260 ;
        RECT 70.690 143.060 71.455 143.200 ;
        RECT 70.690 143.015 70.980 143.060 ;
        RECT 25.250 142.860 25.540 142.905 ;
        RECT 28.370 142.860 28.660 142.905 ;
        RECT 30.260 142.860 30.550 142.905 ;
        RECT 25.250 142.720 30.550 142.860 ;
        RECT 25.250 142.675 25.540 142.720 ;
        RECT 28.370 142.675 28.660 142.720 ;
        RECT 30.260 142.675 30.550 142.720 ;
        RECT 35.715 142.660 36.035 142.920 ;
        RECT 45.375 142.860 45.695 142.920 ;
        RECT 46.385 142.860 46.525 143.015 ;
        RECT 71.135 143.000 71.455 143.060 ;
        RECT 80.350 143.200 80.640 143.245 ;
        RECT 82.635 143.200 82.955 143.260 ;
        RECT 80.350 143.060 82.955 143.200 ;
        RECT 80.350 143.015 80.640 143.060 ;
        RECT 82.635 143.000 82.955 143.060 ;
        RECT 45.375 142.720 46.525 142.860 ;
        RECT 45.375 142.660 45.695 142.720 ;
        RECT 54.575 142.660 54.895 142.920 ;
        RECT 83.185 142.905 83.325 143.400 ;
        RECT 85.410 143.355 85.700 143.400 ;
        RECT 92.295 143.540 92.615 143.600 ;
        RECT 93.690 143.540 93.980 143.585 ;
        RECT 92.295 143.400 93.980 143.540 ;
        RECT 92.295 143.340 92.615 143.400 ;
        RECT 93.690 143.355 93.980 143.400 ;
        RECT 96.435 143.540 96.755 143.600 ;
        RECT 97.445 143.585 97.585 144.080 ;
        RECT 97.815 144.020 98.135 144.080 ;
        RECT 99.195 143.880 99.515 143.940 ;
        RECT 97.905 143.740 101.495 143.880 ;
        RECT 97.905 143.585 98.045 143.740 ;
        RECT 99.195 143.680 99.515 143.740 ;
        RECT 96.910 143.540 97.200 143.585 ;
        RECT 96.435 143.400 97.200 143.540 ;
        RECT 96.435 143.340 96.755 143.400 ;
        RECT 96.910 143.355 97.200 143.400 ;
        RECT 97.370 143.355 97.660 143.585 ;
        RECT 97.830 143.355 98.120 143.585 ;
        RECT 98.275 143.540 98.595 143.600 ;
        RECT 98.750 143.540 99.040 143.585 ;
        RECT 98.275 143.400 99.040 143.540 ;
        RECT 101.355 143.540 101.495 143.740 ;
        RECT 101.955 143.540 102.275 143.600 ;
        RECT 101.355 143.400 102.275 143.540 ;
        RECT 94.595 143.000 94.915 143.260 ;
        RECT 95.515 143.200 95.835 143.260 ;
        RECT 97.445 143.200 97.585 143.355 ;
        RECT 98.275 143.340 98.595 143.400 ;
        RECT 98.750 143.355 99.040 143.400 ;
        RECT 101.955 143.340 102.275 143.400 ;
        RECT 103.795 143.540 104.115 143.600 ;
        RECT 105.190 143.540 105.480 143.585 ;
        RECT 103.795 143.400 105.480 143.540 ;
        RECT 103.795 143.340 104.115 143.400 ;
        RECT 105.190 143.355 105.480 143.400 ;
        RECT 106.555 143.340 106.875 143.600 ;
        RECT 95.515 143.060 97.585 143.200 ;
        RECT 95.515 143.000 95.835 143.060 ;
        RECT 65.585 142.860 65.875 142.905 ;
        RECT 68.365 142.860 68.655 142.905 ;
        RECT 70.225 142.860 70.515 142.905 ;
        RECT 65.585 142.720 70.515 142.860 ;
        RECT 65.585 142.675 65.875 142.720 ;
        RECT 68.365 142.675 68.655 142.720 ;
        RECT 70.225 142.675 70.515 142.720 ;
        RECT 83.110 142.675 83.400 142.905 ;
        RECT 92.770 142.860 93.060 142.905 ;
        RECT 98.735 142.860 99.055 142.920 ;
        RECT 92.770 142.720 99.055 142.860 ;
        RECT 92.770 142.675 93.060 142.720 ;
        RECT 98.735 142.660 99.055 142.720 ;
        RECT 22.375 142.320 22.695 142.580 ;
        RECT 34.335 142.520 34.655 142.580 ;
        RECT 37.570 142.520 37.860 142.565 ;
        RECT 34.335 142.380 37.860 142.520 ;
        RECT 34.335 142.320 34.655 142.380 ;
        RECT 37.570 142.335 37.860 142.380 ;
        RECT 43.535 142.320 43.855 142.580 ;
        RECT 44.915 142.520 45.235 142.580 ;
        RECT 47.215 142.520 47.535 142.580 ;
        RECT 49.515 142.520 49.835 142.580 ;
        RECT 44.915 142.380 49.835 142.520 ;
        RECT 44.915 142.320 45.235 142.380 ;
        RECT 47.215 142.320 47.535 142.380 ;
        RECT 49.515 142.320 49.835 142.380 ;
        RECT 95.070 142.520 95.360 142.565 ;
        RECT 97.815 142.520 98.135 142.580 ;
        RECT 95.070 142.380 98.135 142.520 ;
        RECT 95.070 142.335 95.360 142.380 ;
        RECT 97.815 142.320 98.135 142.380 ;
        RECT 105.650 142.520 105.940 142.565 ;
        RECT 106.095 142.520 106.415 142.580 ;
        RECT 105.650 142.380 106.415 142.520 ;
        RECT 105.650 142.335 105.940 142.380 ;
        RECT 106.095 142.320 106.415 142.380 ;
        RECT 107.490 142.520 107.780 142.565 ;
        RECT 108.855 142.520 109.175 142.580 ;
        RECT 107.490 142.380 109.175 142.520 ;
        RECT 107.490 142.335 107.780 142.380 ;
        RECT 108.855 142.320 109.175 142.380 ;
        RECT 18.165 141.700 112.465 142.180 ;
        RECT 21.915 141.300 22.235 141.560 ;
        RECT 22.835 141.300 23.155 141.560 ;
        RECT 28.355 141.500 28.675 141.560 ;
        RECT 30.670 141.500 30.960 141.545 ;
        RECT 28.355 141.360 30.960 141.500 ;
        RECT 28.355 141.300 28.675 141.360 ;
        RECT 30.670 141.315 30.960 141.360 ;
        RECT 33.415 141.300 33.735 141.560 ;
        RECT 51.355 141.500 51.675 141.560 ;
        RECT 51.830 141.500 52.120 141.545 ;
        RECT 51.355 141.360 52.120 141.500 ;
        RECT 51.355 141.300 51.675 141.360 ;
        RECT 51.830 141.315 52.120 141.360 ;
        RECT 82.635 141.500 82.955 141.560 ;
        RECT 89.995 141.500 90.315 141.560 ;
        RECT 82.635 141.360 90.315 141.500 ;
        RECT 82.635 141.300 82.955 141.360 ;
        RECT 89.995 141.300 90.315 141.360 ;
        RECT 92.755 141.300 93.075 141.560 ;
        RECT 96.435 141.500 96.755 141.560 ;
        RECT 95.145 141.360 96.755 141.500 ;
        RECT 20.535 140.960 20.855 141.220 ;
        RECT 31.115 141.160 31.435 141.220 ;
        RECT 45.345 141.160 45.635 141.205 ;
        RECT 48.125 141.160 48.415 141.205 ;
        RECT 49.985 141.160 50.275 141.205 ;
        RECT 31.115 141.020 38.245 141.160 ;
        RECT 31.115 140.960 31.435 141.020 ;
        RECT 25.135 140.620 25.455 140.880 ;
        RECT 26.070 140.820 26.360 140.865 ;
        RECT 26.975 140.820 27.295 140.880 ;
        RECT 27.450 140.820 27.740 140.865 ;
        RECT 26.070 140.680 27.740 140.820 ;
        RECT 26.070 140.635 26.360 140.680 ;
        RECT 26.975 140.620 27.295 140.680 ;
        RECT 27.450 140.635 27.740 140.680 ;
        RECT 28.370 140.820 28.660 140.865 ;
        RECT 31.575 140.820 31.895 140.880 ;
        RECT 28.370 140.680 31.895 140.820 ;
        RECT 28.370 140.635 28.660 140.680 ;
        RECT 20.995 140.480 21.315 140.540 ;
        RECT 21.470 140.480 21.760 140.525 ;
        RECT 20.995 140.340 21.760 140.480 ;
        RECT 20.995 140.280 21.315 140.340 ;
        RECT 21.470 140.295 21.760 140.340 ;
        RECT 22.375 140.480 22.695 140.540 ;
        RECT 24.690 140.480 24.980 140.525 ;
        RECT 28.445 140.480 28.585 140.635 ;
        RECT 31.575 140.620 31.895 140.680 ;
        RECT 33.875 140.620 34.195 140.880 ;
        RECT 38.105 140.540 38.245 141.020 ;
        RECT 45.345 141.020 50.275 141.160 ;
        RECT 45.345 140.975 45.635 141.020 ;
        RECT 48.125 140.975 48.415 141.020 ;
        RECT 49.985 140.975 50.275 141.020 ;
        RECT 50.910 140.975 51.200 141.205 ;
        RECT 65.125 141.160 65.415 141.205 ;
        RECT 67.905 141.160 68.195 141.205 ;
        RECT 69.765 141.160 70.055 141.205 ;
        RECT 76.900 141.160 77.190 141.205 ;
        RECT 79.875 141.160 80.195 141.220 ;
        RECT 65.125 141.020 70.055 141.160 ;
        RECT 65.125 140.975 65.415 141.020 ;
        RECT 67.905 140.975 68.195 141.020 ;
        RECT 69.765 140.975 70.055 141.020 ;
        RECT 75.365 141.020 80.195 141.160 ;
        RECT 41.480 140.820 41.770 140.865 ;
        RECT 43.075 140.820 43.395 140.880 ;
        RECT 41.480 140.680 43.395 140.820 ;
        RECT 41.480 140.635 41.770 140.680 ;
        RECT 43.075 140.620 43.395 140.680 ;
        RECT 44.915 140.620 45.235 140.880 ;
        RECT 45.835 140.820 46.155 140.880 ;
        RECT 50.985 140.820 51.125 140.975 ;
        RECT 45.835 140.680 51.125 140.820 ;
        RECT 45.835 140.620 46.155 140.680 ;
        RECT 52.275 140.620 52.595 140.880 ;
        RECT 55.955 140.820 56.275 140.880 ;
        RECT 55.955 140.680 59.865 140.820 ;
        RECT 55.955 140.620 56.275 140.680 ;
        RECT 22.375 140.340 28.585 140.480 ;
        RECT 22.375 140.280 22.695 140.340 ;
        RECT 24.690 140.295 24.980 140.340 ;
        RECT 32.955 140.280 33.275 140.540 ;
        RECT 34.335 140.280 34.655 140.540 ;
        RECT 38.015 140.480 38.335 140.540 ;
        RECT 39.870 140.480 40.160 140.525 ;
        RECT 45.005 140.480 45.145 140.620 ;
        RECT 59.725 140.540 59.865 140.680 ;
        RECT 38.015 140.340 45.145 140.480 ;
        RECT 45.345 140.480 45.635 140.525 ;
        RECT 45.345 140.340 47.880 140.480 ;
        RECT 38.015 140.280 38.335 140.340 ;
        RECT 39.870 140.295 40.160 140.340 ;
        RECT 45.345 140.295 45.635 140.340 ;
        RECT 27.895 140.140 28.215 140.200 ;
        RECT 47.665 140.185 47.880 140.340 ;
        RECT 48.595 140.280 48.915 140.540 ;
        RECT 50.435 140.280 50.755 140.540 ;
        RECT 51.815 140.280 52.135 140.540 ;
        RECT 57.795 140.280 58.115 140.540 ;
        RECT 58.255 140.280 58.575 140.540 ;
        RECT 58.715 140.280 59.035 140.540 ;
        RECT 59.635 140.280 59.955 140.540 ;
        RECT 65.125 140.480 65.415 140.525 ;
        RECT 65.125 140.340 67.660 140.480 ;
        RECT 65.125 140.295 65.415 140.340 ;
        RECT 28.830 140.140 29.120 140.185 ;
        RECT 27.895 140.000 29.120 140.140 ;
        RECT 27.895 139.940 28.215 140.000 ;
        RECT 28.830 139.955 29.120 140.000 ;
        RECT 40.330 140.140 40.620 140.185 ;
        RECT 43.485 140.140 43.775 140.185 ;
        RECT 46.745 140.140 47.035 140.185 ;
        RECT 40.330 140.000 47.035 140.140 ;
        RECT 40.330 139.955 40.620 140.000 ;
        RECT 43.485 139.955 43.775 140.000 ;
        RECT 46.745 139.955 47.035 140.000 ;
        RECT 47.665 140.140 47.955 140.185 ;
        RECT 49.525 140.140 49.815 140.185 ;
        RECT 47.665 140.000 49.815 140.140 ;
        RECT 47.665 139.955 47.955 140.000 ;
        RECT 49.525 139.955 49.815 140.000 ;
        RECT 53.210 140.140 53.500 140.185 ;
        RECT 56.430 140.140 56.720 140.185 ;
        RECT 53.210 140.000 56.720 140.140 ;
        RECT 53.210 139.955 53.500 140.000 ;
        RECT 56.430 139.955 56.720 140.000 ;
        RECT 32.050 139.800 32.340 139.845 ;
        RECT 49.975 139.800 50.295 139.860 ;
        RECT 32.050 139.660 50.295 139.800 ;
        RECT 58.805 139.800 58.945 140.280 ;
        RECT 66.535 140.185 66.855 140.200 ;
        RECT 63.265 140.140 63.555 140.185 ;
        RECT 66.525 140.140 66.855 140.185 ;
        RECT 63.265 140.000 66.855 140.140 ;
        RECT 63.265 139.955 63.555 140.000 ;
        RECT 66.525 139.955 66.855 140.000 ;
        RECT 67.445 140.185 67.660 140.340 ;
        RECT 68.375 140.280 68.695 140.540 ;
        RECT 70.230 140.480 70.520 140.525 ;
        RECT 71.135 140.480 71.455 140.540 ;
        RECT 70.230 140.340 71.455 140.480 ;
        RECT 70.230 140.295 70.520 140.340 ;
        RECT 71.135 140.280 71.455 140.340 ;
        RECT 72.055 140.480 72.375 140.540 ;
        RECT 72.975 140.480 73.295 140.540 ;
        RECT 72.055 140.340 73.295 140.480 ;
        RECT 72.055 140.280 72.375 140.340 ;
        RECT 72.975 140.280 73.295 140.340 ;
        RECT 74.355 140.280 74.675 140.540 ;
        RECT 74.815 140.280 75.135 140.540 ;
        RECT 75.365 140.525 75.505 141.020 ;
        RECT 76.900 140.975 77.190 141.020 ;
        RECT 79.875 140.960 80.195 141.020 ;
        RECT 80.765 141.160 81.055 141.205 ;
        RECT 83.545 141.160 83.835 141.205 ;
        RECT 85.405 141.160 85.695 141.205 ;
        RECT 80.765 141.020 85.695 141.160 ;
        RECT 80.765 140.975 81.055 141.020 ;
        RECT 83.545 140.975 83.835 141.020 ;
        RECT 85.405 140.975 85.695 141.020 ;
        RECT 91.375 141.160 91.695 141.220 ;
        RECT 91.375 141.020 92.985 141.160 ;
        RECT 91.375 140.960 91.695 141.020 ;
        RECT 85.855 140.820 86.175 140.880 ;
        RECT 92.295 140.820 92.615 140.880 ;
        RECT 92.845 140.865 92.985 141.020 ;
        RECT 85.855 140.680 92.615 140.820 ;
        RECT 85.855 140.620 86.175 140.680 ;
        RECT 92.295 140.620 92.615 140.680 ;
        RECT 92.770 140.635 93.060 140.865 ;
        RECT 75.290 140.295 75.580 140.525 ;
        RECT 75.735 140.480 76.055 140.540 ;
        RECT 76.210 140.480 76.500 140.525 ;
        RECT 75.735 140.340 76.500 140.480 ;
        RECT 75.735 140.280 76.055 140.340 ;
        RECT 76.210 140.295 76.500 140.340 ;
        RECT 80.765 140.480 81.055 140.525 ;
        RECT 80.765 140.340 83.300 140.480 ;
        RECT 80.765 140.295 81.055 140.340 ;
        RECT 83.085 140.185 83.300 140.340 ;
        RECT 84.015 140.280 84.335 140.540 ;
        RECT 87.695 140.480 88.015 140.540 ;
        RECT 91.375 140.480 91.695 140.540 ;
        RECT 87.695 140.340 91.695 140.480 ;
        RECT 87.695 140.280 88.015 140.340 ;
        RECT 91.375 140.280 91.695 140.340 ;
        RECT 91.835 140.280 92.155 140.540 ;
        RECT 94.595 140.480 94.915 140.540 ;
        RECT 95.145 140.525 95.285 141.360 ;
        RECT 96.435 141.300 96.755 141.360 ;
        RECT 101.050 141.500 101.340 141.545 ;
        RECT 106.555 141.500 106.875 141.560 ;
        RECT 101.050 141.360 106.875 141.500 ;
        RECT 101.050 141.315 101.340 141.360 ;
        RECT 106.555 141.300 106.875 141.360 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 96.895 141.160 97.215 141.220 ;
        RECT 96.065 141.020 97.215 141.160 ;
        RECT 95.070 140.480 95.360 140.525 ;
        RECT 94.595 140.340 95.360 140.480 ;
        RECT 94.595 140.280 94.915 140.340 ;
        RECT 95.070 140.295 95.360 140.340 ;
        RECT 95.515 140.280 95.835 140.540 ;
        RECT 96.065 140.525 96.205 141.020 ;
        RECT 96.895 140.960 97.215 141.020 ;
        RECT 105.605 141.160 105.895 141.205 ;
        RECT 108.385 141.160 108.675 141.205 ;
        RECT 110.245 141.160 110.535 141.205 ;
        RECT 105.605 141.020 110.535 141.160 ;
        RECT 105.605 140.975 105.895 141.020 ;
        RECT 108.385 140.975 108.675 141.020 ;
        RECT 110.245 140.975 110.535 141.020 ;
        RECT 97.830 140.820 98.120 140.865 ;
        RECT 99.655 140.820 99.975 140.880 ;
        RECT 102.415 140.820 102.735 140.880 ;
        RECT 97.830 140.680 102.735 140.820 ;
        RECT 97.830 140.635 98.120 140.680 ;
        RECT 99.655 140.620 99.975 140.680 ;
        RECT 102.415 140.620 102.735 140.680 ;
        RECT 108.855 140.620 109.175 140.880 ;
        RECT 96.985 140.525 97.585 140.530 ;
        RECT 95.990 140.295 96.280 140.525 ;
        RECT 96.790 140.480 97.585 140.525 ;
        RECT 98.275 140.480 98.595 140.540 ;
        RECT 96.790 140.390 98.595 140.480 ;
        RECT 96.790 140.340 97.125 140.390 ;
        RECT 97.445 140.340 98.595 140.390 ;
        RECT 96.790 140.295 97.080 140.340 ;
        RECT 98.275 140.280 98.595 140.340 ;
        RECT 99.195 140.280 99.515 140.540 ;
        RECT 105.605 140.480 105.895 140.525 ;
        RECT 105.605 140.340 108.140 140.480 ;
        RECT 105.605 140.295 105.895 140.340 ;
        RECT 67.445 140.140 67.735 140.185 ;
        RECT 69.305 140.140 69.595 140.185 ;
        RECT 67.445 140.000 69.595 140.140 ;
        RECT 67.445 139.955 67.735 140.000 ;
        RECT 69.305 139.955 69.595 140.000 ;
        RECT 78.905 140.140 79.195 140.185 ;
        RECT 82.165 140.140 82.455 140.185 ;
        RECT 83.085 140.140 83.375 140.185 ;
        RECT 84.945 140.140 85.235 140.185 ;
        RECT 78.905 140.000 82.865 140.140 ;
        RECT 78.905 139.955 79.195 140.000 ;
        RECT 82.165 139.955 82.455 140.000 ;
        RECT 66.535 139.940 66.855 139.955 ;
        RECT 61.260 139.800 61.550 139.845 ;
        RECT 62.395 139.800 62.715 139.860 ;
        RECT 58.805 139.660 62.715 139.800 ;
        RECT 32.050 139.615 32.340 139.660 ;
        RECT 49.975 139.600 50.295 139.660 ;
        RECT 61.260 139.615 61.550 139.660 ;
        RECT 62.395 139.600 62.715 139.660 ;
        RECT 72.975 139.600 73.295 139.860 ;
        RECT 82.725 139.800 82.865 140.000 ;
        RECT 83.085 140.000 85.235 140.140 ;
        RECT 83.085 139.955 83.375 140.000 ;
        RECT 84.945 139.955 85.235 140.000 ;
        RECT 93.230 140.140 93.520 140.185 ;
        RECT 93.690 140.140 93.980 140.185 ;
        RECT 93.230 140.000 93.980 140.140 ;
        RECT 93.230 139.955 93.520 140.000 ;
        RECT 93.690 139.955 93.980 140.000 ;
        RECT 98.750 140.140 99.040 140.185 ;
        RECT 101.740 140.140 102.030 140.185 ;
        RECT 98.750 140.000 102.030 140.140 ;
        RECT 98.750 139.955 99.040 140.000 ;
        RECT 101.740 139.955 102.030 140.000 ;
        RECT 103.745 140.140 104.035 140.185 ;
        RECT 106.095 140.140 106.415 140.200 ;
        RECT 107.925 140.185 108.140 140.340 ;
        RECT 110.695 140.280 111.015 140.540 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 107.005 140.140 107.295 140.185 ;
        RECT 103.745 140.000 107.295 140.140 ;
        RECT 103.745 139.955 104.035 140.000 ;
        RECT 87.250 139.800 87.540 139.845 ;
        RECT 82.725 139.660 87.540 139.800 ;
        RECT 87.250 139.615 87.540 139.660 ;
        RECT 90.455 139.800 90.775 139.860 ;
        RECT 90.930 139.800 91.220 139.845 ;
        RECT 90.455 139.660 91.220 139.800 ;
        RECT 90.455 139.600 90.775 139.660 ;
        RECT 90.930 139.615 91.220 139.660 ;
        RECT 96.895 139.800 97.215 139.860 ;
        RECT 98.825 139.800 98.965 139.955 ;
        RECT 106.095 139.940 106.415 140.000 ;
        RECT 107.005 139.955 107.295 140.000 ;
        RECT 107.925 140.140 108.215 140.185 ;
        RECT 109.785 140.140 110.075 140.185 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 107.925 140.000 110.075 140.140 ;
        RECT 107.925 139.955 108.215 140.000 ;
        RECT 109.785 139.955 110.075 140.000 ;
        RECT 96.895 139.660 98.965 139.800 ;
        RECT 96.895 139.600 97.215 139.660 ;
        RECT 17.370 138.980 112.465 139.460 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 39.395 138.780 39.715 138.840 ;
        RECT 41.235 138.780 41.555 138.840 ;
        RECT 39.395 138.640 41.555 138.780 ;
        RECT 39.395 138.580 39.715 138.640 ;
        RECT 32.510 138.440 32.800 138.485 ;
        RECT 38.030 138.440 38.320 138.485 ;
        RECT 32.510 138.300 38.320 138.440 ;
        RECT 32.510 138.255 32.800 138.300 ;
        RECT 38.030 138.255 38.320 138.300 ;
        RECT 33.890 138.100 34.180 138.145 ;
        RECT 36.175 138.100 36.495 138.160 ;
        RECT 33.890 137.960 36.495 138.100 ;
        RECT 33.890 137.915 34.180 137.960 ;
        RECT 36.175 137.900 36.495 137.960 ;
        RECT 37.095 138.100 37.415 138.160 ;
        RECT 38.935 138.100 39.255 138.160 ;
        RECT 39.945 138.145 40.085 138.640 ;
        RECT 41.235 138.580 41.555 138.640 ;
        RECT 44.470 138.780 44.760 138.825 ;
        RECT 48.595 138.780 48.915 138.840 ;
        RECT 44.470 138.640 48.915 138.780 ;
        RECT 44.470 138.595 44.760 138.640 ;
        RECT 48.595 138.580 48.915 138.640 ;
        RECT 49.975 138.780 50.295 138.840 ;
        RECT 60.095 138.780 60.415 138.840 ;
        RECT 49.975 138.640 60.415 138.780 ;
        RECT 49.975 138.580 50.295 138.640 ;
        RECT 60.095 138.580 60.415 138.640 ;
        RECT 62.395 138.580 62.715 138.840 ;
        RECT 66.535 138.780 66.855 138.840 ;
        RECT 67.010 138.780 67.300 138.825 ;
        RECT 66.535 138.640 67.300 138.780 ;
        RECT 66.535 138.580 66.855 138.640 ;
        RECT 67.010 138.595 67.300 138.640 ;
        RECT 68.375 138.780 68.695 138.840 ;
        RECT 68.850 138.780 69.140 138.825 ;
        RECT 68.375 138.640 69.140 138.780 ;
        RECT 68.375 138.580 68.695 138.640 ;
        RECT 68.850 138.595 69.140 138.640 ;
        RECT 79.875 138.580 80.195 138.840 ;
        RECT 82.190 138.595 82.480 138.825 ;
        RECT 83.570 138.780 83.860 138.825 ;
        RECT 84.015 138.780 84.335 138.840 ;
        RECT 83.570 138.640 84.335 138.780 ;
        RECT 83.570 138.595 83.860 138.640 ;
        RECT 43.075 138.440 43.395 138.500 ;
        RECT 40.405 138.300 43.395 138.440 ;
        RECT 40.405 138.145 40.545 138.300 ;
        RECT 43.075 138.240 43.395 138.300 ;
        RECT 47.230 138.440 47.520 138.485 ;
        RECT 56.430 138.440 56.720 138.485 ;
        RECT 62.870 138.440 63.160 138.485 ;
        RECT 47.230 138.300 56.720 138.440 ;
        RECT 47.230 138.255 47.520 138.300 ;
        RECT 56.430 138.255 56.720 138.300 ;
        RECT 58.805 138.300 63.160 138.440 ;
        RECT 58.805 138.160 58.945 138.300 ;
        RECT 62.870 138.255 63.160 138.300 ;
        RECT 72.975 138.240 73.295 138.500 ;
        RECT 39.410 138.100 39.700 138.145 ;
        RECT 37.095 137.960 39.700 138.100 ;
        RECT 37.095 137.900 37.415 137.960 ;
        RECT 38.935 137.900 39.255 137.960 ;
        RECT 39.410 137.915 39.700 137.960 ;
        RECT 39.870 137.915 40.160 138.145 ;
        RECT 40.330 137.915 40.620 138.145 ;
        RECT 40.775 138.100 41.095 138.160 ;
        RECT 41.250 138.100 41.540 138.145 ;
        RECT 40.775 137.960 41.540 138.100 ;
        RECT 40.775 137.900 41.095 137.960 ;
        RECT 41.250 137.915 41.540 137.960 ;
        RECT 43.535 137.900 43.855 138.160 ;
        RECT 44.455 138.100 44.775 138.160 ;
        RECT 45.850 138.100 46.140 138.145 ;
        RECT 44.455 137.960 46.140 138.100 ;
        RECT 44.455 137.900 44.775 137.960 ;
        RECT 45.850 137.915 46.140 137.960 ;
        RECT 57.795 137.900 58.115 138.160 ;
        RECT 58.255 137.900 58.575 138.160 ;
        RECT 58.715 137.900 59.035 138.160 ;
        RECT 59.635 137.900 59.955 138.160 ;
        RECT 63.315 138.100 63.635 138.160 ;
        RECT 66.090 138.100 66.380 138.145 ;
        RECT 63.315 137.960 66.380 138.100 ;
        RECT 63.315 137.900 63.635 137.960 ;
        RECT 66.090 137.915 66.380 137.960 ;
        RECT 66.995 138.100 67.315 138.160 ;
        RECT 67.470 138.100 67.760 138.145 ;
        RECT 66.995 137.960 67.760 138.100 ;
        RECT 66.995 137.900 67.315 137.960 ;
        RECT 67.470 137.915 67.760 137.960 ;
        RECT 67.930 137.915 68.220 138.145 ;
        RECT 33.430 137.760 33.720 137.805 ;
        RECT 35.715 137.760 36.035 137.820 ;
        RECT 33.430 137.620 36.035 137.760 ;
        RECT 33.430 137.575 33.720 137.620 ;
        RECT 35.715 137.560 36.035 137.620 ;
        RECT 46.770 137.760 47.060 137.805 ;
        RECT 50.895 137.760 51.215 137.820 ;
        RECT 46.770 137.620 51.215 137.760 ;
        RECT 46.770 137.575 47.060 137.620 ;
        RECT 50.895 137.560 51.215 137.620 ;
        RECT 55.495 137.760 55.815 137.820 ;
        RECT 61.490 137.760 61.780 137.805 ;
        RECT 68.005 137.760 68.145 137.915 ;
        RECT 71.595 137.900 71.915 138.160 ;
        RECT 80.335 137.900 80.655 138.160 ;
        RECT 82.265 138.100 82.405 138.595 ;
        RECT 84.015 138.580 84.335 138.640 ;
        RECT 89.995 138.780 90.315 138.840 ;
        RECT 89.995 138.640 96.205 138.780 ;
        RECT 89.995 138.580 90.315 138.640 ;
        RECT 86.330 138.440 86.620 138.485 ;
        RECT 90.470 138.440 90.760 138.485 ;
        RECT 94.595 138.440 94.915 138.500 ;
        RECT 86.330 138.300 90.760 138.440 ;
        RECT 86.330 138.255 86.620 138.300 ;
        RECT 90.470 138.255 90.760 138.300 ;
        RECT 91.925 138.300 94.915 138.440 ;
        RECT 82.650 138.100 82.940 138.145 ;
        RECT 82.265 137.960 82.940 138.100 ;
        RECT 82.650 137.915 82.940 137.960 ;
        RECT 84.935 137.900 85.255 138.160 ;
        RECT 86.775 137.900 87.095 138.160 ;
        RECT 87.695 137.900 88.015 138.160 ;
        RECT 88.155 137.900 88.475 138.160 ;
        RECT 91.925 138.145 92.065 138.300 ;
        RECT 94.595 138.240 94.915 138.300 ;
        RECT 88.630 138.100 88.920 138.145 ;
        RECT 91.850 138.100 92.140 138.145 ;
        RECT 88.630 137.960 92.140 138.100 ;
        RECT 88.630 137.915 88.920 137.960 ;
        RECT 91.850 137.915 92.140 137.960 ;
        RECT 92.310 137.915 92.600 138.145 ;
        RECT 92.770 138.115 93.060 138.145 ;
        RECT 92.770 137.975 93.445 138.115 ;
        RECT 92.770 137.915 93.060 137.975 ;
        RECT 55.495 137.620 61.780 137.760 ;
        RECT 55.495 137.560 55.815 137.620 ;
        RECT 61.490 137.575 61.780 137.620 ;
        RECT 64.785 137.620 68.145 137.760 ;
        RECT 72.530 137.760 72.820 137.805 ;
        RECT 73.435 137.760 73.755 137.820 ;
        RECT 72.530 137.620 73.755 137.760 ;
        RECT 34.810 137.420 35.100 137.465 ;
        RECT 55.035 137.420 55.355 137.480 ;
        RECT 64.785 137.465 64.925 137.620 ;
        RECT 72.530 137.575 72.820 137.620 ;
        RECT 73.435 137.560 73.755 137.620 ;
        RECT 79.430 137.760 79.720 137.805 ;
        RECT 82.175 137.760 82.495 137.820 ;
        RECT 79.430 137.620 82.495 137.760 ;
        RECT 79.430 137.575 79.720 137.620 ;
        RECT 82.175 137.560 82.495 137.620 ;
        RECT 85.870 137.760 86.160 137.805 ;
        RECT 90.915 137.760 91.235 137.820 ;
        RECT 85.870 137.620 91.235 137.760 ;
        RECT 85.870 137.575 86.160 137.620 ;
        RECT 90.915 137.560 91.235 137.620 ;
        RECT 91.375 137.760 91.695 137.820 ;
        RECT 92.385 137.760 92.525 137.915 ;
        RECT 91.375 137.620 92.525 137.760 ;
        RECT 93.305 137.760 93.445 137.975 ;
        RECT 93.690 138.100 93.980 138.145 ;
        RECT 94.135 138.100 94.455 138.160 ;
        RECT 93.690 137.960 94.455 138.100 ;
        RECT 93.690 137.915 93.980 137.960 ;
        RECT 94.135 137.900 94.455 137.960 ;
        RECT 96.065 138.100 96.205 138.640 ;
        RECT 96.895 138.580 97.215 138.840 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 100.590 138.440 100.880 138.485 ;
        RECT 103.745 138.440 104.035 138.485 ;
        RECT 107.005 138.440 107.295 138.485 ;
        RECT 100.590 138.300 107.295 138.440 ;
        RECT 100.590 138.255 100.880 138.300 ;
        RECT 103.745 138.255 104.035 138.300 ;
        RECT 107.005 138.255 107.295 138.300 ;
        RECT 107.925 138.440 108.215 138.485 ;
        RECT 109.785 138.440 110.075 138.485 ;
        RECT 107.925 138.300 110.075 138.440 ;
        RECT 107.925 138.255 108.215 138.300 ;
        RECT 109.785 138.255 110.075 138.300 ;
        RECT 99.655 138.100 99.975 138.160 ;
        RECT 96.065 137.960 99.975 138.100 ;
        RECT 94.595 137.760 94.915 137.820 ;
        RECT 96.065 137.805 96.205 137.960 ;
        RECT 99.655 137.900 99.975 137.960 ;
        RECT 100.130 138.100 100.420 138.145 ;
        RECT 105.605 138.100 105.895 138.145 ;
        RECT 107.925 138.100 108.140 138.255 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 100.130 137.960 101.495 138.100 ;
        RECT 100.130 137.915 100.420 137.960 ;
        RECT 93.305 137.620 94.915 137.760 ;
        RECT 91.375 137.560 91.695 137.620 ;
        RECT 94.595 137.560 94.915 137.620 ;
        RECT 95.990 137.575 96.280 137.805 ;
        RECT 96.450 137.575 96.740 137.805 ;
        RECT 101.355 137.760 101.495 137.960 ;
        RECT 105.605 137.960 108.140 138.100 ;
        RECT 105.605 137.915 105.895 137.960 ;
        RECT 108.855 137.900 109.175 138.160 ;
        RECT 103.795 137.760 104.115 137.820 ;
        RECT 101.355 137.620 104.115 137.760 ;
        RECT 34.810 137.280 55.355 137.420 ;
        RECT 34.810 137.235 35.100 137.280 ;
        RECT 55.035 137.220 55.355 137.280 ;
        RECT 64.710 137.235 65.000 137.465 ;
        RECT 68.835 137.420 69.155 137.480 ;
        RECT 87.695 137.420 88.015 137.480 ;
        RECT 96.525 137.420 96.665 137.575 ;
        RECT 103.795 137.560 104.115 137.620 ;
        RECT 106.095 137.760 106.415 137.820 ;
        RECT 110.695 137.760 111.015 137.820 ;
        RECT 106.095 137.620 111.015 137.760 ;
        RECT 106.095 137.560 106.415 137.620 ;
        RECT 110.695 137.560 111.015 137.620 ;
        RECT 101.955 137.465 102.275 137.480 ;
        RECT 101.740 137.420 102.275 137.465 ;
        RECT 68.835 137.280 71.825 137.420 ;
        RECT 68.835 137.220 69.155 137.280 ;
        RECT 32.955 136.880 33.275 137.140 ;
        RECT 44.455 137.080 44.775 137.140 ;
        RECT 44.930 137.080 45.220 137.125 ;
        RECT 44.455 136.940 45.220 137.080 ;
        RECT 44.455 136.880 44.775 136.940 ;
        RECT 44.930 136.895 45.220 136.940 ;
        RECT 47.215 136.880 47.535 137.140 ;
        RECT 61.475 137.080 61.795 137.140 ;
        RECT 65.170 137.080 65.460 137.125 ;
        RECT 61.475 136.940 65.460 137.080 ;
        RECT 61.475 136.880 61.795 136.940 ;
        RECT 65.170 136.895 65.460 136.940 ;
        RECT 70.215 137.080 70.535 137.140 ;
        RECT 71.685 137.125 71.825 137.280 ;
        RECT 87.695 137.280 102.275 137.420 ;
        RECT 87.695 137.220 88.015 137.280 ;
        RECT 101.740 137.235 102.275 137.280 ;
        RECT 105.605 137.420 105.895 137.465 ;
        RECT 108.385 137.420 108.675 137.465 ;
        RECT 110.245 137.420 110.535 137.465 ;
        RECT 105.605 137.280 110.535 137.420 ;
        RECT 105.605 137.235 105.895 137.280 ;
        RECT 108.385 137.235 108.675 137.280 ;
        RECT 110.245 137.235 110.535 137.280 ;
        RECT 101.955 137.220 102.275 137.235 ;
        RECT 70.690 137.080 70.980 137.125 ;
        RECT 70.215 136.940 70.980 137.080 ;
        RECT 70.215 136.880 70.535 136.940 ;
        RECT 70.690 136.895 70.980 136.940 ;
        RECT 71.610 136.895 71.900 137.125 ;
        RECT 84.015 136.880 84.335 137.140 ;
        RECT 86.330 137.080 86.620 137.125 ;
        RECT 87.235 137.080 87.555 137.140 ;
        RECT 86.330 136.940 87.555 137.080 ;
        RECT 86.330 136.895 86.620 136.940 ;
        RECT 87.235 136.880 87.555 136.940 ;
        RECT 90.010 137.080 90.300 137.125 ;
        RECT 95.515 137.080 95.835 137.140 ;
        RECT 90.010 136.940 95.835 137.080 ;
        RECT 90.010 136.895 90.300 136.940 ;
        RECT 95.515 136.880 95.835 136.940 ;
        RECT 98.750 137.080 99.040 137.125 ;
        RECT 106.555 137.080 106.875 137.140 ;
        RECT 98.750 136.940 106.875 137.080 ;
        RECT 98.750 136.895 99.040 136.940 ;
        RECT 106.555 136.880 106.875 136.940 ;
        RECT 18.165 136.260 112.465 136.740 ;
        RECT 31.575 136.060 31.895 136.120 ;
        RECT 32.510 136.060 32.800 136.105 ;
        RECT 31.575 135.920 32.800 136.060 ;
        RECT 31.575 135.860 31.895 135.920 ;
        RECT 32.510 135.875 32.800 135.920 ;
        RECT 39.855 136.060 40.175 136.120 ;
        RECT 45.835 136.060 46.155 136.120 ;
        RECT 53.655 136.060 53.975 136.120 ;
        RECT 39.855 135.920 46.155 136.060 ;
        RECT 39.855 135.860 40.175 135.920 ;
        RECT 45.835 135.860 46.155 135.920 ;
        RECT 48.225 135.920 53.975 136.060 ;
        RECT 34.350 135.720 34.640 135.765 ;
        RECT 47.675 135.720 47.995 135.780 ;
        RECT 34.350 135.580 47.995 135.720 ;
        RECT 34.350 135.535 34.640 135.580 ;
        RECT 47.675 135.520 47.995 135.580 ;
        RECT 32.970 135.380 33.260 135.425 ;
        RECT 34.795 135.380 35.115 135.440 ;
        RECT 38.015 135.380 38.335 135.440 ;
        RECT 32.970 135.240 35.115 135.380 ;
        RECT 32.970 135.195 33.260 135.240 ;
        RECT 34.795 135.180 35.115 135.240 ;
        RECT 37.645 135.240 38.335 135.380 ;
        RECT 33.430 135.040 33.720 135.085 ;
        RECT 36.635 135.040 36.955 135.100 ;
        RECT 37.645 135.085 37.785 135.240 ;
        RECT 38.015 135.180 38.335 135.240 ;
        RECT 38.935 135.380 39.255 135.440 ;
        RECT 44.915 135.380 45.235 135.440 ;
        RECT 46.080 135.380 46.370 135.425 ;
        RECT 38.935 135.240 41.005 135.380 ;
        RECT 38.935 135.180 39.255 135.240 ;
        RECT 40.865 135.100 41.005 135.240 ;
        RECT 41.325 135.240 46.370 135.380 ;
        RECT 33.430 134.900 36.955 135.040 ;
        RECT 33.430 134.855 33.720 134.900 ;
        RECT 36.635 134.840 36.955 134.900 ;
        RECT 37.570 134.855 37.860 135.085 ;
        RECT 40.315 134.840 40.635 135.100 ;
        RECT 40.775 134.840 41.095 135.100 ;
        RECT 41.325 135.085 41.465 135.240 ;
        RECT 44.915 135.180 45.235 135.240 ;
        RECT 46.080 135.195 46.370 135.240 ;
        RECT 41.250 134.855 41.540 135.085 ;
        RECT 42.170 134.855 42.460 135.085 ;
        RECT 43.075 135.040 43.395 135.100 ;
        RECT 48.225 135.040 48.365 135.920 ;
        RECT 53.655 135.860 53.975 135.920 ;
        RECT 60.095 136.060 60.415 136.120 ;
        RECT 61.935 136.060 62.255 136.120 ;
        RECT 60.095 135.920 62.255 136.060 ;
        RECT 60.095 135.860 60.415 135.920 ;
        RECT 61.935 135.860 62.255 135.920 ;
        RECT 63.315 136.060 63.635 136.120 ;
        RECT 66.535 136.060 66.855 136.120 ;
        RECT 63.315 135.920 66.855 136.060 ;
        RECT 63.315 135.860 63.635 135.920 ;
        RECT 66.535 135.860 66.855 135.920 ;
        RECT 96.435 135.860 96.755 136.120 ;
        RECT 97.140 136.060 97.430 136.105 ;
        RECT 99.195 136.060 99.515 136.120 ;
        RECT 97.140 135.920 99.515 136.060 ;
        RECT 97.140 135.875 97.430 135.920 ;
        RECT 49.945 135.720 50.235 135.765 ;
        RECT 52.725 135.720 53.015 135.765 ;
        RECT 54.585 135.720 54.875 135.765 ;
        RECT 49.945 135.580 54.875 135.720 ;
        RECT 49.945 135.535 50.235 135.580 ;
        RECT 52.725 135.535 53.015 135.580 ;
        RECT 54.585 135.535 54.875 135.580 ;
        RECT 65.125 135.720 65.415 135.765 ;
        RECT 67.905 135.720 68.195 135.765 ;
        RECT 69.765 135.720 70.055 135.765 ;
        RECT 65.125 135.580 70.055 135.720 ;
        RECT 65.125 135.535 65.415 135.580 ;
        RECT 67.905 135.535 68.195 135.580 ;
        RECT 69.765 135.535 70.055 135.580 ;
        RECT 75.735 135.520 76.055 135.780 ;
        RECT 83.110 135.535 83.400 135.765 ;
        RECT 93.215 135.720 93.535 135.780 ;
        RECT 93.690 135.720 93.980 135.765 ;
        RECT 93.215 135.580 93.980 135.720 ;
        RECT 50.435 135.380 50.755 135.440 ;
        RECT 52.275 135.380 52.595 135.440 ;
        RECT 50.435 135.240 52.965 135.380 ;
        RECT 50.435 135.180 50.755 135.240 ;
        RECT 52.275 135.180 52.595 135.240 ;
        RECT 43.075 134.900 48.365 135.040 ;
        RECT 49.945 135.040 50.235 135.085 ;
        RECT 52.825 135.040 52.965 135.240 ;
        RECT 53.195 135.180 53.515 135.440 ;
        RECT 55.495 135.380 55.815 135.440 ;
        RECT 56.890 135.380 57.180 135.425 ;
        RECT 55.495 135.240 57.180 135.380 ;
        RECT 55.495 135.180 55.815 135.240 ;
        RECT 56.890 135.195 57.180 135.240 ;
        RECT 57.810 135.380 58.100 135.425 ;
        RECT 58.715 135.380 59.035 135.440 ;
        RECT 61.260 135.380 61.550 135.425 ;
        RECT 74.355 135.380 74.675 135.440 ;
        RECT 57.810 135.240 61.550 135.380 ;
        RECT 57.810 135.195 58.100 135.240 ;
        RECT 58.715 135.180 59.035 135.240 ;
        RECT 61.260 135.195 61.550 135.240 ;
        RECT 61.795 135.240 74.675 135.380 ;
        RECT 75.825 135.380 75.965 135.520 ;
        RECT 80.350 135.380 80.640 135.425 ;
        RECT 82.635 135.380 82.955 135.440 ;
        RECT 75.825 135.240 77.345 135.380 ;
        RECT 55.050 135.040 55.340 135.085 ;
        RECT 49.945 134.900 52.480 135.040 ;
        RECT 52.825 134.900 55.340 135.040 ;
        RECT 32.050 134.700 32.340 134.745 ;
        RECT 38.950 134.700 39.240 134.745 ;
        RECT 32.050 134.560 39.240 134.700 ;
        RECT 32.050 134.515 32.340 134.560 ;
        RECT 38.950 134.515 39.240 134.560 ;
        RECT 39.395 134.700 39.715 134.760 ;
        RECT 42.245 134.700 42.385 134.855 ;
        RECT 43.075 134.840 43.395 134.900 ;
        RECT 49.945 134.855 50.235 134.900 ;
        RECT 48.085 134.700 48.375 134.745 ;
        RECT 49.515 134.700 49.835 134.760 ;
        RECT 52.265 134.745 52.480 134.900 ;
        RECT 55.050 134.855 55.340 134.900 ;
        RECT 55.955 135.040 56.275 135.100 ;
        RECT 61.795 135.040 61.935 135.240 ;
        RECT 74.355 135.180 74.675 135.240 ;
        RECT 55.955 134.900 61.935 135.040 ;
        RECT 65.125 135.040 65.415 135.085 ;
        RECT 65.125 134.900 67.660 135.040 ;
        RECT 55.955 134.840 56.275 134.900 ;
        RECT 65.125 134.855 65.415 134.900 ;
        RECT 66.535 134.745 66.855 134.760 ;
        RECT 51.345 134.700 51.635 134.745 ;
        RECT 39.395 134.560 46.525 134.700 ;
        RECT 39.395 134.500 39.715 134.560 ;
        RECT 38.015 134.160 38.335 134.420 ;
        RECT 46.385 134.360 46.525 134.560 ;
        RECT 48.085 134.560 51.635 134.700 ;
        RECT 48.085 134.515 48.375 134.560 ;
        RECT 49.515 134.500 49.835 134.560 ;
        RECT 51.345 134.515 51.635 134.560 ;
        RECT 52.265 134.700 52.555 134.745 ;
        RECT 54.125 134.700 54.415 134.745 ;
        RECT 52.265 134.560 54.415 134.700 ;
        RECT 52.265 134.515 52.555 134.560 ;
        RECT 54.125 134.515 54.415 134.560 ;
        RECT 63.265 134.700 63.555 134.745 ;
        RECT 66.525 134.700 66.855 134.745 ;
        RECT 63.265 134.560 66.855 134.700 ;
        RECT 63.265 134.515 63.555 134.560 ;
        RECT 66.525 134.515 66.855 134.560 ;
        RECT 67.445 134.745 67.660 134.900 ;
        RECT 68.375 134.840 68.695 135.100 ;
        RECT 70.230 135.040 70.520 135.085 ;
        RECT 71.135 135.040 71.455 135.100 ;
        RECT 70.230 134.900 71.455 135.040 ;
        RECT 74.445 135.040 74.585 135.180 ;
        RECT 77.205 135.100 77.345 135.240 ;
        RECT 80.350 135.240 82.955 135.380 ;
        RECT 80.350 135.195 80.640 135.240 ;
        RECT 82.635 135.180 82.955 135.240 ;
        RECT 75.290 135.040 75.580 135.085 ;
        RECT 74.445 134.900 75.580 135.040 ;
        RECT 70.230 134.855 70.520 134.900 ;
        RECT 71.135 134.840 71.455 134.900 ;
        RECT 75.290 134.855 75.580 134.900 ;
        RECT 75.750 134.855 76.040 135.085 ;
        RECT 76.210 134.855 76.500 135.085 ;
        RECT 67.445 134.700 67.735 134.745 ;
        RECT 69.305 134.700 69.595 134.745 ;
        RECT 67.445 134.560 69.595 134.700 ;
        RECT 67.445 134.515 67.735 134.560 ;
        RECT 69.305 134.515 69.595 134.560 ;
        RECT 74.815 134.700 75.135 134.760 ;
        RECT 75.825 134.700 75.965 134.855 ;
        RECT 74.815 134.560 75.965 134.700 ;
        RECT 76.285 134.700 76.425 134.855 ;
        RECT 77.115 134.840 77.435 135.100 ;
        RECT 83.185 135.040 83.325 135.535 ;
        RECT 93.215 135.520 93.535 135.580 ;
        RECT 93.690 135.535 93.980 135.580 ;
        RECT 94.135 135.520 94.455 135.780 ;
        RECT 94.595 135.720 94.915 135.780 ;
        RECT 97.215 135.720 97.355 135.875 ;
        RECT 99.195 135.860 99.515 135.920 ;
        RECT 107.490 136.060 107.780 136.105 ;
        RECT 108.855 136.060 109.175 136.120 ;
        RECT 107.490 135.920 109.175 136.060 ;
        RECT 107.490 135.875 107.780 135.920 ;
        RECT 108.855 135.860 109.175 135.920 ;
        RECT 94.595 135.580 97.355 135.720 ;
        RECT 101.005 135.720 101.295 135.765 ;
        RECT 103.785 135.720 104.075 135.765 ;
        RECT 105.645 135.720 105.935 135.765 ;
        RECT 101.005 135.580 105.935 135.720 ;
        RECT 94.595 135.520 94.915 135.580 ;
        RECT 101.005 135.535 101.295 135.580 ;
        RECT 103.785 135.535 104.075 135.580 ;
        RECT 105.645 135.535 105.935 135.580 ;
        RECT 89.995 135.380 90.315 135.440 ;
        RECT 90.470 135.380 90.760 135.425 ;
        RECT 89.995 135.240 90.760 135.380 ;
        RECT 89.995 135.180 90.315 135.240 ;
        RECT 90.470 135.195 90.760 135.240 ;
        RECT 83.570 135.040 83.860 135.085 ;
        RECT 83.185 134.900 83.860 135.040 ;
        RECT 83.570 134.855 83.860 134.900 ;
        RECT 91.850 135.040 92.140 135.085 ;
        RECT 94.685 135.040 94.825 135.520 ;
        RECT 95.990 135.380 96.280 135.425 ;
        RECT 97.355 135.380 97.675 135.440 ;
        RECT 95.990 135.240 97.675 135.380 ;
        RECT 95.990 135.195 96.280 135.240 ;
        RECT 97.355 135.180 97.675 135.240 ;
        RECT 91.850 134.900 94.825 135.040 ;
        RECT 91.850 134.855 92.140 134.900 ;
        RECT 95.055 134.840 95.375 135.100 ;
        RECT 95.515 135.040 95.835 135.100 ;
        RECT 96.450 135.040 96.740 135.085 ;
        RECT 95.515 134.900 96.740 135.040 ;
        RECT 95.515 134.840 95.835 134.900 ;
        RECT 96.450 134.855 96.740 134.900 ;
        RECT 101.005 135.040 101.295 135.085 ;
        RECT 104.270 135.040 104.560 135.085 ;
        RECT 104.715 135.040 105.035 135.100 ;
        RECT 101.005 134.900 103.540 135.040 ;
        RECT 101.005 134.855 101.295 134.900 ;
        RECT 77.575 134.700 77.895 134.760 ;
        RECT 80.335 134.700 80.655 134.760 ;
        RECT 80.810 134.700 81.100 134.745 ;
        RECT 76.285 134.560 81.100 134.700 ;
        RECT 66.535 134.500 66.855 134.515 ;
        RECT 74.815 134.500 75.135 134.560 ;
        RECT 77.575 134.500 77.895 134.560 ;
        RECT 80.335 134.500 80.655 134.560 ;
        RECT 80.810 134.515 81.100 134.560 ;
        RECT 98.275 134.700 98.595 134.760 ;
        RECT 103.325 134.745 103.540 134.900 ;
        RECT 104.270 134.900 105.035 135.040 ;
        RECT 104.270 134.855 104.560 134.900 ;
        RECT 104.715 134.840 105.035 134.900 ;
        RECT 106.095 134.840 106.415 135.100 ;
        RECT 106.555 134.840 106.875 135.100 ;
        RECT 99.145 134.700 99.435 134.745 ;
        RECT 102.405 134.700 102.695 134.745 ;
        RECT 98.275 134.560 102.695 134.700 ;
        RECT 98.275 134.500 98.595 134.560 ;
        RECT 99.145 134.515 99.435 134.560 ;
        RECT 102.405 134.515 102.695 134.560 ;
        RECT 103.325 134.700 103.615 134.745 ;
        RECT 105.185 134.700 105.475 134.745 ;
        RECT 103.325 134.560 105.475 134.700 ;
        RECT 103.325 134.515 103.615 134.560 ;
        RECT 105.185 134.515 105.475 134.560 ;
        RECT 54.575 134.360 54.895 134.420 ;
        RECT 46.385 134.220 54.895 134.360 ;
        RECT 54.575 134.160 54.895 134.220 ;
        RECT 57.335 134.360 57.655 134.420 ;
        RECT 58.270 134.360 58.560 134.405 ;
        RECT 57.335 134.220 58.560 134.360 ;
        RECT 57.335 134.160 57.655 134.220 ;
        RECT 58.270 134.175 58.560 134.220 ;
        RECT 60.095 134.160 60.415 134.420 ;
        RECT 72.975 134.360 73.295 134.420 ;
        RECT 73.910 134.360 74.200 134.405 ;
        RECT 72.975 134.220 74.200 134.360 ;
        RECT 72.975 134.160 73.295 134.220 ;
        RECT 73.910 134.175 74.200 134.220 ;
        RECT 81.255 134.160 81.575 134.420 ;
        RECT 84.490 134.360 84.780 134.405 ;
        RECT 84.935 134.360 85.255 134.420 ;
        RECT 84.490 134.220 85.255 134.360 ;
        RECT 84.490 134.175 84.780 134.220 ;
        RECT 84.935 134.160 85.255 134.220 ;
        RECT 91.375 134.160 91.695 134.420 ;
        RECT 92.295 134.360 92.615 134.420 ;
        RECT 106.185 134.360 106.325 134.840 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 92.295 134.220 106.325 134.360 ;
        RECT 92.295 134.160 92.615 134.220 ;
        RECT 17.370 133.540 112.465 134.020 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 23.295 133.340 23.615 133.400 ;
        RECT 27.895 133.340 28.215 133.400 ;
        RECT 23.295 133.200 27.665 133.340 ;
        RECT 23.295 133.140 23.615 133.200 ;
        RECT 22.850 132.475 23.140 132.705 ;
        RECT 24.675 132.660 24.995 132.720 ;
        RECT 26.990 132.660 27.280 132.705 ;
        RECT 24.675 132.520 27.280 132.660 ;
        RECT 27.525 132.660 27.665 133.200 ;
        RECT 27.895 133.200 32.725 133.340 ;
        RECT 27.895 133.140 28.215 133.200 ;
        RECT 31.590 132.660 31.880 132.705 ;
        RECT 27.525 132.520 31.880 132.660 ;
        RECT 22.925 132.320 23.065 132.475 ;
        RECT 24.675 132.460 24.995 132.520 ;
        RECT 26.990 132.475 27.280 132.520 ;
        RECT 31.590 132.475 31.880 132.520 ;
        RECT 32.035 132.460 32.355 132.720 ;
        RECT 26.055 132.320 26.375 132.380 ;
        RECT 22.925 132.180 26.375 132.320 ;
        RECT 26.055 132.120 26.375 132.180 ;
        RECT 27.450 132.320 27.740 132.365 ;
        RECT 27.895 132.320 28.215 132.380 ;
        RECT 27.450 132.180 28.215 132.320 ;
        RECT 27.450 132.135 27.740 132.180 ;
        RECT 27.895 132.120 28.215 132.180 ;
        RECT 28.370 132.135 28.660 132.365 ;
        RECT 32.585 132.320 32.725 133.200 ;
        RECT 33.415 133.140 33.735 133.400 ;
        RECT 38.935 133.340 39.255 133.400 ;
        RECT 37.645 133.200 39.255 133.340 ;
        RECT 32.970 133.000 33.260 133.045 ;
        RECT 35.730 133.000 36.020 133.045 ;
        RECT 32.970 132.860 36.020 133.000 ;
        RECT 32.970 132.815 33.260 132.860 ;
        RECT 35.730 132.815 36.020 132.860 ;
        RECT 34.335 132.460 34.655 132.720 ;
        RECT 37.095 132.460 37.415 132.720 ;
        RECT 37.645 132.705 37.785 133.200 ;
        RECT 38.935 133.140 39.255 133.200 ;
        RECT 41.250 133.340 41.540 133.385 ;
        RECT 44.915 133.340 45.235 133.400 ;
        RECT 41.250 133.200 45.235 133.340 ;
        RECT 41.250 133.155 41.540 133.200 ;
        RECT 44.915 133.140 45.235 133.200 ;
        RECT 49.515 133.140 49.835 133.400 ;
        RECT 60.095 133.340 60.415 133.400 ;
        RECT 65.630 133.340 65.920 133.385 ;
        RECT 66.535 133.340 66.855 133.400 ;
        RECT 60.095 133.200 64.465 133.340 ;
        RECT 60.095 133.140 60.415 133.200 ;
        RECT 43.535 133.000 43.855 133.060 ;
        RECT 45.390 133.000 45.680 133.045 ;
        RECT 55.955 133.000 56.275 133.060 ;
        RECT 61.015 133.045 61.335 133.060 ;
        RECT 38.105 132.860 39.625 133.000 ;
        RECT 38.105 132.705 38.245 132.860 ;
        RECT 37.570 132.475 37.860 132.705 ;
        RECT 38.030 132.475 38.320 132.705 ;
        RECT 38.935 132.460 39.255 132.720 ;
        RECT 39.485 132.660 39.625 132.860 ;
        RECT 43.535 132.860 45.680 133.000 ;
        RECT 43.535 132.800 43.855 132.860 ;
        RECT 45.390 132.815 45.680 132.860 ;
        RECT 53.285 132.860 56.275 133.000 ;
        RECT 49.070 132.660 49.360 132.705 ;
        RECT 49.975 132.660 50.295 132.720 ;
        RECT 53.285 132.705 53.425 132.860 ;
        RECT 55.955 132.800 56.275 132.860 ;
        RECT 57.745 133.000 58.035 133.045 ;
        RECT 61.005 133.000 61.335 133.045 ;
        RECT 57.745 132.860 61.335 133.000 ;
        RECT 57.745 132.815 58.035 132.860 ;
        RECT 61.005 132.815 61.335 132.860 ;
        RECT 61.015 132.800 61.335 132.815 ;
        RECT 61.925 133.000 62.215 133.045 ;
        RECT 63.785 133.000 64.075 133.045 ;
        RECT 61.925 132.860 64.075 133.000 ;
        RECT 64.325 133.000 64.465 133.200 ;
        RECT 65.630 133.200 66.855 133.340 ;
        RECT 65.630 133.155 65.920 133.200 ;
        RECT 66.535 133.140 66.855 133.200 ;
        RECT 67.470 133.340 67.760 133.385 ;
        RECT 68.375 133.340 68.695 133.400 ;
        RECT 67.470 133.200 68.695 133.340 ;
        RECT 67.470 133.155 67.760 133.200 ;
        RECT 68.375 133.140 68.695 133.200 ;
        RECT 77.575 133.385 77.895 133.400 ;
        RECT 77.575 133.155 78.110 133.385 ;
        RECT 81.255 133.340 81.575 133.400 ;
        RECT 87.480 133.340 87.770 133.385 ;
        RECT 91.375 133.340 91.695 133.400 ;
        RECT 79.505 133.200 91.695 133.340 ;
        RECT 77.575 133.140 77.895 133.155 ;
        RECT 64.325 132.860 66.765 133.000 ;
        RECT 61.925 132.815 62.215 132.860 ;
        RECT 63.785 132.815 64.075 132.860 ;
        RECT 39.485 132.520 41.005 132.660 ;
        RECT 40.865 132.380 41.005 132.520 ;
        RECT 49.070 132.520 50.295 132.660 ;
        RECT 49.070 132.475 49.360 132.520 ;
        RECT 49.975 132.460 50.295 132.520 ;
        RECT 50.450 132.475 50.740 132.705 ;
        RECT 53.210 132.475 53.500 132.705 ;
        RECT 35.270 132.320 35.560 132.365 ;
        RECT 39.395 132.320 39.715 132.380 ;
        RECT 32.585 132.180 39.715 132.320 ;
        RECT 35.270 132.135 35.560 132.180 ;
        RECT 25.595 131.980 25.915 132.040 ;
        RECT 28.445 131.980 28.585 132.135 ;
        RECT 39.395 132.120 39.715 132.180 ;
        RECT 40.330 132.135 40.620 132.365 ;
        RECT 25.595 131.840 28.585 131.980 ;
        RECT 40.405 131.980 40.545 132.135 ;
        RECT 40.775 132.120 41.095 132.380 ;
        RECT 44.010 132.320 44.300 132.365 ;
        RECT 45.375 132.320 45.695 132.380 ;
        RECT 44.010 132.180 45.695 132.320 ;
        RECT 44.010 132.135 44.300 132.180 ;
        RECT 44.085 131.980 44.225 132.135 ;
        RECT 45.375 132.120 45.695 132.180 ;
        RECT 40.405 131.840 44.225 131.980 ;
        RECT 47.230 131.980 47.520 132.025 ;
        RECT 50.525 131.980 50.665 132.475 ;
        RECT 53.655 132.460 53.975 132.720 ;
        RECT 54.115 132.460 54.435 132.720 ;
        RECT 54.575 132.660 54.895 132.720 ;
        RECT 55.050 132.660 55.340 132.705 ;
        RECT 58.255 132.660 58.575 132.720 ;
        RECT 54.575 132.520 58.575 132.660 ;
        RECT 54.575 132.460 54.895 132.520 ;
        RECT 55.050 132.475 55.340 132.520 ;
        RECT 58.255 132.460 58.575 132.520 ;
        RECT 59.605 132.660 59.895 132.705 ;
        RECT 61.925 132.660 62.140 132.815 ;
        RECT 59.605 132.520 62.140 132.660 ;
        RECT 63.315 132.660 63.635 132.720 ;
        RECT 66.625 132.705 66.765 132.860 ;
        RECT 72.975 132.800 73.295 133.060 ;
        RECT 74.815 133.000 75.135 133.060 ;
        RECT 79.505 133.000 79.645 133.200 ;
        RECT 81.255 133.140 81.575 133.200 ;
        RECT 87.480 133.155 87.770 133.200 ;
        RECT 91.375 133.140 91.695 133.200 ;
        RECT 91.835 133.340 92.155 133.400 ;
        RECT 91.835 133.200 98.045 133.340 ;
        RECT 91.835 133.140 92.155 133.200 ;
        RECT 73.525 132.860 75.965 133.000 ;
        RECT 66.090 132.660 66.380 132.705 ;
        RECT 63.315 132.520 66.380 132.660 ;
        RECT 59.605 132.475 59.895 132.520 ;
        RECT 63.315 132.460 63.635 132.520 ;
        RECT 66.090 132.475 66.380 132.520 ;
        RECT 66.550 132.475 66.840 132.705 ;
        RECT 69.295 132.660 69.615 132.720 ;
        RECT 71.610 132.660 71.900 132.705 ;
        RECT 73.525 132.660 73.665 132.860 ;
        RECT 74.815 132.800 75.135 132.860 ;
        RECT 69.295 132.520 71.900 132.660 ;
        RECT 69.295 132.460 69.615 132.520 ;
        RECT 71.610 132.475 71.900 132.520 ;
        RECT 72.145 132.520 73.665 132.660 ;
        RECT 74.355 132.660 74.675 132.720 ;
        RECT 75.825 132.705 75.965 132.860 ;
        RECT 76.285 132.860 79.645 133.000 ;
        RECT 79.825 133.000 80.115 133.045 ;
        RECT 82.175 133.000 82.495 133.060 ;
        RECT 89.535 133.045 89.855 133.060 ;
        RECT 83.085 133.000 83.375 133.045 ;
        RECT 79.825 132.860 83.375 133.000 ;
        RECT 76.285 132.705 76.425 132.860 ;
        RECT 79.825 132.815 80.115 132.860 ;
        RECT 82.175 132.800 82.495 132.860 ;
        RECT 83.085 132.815 83.375 132.860 ;
        RECT 84.005 133.000 84.295 133.045 ;
        RECT 85.865 133.000 86.155 133.045 ;
        RECT 84.005 132.860 86.155 133.000 ;
        RECT 84.005 132.815 84.295 132.860 ;
        RECT 85.865 132.815 86.155 132.860 ;
        RECT 89.485 133.000 89.855 133.045 ;
        RECT 92.745 133.000 93.035 133.045 ;
        RECT 89.485 132.860 93.035 133.000 ;
        RECT 89.485 132.815 89.855 132.860 ;
        RECT 92.745 132.815 93.035 132.860 ;
        RECT 93.665 133.000 93.955 133.045 ;
        RECT 95.525 133.000 95.815 133.045 ;
        RECT 93.665 132.860 95.815 133.000 ;
        RECT 93.665 132.815 93.955 132.860 ;
        RECT 95.525 132.815 95.815 132.860 ;
        RECT 75.290 132.660 75.580 132.705 ;
        RECT 74.355 132.520 75.580 132.660 ;
        RECT 61.935 132.320 62.255 132.380 ;
        RECT 62.870 132.320 63.160 132.365 ;
        RECT 61.935 132.180 63.160 132.320 ;
        RECT 61.935 132.120 62.255 132.180 ;
        RECT 62.870 132.135 63.160 132.180 ;
        RECT 63.775 132.320 64.095 132.380 ;
        RECT 64.710 132.320 65.000 132.365 ;
        RECT 72.145 132.320 72.285 132.520 ;
        RECT 74.355 132.460 74.675 132.520 ;
        RECT 75.290 132.475 75.580 132.520 ;
        RECT 75.750 132.475 76.040 132.705 ;
        RECT 76.210 132.475 76.500 132.705 ;
        RECT 77.115 132.460 77.435 132.720 ;
        RECT 81.685 132.660 81.975 132.705 ;
        RECT 84.005 132.660 84.220 132.815 ;
        RECT 89.535 132.800 89.855 132.815 ;
        RECT 81.685 132.520 84.220 132.660 ;
        RECT 81.685 132.475 81.975 132.520 ;
        RECT 84.935 132.460 85.255 132.720 ;
        RECT 91.345 132.660 91.635 132.705 ;
        RECT 93.665 132.660 93.880 132.815 ;
        RECT 91.345 132.520 93.880 132.660 ;
        RECT 91.345 132.475 91.635 132.520 ;
        RECT 94.595 132.460 94.915 132.720 ;
        RECT 97.905 132.705 98.045 133.200 ;
        RECT 98.275 133.140 98.595 133.400 ;
        RECT 99.195 133.340 99.515 133.400 ;
        RECT 101.050 133.340 101.340 133.385 ;
        RECT 99.195 133.200 101.340 133.340 ;
        RECT 99.195 133.140 99.515 133.200 ;
        RECT 101.050 133.155 101.340 133.200 ;
        RECT 101.510 133.340 101.800 133.385 ;
        RECT 101.955 133.340 102.275 133.400 ;
        RECT 101.510 133.200 102.275 133.340 ;
        RECT 101.510 133.155 101.800 133.200 ;
        RECT 101.955 133.140 102.275 133.200 ;
        RECT 103.350 133.155 103.640 133.385 ;
        RECT 97.830 132.475 98.120 132.705 ;
        RECT 103.425 132.660 103.565 133.155 ;
        RECT 104.715 133.140 105.035 133.400 ;
        RECT 103.810 132.660 104.100 132.705 ;
        RECT 103.425 132.520 104.100 132.660 ;
        RECT 103.810 132.475 104.100 132.520 ;
        RECT 63.775 132.180 65.000 132.320 ;
        RECT 63.775 132.120 64.095 132.180 ;
        RECT 64.710 132.135 65.000 132.180 ;
        RECT 65.245 132.180 72.285 132.320 ;
        RECT 47.230 131.840 50.665 131.980 ;
        RECT 51.370 131.980 51.660 132.025 ;
        RECT 52.735 131.980 53.055 132.040 ;
        RECT 51.370 131.840 53.055 131.980 ;
        RECT 25.595 131.780 25.915 131.840 ;
        RECT 47.230 131.795 47.520 131.840 ;
        RECT 51.370 131.795 51.660 131.840 ;
        RECT 52.735 131.780 53.055 131.840 ;
        RECT 53.655 131.980 53.975 132.040 ;
        RECT 59.605 131.980 59.895 132.025 ;
        RECT 62.385 131.980 62.675 132.025 ;
        RECT 64.245 131.980 64.535 132.025 ;
        RECT 53.655 131.840 58.025 131.980 ;
        RECT 53.655 131.780 53.975 131.840 ;
        RECT 23.295 131.440 23.615 131.700 ;
        RECT 25.135 131.440 25.455 131.700 ;
        RECT 28.355 131.640 28.675 131.700 ;
        RECT 30.670 131.640 30.960 131.685 ;
        RECT 28.355 131.500 30.960 131.640 ;
        RECT 28.355 131.440 28.675 131.500 ;
        RECT 30.670 131.455 30.960 131.500 ;
        RECT 31.575 131.640 31.895 131.700 ;
        RECT 32.510 131.640 32.800 131.685 ;
        RECT 31.575 131.500 32.800 131.640 ;
        RECT 31.575 131.440 31.895 131.500 ;
        RECT 32.510 131.455 32.800 131.500 ;
        RECT 43.075 131.440 43.395 131.700 ;
        RECT 43.535 131.640 43.855 131.700 ;
        RECT 49.515 131.640 49.835 131.700 ;
        RECT 43.535 131.500 49.835 131.640 ;
        RECT 43.535 131.440 43.855 131.500 ;
        RECT 49.515 131.440 49.835 131.500 ;
        RECT 51.815 131.440 52.135 131.700 ;
        RECT 54.115 131.640 54.435 131.700 ;
        RECT 55.740 131.640 56.030 131.685 ;
        RECT 57.335 131.640 57.655 131.700 ;
        RECT 54.115 131.500 57.655 131.640 ;
        RECT 57.885 131.640 58.025 131.840 ;
        RECT 59.605 131.840 64.535 131.980 ;
        RECT 59.605 131.795 59.895 131.840 ;
        RECT 62.385 131.795 62.675 131.840 ;
        RECT 64.245 131.795 64.535 131.840 ;
        RECT 65.245 131.640 65.385 132.180 ;
        RECT 72.515 132.120 72.835 132.380 ;
        RECT 73.895 132.320 74.215 132.380 ;
        RECT 77.205 132.320 77.345 132.460 ;
        RECT 73.895 132.180 77.345 132.320 ;
        RECT 83.095 132.320 83.415 132.380 ;
        RECT 86.790 132.320 87.080 132.365 ;
        RECT 83.095 132.180 87.080 132.320 ;
        RECT 73.895 132.120 74.215 132.180 ;
        RECT 83.095 132.120 83.415 132.180 ;
        RECT 86.790 132.135 87.080 132.180 ;
        RECT 92.295 132.320 92.615 132.380 ;
        RECT 96.450 132.320 96.740 132.365 ;
        RECT 92.295 132.180 96.740 132.320 ;
        RECT 92.295 132.120 92.615 132.180 ;
        RECT 96.450 132.135 96.740 132.180 ;
        RECT 100.590 132.320 100.880 132.365 ;
        RECT 102.415 132.320 102.735 132.380 ;
        RECT 100.590 132.180 102.735 132.320 ;
        RECT 100.590 132.135 100.880 132.180 ;
        RECT 102.415 132.120 102.735 132.180 ;
        RECT 70.690 131.980 70.980 132.025 ;
        RECT 74.355 131.980 74.675 132.040 ;
        RECT 70.690 131.840 74.675 131.980 ;
        RECT 70.690 131.795 70.980 131.840 ;
        RECT 74.355 131.780 74.675 131.840 ;
        RECT 81.685 131.980 81.975 132.025 ;
        RECT 84.465 131.980 84.755 132.025 ;
        RECT 86.325 131.980 86.615 132.025 ;
        RECT 81.685 131.840 86.615 131.980 ;
        RECT 81.685 131.795 81.975 131.840 ;
        RECT 84.465 131.795 84.755 131.840 ;
        RECT 86.325 131.795 86.615 131.840 ;
        RECT 91.345 131.980 91.635 132.025 ;
        RECT 94.125 131.980 94.415 132.025 ;
        RECT 95.985 131.980 96.275 132.025 ;
        RECT 91.345 131.840 96.275 131.980 ;
        RECT 91.345 131.795 91.635 131.840 ;
        RECT 94.125 131.795 94.415 131.840 ;
        RECT 95.985 131.795 96.275 131.840 ;
        RECT 57.885 131.500 65.385 131.640 ;
        RECT 54.115 131.440 54.435 131.500 ;
        RECT 55.740 131.455 56.030 131.500 ;
        RECT 57.335 131.440 57.655 131.500 ;
        RECT 72.975 131.440 73.295 131.700 ;
        RECT 73.435 131.640 73.755 131.700 ;
        RECT 73.910 131.640 74.200 131.685 ;
        RECT 73.435 131.500 74.200 131.640 ;
        RECT 73.435 131.440 73.755 131.500 ;
        RECT 73.910 131.455 74.200 131.500 ;
        RECT 18.165 130.820 112.465 131.300 ;
        RECT 26.055 130.620 26.375 130.680 ;
        RECT 29.735 130.620 30.055 130.680 ;
        RECT 26.055 130.480 30.055 130.620 ;
        RECT 26.055 130.420 26.375 130.480 ;
        RECT 29.735 130.420 30.055 130.480 ;
        RECT 32.955 130.420 33.275 130.680 ;
        RECT 35.255 130.620 35.575 130.680 ;
        RECT 35.730 130.620 36.020 130.665 ;
        RECT 35.255 130.480 36.020 130.620 ;
        RECT 35.255 130.420 35.575 130.480 ;
        RECT 35.730 130.435 36.020 130.480 ;
        RECT 38.260 130.620 38.550 130.665 ;
        RECT 40.775 130.620 41.095 130.680 ;
        RECT 43.535 130.620 43.855 130.680 ;
        RECT 38.260 130.480 43.855 130.620 ;
        RECT 38.260 130.435 38.550 130.480 ;
        RECT 40.775 130.420 41.095 130.480 ;
        RECT 43.535 130.420 43.855 130.480 ;
        RECT 45.375 130.620 45.695 130.680 ;
        RECT 48.610 130.620 48.900 130.665 ;
        RECT 45.375 130.480 48.900 130.620 ;
        RECT 45.375 130.420 45.695 130.480 ;
        RECT 48.610 130.435 48.900 130.480 ;
        RECT 61.935 130.420 62.255 130.680 ;
        RECT 70.230 130.620 70.520 130.665 ;
        RECT 70.675 130.620 70.995 130.680 ;
        RECT 70.230 130.480 70.995 130.620 ;
        RECT 70.230 130.435 70.520 130.480 ;
        RECT 70.675 130.420 70.995 130.480 ;
        RECT 82.175 130.620 82.495 130.680 ;
        RECT 82.650 130.620 82.940 130.665 ;
        RECT 82.175 130.480 82.940 130.620 ;
        RECT 82.175 130.420 82.495 130.480 ;
        RECT 82.650 130.435 82.940 130.480 ;
        RECT 85.410 130.620 85.700 130.665 ;
        RECT 89.535 130.620 89.855 130.680 ;
        RECT 85.410 130.480 89.855 130.620 ;
        RECT 85.410 130.435 85.700 130.480 ;
        RECT 89.535 130.420 89.855 130.480 ;
        RECT 92.295 130.620 92.615 130.680 ;
        RECT 93.230 130.620 93.520 130.665 ;
        RECT 92.295 130.480 93.520 130.620 ;
        RECT 92.295 130.420 92.615 130.480 ;
        RECT 93.230 130.435 93.520 130.480 ;
        RECT 94.595 130.620 94.915 130.680 ;
        RECT 95.990 130.620 96.280 130.665 ;
        RECT 94.595 130.480 96.280 130.620 ;
        RECT 94.595 130.420 94.915 130.480 ;
        RECT 95.990 130.435 96.280 130.480 ;
        RECT 23.725 130.280 24.015 130.325 ;
        RECT 26.505 130.280 26.795 130.325 ;
        RECT 28.365 130.280 28.655 130.325 ;
        RECT 23.725 130.140 28.655 130.280 ;
        RECT 23.725 130.095 24.015 130.140 ;
        RECT 26.505 130.095 26.795 130.140 ;
        RECT 28.365 130.095 28.655 130.140 ;
        RECT 42.125 130.280 42.415 130.325 ;
        RECT 44.905 130.280 45.195 130.325 ;
        RECT 46.765 130.280 47.055 130.325 ;
        RECT 42.125 130.140 47.055 130.280 ;
        RECT 42.125 130.095 42.415 130.140 ;
        RECT 44.905 130.095 45.195 130.140 ;
        RECT 46.765 130.095 47.055 130.140 ;
        RECT 61.015 130.280 61.335 130.340 ;
        RECT 62.870 130.280 63.160 130.325 ;
        RECT 73.895 130.280 74.215 130.340 ;
        RECT 61.015 130.140 63.160 130.280 ;
        RECT 61.015 130.080 61.335 130.140 ;
        RECT 62.870 130.095 63.160 130.140 ;
        RECT 66.855 130.140 74.215 130.280 ;
        RECT 24.675 129.940 24.995 130.000 ;
        RECT 31.130 129.940 31.420 129.985 ;
        RECT 24.675 129.800 31.420 129.940 ;
        RECT 24.675 129.740 24.995 129.800 ;
        RECT 31.130 129.755 31.420 129.800 ;
        RECT 42.615 129.940 42.935 130.000 ;
        RECT 45.390 129.940 45.680 129.985 ;
        RECT 42.615 129.800 45.680 129.940 ;
        RECT 42.615 129.740 42.935 129.800 ;
        RECT 45.390 129.755 45.680 129.800 ;
        RECT 49.055 129.740 49.375 130.000 ;
        RECT 49.515 129.940 49.835 130.000 ;
        RECT 55.495 129.940 55.815 130.000 ;
        RECT 56.430 129.940 56.720 129.985 ;
        RECT 49.515 129.800 52.505 129.940 ;
        RECT 49.515 129.740 49.835 129.800 ;
        RECT 23.725 129.600 24.015 129.645 ;
        RECT 26.990 129.600 27.280 129.645 ;
        RECT 27.435 129.600 27.755 129.660 ;
        RECT 23.725 129.460 26.260 129.600 ;
        RECT 23.725 129.415 24.015 129.460 ;
        RECT 21.865 129.260 22.155 129.305 ;
        RECT 23.295 129.260 23.615 129.320 ;
        RECT 26.045 129.305 26.260 129.460 ;
        RECT 26.990 129.460 27.755 129.600 ;
        RECT 26.990 129.415 27.280 129.460 ;
        RECT 27.435 129.400 27.755 129.460 ;
        RECT 28.815 129.400 29.135 129.660 ;
        RECT 29.735 129.400 30.055 129.660 ;
        RECT 32.050 129.600 32.340 129.645 ;
        RECT 34.335 129.600 34.655 129.660 ;
        RECT 36.635 129.600 36.955 129.660 ;
        RECT 32.050 129.460 36.955 129.600 ;
        RECT 32.050 129.415 32.340 129.460 ;
        RECT 34.335 129.400 34.655 129.460 ;
        RECT 36.635 129.400 36.955 129.460 ;
        RECT 37.570 129.600 37.860 129.645 ;
        RECT 38.935 129.600 39.255 129.660 ;
        RECT 37.570 129.460 39.255 129.600 ;
        RECT 37.570 129.415 37.860 129.460 ;
        RECT 38.935 129.400 39.255 129.460 ;
        RECT 42.125 129.600 42.415 129.645 ;
        RECT 42.125 129.460 44.660 129.600 ;
        RECT 42.125 129.415 42.415 129.460 ;
        RECT 25.125 129.260 25.415 129.305 ;
        RECT 21.865 129.120 25.415 129.260 ;
        RECT 21.865 129.075 22.155 129.120 ;
        RECT 23.295 129.060 23.615 129.120 ;
        RECT 25.125 129.075 25.415 129.120 ;
        RECT 26.045 129.260 26.335 129.305 ;
        RECT 27.905 129.260 28.195 129.305 ;
        RECT 26.045 129.120 28.195 129.260 ;
        RECT 26.045 129.075 26.335 129.120 ;
        RECT 27.905 129.075 28.195 129.120 ;
        RECT 38.015 129.260 38.335 129.320 ;
        RECT 44.445 129.305 44.660 129.460 ;
        RECT 47.230 129.415 47.520 129.645 ;
        RECT 40.265 129.260 40.555 129.305 ;
        RECT 43.525 129.260 43.815 129.305 ;
        RECT 38.015 129.120 43.815 129.260 ;
        RECT 38.015 129.060 38.335 129.120 ;
        RECT 40.265 129.075 40.555 129.120 ;
        RECT 43.525 129.075 43.815 129.120 ;
        RECT 44.445 129.260 44.735 129.305 ;
        RECT 46.305 129.260 46.595 129.305 ;
        RECT 44.445 129.120 46.595 129.260 ;
        RECT 47.305 129.260 47.445 129.415 ;
        RECT 48.595 129.400 48.915 129.660 ;
        RECT 49.990 129.600 50.280 129.645 ;
        RECT 51.815 129.600 52.135 129.660 ;
        RECT 49.990 129.460 52.135 129.600 ;
        RECT 52.365 129.600 52.505 129.800 ;
        RECT 55.495 129.800 56.720 129.940 ;
        RECT 55.495 129.740 55.815 129.800 ;
        RECT 56.430 129.755 56.720 129.800 ;
        RECT 57.335 129.740 57.655 130.000 ;
        RECT 58.255 129.940 58.575 130.000 ;
        RECT 66.855 129.940 66.995 130.140 ;
        RECT 73.895 130.080 74.215 130.140 ;
        RECT 58.255 129.800 66.995 129.940 ;
        RECT 58.255 129.740 58.575 129.800 ;
        RECT 71.135 129.740 71.455 130.000 ;
        RECT 57.810 129.600 58.100 129.645 ;
        RECT 61.030 129.600 61.320 129.645 ;
        RECT 52.365 129.460 58.100 129.600 ;
        RECT 49.990 129.415 50.280 129.460 ;
        RECT 51.815 129.400 52.135 129.460 ;
        RECT 57.810 129.415 58.100 129.460 ;
        RECT 59.725 129.460 61.320 129.600 ;
        RECT 52.275 129.260 52.595 129.320 ;
        RECT 47.305 129.120 52.595 129.260 ;
        RECT 44.445 129.075 44.735 129.120 ;
        RECT 46.305 129.075 46.595 129.120 ;
        RECT 52.275 129.060 52.595 129.120 ;
        RECT 19.860 128.920 20.150 128.965 ;
        RECT 24.675 128.920 24.995 128.980 ;
        RECT 19.860 128.780 24.995 128.920 ;
        RECT 19.860 128.735 20.150 128.780 ;
        RECT 24.675 128.720 24.995 128.780 ;
        RECT 30.195 128.720 30.515 128.980 ;
        RECT 45.375 128.920 45.695 128.980 ;
        RECT 59.725 128.965 59.865 129.460 ;
        RECT 61.030 129.415 61.320 129.460 ;
        RECT 63.315 129.400 63.635 129.660 ;
        RECT 68.850 129.415 69.140 129.645 ;
        RECT 68.925 129.260 69.065 129.415 ;
        RECT 69.295 129.400 69.615 129.660 ;
        RECT 79.415 129.400 79.735 129.660 ;
        RECT 83.110 129.600 83.400 129.645 ;
        RECT 84.950 129.600 85.240 129.645 ;
        RECT 87.695 129.600 88.015 129.660 ;
        RECT 91.835 129.600 92.155 129.660 ;
        RECT 83.110 129.460 92.155 129.600 ;
        RECT 83.110 129.415 83.400 129.460 ;
        RECT 84.950 129.415 85.240 129.460 ;
        RECT 87.695 129.400 88.015 129.460 ;
        RECT 91.835 129.400 92.155 129.460 ;
        RECT 93.215 129.600 93.535 129.660 ;
        RECT 96.910 129.600 97.200 129.645 ;
        RECT 93.215 129.460 97.200 129.600 ;
        RECT 93.215 129.400 93.535 129.460 ;
        RECT 96.910 129.415 97.200 129.460 ;
        RECT 74.815 129.260 75.135 129.320 ;
        RECT 68.925 129.120 75.135 129.260 ;
        RECT 79.505 129.260 79.645 129.400 ;
        RECT 86.790 129.260 87.080 129.305 ;
        RECT 79.505 129.120 87.080 129.260 ;
        RECT 74.815 129.060 75.135 129.120 ;
        RECT 86.790 129.075 87.080 129.120 ;
        RECT 47.690 128.920 47.980 128.965 ;
        RECT 45.375 128.780 47.980 128.920 ;
        RECT 45.375 128.720 45.695 128.780 ;
        RECT 47.690 128.735 47.980 128.780 ;
        RECT 59.650 128.735 59.940 128.965 ;
        RECT 17.370 128.100 112.465 128.580 ;
        RECT 24.675 127.700 24.995 127.960 ;
        RECT 27.435 127.700 27.755 127.960 ;
        RECT 27.895 127.945 28.215 127.960 ;
        RECT 27.895 127.715 28.430 127.945 ;
        RECT 37.570 127.715 37.860 127.945 ;
        RECT 27.895 127.700 28.215 127.715 ;
        RECT 30.195 127.605 30.515 127.620 ;
        RECT 30.145 127.560 30.515 127.605 ;
        RECT 33.405 127.560 33.695 127.605 ;
        RECT 30.145 127.420 33.695 127.560 ;
        RECT 30.145 127.375 30.515 127.420 ;
        RECT 33.405 127.375 33.695 127.420 ;
        RECT 34.325 127.560 34.615 127.605 ;
        RECT 36.185 127.560 36.475 127.605 ;
        RECT 34.325 127.420 36.475 127.560 ;
        RECT 34.325 127.375 34.615 127.420 ;
        RECT 36.185 127.375 36.475 127.420 ;
        RECT 30.195 127.360 30.515 127.375 ;
        RECT 20.550 127.220 20.840 127.265 ;
        RECT 20.550 127.080 22.605 127.220 ;
        RECT 20.550 127.035 20.840 127.080 ;
        RECT 22.465 126.585 22.605 127.080 ;
        RECT 24.215 127.020 24.535 127.280 ;
        RECT 25.135 127.220 25.455 127.280 ;
        RECT 26.530 127.220 26.820 127.265 ;
        RECT 25.135 127.080 26.820 127.220 ;
        RECT 25.135 127.020 25.455 127.080 ;
        RECT 26.530 127.035 26.820 127.080 ;
        RECT 32.005 127.220 32.295 127.265 ;
        RECT 34.325 127.220 34.540 127.375 ;
        RECT 32.005 127.080 34.540 127.220 ;
        RECT 37.645 127.220 37.785 127.715 ;
        RECT 39.395 127.700 39.715 127.960 ;
        RECT 42.615 127.700 42.935 127.960 ;
        RECT 71.135 127.900 71.455 127.960 ;
        RECT 75.735 127.900 76.055 127.960 ;
        RECT 76.210 127.900 76.500 127.945 ;
        RECT 71.135 127.760 75.505 127.900 ;
        RECT 71.135 127.700 71.455 127.760 ;
        RECT 60.555 127.560 60.875 127.620 ;
        RECT 61.490 127.560 61.780 127.605 ;
        RECT 58.805 127.420 61.780 127.560 ;
        RECT 38.015 127.220 38.335 127.280 ;
        RECT 37.645 127.080 38.335 127.220 ;
        RECT 32.005 127.035 32.295 127.080 ;
        RECT 38.015 127.020 38.335 127.080 ;
        RECT 41.710 127.220 42.000 127.265 ;
        RECT 42.615 127.220 42.935 127.280 ;
        RECT 41.710 127.080 42.935 127.220 ;
        RECT 41.710 127.035 42.000 127.080 ;
        RECT 42.615 127.020 42.935 127.080 ;
        RECT 43.535 127.020 43.855 127.280 ;
        RECT 44.010 127.220 44.300 127.265 ;
        RECT 46.310 127.220 46.600 127.265 ;
        RECT 44.010 127.080 46.600 127.220 ;
        RECT 44.010 127.035 44.300 127.080 ;
        RECT 46.310 127.035 46.600 127.080 ;
        RECT 24.675 126.880 24.995 126.940 ;
        RECT 25.595 126.880 25.915 126.940 ;
        RECT 24.675 126.740 25.915 126.880 ;
        RECT 24.675 126.680 24.995 126.740 ;
        RECT 25.595 126.680 25.915 126.740 ;
        RECT 35.255 126.680 35.575 126.940 ;
        RECT 37.110 126.695 37.400 126.925 ;
        RECT 38.935 126.880 39.255 126.940 ;
        RECT 39.870 126.880 40.160 126.925 ;
        RECT 38.935 126.740 40.160 126.880 ;
        RECT 22.390 126.355 22.680 126.585 ;
        RECT 32.005 126.540 32.295 126.585 ;
        RECT 34.785 126.540 35.075 126.585 ;
        RECT 36.645 126.540 36.935 126.585 ;
        RECT 32.005 126.400 36.935 126.540 ;
        RECT 37.185 126.540 37.325 126.695 ;
        RECT 38.935 126.680 39.255 126.740 ;
        RECT 39.870 126.695 40.160 126.740 ;
        RECT 40.775 126.680 41.095 126.940 ;
        RECT 42.155 126.880 42.475 126.940 ;
        RECT 45.390 126.880 45.680 126.925 ;
        RECT 42.155 126.740 45.680 126.880 ;
        RECT 46.385 126.880 46.525 127.035 ;
        RECT 47.215 127.020 47.535 127.280 ;
        RECT 48.135 127.220 48.455 127.280 ;
        RECT 48.610 127.220 48.900 127.265 ;
        RECT 48.135 127.080 48.900 127.220 ;
        RECT 48.135 127.020 48.455 127.080 ;
        RECT 48.610 127.035 48.900 127.080 ;
        RECT 49.530 127.035 49.820 127.265 ;
        RECT 52.275 127.220 52.595 127.280 ;
        RECT 52.750 127.220 53.040 127.265 ;
        RECT 52.275 127.080 53.040 127.220 ;
        RECT 49.605 126.880 49.745 127.035 ;
        RECT 52.275 127.020 52.595 127.080 ;
        RECT 52.750 127.035 53.040 127.080 ;
        RECT 57.350 127.220 57.640 127.265 ;
        RECT 58.805 127.220 58.945 127.420 ;
        RECT 60.555 127.360 60.875 127.420 ;
        RECT 61.490 127.375 61.780 127.420 ;
        RECT 72.990 127.560 73.280 127.605 ;
        RECT 73.435 127.560 73.755 127.620 ;
        RECT 72.990 127.420 73.755 127.560 ;
        RECT 75.365 127.560 75.505 127.760 ;
        RECT 75.735 127.760 76.500 127.900 ;
        RECT 75.735 127.700 76.055 127.760 ;
        RECT 76.210 127.715 76.500 127.760 ;
        RECT 86.775 127.605 87.095 127.620 ;
        RECT 80.810 127.560 81.100 127.605 ;
        RECT 84.035 127.560 84.325 127.605 ;
        RECT 85.895 127.560 86.185 127.605 ;
        RECT 75.365 127.420 83.325 127.560 ;
        RECT 72.990 127.375 73.280 127.420 ;
        RECT 73.435 127.360 73.755 127.420 ;
        RECT 80.810 127.375 81.100 127.420 ;
        RECT 83.185 127.280 83.325 127.420 ;
        RECT 84.035 127.420 86.185 127.560 ;
        RECT 84.035 127.375 84.325 127.420 ;
        RECT 85.895 127.375 86.185 127.420 ;
        RECT 57.350 127.080 58.945 127.220 ;
        RECT 59.190 127.220 59.480 127.265 ;
        RECT 63.330 127.220 63.620 127.265 ;
        RECT 59.190 127.080 63.620 127.220 ;
        RECT 57.350 127.035 57.640 127.080 ;
        RECT 59.190 127.035 59.480 127.080 ;
        RECT 63.330 127.035 63.620 127.080 ;
        RECT 46.385 126.740 49.745 126.880 ;
        RECT 42.155 126.680 42.475 126.740 ;
        RECT 45.390 126.695 45.680 126.740 ;
        RECT 37.555 126.540 37.875 126.600 ;
        RECT 45.835 126.540 46.155 126.600 ;
        RECT 37.185 126.400 46.155 126.540 ;
        RECT 32.005 126.355 32.295 126.400 ;
        RECT 34.785 126.355 35.075 126.400 ;
        RECT 36.645 126.355 36.935 126.400 ;
        RECT 37.555 126.340 37.875 126.400 ;
        RECT 45.835 126.340 46.155 126.400 ;
        RECT 21.455 126.000 21.775 126.260 ;
        RECT 43.995 126.200 44.315 126.260 ;
        RECT 44.930 126.200 45.220 126.245 ;
        RECT 43.995 126.060 45.220 126.200 ;
        RECT 49.605 126.200 49.745 126.740 ;
        RECT 50.450 126.880 50.740 126.925 ;
        RECT 51.815 126.880 52.135 126.940 ;
        RECT 50.450 126.740 52.135 126.880 ;
        RECT 50.450 126.695 50.740 126.740 ;
        RECT 51.815 126.680 52.135 126.740 ;
        RECT 58.270 126.540 58.560 126.585 ;
        RECT 59.265 126.540 59.405 127.035 ;
        RECT 69.295 127.020 69.615 127.280 ;
        RECT 69.755 127.220 70.075 127.280 ;
        RECT 71.610 127.220 71.900 127.265 ;
        RECT 69.755 127.080 71.900 127.220 ;
        RECT 69.755 127.020 70.075 127.080 ;
        RECT 71.610 127.035 71.900 127.080 ;
        RECT 72.055 127.020 72.375 127.280 ;
        RECT 72.515 127.220 72.835 127.280 ;
        RECT 82.190 127.220 82.480 127.265 ;
        RECT 72.515 127.080 82.480 127.220 ;
        RECT 72.515 127.020 72.835 127.080 ;
        RECT 82.190 127.035 82.480 127.080 ;
        RECT 83.095 127.020 83.415 127.280 ;
        RECT 85.970 127.220 86.185 127.375 ;
        RECT 86.775 127.560 87.105 127.605 ;
        RECT 90.075 127.560 90.365 127.605 ;
        RECT 86.775 127.420 90.365 127.560 ;
        RECT 86.775 127.375 87.105 127.420 ;
        RECT 90.075 127.375 90.365 127.420 ;
        RECT 91.835 127.560 92.155 127.620 ;
        RECT 100.590 127.560 100.880 127.605 ;
        RECT 103.745 127.560 104.035 127.605 ;
        RECT 107.005 127.560 107.295 127.605 ;
        RECT 91.835 127.420 100.345 127.560 ;
        RECT 86.775 127.360 87.095 127.375 ;
        RECT 91.835 127.360 92.155 127.420 ;
        RECT 88.215 127.220 88.505 127.265 ;
        RECT 85.970 127.080 88.505 127.220 ;
        RECT 88.215 127.035 88.505 127.080 ;
        RECT 93.675 127.020 93.995 127.280 ;
        RECT 94.595 127.220 94.915 127.280 ;
        RECT 96.435 127.220 96.755 127.280 ;
        RECT 100.205 127.265 100.345 127.420 ;
        RECT 100.590 127.420 107.295 127.560 ;
        RECT 100.590 127.375 100.880 127.420 ;
        RECT 103.745 127.375 104.035 127.420 ;
        RECT 107.005 127.375 107.295 127.420 ;
        RECT 107.925 127.560 108.215 127.605 ;
        RECT 109.785 127.560 110.075 127.605 ;
        RECT 107.925 127.420 110.075 127.560 ;
        RECT 107.925 127.375 108.215 127.420 ;
        RECT 109.785 127.375 110.075 127.420 ;
        RECT 96.910 127.220 97.200 127.265 ;
        RECT 94.595 127.080 96.205 127.220 ;
        RECT 94.595 127.020 94.915 127.080 ;
        RECT 64.250 126.880 64.540 126.925 ;
        RECT 64.250 126.740 65.385 126.880 ;
        RECT 64.250 126.695 64.540 126.740 ;
        RECT 58.270 126.400 59.405 126.540 ;
        RECT 58.270 126.355 58.560 126.400 ;
        RECT 50.895 126.200 51.215 126.260 ;
        RECT 59.635 126.200 59.955 126.260 ;
        RECT 49.605 126.060 59.955 126.200 ;
        RECT 43.995 126.000 44.315 126.060 ;
        RECT 44.930 126.015 45.220 126.060 ;
        RECT 50.895 126.000 51.215 126.060 ;
        RECT 59.635 126.000 59.955 126.060 ;
        RECT 61.015 126.000 61.335 126.260 ;
        RECT 62.395 126.000 62.715 126.260 ;
        RECT 65.245 126.200 65.385 126.740 ;
        RECT 68.390 126.695 68.680 126.925 ;
        RECT 68.835 126.880 69.155 126.940 ;
        RECT 70.230 126.880 70.520 126.925 ;
        RECT 68.835 126.740 70.520 126.880 ;
        RECT 67.915 126.540 68.235 126.600 ;
        RECT 68.465 126.540 68.605 126.695 ;
        RECT 68.835 126.680 69.155 126.740 ;
        RECT 70.230 126.695 70.520 126.740 ;
        RECT 75.275 126.680 75.595 126.940 ;
        RECT 75.750 126.695 76.040 126.925 ;
        RECT 84.950 126.880 85.240 126.925 ;
        RECT 86.775 126.880 87.095 126.940 ;
        RECT 84.950 126.740 87.095 126.880 ;
        RECT 84.950 126.695 85.240 126.740 ;
        RECT 75.825 126.540 75.965 126.695 ;
        RECT 86.775 126.680 87.095 126.740 ;
        RECT 95.530 126.695 95.820 126.925 ;
        RECT 96.065 126.880 96.205 127.080 ;
        RECT 96.435 127.080 97.200 127.220 ;
        RECT 96.435 127.020 96.755 127.080 ;
        RECT 96.910 127.035 97.200 127.080 ;
        RECT 97.830 127.035 98.120 127.265 ;
        RECT 100.130 127.220 100.420 127.265 ;
        RECT 104.715 127.220 105.035 127.280 ;
        RECT 100.130 127.080 105.035 127.220 ;
        RECT 100.130 127.035 100.420 127.080 ;
        RECT 97.905 126.880 98.045 127.035 ;
        RECT 104.715 127.020 105.035 127.080 ;
        RECT 105.605 127.220 105.895 127.265 ;
        RECT 107.925 127.220 108.140 127.375 ;
        RECT 105.605 127.080 108.140 127.220 ;
        RECT 105.605 127.035 105.895 127.080 ;
        RECT 110.695 127.020 111.015 127.280 ;
        RECT 96.065 126.740 98.045 126.880 ;
        RECT 98.750 126.880 99.040 126.925 ;
        RECT 99.195 126.880 99.515 126.940 ;
        RECT 101.740 126.880 102.030 126.925 ;
        RECT 98.750 126.740 102.030 126.880 ;
        RECT 98.750 126.695 99.040 126.740 ;
        RECT 67.915 126.400 75.965 126.540 ;
        RECT 83.575 126.540 83.865 126.585 ;
        RECT 85.435 126.540 85.725 126.585 ;
        RECT 88.215 126.540 88.505 126.585 ;
        RECT 83.575 126.400 88.505 126.540 ;
        RECT 67.915 126.340 68.235 126.400 ;
        RECT 83.575 126.355 83.865 126.400 ;
        RECT 85.435 126.355 85.725 126.400 ;
        RECT 88.215 126.355 88.505 126.400 ;
        RECT 95.605 126.260 95.745 126.695 ;
        RECT 99.195 126.680 99.515 126.740 ;
        RECT 101.740 126.695 102.030 126.740 ;
        RECT 108.855 126.680 109.175 126.940 ;
        RECT 105.605 126.540 105.895 126.585 ;
        RECT 108.385 126.540 108.675 126.585 ;
        RECT 110.245 126.540 110.535 126.585 ;
        RECT 105.605 126.400 110.535 126.540 ;
        RECT 105.605 126.355 105.895 126.400 ;
        RECT 108.385 126.355 108.675 126.400 ;
        RECT 110.245 126.355 110.535 126.400 ;
        RECT 67.455 126.200 67.775 126.260 ;
        RECT 68.835 126.200 69.155 126.260 ;
        RECT 65.245 126.060 69.155 126.200 ;
        RECT 67.455 126.000 67.775 126.060 ;
        RECT 68.835 126.000 69.155 126.060 ;
        RECT 70.690 126.200 70.980 126.245 ;
        RECT 71.595 126.200 71.915 126.260 ;
        RECT 70.690 126.060 71.915 126.200 ;
        RECT 70.690 126.015 70.980 126.060 ;
        RECT 71.595 126.000 71.915 126.060 ;
        RECT 72.055 126.000 72.375 126.260 ;
        RECT 78.035 126.000 78.355 126.260 ;
        RECT 79.415 126.200 79.735 126.260 ;
        RECT 81.730 126.200 82.020 126.245 ;
        RECT 79.415 126.060 82.020 126.200 ;
        RECT 79.415 126.000 79.735 126.060 ;
        RECT 81.730 126.015 82.020 126.060 ;
        RECT 85.855 126.200 86.175 126.260 ;
        RECT 92.080 126.200 92.370 126.245 ;
        RECT 95.515 126.200 95.835 126.260 ;
        RECT 85.855 126.060 95.835 126.200 ;
        RECT 85.855 126.000 86.175 126.060 ;
        RECT 92.080 126.015 92.370 126.060 ;
        RECT 95.515 126.000 95.835 126.060 ;
        RECT 18.165 125.380 112.465 125.860 ;
        RECT 19.860 125.180 20.150 125.225 ;
        RECT 24.215 125.180 24.535 125.240 ;
        RECT 19.860 125.040 29.045 125.180 ;
        RECT 19.860 124.995 20.150 125.040 ;
        RECT 24.215 124.980 24.535 125.040 ;
        RECT 23.725 124.840 24.015 124.885 ;
        RECT 26.505 124.840 26.795 124.885 ;
        RECT 28.365 124.840 28.655 124.885 ;
        RECT 23.725 124.700 28.655 124.840 ;
        RECT 28.905 124.840 29.045 125.040 ;
        RECT 31.575 124.980 31.895 125.240 ;
        RECT 32.035 124.980 32.355 125.240 ;
        RECT 37.555 124.980 37.875 125.240 ;
        RECT 43.075 125.180 43.395 125.240 ;
        RECT 44.915 125.180 45.235 125.240 ;
        RECT 43.075 125.040 45.235 125.180 ;
        RECT 43.075 124.980 43.395 125.040 ;
        RECT 44.915 124.980 45.235 125.040 ;
        RECT 52.275 125.180 52.595 125.240 ;
        RECT 52.750 125.180 53.040 125.225 ;
        RECT 52.275 125.040 53.040 125.180 ;
        RECT 52.275 124.980 52.595 125.040 ;
        RECT 52.750 124.995 53.040 125.040 ;
        RECT 59.635 125.180 59.955 125.240 ;
        RECT 70.690 125.180 70.980 125.225 ;
        RECT 72.055 125.180 72.375 125.240 ;
        RECT 59.635 125.040 70.445 125.180 ;
        RECT 59.635 124.980 59.955 125.040 ;
        RECT 36.635 124.840 36.955 124.900 ;
        RECT 28.905 124.700 34.105 124.840 ;
        RECT 23.725 124.655 24.015 124.700 ;
        RECT 26.505 124.655 26.795 124.700 ;
        RECT 28.365 124.655 28.655 124.700 ;
        RECT 21.455 124.500 21.775 124.560 ;
        RECT 26.990 124.500 27.280 124.545 ;
        RECT 21.455 124.360 27.280 124.500 ;
        RECT 21.455 124.300 21.775 124.360 ;
        RECT 26.990 124.315 27.280 124.360 ;
        RECT 28.815 124.300 29.135 124.560 ;
        RECT 23.725 124.160 24.015 124.205 ;
        RECT 27.435 124.160 27.755 124.220 ;
        RECT 33.965 124.205 34.105 124.700 ;
        RECT 36.635 124.700 47.905 124.840 ;
        RECT 36.635 124.640 36.955 124.700 ;
        RECT 47.765 124.560 47.905 124.700 ;
        RECT 69.295 124.640 69.615 124.900 ;
        RECT 70.305 124.840 70.445 125.040 ;
        RECT 70.690 125.040 72.375 125.180 ;
        RECT 70.690 124.995 70.980 125.040 ;
        RECT 72.055 124.980 72.375 125.040 ;
        RECT 72.975 124.980 73.295 125.240 ;
        RECT 85.410 125.180 85.700 125.225 ;
        RECT 86.315 125.180 86.635 125.240 ;
        RECT 85.410 125.040 86.635 125.180 ;
        RECT 85.410 124.995 85.700 125.040 ;
        RECT 86.315 124.980 86.635 125.040 ;
        RECT 86.775 124.980 87.095 125.240 ;
        RECT 87.235 125.180 87.555 125.240 ;
        RECT 88.170 125.180 88.460 125.225 ;
        RECT 87.235 125.040 88.460 125.180 ;
        RECT 87.235 124.980 87.555 125.040 ;
        RECT 88.170 124.995 88.460 125.040 ;
        RECT 92.755 125.180 93.075 125.240 ;
        RECT 94.610 125.180 94.900 125.225 ;
        RECT 92.755 125.040 94.900 125.180 ;
        RECT 92.755 124.980 93.075 125.040 ;
        RECT 94.610 124.995 94.900 125.040 ;
        RECT 96.910 125.180 97.200 125.225 ;
        RECT 97.355 125.180 97.675 125.240 ;
        RECT 96.910 125.040 97.675 125.180 ;
        RECT 96.910 124.995 97.200 125.040 ;
        RECT 97.355 124.980 97.675 125.040 ;
        RECT 107.030 125.180 107.320 125.225 ;
        RECT 108.855 125.180 109.175 125.240 ;
        RECT 107.030 125.040 109.175 125.180 ;
        RECT 107.030 124.995 107.320 125.040 ;
        RECT 108.855 124.980 109.175 125.040 ;
        RECT 78.005 124.840 78.295 124.885 ;
        RECT 80.785 124.840 81.075 124.885 ;
        RECT 82.645 124.840 82.935 124.885 ;
        RECT 87.695 124.840 88.015 124.900 ;
        RECT 70.305 124.700 77.805 124.840 ;
        RECT 40.775 124.500 41.095 124.560 ;
        RECT 47.675 124.500 47.995 124.560 ;
        RECT 61.015 124.500 61.335 124.560 ;
        RECT 69.385 124.500 69.525 124.640 ;
        RECT 77.665 124.500 77.805 124.700 ;
        RECT 78.005 124.700 82.935 124.840 ;
        RECT 78.005 124.655 78.295 124.700 ;
        RECT 80.785 124.655 81.075 124.700 ;
        RECT 82.645 124.655 82.935 124.700 ;
        RECT 85.025 124.700 88.015 124.840 ;
        RECT 40.775 124.360 47.445 124.500 ;
        RECT 40.775 124.300 41.095 124.360 ;
        RECT 29.750 124.160 30.040 124.205 ;
        RECT 23.725 124.020 26.260 124.160 ;
        RECT 23.725 123.975 24.015 124.020 ;
        RECT 20.995 123.820 21.315 123.880 ;
        RECT 26.045 123.865 26.260 124.020 ;
        RECT 27.435 124.020 30.040 124.160 ;
        RECT 27.435 123.960 27.755 124.020 ;
        RECT 29.750 123.975 30.040 124.020 ;
        RECT 30.670 124.160 30.960 124.205 ;
        RECT 32.970 124.160 33.260 124.205 ;
        RECT 30.670 124.020 33.260 124.160 ;
        RECT 30.670 123.975 30.960 124.020 ;
        RECT 32.970 123.975 33.260 124.020 ;
        RECT 33.890 124.160 34.180 124.205 ;
        RECT 34.335 124.160 34.655 124.220 ;
        RECT 33.890 124.020 34.655 124.160 ;
        RECT 33.890 123.975 34.180 124.020 ;
        RECT 21.865 123.820 22.155 123.865 ;
        RECT 25.125 123.820 25.415 123.865 ;
        RECT 20.995 123.680 25.415 123.820 ;
        RECT 20.995 123.620 21.315 123.680 ;
        RECT 21.865 123.635 22.155 123.680 ;
        RECT 25.125 123.635 25.415 123.680 ;
        RECT 26.045 123.820 26.335 123.865 ;
        RECT 27.905 123.820 28.195 123.865 ;
        RECT 26.045 123.680 28.195 123.820 ;
        RECT 29.825 123.820 29.965 123.975 ;
        RECT 32.035 123.820 32.355 123.880 ;
        RECT 29.825 123.680 32.355 123.820 ;
        RECT 33.045 123.820 33.185 123.975 ;
        RECT 34.335 123.960 34.655 124.020 ;
        RECT 44.915 123.960 45.235 124.220 ;
        RECT 46.310 124.160 46.600 124.205 ;
        RECT 46.755 124.160 47.075 124.220 ;
        RECT 46.310 124.020 47.075 124.160 ;
        RECT 46.310 123.975 46.600 124.020 ;
        RECT 36.635 123.820 36.955 123.880 ;
        RECT 33.045 123.680 36.955 123.820 ;
        RECT 26.045 123.635 26.335 123.680 ;
        RECT 27.905 123.635 28.195 123.680 ;
        RECT 32.035 123.620 32.355 123.680 ;
        RECT 36.635 123.620 36.955 123.680 ;
        RECT 44.010 123.820 44.300 123.865 ;
        RECT 46.385 123.820 46.525 123.975 ;
        RECT 46.755 123.960 47.075 124.020 ;
        RECT 44.010 123.680 46.525 123.820 ;
        RECT 44.010 123.635 44.300 123.680 ;
        RECT 24.675 123.480 24.995 123.540 ;
        RECT 30.195 123.480 30.515 123.540 ;
        RECT 24.675 123.340 30.515 123.480 ;
        RECT 24.675 123.280 24.995 123.340 ;
        RECT 30.195 123.280 30.515 123.340 ;
        RECT 45.835 123.280 46.155 123.540 ;
        RECT 46.755 123.480 47.075 123.540 ;
        RECT 47.305 123.480 47.445 124.360 ;
        RECT 47.675 124.360 72.285 124.500 ;
        RECT 77.665 124.360 82.865 124.500 ;
        RECT 47.675 124.300 47.995 124.360 ;
        RECT 61.015 124.300 61.335 124.360 ;
        RECT 58.730 124.160 59.020 124.205 ;
        RECT 62.395 124.160 62.715 124.220 ;
        RECT 63.330 124.160 63.620 124.205 ;
        RECT 58.730 124.020 63.620 124.160 ;
        RECT 58.730 123.975 59.020 124.020 ;
        RECT 62.395 123.960 62.715 124.020 ;
        RECT 63.330 123.975 63.620 124.020 ;
        RECT 66.995 124.160 67.315 124.220 ;
        RECT 69.845 124.205 69.985 124.360 ;
        RECT 67.470 124.160 67.760 124.205 ;
        RECT 66.995 124.020 69.065 124.160 ;
        RECT 66.995 123.960 67.315 124.020 ;
        RECT 67.470 123.975 67.760 124.020 ;
        RECT 53.195 123.820 53.515 123.880 ;
        RECT 57.795 123.820 58.115 123.880 ;
        RECT 53.195 123.680 58.115 123.820 ;
        RECT 53.195 123.620 53.515 123.680 ;
        RECT 57.795 123.620 58.115 123.680 ;
        RECT 53.655 123.480 53.975 123.540 ;
        RECT 57.350 123.480 57.640 123.525 ;
        RECT 46.755 123.340 57.640 123.480 ;
        RECT 46.755 123.280 47.075 123.340 ;
        RECT 53.655 123.280 53.975 123.340 ;
        RECT 57.350 123.295 57.640 123.340 ;
        RECT 64.710 123.480 65.000 123.525 ;
        RECT 67.455 123.480 67.775 123.540 ;
        RECT 64.710 123.340 67.775 123.480 ;
        RECT 64.710 123.295 65.000 123.340 ;
        RECT 67.455 123.280 67.775 123.340 ;
        RECT 67.930 123.480 68.220 123.525 ;
        RECT 68.375 123.480 68.695 123.540 ;
        RECT 67.930 123.340 68.695 123.480 ;
        RECT 68.925 123.480 69.065 124.020 ;
        RECT 69.310 123.975 69.600 124.205 ;
        RECT 69.770 123.975 70.060 124.205 ;
        RECT 70.675 124.160 70.995 124.220 ;
        RECT 72.145 124.205 72.285 124.360 ;
        RECT 71.150 124.160 71.440 124.205 ;
        RECT 70.675 124.020 71.440 124.160 ;
        RECT 69.385 123.820 69.525 123.975 ;
        RECT 70.675 123.960 70.995 124.020 ;
        RECT 71.150 123.975 71.440 124.020 ;
        RECT 72.070 123.975 72.360 124.205 ;
        RECT 78.005 124.160 78.295 124.205 ;
        RECT 78.005 124.020 80.540 124.160 ;
        RECT 78.005 123.975 78.295 124.020 ;
        RECT 73.435 123.820 73.755 123.880 ;
        RECT 79.415 123.865 79.735 123.880 ;
        RECT 69.385 123.680 73.755 123.820 ;
        RECT 73.435 123.620 73.755 123.680 ;
        RECT 76.145 123.820 76.435 123.865 ;
        RECT 79.405 123.820 79.735 123.865 ;
        RECT 76.145 123.680 79.735 123.820 ;
        RECT 76.145 123.635 76.435 123.680 ;
        RECT 79.405 123.635 79.735 123.680 ;
        RECT 80.325 123.865 80.540 124.020 ;
        RECT 81.255 123.960 81.575 124.220 ;
        RECT 80.325 123.820 80.615 123.865 ;
        RECT 82.185 123.820 82.475 123.865 ;
        RECT 80.325 123.680 82.475 123.820 ;
        RECT 82.725 123.820 82.865 124.360 ;
        RECT 83.095 124.300 83.415 124.560 ;
        RECT 85.025 124.205 85.165 124.700 ;
        RECT 87.695 124.640 88.015 124.700 ;
        RECT 95.515 124.840 95.835 124.900 ;
        RECT 95.515 124.700 100.805 124.840 ;
        RECT 95.515 124.640 95.835 124.700 ;
        RECT 92.755 124.500 93.075 124.560 ;
        RECT 94.595 124.500 94.915 124.560 ;
        RECT 98.275 124.500 98.595 124.560 ;
        RECT 86.405 124.360 96.665 124.500 ;
        RECT 84.950 123.975 85.240 124.205 ;
        RECT 86.405 123.820 86.545 124.360 ;
        RECT 87.235 124.160 87.555 124.220 ;
        RECT 89.165 124.205 89.305 124.360 ;
        RECT 92.755 124.300 93.075 124.360 ;
        RECT 94.595 124.300 94.915 124.360 ;
        RECT 95.605 124.205 95.745 124.360 ;
        RECT 87.710 124.160 88.000 124.205 ;
        RECT 87.235 124.020 88.000 124.160 ;
        RECT 87.235 123.960 87.555 124.020 ;
        RECT 87.710 123.975 88.000 124.020 ;
        RECT 89.090 123.975 89.380 124.205 ;
        RECT 89.550 123.975 89.840 124.205 ;
        RECT 95.530 123.975 95.820 124.205 ;
        RECT 82.725 123.680 86.545 123.820 ;
        RECT 86.775 123.820 87.095 123.880 ;
        RECT 89.625 123.820 89.765 123.975 ;
        RECT 95.975 123.960 96.295 124.220 ;
        RECT 96.525 124.160 96.665 124.360 ;
        RECT 98.275 124.360 99.885 124.500 ;
        RECT 98.275 124.300 98.595 124.360 ;
        RECT 97.730 124.160 98.020 124.205 ;
        RECT 96.525 124.020 98.020 124.160 ;
        RECT 97.730 123.975 98.020 124.020 ;
        RECT 98.750 123.975 99.040 124.205 ;
        RECT 99.745 124.160 99.885 124.360 ;
        RECT 100.115 124.300 100.435 124.560 ;
        RECT 100.665 124.545 100.805 124.700 ;
        RECT 100.590 124.315 100.880 124.545 ;
        RECT 104.270 124.160 104.560 124.205 ;
        RECT 99.745 124.020 104.560 124.160 ;
        RECT 104.270 123.975 104.560 124.020 ;
        RECT 106.110 123.975 106.400 124.205 ;
        RECT 86.775 123.680 89.765 123.820 ;
        RECT 98.825 123.820 98.965 123.975 ;
        RECT 102.415 123.820 102.735 123.880 ;
        RECT 106.185 123.820 106.325 123.975 ;
        RECT 98.825 123.680 102.735 123.820 ;
        RECT 80.325 123.635 80.615 123.680 ;
        RECT 82.185 123.635 82.475 123.680 ;
        RECT 79.415 123.620 79.735 123.635 ;
        RECT 86.775 123.620 87.095 123.680 ;
        RECT 102.415 123.620 102.735 123.680 ;
        RECT 102.965 123.680 106.325 123.820 ;
        RECT 72.515 123.480 72.835 123.540 ;
        RECT 68.925 123.340 72.835 123.480 ;
        RECT 67.930 123.295 68.220 123.340 ;
        RECT 68.375 123.280 68.695 123.340 ;
        RECT 72.515 123.280 72.835 123.340 ;
        RECT 74.140 123.480 74.430 123.525 ;
        RECT 74.815 123.480 75.135 123.540 ;
        RECT 74.140 123.340 75.135 123.480 ;
        RECT 74.140 123.295 74.430 123.340 ;
        RECT 74.815 123.280 75.135 123.340 ;
        RECT 99.195 123.480 99.515 123.540 ;
        RECT 102.965 123.525 103.105 123.680 ;
        RECT 101.050 123.480 101.340 123.525 ;
        RECT 99.195 123.340 101.340 123.480 ;
        RECT 99.195 123.280 99.515 123.340 ;
        RECT 101.050 123.295 101.340 123.340 ;
        RECT 102.890 123.295 103.180 123.525 ;
        RECT 105.190 123.480 105.480 123.525 ;
        RECT 107.015 123.480 107.335 123.540 ;
        RECT 105.190 123.340 107.335 123.480 ;
        RECT 105.190 123.295 105.480 123.340 ;
        RECT 107.015 123.280 107.335 123.340 ;
        RECT 17.370 122.660 112.465 123.140 ;
        RECT 20.995 122.260 21.315 122.520 ;
        RECT 22.835 122.505 23.155 122.520 ;
        RECT 22.620 122.460 23.155 122.505 ;
        RECT 31.575 122.460 31.895 122.520 ;
        RECT 22.620 122.320 31.895 122.460 ;
        RECT 22.620 122.275 23.155 122.320 ;
        RECT 22.835 122.260 23.155 122.275 ;
        RECT 31.575 122.260 31.895 122.320 ;
        RECT 32.035 122.460 32.355 122.520 ;
        RECT 33.890 122.460 34.180 122.505 ;
        RECT 32.035 122.320 34.180 122.460 ;
        RECT 32.035 122.260 32.355 122.320 ;
        RECT 33.890 122.275 34.180 122.320 ;
        RECT 34.335 122.260 34.655 122.520 ;
        RECT 35.255 122.460 35.575 122.520 ;
        RECT 36.190 122.460 36.480 122.505 ;
        RECT 35.255 122.320 36.480 122.460 ;
        RECT 35.255 122.260 35.575 122.320 ;
        RECT 36.190 122.275 36.480 122.320 ;
        RECT 43.075 122.260 43.395 122.520 ;
        RECT 43.550 122.460 43.840 122.505 ;
        RECT 44.915 122.460 45.235 122.520 ;
        RECT 43.550 122.320 45.235 122.460 ;
        RECT 43.550 122.275 43.840 122.320 ;
        RECT 44.915 122.260 45.235 122.320 ;
        RECT 51.355 122.460 51.675 122.520 ;
        RECT 52.290 122.460 52.580 122.505 ;
        RECT 51.355 122.320 52.580 122.460 ;
        RECT 51.355 122.260 51.675 122.320 ;
        RECT 52.290 122.275 52.580 122.320 ;
        RECT 52.735 122.460 53.055 122.520 ;
        RECT 54.130 122.460 54.420 122.505 ;
        RECT 55.035 122.460 55.355 122.520 ;
        RECT 52.735 122.320 53.885 122.460 ;
        RECT 52.735 122.260 53.055 122.320 ;
        RECT 23.755 122.120 24.075 122.180 ;
        RECT 24.625 122.120 24.915 122.165 ;
        RECT 27.885 122.120 28.175 122.165 ;
        RECT 23.755 121.980 28.175 122.120 ;
        RECT 23.755 121.920 24.075 121.980 ;
        RECT 24.625 121.935 24.915 121.980 ;
        RECT 27.885 121.935 28.175 121.980 ;
        RECT 28.805 122.120 29.095 122.165 ;
        RECT 30.665 122.120 30.955 122.165 ;
        RECT 28.805 121.980 30.955 122.120 ;
        RECT 28.805 121.935 29.095 121.980 ;
        RECT 30.665 121.935 30.955 121.980 ;
        RECT 31.115 122.120 31.435 122.180 ;
        RECT 34.795 122.120 35.115 122.180 ;
        RECT 37.555 122.120 37.875 122.180 ;
        RECT 40.790 122.120 41.080 122.165 ;
        RECT 49.530 122.120 49.820 122.165 ;
        RECT 53.745 122.120 53.885 122.320 ;
        RECT 54.130 122.320 55.355 122.460 ;
        RECT 54.130 122.275 54.420 122.320 ;
        RECT 55.035 122.260 55.355 122.320 ;
        RECT 79.890 122.460 80.180 122.505 ;
        RECT 81.255 122.460 81.575 122.520 ;
        RECT 79.890 122.320 81.575 122.460 ;
        RECT 79.890 122.275 80.180 122.320 ;
        RECT 81.255 122.260 81.575 122.320 ;
        RECT 85.410 122.460 85.700 122.505 ;
        RECT 85.855 122.460 86.175 122.520 ;
        RECT 85.410 122.320 86.175 122.460 ;
        RECT 85.410 122.275 85.700 122.320 ;
        RECT 85.855 122.260 86.175 122.320 ;
        RECT 87.235 122.260 87.555 122.520 ;
        RECT 93.690 122.460 93.980 122.505 ;
        RECT 96.895 122.460 97.215 122.520 ;
        RECT 93.690 122.320 97.215 122.460 ;
        RECT 93.690 122.275 93.980 122.320 ;
        RECT 96.895 122.260 97.215 122.320 ;
        RECT 99.195 122.460 99.515 122.520 ;
        RECT 101.970 122.460 102.260 122.505 ;
        RECT 99.195 122.320 102.260 122.460 ;
        RECT 99.195 122.260 99.515 122.320 ;
        RECT 101.970 122.275 102.260 122.320 ;
        RECT 54.590 122.120 54.880 122.165 ;
        RECT 31.115 121.980 41.080 122.120 ;
        RECT 21.470 121.780 21.760 121.825 ;
        RECT 25.595 121.780 25.915 121.840 ;
        RECT 21.470 121.640 25.915 121.780 ;
        RECT 21.470 121.595 21.760 121.640 ;
        RECT 25.595 121.580 25.915 121.640 ;
        RECT 26.485 121.780 26.775 121.825 ;
        RECT 28.805 121.780 29.020 121.935 ;
        RECT 31.115 121.920 31.435 121.980 ;
        RECT 34.795 121.920 35.115 121.980 ;
        RECT 37.555 121.920 37.875 121.980 ;
        RECT 40.790 121.935 41.080 121.980 ;
        RECT 41.785 121.980 49.285 122.120 ;
        RECT 26.485 121.640 29.020 121.780 ;
        RECT 26.485 121.595 26.775 121.640 ;
        RECT 29.735 121.580 30.055 121.840 ;
        RECT 30.195 121.780 30.515 121.840 ;
        RECT 37.110 121.780 37.400 121.825 ;
        RECT 38.015 121.780 38.335 121.840 ;
        RECT 30.195 121.770 31.345 121.780 ;
        RECT 31.665 121.770 32.495 121.780 ;
        RECT 30.195 121.640 32.495 121.770 ;
        RECT 30.195 121.580 30.515 121.640 ;
        RECT 31.205 121.630 31.805 121.640 ;
        RECT 28.815 121.440 29.135 121.500 ;
        RECT 30.655 121.440 30.975 121.500 ;
        RECT 31.590 121.440 31.880 121.485 ;
        RECT 28.815 121.300 31.880 121.440 ;
        RECT 32.355 121.440 32.495 121.640 ;
        RECT 37.110 121.640 38.335 121.780 ;
        RECT 37.110 121.595 37.400 121.640 ;
        RECT 38.015 121.580 38.335 121.640 ;
        RECT 38.490 121.780 38.780 121.825 ;
        RECT 41.785 121.780 41.925 121.980 ;
        RECT 38.490 121.640 41.925 121.780 ;
        RECT 38.490 121.595 38.780 121.640 ;
        RECT 42.170 121.595 42.460 121.825 ;
        RECT 43.995 121.780 44.315 121.840 ;
        RECT 45.390 121.780 45.680 121.825 ;
        RECT 43.995 121.640 45.680 121.780 ;
        RECT 35.255 121.440 35.575 121.500 ;
        RECT 32.355 121.300 35.575 121.440 ;
        RECT 28.815 121.240 29.135 121.300 ;
        RECT 30.655 121.240 30.975 121.300 ;
        RECT 31.590 121.255 31.880 121.300 ;
        RECT 35.255 121.240 35.575 121.300 ;
        RECT 36.635 121.440 36.955 121.500 ;
        RECT 38.565 121.440 38.705 121.595 ;
        RECT 36.635 121.300 38.705 121.440 ;
        RECT 36.635 121.240 36.955 121.300 ;
        RECT 41.250 121.255 41.540 121.485 ;
        RECT 42.245 121.440 42.385 121.595 ;
        RECT 43.995 121.580 44.315 121.640 ;
        RECT 45.390 121.595 45.680 121.640 ;
        RECT 45.850 121.780 46.140 121.825 ;
        RECT 48.595 121.780 48.915 121.840 ;
        RECT 49.145 121.825 49.285 121.980 ;
        RECT 49.530 121.980 53.425 122.120 ;
        RECT 53.745 121.980 54.880 122.120 ;
        RECT 49.530 121.935 49.820 121.980 ;
        RECT 45.850 121.640 48.915 121.780 ;
        RECT 45.850 121.595 46.140 121.640 ;
        RECT 48.595 121.580 48.915 121.640 ;
        RECT 49.070 121.780 49.360 121.825 ;
        RECT 49.070 121.640 51.125 121.780 ;
        RECT 49.070 121.595 49.360 121.640 ;
        RECT 42.245 121.300 44.225 121.440 ;
        RECT 26.485 121.100 26.775 121.145 ;
        RECT 29.265 121.100 29.555 121.145 ;
        RECT 31.125 121.100 31.415 121.145 ;
        RECT 41.325 121.100 41.465 121.255 ;
        RECT 43.535 121.100 43.855 121.160 ;
        RECT 26.485 120.960 31.415 121.100 ;
        RECT 26.485 120.915 26.775 120.960 ;
        RECT 29.265 120.915 29.555 120.960 ;
        RECT 31.125 120.915 31.415 120.960 ;
        RECT 31.665 120.960 43.855 121.100 ;
        RECT 44.085 121.100 44.225 121.300 ;
        RECT 46.755 121.240 47.075 121.500 ;
        RECT 50.450 121.255 50.740 121.485 ;
        RECT 50.985 121.440 51.125 121.640 ;
        RECT 51.355 121.580 51.675 121.840 ;
        RECT 51.815 121.780 52.135 121.840 ;
        RECT 52.735 121.780 53.055 121.840 ;
        RECT 51.815 121.640 53.055 121.780 ;
        RECT 53.285 121.780 53.425 121.980 ;
        RECT 54.590 121.935 54.880 121.980 ;
        RECT 57.795 121.920 58.115 122.180 ;
        RECT 64.715 122.120 65.005 122.165 ;
        RECT 66.575 122.120 66.865 122.165 ;
        RECT 64.715 121.980 66.865 122.120 ;
        RECT 64.715 121.935 65.005 121.980 ;
        RECT 66.575 121.935 66.865 121.980 ;
        RECT 67.495 122.120 67.785 122.165 ;
        RECT 68.375 122.120 68.695 122.180 ;
        RECT 70.755 122.120 71.045 122.165 ;
        RECT 67.495 121.980 71.045 122.120 ;
        RECT 67.495 121.935 67.785 121.980 ;
        RECT 59.190 121.780 59.480 121.825 ;
        RECT 61.015 121.780 61.335 121.840 ;
        RECT 63.315 121.780 63.635 121.840 ;
        RECT 53.285 121.640 54.345 121.780 ;
        RECT 51.815 121.580 52.135 121.640 ;
        RECT 52.735 121.580 53.055 121.640 ;
        RECT 53.195 121.440 53.515 121.500 ;
        RECT 50.985 121.300 53.515 121.440 ;
        RECT 47.675 121.100 47.995 121.160 ;
        RECT 44.085 120.960 47.995 121.100 ;
        RECT 50.525 121.100 50.665 121.255 ;
        RECT 53.195 121.240 53.515 121.300 ;
        RECT 53.655 121.240 53.975 121.500 ;
        RECT 54.205 121.440 54.345 121.640 ;
        RECT 59.190 121.640 63.635 121.780 ;
        RECT 59.190 121.595 59.480 121.640 ;
        RECT 61.015 121.580 61.335 121.640 ;
        RECT 63.315 121.580 63.635 121.640 ;
        RECT 63.775 121.580 64.095 121.840 ;
        RECT 66.650 121.780 66.865 121.935 ;
        RECT 68.375 121.920 68.695 121.980 ;
        RECT 70.755 121.935 71.045 121.980 ;
        RECT 74.815 122.120 75.135 122.180 ;
        RECT 84.950 122.120 85.240 122.165 ;
        RECT 95.990 122.120 96.280 122.165 ;
        RECT 74.815 121.980 85.240 122.120 ;
        RECT 74.815 121.920 75.135 121.980 ;
        RECT 84.950 121.935 85.240 121.980 ;
        RECT 91.925 121.980 96.280 122.120 ;
        RECT 68.895 121.780 69.185 121.825 ;
        RECT 66.650 121.640 69.185 121.780 ;
        RECT 68.895 121.595 69.185 121.640 ;
        RECT 72.975 121.780 73.295 121.840 ;
        RECT 75.290 121.780 75.580 121.825 ;
        RECT 72.975 121.640 75.580 121.780 ;
        RECT 72.975 121.580 73.295 121.640 ;
        RECT 75.290 121.595 75.580 121.640 ;
        RECT 78.035 121.780 78.355 121.840 ;
        RECT 78.970 121.780 79.260 121.825 ;
        RECT 78.035 121.640 79.260 121.780 ;
        RECT 78.035 121.580 78.355 121.640 ;
        RECT 78.970 121.595 79.260 121.640 ;
        RECT 87.235 121.780 87.555 121.840 ;
        RECT 91.925 121.825 92.065 121.980 ;
        RECT 95.990 121.935 96.280 121.980 ;
        RECT 89.550 121.780 89.840 121.825 ;
        RECT 91.850 121.780 92.140 121.825 ;
        RECT 87.235 121.640 89.840 121.780 ;
        RECT 87.235 121.580 87.555 121.640 ;
        RECT 89.550 121.595 89.840 121.640 ;
        RECT 90.085 121.640 92.140 121.780 ;
        RECT 90.085 121.500 90.225 121.640 ;
        RECT 91.850 121.595 92.140 121.640 ;
        RECT 92.755 121.580 93.075 121.840 ;
        RECT 102.415 121.580 102.735 121.840 ;
        RECT 104.715 121.580 105.035 121.840 ;
        RECT 106.570 121.595 106.860 121.825 ;
        RECT 54.575 121.440 54.895 121.500 ;
        RECT 54.205 121.300 54.895 121.440 ;
        RECT 54.575 121.240 54.895 121.300 ;
        RECT 65.630 121.440 65.920 121.485 ;
        RECT 75.735 121.440 76.055 121.500 ;
        RECT 84.030 121.440 84.320 121.485 ;
        RECT 65.630 121.300 74.585 121.440 ;
        RECT 65.630 121.255 65.920 121.300 ;
        RECT 55.035 121.100 55.355 121.160 ;
        RECT 50.525 120.960 55.355 121.100 ;
        RECT 31.665 120.820 31.805 120.960 ;
        RECT 43.535 120.900 43.855 120.960 ;
        RECT 47.675 120.900 47.995 120.960 ;
        RECT 55.035 120.900 55.355 120.960 ;
        RECT 56.430 121.100 56.720 121.145 ;
        RECT 59.635 121.100 59.955 121.160 ;
        RECT 56.430 120.960 59.955 121.100 ;
        RECT 56.430 120.915 56.720 120.960 ;
        RECT 59.635 120.900 59.955 120.960 ;
        RECT 64.255 121.100 64.545 121.145 ;
        RECT 66.115 121.100 66.405 121.145 ;
        RECT 68.895 121.100 69.185 121.145 ;
        RECT 64.255 120.960 69.185 121.100 ;
        RECT 64.255 120.915 64.545 120.960 ;
        RECT 66.115 120.915 66.405 120.960 ;
        RECT 68.895 120.915 69.185 120.960 ;
        RECT 71.595 121.100 71.915 121.160 ;
        RECT 74.445 121.145 74.585 121.300 ;
        RECT 75.735 121.300 84.320 121.440 ;
        RECT 75.735 121.240 76.055 121.300 ;
        RECT 84.030 121.255 84.320 121.300 ;
        RECT 71.595 120.960 73.665 121.100 ;
        RECT 71.595 120.900 71.915 120.960 ;
        RECT 26.975 120.760 27.295 120.820 ;
        RECT 29.735 120.760 30.055 120.820 ;
        RECT 26.975 120.620 30.055 120.760 ;
        RECT 26.975 120.560 27.295 120.620 ;
        RECT 29.735 120.560 30.055 120.620 ;
        RECT 31.575 120.560 31.895 120.820 ;
        RECT 32.035 120.560 32.355 120.820 ;
        RECT 38.475 120.760 38.795 120.820 ;
        RECT 38.950 120.760 39.240 120.805 ;
        RECT 38.475 120.620 39.240 120.760 ;
        RECT 38.475 120.560 38.795 120.620 ;
        RECT 38.950 120.575 39.240 120.620 ;
        RECT 52.275 120.760 52.595 120.820 ;
        RECT 63.775 120.760 64.095 120.820 ;
        RECT 52.275 120.620 64.095 120.760 ;
        RECT 52.275 120.560 52.595 120.620 ;
        RECT 63.775 120.560 64.095 120.620 ;
        RECT 70.675 120.760 70.995 120.820 ;
        RECT 72.760 120.760 73.050 120.805 ;
        RECT 70.675 120.620 73.050 120.760 ;
        RECT 73.525 120.760 73.665 120.960 ;
        RECT 74.370 120.915 74.660 121.145 ;
        RECT 84.105 121.100 84.245 121.255 ;
        RECT 89.995 121.240 90.315 121.500 ;
        RECT 90.470 121.440 90.760 121.485 ;
        RECT 94.595 121.440 94.915 121.500 ;
        RECT 90.470 121.300 94.915 121.440 ;
        RECT 90.470 121.255 90.760 121.300 ;
        RECT 90.545 121.100 90.685 121.255 ;
        RECT 94.595 121.240 94.915 121.300 ;
        RECT 95.530 121.440 95.820 121.485 ;
        RECT 95.975 121.440 96.295 121.500 ;
        RECT 95.530 121.300 96.295 121.440 ;
        RECT 95.530 121.255 95.820 121.300 ;
        RECT 95.975 121.240 96.295 121.300 ;
        RECT 101.050 121.255 101.340 121.485 ;
        RECT 106.645 121.440 106.785 121.595 ;
        RECT 104.345 121.300 106.785 121.440 ;
        RECT 84.105 120.960 90.685 121.100 ;
        RECT 94.685 121.100 94.825 121.240 ;
        RECT 100.115 121.100 100.435 121.160 ;
        RECT 101.125 121.100 101.265 121.255 ;
        RECT 104.345 121.145 104.485 121.300 ;
        RECT 94.685 120.960 101.265 121.100 ;
        RECT 100.115 120.900 100.435 120.960 ;
        RECT 104.270 120.915 104.560 121.145 ;
        RECT 81.255 120.760 81.575 120.820 ;
        RECT 73.525 120.620 81.575 120.760 ;
        RECT 70.675 120.560 70.995 120.620 ;
        RECT 72.760 120.575 73.050 120.620 ;
        RECT 81.255 120.560 81.575 120.620 ;
        RECT 87.695 120.560 88.015 120.820 ;
        RECT 97.355 120.760 97.675 120.820 ;
        RECT 97.830 120.760 98.120 120.805 ;
        RECT 97.355 120.620 98.120 120.760 ;
        RECT 97.355 120.560 97.675 120.620 ;
        RECT 97.830 120.575 98.120 120.620 ;
        RECT 105.175 120.560 105.495 120.820 ;
        RECT 107.490 120.760 107.780 120.805 ;
        RECT 108.855 120.760 109.175 120.820 ;
        RECT 107.490 120.620 109.175 120.760 ;
        RECT 107.490 120.575 107.780 120.620 ;
        RECT 108.855 120.560 109.175 120.620 ;
        RECT 18.165 119.940 112.465 120.420 ;
        RECT 46.755 119.740 47.075 119.800 ;
        RECT 44.545 119.600 47.075 119.740 ;
        RECT 24.675 119.400 24.995 119.460 ;
        RECT 22.005 119.260 24.995 119.400 ;
        RECT 22.005 119.105 22.145 119.260 ;
        RECT 24.675 119.200 24.995 119.260 ;
        RECT 26.055 119.400 26.375 119.460 ;
        RECT 29.245 119.400 29.535 119.445 ;
        RECT 32.025 119.400 32.315 119.445 ;
        RECT 33.885 119.400 34.175 119.445 ;
        RECT 26.055 119.260 28.125 119.400 ;
        RECT 26.055 119.200 26.375 119.260 ;
        RECT 21.930 118.875 22.220 119.105 ;
        RECT 22.390 119.060 22.680 119.105 ;
        RECT 25.380 119.060 25.670 119.105 ;
        RECT 27.435 119.060 27.755 119.120 ;
        RECT 22.390 118.920 27.755 119.060 ;
        RECT 27.985 119.060 28.125 119.260 ;
        RECT 29.245 119.260 34.175 119.400 ;
        RECT 29.245 119.215 29.535 119.260 ;
        RECT 32.025 119.215 32.315 119.260 ;
        RECT 33.885 119.215 34.175 119.260 ;
        RECT 34.350 119.060 34.640 119.105 ;
        RECT 34.795 119.060 35.115 119.120 ;
        RECT 27.985 118.920 34.105 119.060 ;
        RECT 22.390 118.875 22.680 118.920 ;
        RECT 25.380 118.875 25.670 118.920 ;
        RECT 27.435 118.860 27.755 118.920 ;
        RECT 22.835 118.520 23.155 118.780 ;
        RECT 29.245 118.720 29.535 118.765 ;
        RECT 32.510 118.720 32.800 118.765 ;
        RECT 32.955 118.720 33.275 118.780 ;
        RECT 29.245 118.580 31.780 118.720 ;
        RECT 29.245 118.535 29.535 118.580 ;
        RECT 27.435 118.425 27.755 118.440 ;
        RECT 31.565 118.425 31.780 118.580 ;
        RECT 32.510 118.580 33.275 118.720 ;
        RECT 33.965 118.720 34.105 118.920 ;
        RECT 34.350 118.920 35.115 119.060 ;
        RECT 34.350 118.875 34.640 118.920 ;
        RECT 34.795 118.860 35.115 118.920 ;
        RECT 35.255 119.060 35.575 119.120 ;
        RECT 40.330 119.060 40.620 119.105 ;
        RECT 44.545 119.060 44.685 119.600 ;
        RECT 46.755 119.540 47.075 119.600 ;
        RECT 48.595 119.740 48.915 119.800 ;
        RECT 51.140 119.740 51.430 119.785 ;
        RECT 51.815 119.740 52.135 119.800 ;
        RECT 48.595 119.600 52.135 119.740 ;
        RECT 48.595 119.540 48.915 119.600 ;
        RECT 51.140 119.555 51.430 119.600 ;
        RECT 51.815 119.540 52.135 119.600 ;
        RECT 63.560 119.740 63.850 119.785 ;
        RECT 67.915 119.740 68.235 119.800 ;
        RECT 63.560 119.600 68.235 119.740 ;
        RECT 63.560 119.555 63.850 119.600 ;
        RECT 67.915 119.540 68.235 119.600 ;
        RECT 72.975 119.540 73.295 119.800 ;
        RECT 89.995 119.785 90.315 119.800 ;
        RECT 89.780 119.555 90.315 119.785 ;
        RECT 101.740 119.740 102.030 119.785 ;
        RECT 102.415 119.740 102.735 119.800 ;
        RECT 101.740 119.600 102.735 119.740 ;
        RECT 101.740 119.555 102.030 119.600 ;
        RECT 89.995 119.540 90.315 119.555 ;
        RECT 102.415 119.540 102.735 119.600 ;
        RECT 45.345 119.400 45.635 119.445 ;
        RECT 48.125 119.400 48.415 119.445 ;
        RECT 49.985 119.400 50.275 119.445 ;
        RECT 45.345 119.260 50.275 119.400 ;
        RECT 45.345 119.215 45.635 119.260 ;
        RECT 48.125 119.215 48.415 119.260 ;
        RECT 49.985 119.215 50.275 119.260 ;
        RECT 55.005 119.400 55.295 119.445 ;
        RECT 57.785 119.400 58.075 119.445 ;
        RECT 59.645 119.400 59.935 119.445 ;
        RECT 61.030 119.400 61.320 119.445 ;
        RECT 55.005 119.260 59.935 119.400 ;
        RECT 55.005 119.215 55.295 119.260 ;
        RECT 57.785 119.215 58.075 119.260 ;
        RECT 59.645 119.215 59.935 119.260 ;
        RECT 60.185 119.260 61.320 119.400 ;
        RECT 35.255 118.920 44.685 119.060 ;
        RECT 45.835 119.060 46.155 119.120 ;
        RECT 48.610 119.060 48.900 119.105 ;
        RECT 45.835 118.920 48.900 119.060 ;
        RECT 35.255 118.860 35.575 118.920 ;
        RECT 40.330 118.875 40.620 118.920 ;
        RECT 45.835 118.860 46.155 118.920 ;
        RECT 48.610 118.875 48.900 118.920 ;
        RECT 50.450 119.060 50.740 119.105 ;
        RECT 52.275 119.060 52.595 119.120 ;
        RECT 60.185 119.060 60.325 119.260 ;
        RECT 61.030 119.215 61.320 119.260 ;
        RECT 67.425 119.400 67.715 119.445 ;
        RECT 70.205 119.400 70.495 119.445 ;
        RECT 72.065 119.400 72.355 119.445 ;
        RECT 67.425 119.260 72.355 119.400 ;
        RECT 67.425 119.215 67.715 119.260 ;
        RECT 70.205 119.215 70.495 119.260 ;
        RECT 72.065 119.215 72.355 119.260 ;
        RECT 93.645 119.400 93.935 119.445 ;
        RECT 96.425 119.400 96.715 119.445 ;
        RECT 98.285 119.400 98.575 119.445 ;
        RECT 93.645 119.260 98.575 119.400 ;
        RECT 93.645 119.215 93.935 119.260 ;
        RECT 96.425 119.215 96.715 119.260 ;
        RECT 98.285 119.215 98.575 119.260 ;
        RECT 105.605 119.400 105.895 119.445 ;
        RECT 108.385 119.400 108.675 119.445 ;
        RECT 110.245 119.400 110.535 119.445 ;
        RECT 105.605 119.260 110.535 119.400 ;
        RECT 105.605 119.215 105.895 119.260 ;
        RECT 108.385 119.215 108.675 119.260 ;
        RECT 110.245 119.215 110.535 119.260 ;
        RECT 63.775 119.060 64.095 119.120 ;
        RECT 50.450 118.920 52.595 119.060 ;
        RECT 50.450 118.875 50.740 118.920 ;
        RECT 52.275 118.860 52.595 118.920 ;
        RECT 58.345 118.920 60.325 119.060 ;
        RECT 61.565 118.920 64.095 119.060 ;
        RECT 36.635 118.720 36.955 118.780 ;
        RECT 33.965 118.580 36.955 118.720 ;
        RECT 32.510 118.535 32.800 118.580 ;
        RECT 32.955 118.520 33.275 118.580 ;
        RECT 36.635 118.520 36.955 118.580 ;
        RECT 39.410 118.720 39.700 118.765 ;
        RECT 41.480 118.720 41.770 118.765 ;
        RECT 43.995 118.720 44.315 118.780 ;
        RECT 58.345 118.765 58.485 118.920 ;
        RECT 39.410 118.580 44.315 118.720 ;
        RECT 39.410 118.535 39.700 118.580 ;
        RECT 41.480 118.535 41.770 118.580 ;
        RECT 43.995 118.520 44.315 118.580 ;
        RECT 45.345 118.720 45.635 118.765 ;
        RECT 55.005 118.720 55.295 118.765 ;
        RECT 45.345 118.580 47.880 118.720 ;
        RECT 45.345 118.535 45.635 118.580 ;
        RECT 27.385 118.380 27.755 118.425 ;
        RECT 30.645 118.380 30.935 118.425 ;
        RECT 27.385 118.240 30.935 118.380 ;
        RECT 27.385 118.195 27.755 118.240 ;
        RECT 30.645 118.195 30.935 118.240 ;
        RECT 31.565 118.380 31.855 118.425 ;
        RECT 33.425 118.380 33.715 118.425 ;
        RECT 31.565 118.240 33.715 118.380 ;
        RECT 31.565 118.195 31.855 118.240 ;
        RECT 33.425 118.195 33.715 118.240 ;
        RECT 38.475 118.380 38.795 118.440 ;
        RECT 47.665 118.425 47.880 118.580 ;
        RECT 55.005 118.580 57.540 118.720 ;
        RECT 55.005 118.535 55.295 118.580 ;
        RECT 43.485 118.380 43.775 118.425 ;
        RECT 46.745 118.380 47.035 118.425 ;
        RECT 38.475 118.240 47.035 118.380 ;
        RECT 27.435 118.180 27.755 118.195 ;
        RECT 38.475 118.180 38.795 118.240 ;
        RECT 43.485 118.195 43.775 118.240 ;
        RECT 46.745 118.195 47.035 118.240 ;
        RECT 47.665 118.380 47.955 118.425 ;
        RECT 49.525 118.380 49.815 118.425 ;
        RECT 47.665 118.240 49.815 118.380 ;
        RECT 47.665 118.195 47.955 118.240 ;
        RECT 49.525 118.195 49.815 118.240 ;
        RECT 53.145 118.380 53.435 118.425 ;
        RECT 54.575 118.380 54.895 118.440 ;
        RECT 57.325 118.425 57.540 118.580 ;
        RECT 58.270 118.535 58.560 118.765 ;
        RECT 60.110 118.720 60.400 118.765 ;
        RECT 61.565 118.720 61.705 118.920 ;
        RECT 63.775 118.860 64.095 118.920 ;
        RECT 71.135 119.060 71.455 119.120 ;
        RECT 72.530 119.060 72.820 119.105 ;
        RECT 71.135 118.920 72.820 119.060 ;
        RECT 71.135 118.860 71.455 118.920 ;
        RECT 72.530 118.875 72.820 118.920 ;
        RECT 73.435 119.060 73.755 119.120 ;
        RECT 75.290 119.060 75.580 119.105 ;
        RECT 73.435 118.920 75.580 119.060 ;
        RECT 73.435 118.860 73.755 118.920 ;
        RECT 75.290 118.875 75.580 118.920 ;
        RECT 75.735 119.060 76.055 119.120 ;
        RECT 81.270 119.060 81.560 119.105 ;
        RECT 75.735 118.920 81.560 119.060 ;
        RECT 60.110 118.580 61.705 118.720 ;
        RECT 60.110 118.535 60.400 118.580 ;
        RECT 61.950 118.535 62.240 118.765 ;
        RECT 67.425 118.720 67.715 118.765 ;
        RECT 70.690 118.720 70.980 118.765 ;
        RECT 72.055 118.720 72.375 118.780 ;
        RECT 67.425 118.580 69.960 118.720 ;
        RECT 67.425 118.535 67.715 118.580 ;
        RECT 56.405 118.380 56.695 118.425 ;
        RECT 53.145 118.240 56.695 118.380 ;
        RECT 53.145 118.195 53.435 118.240 ;
        RECT 54.575 118.180 54.895 118.240 ;
        RECT 56.405 118.195 56.695 118.240 ;
        RECT 57.325 118.380 57.615 118.425 ;
        RECT 59.185 118.380 59.475 118.425 ;
        RECT 57.325 118.240 59.475 118.380 ;
        RECT 57.325 118.195 57.615 118.240 ;
        RECT 59.185 118.195 59.475 118.240 ;
        RECT 59.635 118.380 59.955 118.440 ;
        RECT 62.025 118.380 62.165 118.535 ;
        RECT 59.635 118.240 62.165 118.380 ;
        RECT 65.565 118.380 65.855 118.425 ;
        RECT 66.535 118.380 66.855 118.440 ;
        RECT 69.745 118.425 69.960 118.580 ;
        RECT 70.690 118.580 72.375 118.720 ;
        RECT 75.365 118.720 75.505 118.875 ;
        RECT 75.735 118.860 76.055 118.920 ;
        RECT 81.270 118.875 81.560 118.920 ;
        RECT 88.245 118.920 96.665 119.060 ;
        RECT 88.245 118.765 88.385 118.920 ;
        RECT 80.350 118.720 80.640 118.765 ;
        RECT 75.365 118.580 80.640 118.720 ;
        RECT 70.690 118.535 70.980 118.580 ;
        RECT 72.055 118.520 72.375 118.580 ;
        RECT 80.350 118.535 80.640 118.580 ;
        RECT 88.170 118.535 88.460 118.765 ;
        RECT 93.645 118.720 93.935 118.765 ;
        RECT 96.525 118.720 96.665 118.920 ;
        RECT 96.895 118.860 97.215 119.120 ;
        RECT 98.735 119.060 99.055 119.120 ;
        RECT 98.735 118.920 108.625 119.060 ;
        RECT 98.735 118.860 99.055 118.920 ;
        RECT 100.130 118.720 100.420 118.765 ;
        RECT 104.715 118.720 105.035 118.780 ;
        RECT 93.645 118.580 96.180 118.720 ;
        RECT 96.525 118.580 105.035 118.720 ;
        RECT 93.645 118.535 93.935 118.580 ;
        RECT 95.965 118.425 96.180 118.580 ;
        RECT 100.130 118.535 100.420 118.580 ;
        RECT 104.715 118.520 105.035 118.580 ;
        RECT 105.605 118.720 105.895 118.765 ;
        RECT 108.485 118.720 108.625 118.920 ;
        RECT 108.855 118.860 109.175 119.120 ;
        RECT 110.695 118.860 111.015 119.120 ;
        RECT 110.785 118.720 110.925 118.860 ;
        RECT 105.605 118.580 108.140 118.720 ;
        RECT 108.485 118.580 110.925 118.720 ;
        RECT 105.605 118.535 105.895 118.580 ;
        RECT 68.825 118.380 69.115 118.425 ;
        RECT 65.565 118.240 69.115 118.380 ;
        RECT 59.635 118.180 59.955 118.240 ;
        RECT 65.565 118.195 65.855 118.240 ;
        RECT 66.535 118.180 66.855 118.240 ;
        RECT 68.825 118.195 69.115 118.240 ;
        RECT 69.745 118.380 70.035 118.425 ;
        RECT 71.605 118.380 71.895 118.425 ;
        RECT 69.745 118.240 71.895 118.380 ;
        RECT 69.745 118.195 70.035 118.240 ;
        RECT 71.605 118.195 71.895 118.240 ;
        RECT 88.630 118.380 88.920 118.425 ;
        RECT 91.785 118.380 92.075 118.425 ;
        RECT 95.045 118.380 95.335 118.425 ;
        RECT 88.630 118.240 95.335 118.380 ;
        RECT 88.630 118.195 88.920 118.240 ;
        RECT 91.785 118.195 92.075 118.240 ;
        RECT 95.045 118.195 95.335 118.240 ;
        RECT 95.965 118.380 96.255 118.425 ;
        RECT 97.825 118.380 98.115 118.425 ;
        RECT 95.965 118.240 98.115 118.380 ;
        RECT 95.965 118.195 96.255 118.240 ;
        RECT 97.825 118.195 98.115 118.240 ;
        RECT 103.745 118.380 104.035 118.425 ;
        RECT 105.175 118.380 105.495 118.440 ;
        RECT 107.925 118.425 108.140 118.580 ;
        RECT 107.005 118.380 107.295 118.425 ;
        RECT 103.745 118.240 107.295 118.380 ;
        RECT 103.745 118.195 104.035 118.240 ;
        RECT 105.175 118.180 105.495 118.240 ;
        RECT 107.005 118.195 107.295 118.240 ;
        RECT 107.925 118.380 108.215 118.425 ;
        RECT 109.785 118.380 110.075 118.425 ;
        RECT 107.925 118.240 110.075 118.380 ;
        RECT 107.925 118.195 108.215 118.240 ;
        RECT 109.785 118.195 110.075 118.240 ;
        RECT 24.675 117.840 24.995 118.100 ;
        RECT 36.175 117.840 36.495 118.100 ;
        RECT 36.635 118.040 36.955 118.100 ;
        RECT 37.110 118.040 37.400 118.085 ;
        RECT 36.635 117.900 37.400 118.040 ;
        RECT 36.635 117.840 36.955 117.900 ;
        RECT 37.110 117.855 37.400 117.900 ;
        RECT 37.555 118.040 37.875 118.100 ;
        RECT 38.935 118.040 39.255 118.100 ;
        RECT 37.555 117.900 39.255 118.040 ;
        RECT 37.555 117.840 37.875 117.900 ;
        RECT 38.935 117.840 39.255 117.900 ;
        RECT 70.675 118.040 70.995 118.100 ;
        RECT 74.830 118.040 75.120 118.085 ;
        RECT 70.675 117.900 75.120 118.040 ;
        RECT 70.675 117.840 70.995 117.900 ;
        RECT 74.830 117.855 75.120 117.900 ;
        RECT 78.510 118.040 78.800 118.085 ;
        RECT 79.875 118.040 80.195 118.100 ;
        RECT 78.510 117.900 80.195 118.040 ;
        RECT 78.510 117.855 78.800 117.900 ;
        RECT 79.875 117.840 80.195 117.900 ;
        RECT 80.795 117.840 81.115 118.100 ;
        RECT 100.575 117.840 100.895 118.100 ;
        RECT 17.370 117.220 112.465 117.700 ;
        RECT 23.755 116.820 24.075 117.080 ;
        RECT 26.530 117.020 26.820 117.065 ;
        RECT 26.975 117.020 27.295 117.080 ;
        RECT 26.530 116.880 27.295 117.020 ;
        RECT 26.530 116.835 26.820 116.880 ;
        RECT 26.975 116.820 27.295 116.880 ;
        RECT 27.435 116.820 27.755 117.080 ;
        RECT 37.555 117.065 37.875 117.080 ;
        RECT 37.340 116.835 37.875 117.065 ;
        RECT 38.260 117.020 38.550 117.065 ;
        RECT 42.615 117.020 42.935 117.080 ;
        RECT 50.450 117.020 50.740 117.065 ;
        RECT 38.260 116.880 50.740 117.020 ;
        RECT 38.260 116.835 38.550 116.880 ;
        RECT 37.555 116.820 37.875 116.835 ;
        RECT 42.615 116.820 42.935 116.880 ;
        RECT 50.450 116.835 50.740 116.880 ;
        RECT 50.910 117.020 51.200 117.065 ;
        RECT 53.440 117.020 53.730 117.065 ;
        RECT 54.575 117.020 54.895 117.080 ;
        RECT 50.910 116.880 54.895 117.020 ;
        RECT 50.910 116.835 51.200 116.880 ;
        RECT 53.440 116.835 53.730 116.880 ;
        RECT 54.575 116.820 54.895 116.880 ;
        RECT 66.535 116.820 66.855 117.080 ;
        RECT 67.915 117.020 68.235 117.080 ;
        RECT 69.310 117.020 69.600 117.065 ;
        RECT 67.915 116.880 69.600 117.020 ;
        RECT 67.915 116.820 68.235 116.880 ;
        RECT 69.310 116.835 69.600 116.880 ;
        RECT 71.150 116.835 71.440 117.065 ;
        RECT 71.610 117.020 71.900 117.065 ;
        RECT 72.055 117.020 72.375 117.080 ;
        RECT 71.610 116.880 72.375 117.020 ;
        RECT 71.610 116.835 71.900 116.880 ;
        RECT 29.295 116.680 29.585 116.725 ;
        RECT 31.155 116.680 31.445 116.725 ;
        RECT 23.385 116.540 26.285 116.680 ;
        RECT 23.385 116.385 23.525 116.540 ;
        RECT 26.145 116.400 26.285 116.540 ;
        RECT 29.295 116.540 31.445 116.680 ;
        RECT 29.295 116.495 29.585 116.540 ;
        RECT 31.155 116.495 31.445 116.540 ;
        RECT 32.075 116.680 32.365 116.725 ;
        RECT 35.335 116.680 35.625 116.725 ;
        RECT 36.175 116.680 36.495 116.740 ;
        RECT 32.075 116.540 36.495 116.680 ;
        RECT 32.075 116.495 32.365 116.540 ;
        RECT 35.335 116.495 35.625 116.540 ;
        RECT 23.310 116.155 23.600 116.385 ;
        RECT 24.675 116.340 24.995 116.400 ;
        RECT 25.610 116.340 25.900 116.385 ;
        RECT 24.675 116.200 25.900 116.340 ;
        RECT 24.675 116.140 24.995 116.200 ;
        RECT 25.610 116.155 25.900 116.200 ;
        RECT 26.055 116.340 26.375 116.400 ;
        RECT 26.990 116.340 27.280 116.385 ;
        RECT 26.055 116.200 27.280 116.340 ;
        RECT 26.055 116.140 26.375 116.200 ;
        RECT 26.990 116.155 27.280 116.200 ;
        RECT 30.210 116.340 30.500 116.385 ;
        RECT 30.655 116.340 30.975 116.400 ;
        RECT 30.210 116.200 30.975 116.340 ;
        RECT 31.230 116.340 31.445 116.495 ;
        RECT 36.175 116.480 36.495 116.540 ;
        RECT 40.265 116.680 40.555 116.725 ;
        RECT 41.235 116.680 41.555 116.740 ;
        RECT 43.525 116.680 43.815 116.725 ;
        RECT 40.265 116.540 43.815 116.680 ;
        RECT 40.265 116.495 40.555 116.540 ;
        RECT 41.235 116.480 41.555 116.540 ;
        RECT 43.525 116.495 43.815 116.540 ;
        RECT 44.445 116.680 44.735 116.725 ;
        RECT 46.305 116.680 46.595 116.725 ;
        RECT 44.445 116.540 46.595 116.680 ;
        RECT 44.445 116.495 44.735 116.540 ;
        RECT 46.305 116.495 46.595 116.540 ;
        RECT 55.445 116.680 55.735 116.725 ;
        RECT 56.875 116.680 57.195 116.740 ;
        RECT 58.705 116.680 58.995 116.725 ;
        RECT 55.445 116.540 58.995 116.680 ;
        RECT 55.445 116.495 55.735 116.540 ;
        RECT 33.475 116.340 33.765 116.385 ;
        RECT 31.230 116.200 33.765 116.340 ;
        RECT 30.210 116.155 30.500 116.200 ;
        RECT 30.655 116.140 30.975 116.200 ;
        RECT 33.475 116.155 33.765 116.200 ;
        RECT 42.125 116.340 42.415 116.385 ;
        RECT 44.445 116.340 44.660 116.495 ;
        RECT 56.875 116.480 57.195 116.540 ;
        RECT 58.705 116.495 58.995 116.540 ;
        RECT 59.625 116.680 59.915 116.725 ;
        RECT 61.485 116.680 61.775 116.725 ;
        RECT 59.625 116.540 61.775 116.680 ;
        RECT 59.625 116.495 59.915 116.540 ;
        RECT 61.485 116.495 61.775 116.540 ;
        RECT 68.850 116.680 69.140 116.725 ;
        RECT 70.675 116.680 70.995 116.740 ;
        RECT 68.850 116.540 70.995 116.680 ;
        RECT 68.850 116.495 69.140 116.540 ;
        RECT 42.125 116.200 44.660 116.340 ;
        RECT 46.755 116.340 47.075 116.400 ;
        RECT 57.305 116.340 57.595 116.385 ;
        RECT 59.625 116.340 59.840 116.495 ;
        RECT 70.675 116.480 70.995 116.540 ;
        RECT 46.755 116.200 49.745 116.340 ;
        RECT 42.125 116.155 42.415 116.200 ;
        RECT 46.755 116.140 47.075 116.200 ;
        RECT 28.370 116.000 28.660 116.045 ;
        RECT 32.495 116.000 32.815 116.060 ;
        RECT 34.795 116.000 35.115 116.060 ;
        RECT 28.370 115.860 35.115 116.000 ;
        RECT 28.370 115.815 28.660 115.860 ;
        RECT 32.495 115.800 32.815 115.860 ;
        RECT 34.795 115.800 35.115 115.860 ;
        RECT 45.375 115.800 45.695 116.060 ;
        RECT 46.295 116.000 46.615 116.060 ;
        RECT 47.230 116.000 47.520 116.045 ;
        RECT 47.675 116.000 47.995 116.060 ;
        RECT 49.605 116.045 49.745 116.200 ;
        RECT 57.305 116.200 59.840 116.340 ;
        RECT 60.095 116.340 60.415 116.400 ;
        RECT 62.410 116.340 62.700 116.385 ;
        RECT 63.775 116.340 64.095 116.400 ;
        RECT 60.095 116.200 64.095 116.340 ;
        RECT 57.305 116.155 57.595 116.200 ;
        RECT 60.095 116.140 60.415 116.200 ;
        RECT 62.410 116.155 62.700 116.200 ;
        RECT 63.775 116.140 64.095 116.200 ;
        RECT 66.090 116.340 66.380 116.385 ;
        RECT 66.995 116.340 67.315 116.400 ;
        RECT 66.090 116.200 67.315 116.340 ;
        RECT 71.225 116.340 71.365 116.835 ;
        RECT 72.055 116.820 72.375 116.880 ;
        RECT 73.435 117.020 73.755 117.080 ;
        RECT 75.060 117.020 75.350 117.065 ;
        RECT 73.435 116.880 75.350 117.020 ;
        RECT 73.435 116.820 73.755 116.880 ;
        RECT 75.060 116.835 75.350 116.880 ;
        RECT 80.795 117.020 81.115 117.080 ;
        RECT 84.720 117.020 85.010 117.065 ;
        RECT 87.235 117.020 87.555 117.080 ;
        RECT 80.795 116.880 87.555 117.020 ;
        RECT 80.795 116.820 81.115 116.880 ;
        RECT 84.720 116.835 85.010 116.880 ;
        RECT 87.235 116.820 87.555 116.880 ;
        RECT 95.975 117.020 96.295 117.080 ;
        RECT 96.910 117.020 97.200 117.065 ;
        RECT 95.975 116.880 97.200 117.020 ;
        RECT 95.975 116.820 96.295 116.880 ;
        RECT 96.910 116.835 97.200 116.880 ;
        RECT 98.275 117.020 98.595 117.080 ;
        RECT 98.750 117.020 99.040 117.065 ;
        RECT 98.275 116.880 99.040 117.020 ;
        RECT 77.065 116.680 77.355 116.725 ;
        RECT 78.495 116.680 78.815 116.740 ;
        RECT 86.775 116.725 87.095 116.740 ;
        RECT 80.325 116.680 80.615 116.725 ;
        RECT 77.065 116.540 80.615 116.680 ;
        RECT 77.065 116.495 77.355 116.540 ;
        RECT 78.495 116.480 78.815 116.540 ;
        RECT 80.325 116.495 80.615 116.540 ;
        RECT 81.245 116.680 81.535 116.725 ;
        RECT 83.105 116.680 83.395 116.725 ;
        RECT 81.245 116.540 83.395 116.680 ;
        RECT 81.245 116.495 81.535 116.540 ;
        RECT 83.105 116.495 83.395 116.540 ;
        RECT 86.725 116.680 87.095 116.725 ;
        RECT 89.985 116.680 90.275 116.725 ;
        RECT 86.725 116.540 90.275 116.680 ;
        RECT 86.725 116.495 87.095 116.540 ;
        RECT 89.985 116.495 90.275 116.540 ;
        RECT 90.905 116.680 91.195 116.725 ;
        RECT 92.765 116.680 93.055 116.725 ;
        RECT 90.905 116.540 93.055 116.680 ;
        RECT 96.985 116.680 97.125 116.835 ;
        RECT 98.275 116.820 98.595 116.880 ;
        RECT 98.750 116.835 99.040 116.880 ;
        RECT 99.900 116.680 100.190 116.725 ;
        RECT 96.985 116.540 100.190 116.680 ;
        RECT 90.905 116.495 91.195 116.540 ;
        RECT 92.765 116.495 93.055 116.540 ;
        RECT 99.900 116.495 100.190 116.540 ;
        RECT 100.575 116.680 100.895 116.740 ;
        RECT 101.905 116.680 102.195 116.725 ;
        RECT 105.165 116.680 105.455 116.725 ;
        RECT 100.575 116.540 105.455 116.680 ;
        RECT 72.530 116.340 72.820 116.385 ;
        RECT 71.225 116.200 72.820 116.340 ;
        RECT 66.090 116.155 66.380 116.200 ;
        RECT 66.995 116.140 67.315 116.200 ;
        RECT 72.530 116.155 72.820 116.200 ;
        RECT 78.925 116.340 79.215 116.385 ;
        RECT 81.245 116.340 81.460 116.495 ;
        RECT 86.775 116.480 87.095 116.495 ;
        RECT 78.925 116.200 81.460 116.340 ;
        RECT 88.585 116.340 88.875 116.385 ;
        RECT 90.905 116.340 91.120 116.495 ;
        RECT 100.575 116.480 100.895 116.540 ;
        RECT 101.905 116.495 102.195 116.540 ;
        RECT 105.165 116.495 105.455 116.540 ;
        RECT 106.085 116.680 106.375 116.725 ;
        RECT 107.945 116.680 108.235 116.725 ;
        RECT 106.085 116.540 108.235 116.680 ;
        RECT 106.085 116.495 106.375 116.540 ;
        RECT 107.945 116.495 108.235 116.540 ;
        RECT 88.585 116.200 91.120 116.340 ;
        RECT 93.690 116.340 93.980 116.385 ;
        RECT 96.895 116.340 97.215 116.400 ;
        RECT 98.735 116.340 99.055 116.400 ;
        RECT 93.690 116.200 99.055 116.340 ;
        RECT 78.925 116.155 79.215 116.200 ;
        RECT 88.585 116.155 88.875 116.200 ;
        RECT 93.690 116.155 93.980 116.200 ;
        RECT 96.895 116.140 97.215 116.200 ;
        RECT 98.735 116.140 99.055 116.200 ;
        RECT 103.765 116.340 104.055 116.385 ;
        RECT 106.085 116.340 106.300 116.495 ;
        RECT 103.765 116.200 106.300 116.340 ;
        RECT 103.765 116.155 104.055 116.200 ;
        RECT 107.015 116.140 107.335 116.400 ;
        RECT 108.870 116.340 109.160 116.385 ;
        RECT 110.695 116.340 111.015 116.400 ;
        RECT 108.870 116.200 111.015 116.340 ;
        RECT 108.870 116.155 109.160 116.200 ;
        RECT 110.695 116.140 111.015 116.200 ;
        RECT 46.295 115.860 47.995 116.000 ;
        RECT 46.295 115.800 46.615 115.860 ;
        RECT 47.230 115.815 47.520 115.860 ;
        RECT 47.675 115.800 47.995 115.860 ;
        RECT 49.530 115.815 49.820 116.045 ;
        RECT 59.175 116.000 59.495 116.060 ;
        RECT 60.570 116.000 60.860 116.045 ;
        RECT 59.175 115.860 60.860 116.000 ;
        RECT 59.175 115.800 59.495 115.860 ;
        RECT 60.570 115.815 60.860 115.860 ;
        RECT 67.455 116.000 67.775 116.060 ;
        RECT 67.930 116.000 68.220 116.045 ;
        RECT 75.735 116.000 76.055 116.060 ;
        RECT 67.455 115.860 76.055 116.000 ;
        RECT 67.455 115.800 67.775 115.860 ;
        RECT 67.930 115.815 68.220 115.860 ;
        RECT 75.735 115.800 76.055 115.860 ;
        RECT 80.795 116.000 81.115 116.060 ;
        RECT 82.190 116.000 82.480 116.045 ;
        RECT 80.795 115.860 82.480 116.000 ;
        RECT 80.795 115.800 81.115 115.860 ;
        RECT 82.190 115.815 82.480 115.860 ;
        RECT 83.095 116.000 83.415 116.060 ;
        RECT 84.030 116.000 84.320 116.045 ;
        RECT 85.855 116.000 86.175 116.060 ;
        RECT 83.095 115.860 86.175 116.000 ;
        RECT 83.095 115.800 83.415 115.860 ;
        RECT 84.030 115.815 84.320 115.860 ;
        RECT 85.855 115.800 86.175 115.860 ;
        RECT 89.535 116.000 89.855 116.060 ;
        RECT 91.850 116.000 92.140 116.045 ;
        RECT 89.535 115.860 92.140 116.000 ;
        RECT 89.535 115.800 89.855 115.860 ;
        RECT 91.850 115.815 92.140 115.860 ;
        RECT 94.595 116.000 94.915 116.060 ;
        RECT 95.530 116.000 95.820 116.045 ;
        RECT 94.595 115.860 95.820 116.000 ;
        RECT 94.595 115.800 94.915 115.860 ;
        RECT 95.530 115.815 95.820 115.860 ;
        RECT 96.450 116.000 96.740 116.045 ;
        RECT 102.415 116.000 102.735 116.060 ;
        RECT 96.450 115.860 102.735 116.000 ;
        RECT 96.450 115.815 96.740 115.860 ;
        RECT 102.415 115.800 102.735 115.860 ;
        RECT 28.835 115.660 29.125 115.705 ;
        RECT 30.695 115.660 30.985 115.705 ;
        RECT 33.475 115.660 33.765 115.705 ;
        RECT 28.835 115.520 33.765 115.660 ;
        RECT 28.835 115.475 29.125 115.520 ;
        RECT 30.695 115.475 30.985 115.520 ;
        RECT 33.475 115.475 33.765 115.520 ;
        RECT 42.125 115.660 42.415 115.705 ;
        RECT 44.905 115.660 45.195 115.705 ;
        RECT 46.765 115.660 47.055 115.705 ;
        RECT 42.125 115.520 47.055 115.660 ;
        RECT 42.125 115.475 42.415 115.520 ;
        RECT 44.905 115.475 45.195 115.520 ;
        RECT 46.765 115.475 47.055 115.520 ;
        RECT 57.305 115.660 57.595 115.705 ;
        RECT 60.085 115.660 60.375 115.705 ;
        RECT 61.945 115.660 62.235 115.705 ;
        RECT 57.305 115.520 62.235 115.660 ;
        RECT 57.305 115.475 57.595 115.520 ;
        RECT 60.085 115.475 60.375 115.520 ;
        RECT 61.945 115.475 62.235 115.520 ;
        RECT 78.925 115.660 79.215 115.705 ;
        RECT 81.705 115.660 81.995 115.705 ;
        RECT 83.565 115.660 83.855 115.705 ;
        RECT 78.925 115.520 83.855 115.660 ;
        RECT 78.925 115.475 79.215 115.520 ;
        RECT 81.705 115.475 81.995 115.520 ;
        RECT 83.565 115.475 83.855 115.520 ;
        RECT 88.585 115.660 88.875 115.705 ;
        RECT 91.365 115.660 91.655 115.705 ;
        RECT 93.225 115.660 93.515 115.705 ;
        RECT 88.585 115.520 93.515 115.660 ;
        RECT 88.585 115.475 88.875 115.520 ;
        RECT 91.365 115.475 91.655 115.520 ;
        RECT 93.225 115.475 93.515 115.520 ;
        RECT 103.765 115.660 104.055 115.705 ;
        RECT 106.545 115.660 106.835 115.705 ;
        RECT 108.405 115.660 108.695 115.705 ;
        RECT 103.765 115.520 108.695 115.660 ;
        RECT 103.765 115.475 104.055 115.520 ;
        RECT 106.545 115.475 106.835 115.520 ;
        RECT 108.405 115.475 108.695 115.520 ;
        RECT 52.275 115.320 52.595 115.380 ;
        RECT 52.750 115.320 53.040 115.365 ;
        RECT 52.275 115.180 53.040 115.320 ;
        RECT 52.275 115.120 52.595 115.180 ;
        RECT 52.750 115.135 53.040 115.180 ;
        RECT 18.165 114.500 112.465 114.980 ;
        RECT 32.955 114.100 33.275 114.360 ;
        RECT 41.235 114.100 41.555 114.360 ;
        RECT 45.850 114.300 46.140 114.345 ;
        RECT 45.850 114.160 47.445 114.300 ;
        RECT 45.850 114.115 46.140 114.160 ;
        RECT 23.870 113.960 24.160 114.005 ;
        RECT 26.990 113.960 27.280 114.005 ;
        RECT 28.880 113.960 29.170 114.005 ;
        RECT 43.995 113.960 44.315 114.020 ;
        RECT 23.870 113.820 29.170 113.960 ;
        RECT 23.870 113.775 24.160 113.820 ;
        RECT 26.990 113.775 27.280 113.820 ;
        RECT 28.880 113.775 29.170 113.820 ;
        RECT 29.365 113.820 44.315 113.960 ;
        RECT 29.365 113.620 29.505 113.820 ;
        RECT 43.995 113.760 44.315 113.820 ;
        RECT 45.375 113.960 45.695 114.020 ;
        RECT 46.310 113.960 46.600 114.005 ;
        RECT 45.375 113.820 46.600 113.960 ;
        RECT 45.375 113.760 45.695 113.820 ;
        RECT 46.310 113.775 46.600 113.820 ;
        RECT 19.705 113.480 29.505 113.620 ;
        RECT 29.750 113.620 30.040 113.665 ;
        RECT 32.495 113.620 32.815 113.680 ;
        RECT 34.335 113.620 34.655 113.680 ;
        RECT 29.750 113.480 34.655 113.620 ;
        RECT 19.705 113.325 19.845 113.480 ;
        RECT 29.750 113.435 30.040 113.480 ;
        RECT 32.495 113.420 32.815 113.480 ;
        RECT 34.335 113.420 34.655 113.480 ;
        RECT 43.090 113.620 43.380 113.665 ;
        RECT 46.755 113.620 47.075 113.680 ;
        RECT 43.090 113.480 47.075 113.620 ;
        RECT 43.090 113.435 43.380 113.480 ;
        RECT 46.755 113.420 47.075 113.480 ;
        RECT 19.630 113.095 19.920 113.325 ;
        RECT 22.790 112.985 23.080 113.300 ;
        RECT 23.870 113.280 24.160 113.325 ;
        RECT 27.450 113.280 27.740 113.325 ;
        RECT 29.285 113.280 29.575 113.325 ;
        RECT 23.870 113.140 29.575 113.280 ;
        RECT 23.870 113.095 24.160 113.140 ;
        RECT 27.450 113.095 27.740 113.140 ;
        RECT 29.285 113.095 29.575 113.140 ;
        RECT 32.035 113.080 32.355 113.340 ;
        RECT 33.415 113.080 33.735 113.340 ;
        RECT 36.635 113.080 36.955 113.340 ;
        RECT 40.790 113.095 41.080 113.325 ;
        RECT 22.490 112.940 23.080 112.985 ;
        RECT 23.295 112.940 23.615 113.000 ;
        RECT 25.730 112.940 26.380 112.985 ;
        RECT 22.490 112.800 26.380 112.940 ;
        RECT 22.490 112.755 22.780 112.800 ;
        RECT 23.295 112.740 23.615 112.800 ;
        RECT 25.730 112.755 26.380 112.800 ;
        RECT 28.355 112.740 28.675 113.000 ;
        RECT 31.115 112.940 31.435 113.000 ;
        RECT 31.115 112.800 35.945 112.940 ;
        RECT 31.115 112.740 31.435 112.800 ;
        RECT 33.890 112.600 34.180 112.645 ;
        RECT 34.795 112.600 35.115 112.660 ;
        RECT 35.805 112.645 35.945 112.800 ;
        RECT 33.890 112.460 35.115 112.600 ;
        RECT 33.890 112.415 34.180 112.460 ;
        RECT 34.795 112.400 35.115 112.460 ;
        RECT 35.730 112.415 36.020 112.645 ;
        RECT 40.865 112.600 41.005 113.095 ;
        RECT 43.535 113.080 43.855 113.340 ;
        RECT 47.305 113.325 47.445 114.160 ;
        RECT 56.875 114.100 57.195 114.360 ;
        RECT 59.175 114.100 59.495 114.360 ;
        RECT 68.835 114.300 69.155 114.360 ;
        RECT 69.310 114.300 69.600 114.345 ;
        RECT 68.835 114.160 69.600 114.300 ;
        RECT 68.835 114.100 69.155 114.160 ;
        RECT 69.310 114.115 69.600 114.160 ;
        RECT 78.495 114.100 78.815 114.360 ;
        RECT 80.795 114.100 81.115 114.360 ;
        RECT 81.730 114.300 82.020 114.345 ;
        RECT 86.775 114.300 87.095 114.360 ;
        RECT 81.730 114.160 87.095 114.300 ;
        RECT 81.730 114.115 82.020 114.160 ;
        RECT 86.775 114.100 87.095 114.160 ;
        RECT 89.535 114.100 89.855 114.360 ;
        RECT 96.435 114.100 96.755 114.360 ;
        RECT 47.230 113.095 47.520 113.325 ;
        RECT 56.430 113.280 56.720 113.325 ;
        RECT 57.795 113.280 58.115 113.340 ;
        RECT 51.905 113.140 58.115 113.280 ;
        RECT 42.615 112.940 42.935 113.000 ;
        RECT 44.010 112.940 44.300 112.985 ;
        RECT 42.615 112.800 44.300 112.940 ;
        RECT 42.615 112.740 42.935 112.800 ;
        RECT 44.010 112.755 44.300 112.800 ;
        RECT 51.905 112.600 52.045 113.140 ;
        RECT 56.430 113.095 56.720 113.140 ;
        RECT 57.795 113.080 58.115 113.140 ;
        RECT 58.270 113.095 58.560 113.325 ;
        RECT 69.770 113.280 70.060 113.325 ;
        RECT 77.115 113.280 77.435 113.340 ;
        RECT 69.770 113.140 77.435 113.280 ;
        RECT 69.770 113.095 70.060 113.140 ;
        RECT 52.275 112.940 52.595 113.000 ;
        RECT 58.345 112.940 58.485 113.095 ;
        RECT 77.115 113.080 77.435 113.140 ;
        RECT 78.050 113.095 78.340 113.325 ;
        RECT 52.275 112.800 58.485 112.940 ;
        RECT 66.995 112.940 67.315 113.000 ;
        RECT 78.125 112.940 78.265 113.095 ;
        RECT 79.875 113.080 80.195 113.340 ;
        RECT 81.270 113.095 81.560 113.325 ;
        RECT 87.695 113.280 88.015 113.340 ;
        RECT 88.630 113.280 88.920 113.325 ;
        RECT 87.695 113.140 88.920 113.280 ;
        RECT 81.345 112.940 81.485 113.095 ;
        RECT 87.695 113.080 88.015 113.140 ;
        RECT 88.630 113.095 88.920 113.140 ;
        RECT 97.355 113.080 97.675 113.340 ;
        RECT 66.995 112.800 81.485 112.940 ;
        RECT 52.275 112.740 52.595 112.800 ;
        RECT 66.995 112.740 67.315 112.800 ;
        RECT 40.865 112.460 52.045 112.600 ;
        RECT 17.370 111.780 112.465 112.260 ;
        RECT 27.910 111.580 28.200 111.625 ;
        RECT 28.355 111.580 28.675 111.640 ;
        RECT 42.630 111.580 42.920 111.625 ;
        RECT 61.015 111.580 61.335 111.640 ;
        RECT 27.910 111.440 28.675 111.580 ;
        RECT 27.910 111.395 28.200 111.440 ;
        RECT 28.355 111.380 28.675 111.440 ;
        RECT 39.945 111.440 42.920 111.580 ;
        RECT 26.515 111.240 26.835 111.300 ;
        RECT 33.990 111.240 34.280 111.285 ;
        RECT 34.795 111.240 35.115 111.300 ;
        RECT 39.945 111.285 40.085 111.440 ;
        RECT 42.630 111.395 42.920 111.440 ;
        RECT 59.265 111.440 70.905 111.580 ;
        RECT 37.230 111.240 37.880 111.285 ;
        RECT 26.515 111.100 29.965 111.240 ;
        RECT 26.515 111.040 26.835 111.100 ;
        RECT 28.815 110.700 29.135 110.960 ;
        RECT 29.825 110.945 29.965 111.100 ;
        RECT 33.990 111.100 37.880 111.240 ;
        RECT 33.990 111.055 34.580 111.100 ;
        RECT 29.750 110.715 30.040 110.945 ;
        RECT 34.290 110.740 34.580 111.055 ;
        RECT 34.795 111.040 35.115 111.100 ;
        RECT 37.230 111.055 37.880 111.100 ;
        RECT 39.870 111.055 40.160 111.285 ;
        RECT 40.315 111.240 40.635 111.300 ;
        RECT 40.315 111.100 43.765 111.240 ;
        RECT 40.315 111.040 40.635 111.100 ;
        RECT 43.625 110.945 43.765 111.100 ;
        RECT 35.370 110.900 35.660 110.945 ;
        RECT 38.950 110.900 39.240 110.945 ;
        RECT 40.785 110.900 41.075 110.945 ;
        RECT 35.370 110.760 41.075 110.900 ;
        RECT 35.370 110.715 35.660 110.760 ;
        RECT 38.950 110.715 39.240 110.760 ;
        RECT 40.785 110.715 41.075 110.760 ;
        RECT 43.550 110.715 43.840 110.945 ;
        RECT 44.455 110.900 44.775 110.960 ;
        RECT 44.930 110.900 45.220 110.945 ;
        RECT 44.455 110.760 45.220 110.900 ;
        RECT 44.455 110.700 44.775 110.760 ;
        RECT 44.930 110.715 45.220 110.760 ;
        RECT 45.390 110.900 45.680 110.945 ;
        RECT 45.835 110.900 46.155 110.960 ;
        RECT 45.390 110.760 46.155 110.900 ;
        RECT 45.390 110.715 45.680 110.760 ;
        RECT 45.835 110.700 46.155 110.760 ;
        RECT 49.055 110.900 49.375 110.960 ;
        RECT 51.830 110.900 52.120 110.945 ;
        RECT 49.055 110.760 52.120 110.900 ;
        RECT 49.055 110.700 49.375 110.760 ;
        RECT 51.830 110.715 52.120 110.760 ;
        RECT 56.890 110.900 57.180 110.945 ;
        RECT 59.265 110.900 59.405 111.440 ;
        RECT 61.015 111.380 61.335 111.440 ;
        RECT 59.635 111.240 59.955 111.300 ;
        RECT 60.210 111.240 60.500 111.285 ;
        RECT 63.450 111.240 64.100 111.285 ;
        RECT 59.635 111.100 64.100 111.240 ;
        RECT 59.635 111.040 59.955 111.100 ;
        RECT 60.210 111.055 60.800 111.100 ;
        RECT 63.450 111.055 64.100 111.100 ;
        RECT 56.890 110.760 59.405 110.900 ;
        RECT 56.890 110.715 57.180 110.760 ;
        RECT 60.510 110.740 60.800 111.055 ;
        RECT 61.590 110.900 61.880 110.945 ;
        RECT 65.170 110.900 65.460 110.945 ;
        RECT 67.005 110.900 67.295 110.945 ;
        RECT 61.590 110.760 67.295 110.900 ;
        RECT 61.590 110.715 61.880 110.760 ;
        RECT 65.170 110.715 65.460 110.760 ;
        RECT 67.005 110.715 67.295 110.760 ;
        RECT 70.215 110.700 70.535 110.960 ;
        RECT 70.765 110.945 70.905 111.440 ;
        RECT 109.790 111.395 110.080 111.625 ;
        RECT 77.115 111.240 77.435 111.300 ;
        RECT 109.865 111.240 110.005 111.395 ;
        RECT 77.115 111.100 110.005 111.240 ;
        RECT 77.115 111.040 77.435 111.100 ;
        RECT 70.690 110.715 70.980 110.945 ;
        RECT 74.355 110.900 74.675 110.960 ;
        RECT 77.590 110.900 77.880 110.945 ;
        RECT 74.355 110.760 77.880 110.900 ;
        RECT 74.355 110.700 74.675 110.760 ;
        RECT 77.590 110.715 77.880 110.760 ;
        RECT 81.255 110.900 81.575 110.960 ;
        RECT 83.110 110.900 83.400 110.945 ;
        RECT 81.255 110.760 83.400 110.900 ;
        RECT 81.255 110.700 81.575 110.760 ;
        RECT 83.110 110.715 83.400 110.760 ;
        RECT 86.315 110.700 86.635 110.960 ;
        RECT 89.090 110.715 89.380 110.945 ;
        RECT 92.310 110.715 92.600 110.945 ;
        RECT 93.690 110.900 93.980 110.945 ;
        RECT 94.135 110.900 94.455 110.960 ;
        RECT 93.690 110.760 94.455 110.900 ;
        RECT 93.690 110.715 93.980 110.760 ;
        RECT 31.130 110.560 31.420 110.605 ;
        RECT 31.575 110.560 31.895 110.620 ;
        RECT 31.130 110.420 31.895 110.560 ;
        RECT 31.130 110.375 31.420 110.420 ;
        RECT 31.575 110.360 31.895 110.420 ;
        RECT 34.795 110.560 35.115 110.620 ;
        RECT 41.250 110.560 41.540 110.605 ;
        RECT 34.795 110.420 41.540 110.560 ;
        RECT 34.795 110.360 35.115 110.420 ;
        RECT 41.250 110.375 41.540 110.420 ;
        RECT 55.035 110.560 55.355 110.620 ;
        RECT 55.510 110.560 55.800 110.605 ;
        RECT 55.035 110.420 55.800 110.560 ;
        RECT 55.035 110.360 55.355 110.420 ;
        RECT 55.510 110.375 55.800 110.420 ;
        RECT 57.350 110.560 57.640 110.605 ;
        RECT 62.855 110.560 63.175 110.620 ;
        RECT 57.350 110.420 63.175 110.560 ;
        RECT 57.350 110.375 57.640 110.420 ;
        RECT 62.855 110.360 63.175 110.420 ;
        RECT 66.075 110.360 66.395 110.620 ;
        RECT 67.455 110.360 67.775 110.620 ;
        RECT 72.070 110.560 72.360 110.605 ;
        RECT 72.515 110.560 72.835 110.620 ;
        RECT 72.070 110.420 72.835 110.560 ;
        RECT 72.070 110.375 72.360 110.420 ;
        RECT 72.515 110.360 72.835 110.420 ;
        RECT 84.015 110.560 84.335 110.620 ;
        RECT 89.165 110.560 89.305 110.715 ;
        RECT 92.385 110.560 92.525 110.715 ;
        RECT 94.135 110.700 94.455 110.760 ;
        RECT 97.830 110.715 98.120 110.945 ;
        RECT 99.195 110.900 99.515 110.960 ;
        RECT 100.130 110.900 100.420 110.945 ;
        RECT 104.730 110.900 105.020 110.945 ;
        RECT 99.195 110.760 100.420 110.900 ;
        RECT 97.905 110.560 98.045 110.715 ;
        RECT 99.195 110.700 99.515 110.760 ;
        RECT 100.130 110.715 100.420 110.760 ;
        RECT 100.665 110.760 105.020 110.900 ;
        RECT 98.735 110.560 99.055 110.620 ;
        RECT 100.665 110.560 100.805 110.760 ;
        RECT 104.730 110.715 105.020 110.760 ;
        RECT 105.635 110.900 105.955 110.960 ;
        RECT 106.110 110.900 106.400 110.945 ;
        RECT 105.635 110.760 106.400 110.900 ;
        RECT 105.635 110.700 105.955 110.760 ;
        RECT 106.110 110.715 106.400 110.760 ;
        RECT 107.475 110.700 107.795 110.960 ;
        RECT 110.710 110.900 111.000 110.945 ;
        RECT 112.535 110.900 112.855 110.960 ;
        RECT 110.710 110.760 112.855 110.900 ;
        RECT 110.710 110.715 111.000 110.760 ;
        RECT 112.535 110.700 112.855 110.760 ;
        RECT 109.775 110.560 110.095 110.620 ;
        RECT 84.015 110.420 89.305 110.560 ;
        RECT 89.625 110.420 100.805 110.560 ;
        RECT 101.125 110.420 110.095 110.560 ;
        RECT 84.015 110.360 84.335 110.420 ;
        RECT 35.370 110.220 35.660 110.265 ;
        RECT 38.490 110.220 38.780 110.265 ;
        RECT 40.380 110.220 40.670 110.265 ;
        RECT 35.370 110.080 40.670 110.220 ;
        RECT 35.370 110.035 35.660 110.080 ;
        RECT 38.490 110.035 38.780 110.080 ;
        RECT 40.380 110.035 40.670 110.080 ;
        RECT 45.835 110.220 46.155 110.280 ;
        RECT 50.910 110.220 51.200 110.265 ;
        RECT 45.835 110.080 51.200 110.220 ;
        RECT 45.835 110.020 46.155 110.080 ;
        RECT 50.910 110.035 51.200 110.080 ;
        RECT 61.590 110.220 61.880 110.265 ;
        RECT 64.710 110.220 65.000 110.265 ;
        RECT 66.600 110.220 66.890 110.265 ;
        RECT 61.590 110.080 66.890 110.220 ;
        RECT 61.590 110.035 61.880 110.080 ;
        RECT 64.710 110.035 65.000 110.080 ;
        RECT 66.600 110.035 66.890 110.080 ;
        RECT 86.315 110.220 86.635 110.280 ;
        RECT 89.625 110.220 89.765 110.420 ;
        RECT 98.735 110.360 99.055 110.420 ;
        RECT 86.315 110.080 89.765 110.220 ;
        RECT 90.010 110.220 90.300 110.265 ;
        RECT 93.215 110.220 93.535 110.280 ;
        RECT 101.125 110.265 101.265 110.420 ;
        RECT 109.775 110.360 110.095 110.420 ;
        RECT 90.010 110.080 93.535 110.220 ;
        RECT 86.315 110.020 86.635 110.080 ;
        RECT 90.010 110.035 90.300 110.080 ;
        RECT 93.215 110.020 93.535 110.080 ;
        RECT 101.050 110.035 101.340 110.265 ;
        RECT 107.030 110.220 107.320 110.265 ;
        RECT 108.855 110.220 109.175 110.280 ;
        RECT 107.030 110.080 109.175 110.220 ;
        RECT 107.030 110.035 107.320 110.080 ;
        RECT 108.855 110.020 109.175 110.080 ;
        RECT 30.670 109.880 30.960 109.925 ;
        RECT 31.115 109.880 31.435 109.940 ;
        RECT 30.670 109.740 31.435 109.880 ;
        RECT 30.670 109.695 30.960 109.740 ;
        RECT 31.115 109.680 31.435 109.740 ;
        RECT 38.015 109.880 38.335 109.940 ;
        RECT 44.010 109.880 44.300 109.925 ;
        RECT 38.015 109.740 44.300 109.880 ;
        RECT 38.015 109.680 38.335 109.740 ;
        RECT 44.010 109.695 44.300 109.740 ;
        RECT 46.295 109.680 46.615 109.940 ;
        RECT 66.995 109.880 67.315 109.940 ;
        RECT 69.310 109.880 69.600 109.925 ;
        RECT 66.995 109.740 69.600 109.880 ;
        RECT 66.995 109.680 67.315 109.740 ;
        RECT 69.310 109.695 69.600 109.740 ;
        RECT 78.495 109.680 78.815 109.940 ;
        RECT 84.015 109.680 84.335 109.940 ;
        RECT 86.775 109.680 87.095 109.940 ;
        RECT 91.835 109.680 92.155 109.940 ;
        RECT 94.610 109.880 94.900 109.925 ;
        RECT 95.515 109.880 95.835 109.940 ;
        RECT 94.610 109.740 95.835 109.880 ;
        RECT 94.610 109.695 94.900 109.740 ;
        RECT 95.515 109.680 95.835 109.740 ;
        RECT 98.290 109.880 98.580 109.925 ;
        RECT 101.955 109.880 102.275 109.940 ;
        RECT 98.290 109.740 102.275 109.880 ;
        RECT 98.290 109.695 98.580 109.740 ;
        RECT 101.955 109.680 102.275 109.740 ;
        RECT 105.190 109.880 105.480 109.925 ;
        RECT 105.635 109.880 105.955 109.940 ;
        RECT 105.190 109.740 105.955 109.880 ;
        RECT 105.190 109.695 105.480 109.740 ;
        RECT 105.635 109.680 105.955 109.740 ;
        RECT 108.410 109.880 108.700 109.925 ;
        RECT 109.315 109.880 109.635 109.940 ;
        RECT 108.410 109.740 109.635 109.880 ;
        RECT 108.410 109.695 108.700 109.740 ;
        RECT 109.315 109.680 109.635 109.740 ;
        RECT 18.165 109.060 112.465 109.540 ;
        RECT 23.295 108.660 23.615 108.920 ;
        RECT 64.250 108.860 64.540 108.905 ;
        RECT 66.075 108.860 66.395 108.920 ;
        RECT 64.250 108.720 66.395 108.860 ;
        RECT 64.250 108.675 64.540 108.720 ;
        RECT 66.075 108.660 66.395 108.720 ;
        RECT 67.455 108.860 67.775 108.920 ;
        RECT 85.855 108.860 86.175 108.920 ;
        RECT 67.455 108.720 86.175 108.860 ;
        RECT 67.455 108.660 67.775 108.720 ;
        RECT 28.470 108.520 28.760 108.565 ;
        RECT 31.590 108.520 31.880 108.565 ;
        RECT 33.480 108.520 33.770 108.565 ;
        RECT 28.470 108.380 33.770 108.520 ;
        RECT 28.470 108.335 28.760 108.380 ;
        RECT 31.590 108.335 31.880 108.380 ;
        RECT 33.480 108.335 33.770 108.380 ;
        RECT 41.810 108.520 42.100 108.565 ;
        RECT 44.930 108.520 45.220 108.565 ;
        RECT 46.820 108.520 47.110 108.565 ;
        RECT 41.810 108.380 47.110 108.520 ;
        RECT 41.810 108.335 42.100 108.380 ;
        RECT 44.930 108.335 45.220 108.380 ;
        RECT 46.820 108.335 47.110 108.380 ;
        RECT 53.310 108.520 53.600 108.565 ;
        RECT 56.430 108.520 56.720 108.565 ;
        RECT 58.320 108.520 58.610 108.565 ;
        RECT 53.310 108.380 58.610 108.520 ;
        RECT 53.310 108.335 53.600 108.380 ;
        RECT 56.430 108.335 56.720 108.380 ;
        RECT 58.320 108.335 58.610 108.380 ;
        RECT 68.950 108.520 69.240 108.565 ;
        RECT 72.070 108.520 72.360 108.565 ;
        RECT 73.960 108.520 74.250 108.565 ;
        RECT 68.950 108.380 74.250 108.520 ;
        RECT 68.950 108.335 69.240 108.380 ;
        RECT 72.070 108.335 72.360 108.380 ;
        RECT 73.960 108.335 74.250 108.380 ;
        RECT 34.335 107.980 34.655 108.240 ;
        RECT 46.295 107.980 46.615 108.240 ;
        RECT 47.675 107.980 47.995 108.240 ;
        RECT 49.070 108.180 49.360 108.225 ;
        RECT 54.575 108.180 54.895 108.240 ;
        RECT 49.070 108.040 54.895 108.180 ;
        RECT 49.070 107.995 49.360 108.040 ;
        RECT 54.575 107.980 54.895 108.040 ;
        RECT 59.190 108.180 59.480 108.225 ;
        RECT 60.095 108.180 60.415 108.240 ;
        RECT 59.190 108.040 60.415 108.180 ;
        RECT 59.190 107.995 59.480 108.040 ;
        RECT 60.095 107.980 60.415 108.040 ;
        RECT 64.710 108.180 65.000 108.225 ;
        RECT 67.455 108.180 67.775 108.240 ;
        RECT 74.905 108.225 75.045 108.720 ;
        RECT 85.855 108.660 86.175 108.720 ;
        RECT 90.455 108.860 90.775 108.920 ;
        RECT 90.455 108.720 98.505 108.860 ;
        RECT 90.455 108.660 90.775 108.720 ;
        RECT 79.990 108.520 80.280 108.565 ;
        RECT 83.110 108.520 83.400 108.565 ;
        RECT 85.000 108.520 85.290 108.565 ;
        RECT 79.990 108.380 85.290 108.520 ;
        RECT 79.990 108.335 80.280 108.380 ;
        RECT 83.110 108.335 83.400 108.380 ;
        RECT 85.000 108.335 85.290 108.380 ;
        RECT 91.030 108.520 91.320 108.565 ;
        RECT 94.150 108.520 94.440 108.565 ;
        RECT 96.040 108.520 96.330 108.565 ;
        RECT 91.030 108.380 96.330 108.520 ;
        RECT 91.030 108.335 91.320 108.380 ;
        RECT 94.150 108.335 94.440 108.380 ;
        RECT 96.040 108.335 96.330 108.380 ;
        RECT 64.710 108.040 67.775 108.180 ;
        RECT 64.710 107.995 65.000 108.040 ;
        RECT 67.455 107.980 67.775 108.040 ;
        RECT 74.830 107.995 75.120 108.225 ;
        RECT 75.750 108.180 76.040 108.225 ;
        RECT 81.255 108.180 81.575 108.240 ;
        RECT 75.750 108.040 81.575 108.180 ;
        RECT 75.750 107.995 76.040 108.040 ;
        RECT 81.255 107.980 81.575 108.040 ;
        RECT 84.015 108.180 84.335 108.240 ;
        RECT 84.490 108.180 84.780 108.225 ;
        RECT 84.015 108.040 84.780 108.180 ;
        RECT 84.015 107.980 84.335 108.040 ;
        RECT 84.490 107.995 84.780 108.040 ;
        RECT 85.855 107.980 86.175 108.240 ;
        RECT 86.790 108.180 87.080 108.225 ;
        RECT 90.455 108.180 90.775 108.240 ;
        RECT 86.790 108.040 90.775 108.180 ;
        RECT 86.790 107.995 87.080 108.040 ;
        RECT 90.455 107.980 90.775 108.040 ;
        RECT 95.515 107.980 95.835 108.240 ;
        RECT 96.895 107.980 97.215 108.240 ;
        RECT 23.755 107.640 24.075 107.900 ;
        RECT 24.230 107.840 24.520 107.885 ;
        RECT 26.055 107.840 26.375 107.900 ;
        RECT 24.230 107.700 26.375 107.840 ;
        RECT 24.230 107.655 24.520 107.700 ;
        RECT 26.055 107.640 26.375 107.700 ;
        RECT 25.595 107.500 25.915 107.560 ;
        RECT 27.390 107.545 27.680 107.860 ;
        RECT 28.470 107.840 28.760 107.885 ;
        RECT 32.050 107.840 32.340 107.885 ;
        RECT 33.885 107.840 34.175 107.885 ;
        RECT 28.470 107.700 34.175 107.840 ;
        RECT 28.470 107.655 28.760 107.700 ;
        RECT 32.050 107.655 32.340 107.700 ;
        RECT 33.885 107.655 34.175 107.700 ;
        RECT 37.095 107.640 37.415 107.900 ;
        RECT 27.090 107.500 27.680 107.545 ;
        RECT 30.330 107.500 30.980 107.545 ;
        RECT 25.595 107.360 30.980 107.500 ;
        RECT 25.595 107.300 25.915 107.360 ;
        RECT 27.090 107.315 27.380 107.360 ;
        RECT 30.330 107.315 30.980 107.360 ;
        RECT 32.970 107.315 33.260 107.545 ;
        RECT 37.570 107.500 37.860 107.545 ;
        RECT 39.855 107.500 40.175 107.560 ;
        RECT 40.730 107.545 41.020 107.860 ;
        RECT 41.810 107.840 42.100 107.885 ;
        RECT 45.390 107.840 45.680 107.885 ;
        RECT 47.225 107.840 47.515 107.885 ;
        RECT 41.810 107.700 47.515 107.840 ;
        RECT 41.810 107.655 42.100 107.700 ;
        RECT 45.390 107.655 45.680 107.700 ;
        RECT 47.225 107.655 47.515 107.700 ;
        RECT 37.570 107.360 40.175 107.500 ;
        RECT 37.570 107.315 37.860 107.360 ;
        RECT 33.045 107.160 33.185 107.315 ;
        RECT 39.855 107.300 40.175 107.360 ;
        RECT 40.430 107.500 41.020 107.545 ;
        RECT 42.615 107.500 42.935 107.560 ;
        RECT 52.230 107.545 52.520 107.860 ;
        RECT 53.310 107.840 53.600 107.885 ;
        RECT 56.890 107.840 57.180 107.885 ;
        RECT 58.725 107.840 59.015 107.885 ;
        RECT 53.310 107.700 59.015 107.840 ;
        RECT 53.310 107.655 53.600 107.700 ;
        RECT 56.890 107.655 57.180 107.700 ;
        RECT 58.725 107.655 59.015 107.700 ;
        RECT 61.030 107.840 61.320 107.885 ;
        RECT 61.475 107.840 61.795 107.900 ;
        RECT 61.030 107.700 61.795 107.840 ;
        RECT 61.030 107.655 61.320 107.700 ;
        RECT 61.475 107.640 61.795 107.700 ;
        RECT 61.935 107.840 62.255 107.900 ;
        RECT 98.365 107.885 98.505 108.720 ;
        RECT 104.830 108.520 105.120 108.565 ;
        RECT 107.950 108.520 108.240 108.565 ;
        RECT 109.840 108.520 110.130 108.565 ;
        RECT 104.830 108.380 110.130 108.520 ;
        RECT 104.830 108.335 105.120 108.380 ;
        RECT 107.950 108.335 108.240 108.380 ;
        RECT 109.840 108.335 110.130 108.380 ;
        RECT 109.315 107.980 109.635 108.240 ;
        RECT 110.695 107.980 111.015 108.240 ;
        RECT 63.330 107.840 63.620 107.885 ;
        RECT 61.935 107.700 63.620 107.840 ;
        RECT 61.935 107.640 62.255 107.700 ;
        RECT 63.330 107.655 63.620 107.700 ;
        RECT 43.670 107.500 44.320 107.545 ;
        RECT 40.430 107.360 44.320 107.500 ;
        RECT 40.430 107.315 40.720 107.360 ;
        RECT 42.615 107.300 42.935 107.360 ;
        RECT 43.670 107.315 44.320 107.360 ;
        RECT 51.930 107.500 52.520 107.545 ;
        RECT 52.735 107.500 53.055 107.560 ;
        RECT 55.170 107.500 55.820 107.545 ;
        RECT 51.930 107.360 55.820 107.500 ;
        RECT 51.930 107.315 52.220 107.360 ;
        RECT 52.735 107.300 53.055 107.360 ;
        RECT 55.170 107.315 55.820 107.360 ;
        RECT 57.335 107.500 57.655 107.560 ;
        RECT 67.870 107.545 68.160 107.860 ;
        RECT 68.950 107.840 69.240 107.885 ;
        RECT 72.530 107.840 72.820 107.885 ;
        RECT 74.365 107.840 74.655 107.885 ;
        RECT 68.950 107.700 74.655 107.840 ;
        RECT 68.950 107.655 69.240 107.700 ;
        RECT 72.530 107.655 72.820 107.700 ;
        RECT 74.365 107.655 74.655 107.700 ;
        RECT 57.810 107.500 58.100 107.545 ;
        RECT 57.335 107.360 58.100 107.500 ;
        RECT 57.335 107.300 57.655 107.360 ;
        RECT 57.810 107.315 58.100 107.360 ;
        RECT 67.570 107.500 68.160 107.545 ;
        RECT 70.675 107.545 70.995 107.560 ;
        RECT 70.675 107.500 71.460 107.545 ;
        RECT 67.570 107.360 71.460 107.500 ;
        RECT 67.570 107.315 67.860 107.360 ;
        RECT 70.675 107.315 71.460 107.360 ;
        RECT 72.975 107.500 73.295 107.560 ;
        RECT 78.910 107.545 79.200 107.860 ;
        RECT 79.990 107.840 80.280 107.885 ;
        RECT 83.570 107.840 83.860 107.885 ;
        RECT 85.405 107.840 85.695 107.885 ;
        RECT 79.990 107.700 85.695 107.840 ;
        RECT 79.990 107.655 80.280 107.700 ;
        RECT 83.570 107.655 83.860 107.700 ;
        RECT 85.405 107.655 85.695 107.700 ;
        RECT 73.450 107.500 73.740 107.545 ;
        RECT 72.975 107.360 73.740 107.500 ;
        RECT 70.675 107.300 70.995 107.315 ;
        RECT 72.975 107.300 73.295 107.360 ;
        RECT 73.450 107.315 73.740 107.360 ;
        RECT 78.610 107.500 79.200 107.545 ;
        RECT 79.415 107.500 79.735 107.560 ;
        RECT 89.950 107.545 90.240 107.860 ;
        RECT 91.030 107.840 91.320 107.885 ;
        RECT 94.610 107.840 94.900 107.885 ;
        RECT 96.445 107.840 96.735 107.885 ;
        RECT 91.030 107.700 96.735 107.840 ;
        RECT 91.030 107.655 91.320 107.700 ;
        RECT 94.610 107.655 94.900 107.700 ;
        RECT 96.445 107.655 96.735 107.700 ;
        RECT 98.290 107.655 98.580 107.885 ;
        RECT 98.735 107.840 99.055 107.900 ;
        RECT 99.670 107.840 99.960 107.885 ;
        RECT 98.735 107.700 99.960 107.840 ;
        RECT 98.735 107.640 99.055 107.700 ;
        RECT 99.670 107.655 99.960 107.700 ;
        RECT 81.850 107.500 82.500 107.545 ;
        RECT 78.610 107.360 82.500 107.500 ;
        RECT 78.610 107.315 78.900 107.360 ;
        RECT 79.415 107.300 79.735 107.360 ;
        RECT 81.850 107.315 82.500 107.360 ;
        RECT 89.650 107.500 90.240 107.545 ;
        RECT 91.835 107.500 92.155 107.560 ;
        RECT 92.890 107.500 93.540 107.545 ;
        RECT 89.650 107.360 93.540 107.500 ;
        RECT 89.650 107.315 89.940 107.360 ;
        RECT 91.835 107.300 92.155 107.360 ;
        RECT 92.890 107.315 93.540 107.360 ;
        RECT 94.135 107.500 94.455 107.560 ;
        RECT 103.750 107.545 104.040 107.860 ;
        RECT 104.830 107.840 105.120 107.885 ;
        RECT 108.410 107.840 108.700 107.885 ;
        RECT 110.245 107.840 110.535 107.885 ;
        RECT 104.830 107.700 110.535 107.840 ;
        RECT 104.830 107.655 105.120 107.700 ;
        RECT 108.410 107.655 108.700 107.700 ;
        RECT 110.245 107.655 110.535 107.700 ;
        RECT 99.210 107.500 99.500 107.545 ;
        RECT 94.135 107.360 99.500 107.500 ;
        RECT 94.135 107.300 94.455 107.360 ;
        RECT 99.210 107.315 99.500 107.360 ;
        RECT 100.590 107.500 100.880 107.545 ;
        RECT 103.450 107.500 104.040 107.545 ;
        RECT 105.635 107.500 105.955 107.560 ;
        RECT 106.690 107.500 107.340 107.545 ;
        RECT 100.590 107.360 103.105 107.500 ;
        RECT 100.590 107.315 100.880 107.360 ;
        RECT 36.190 107.160 36.480 107.205 ;
        RECT 33.045 107.020 36.480 107.160 ;
        RECT 36.190 106.975 36.480 107.020 ;
        RECT 61.950 107.160 62.240 107.205 ;
        RECT 63.775 107.160 64.095 107.220 ;
        RECT 61.950 107.020 64.095 107.160 ;
        RECT 61.950 106.975 62.240 107.020 ;
        RECT 63.775 106.960 64.095 107.020 ;
        RECT 97.355 106.960 97.675 107.220 ;
        RECT 102.965 107.160 103.105 107.360 ;
        RECT 103.450 107.360 107.340 107.500 ;
        RECT 103.450 107.315 103.740 107.360 ;
        RECT 105.635 107.300 105.955 107.360 ;
        RECT 106.690 107.315 107.340 107.360 ;
        RECT 108.395 107.160 108.715 107.220 ;
        RECT 102.965 107.020 108.715 107.160 ;
        RECT 108.395 106.960 108.715 107.020 ;
        RECT 17.370 106.340 112.465 106.820 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 25.595 105.940 25.915 106.200 ;
        RECT 33.415 106.140 33.735 106.200 ;
        RECT 26.605 106.000 50.665 106.140 ;
        RECT 23.755 105.460 24.075 105.520 ;
        RECT 25.150 105.460 25.440 105.505 ;
        RECT 26.605 105.460 26.745 106.000 ;
        RECT 33.415 105.940 33.735 106.000 ;
        RECT 32.955 105.845 33.275 105.860 ;
        RECT 29.390 105.800 29.680 105.845 ;
        RECT 32.630 105.800 33.280 105.845 ;
        RECT 29.390 105.660 33.280 105.800 ;
        RECT 29.390 105.615 29.980 105.660 ;
        RECT 32.630 105.615 33.280 105.660 ;
        RECT 35.270 105.800 35.560 105.845 ;
        RECT 38.015 105.800 38.335 105.860 ;
        RECT 35.270 105.660 38.335 105.800 ;
        RECT 35.270 105.615 35.560 105.660 ;
        RECT 23.755 105.320 26.745 105.460 ;
        RECT 23.755 105.260 24.075 105.320 ;
        RECT 25.150 105.275 25.440 105.320 ;
        RECT 29.690 105.300 29.980 105.615 ;
        RECT 32.955 105.600 33.275 105.615 ;
        RECT 38.015 105.600 38.335 105.660 ;
        RECT 40.770 105.800 41.420 105.845 ;
        RECT 44.370 105.800 44.660 105.845 ;
        RECT 49.990 105.800 50.280 105.845 ;
        RECT 40.770 105.660 50.280 105.800 ;
        RECT 40.770 105.615 41.420 105.660 ;
        RECT 44.070 105.615 44.660 105.660 ;
        RECT 49.990 105.615 50.280 105.660 ;
        RECT 30.770 105.460 31.060 105.505 ;
        RECT 34.350 105.460 34.640 105.505 ;
        RECT 36.185 105.460 36.475 105.505 ;
        RECT 30.770 105.320 36.475 105.460 ;
        RECT 30.770 105.275 31.060 105.320 ;
        RECT 34.350 105.275 34.640 105.320 ;
        RECT 36.185 105.275 36.475 105.320 ;
        RECT 37.575 105.460 37.865 105.505 ;
        RECT 39.410 105.460 39.700 105.505 ;
        RECT 42.990 105.460 43.280 105.505 ;
        RECT 37.575 105.320 43.280 105.460 ;
        RECT 37.575 105.275 37.865 105.320 ;
        RECT 39.410 105.275 39.700 105.320 ;
        RECT 42.990 105.275 43.280 105.320 ;
        RECT 44.070 105.300 44.360 105.615 ;
        RECT 50.525 105.505 50.665 106.000 ;
        RECT 52.735 105.940 53.055 106.200 ;
        RECT 54.590 106.140 54.880 106.185 ;
        RECT 57.335 106.140 57.655 106.200 ;
        RECT 54.590 106.000 57.655 106.140 ;
        RECT 54.590 105.955 54.880 106.000 ;
        RECT 57.335 105.940 57.655 106.000 ;
        RECT 70.675 105.940 70.995 106.200 ;
        RECT 72.975 105.940 73.295 106.200 ;
        RECT 78.495 106.140 78.815 106.200 ;
        RECT 109.775 106.140 110.095 106.200 ;
        RECT 78.495 106.000 82.865 106.140 ;
        RECT 78.495 105.940 78.815 106.000 ;
        RECT 55.035 105.800 55.355 105.860 ;
        RECT 52.365 105.660 55.355 105.800 ;
        RECT 52.365 105.505 52.505 105.660 ;
        RECT 55.035 105.600 55.355 105.660 ;
        RECT 57.910 105.800 58.200 105.845 ;
        RECT 61.150 105.800 61.800 105.845 ;
        RECT 57.910 105.660 61.800 105.800 ;
        RECT 57.910 105.615 58.500 105.660 ;
        RECT 61.150 105.615 61.800 105.660 ;
        RECT 58.210 105.520 58.500 105.615 ;
        RECT 63.775 105.600 64.095 105.860 ;
        RECT 76.770 105.800 77.060 105.845 ;
        RECT 78.955 105.800 79.275 105.860 ;
        RECT 82.725 105.845 82.865 106.000 ;
        RECT 108.485 106.000 110.095 106.140 ;
        RECT 80.010 105.800 80.660 105.845 ;
        RECT 76.770 105.660 80.660 105.800 ;
        RECT 76.770 105.615 77.360 105.660 ;
        RECT 50.450 105.460 50.740 105.505 ;
        RECT 52.290 105.460 52.580 105.505 ;
        RECT 50.450 105.320 52.580 105.460 ;
        RECT 50.450 105.275 50.740 105.320 ;
        RECT 52.290 105.275 52.580 105.320 ;
        RECT 53.670 105.460 53.960 105.505 ;
        RECT 55.495 105.460 55.815 105.520 ;
        RECT 53.670 105.320 55.815 105.460 ;
        RECT 53.670 105.275 53.960 105.320 ;
        RECT 55.495 105.260 55.815 105.320 ;
        RECT 58.210 105.300 58.575 105.520 ;
        RECT 58.255 105.260 58.575 105.300 ;
        RECT 59.290 105.460 59.580 105.505 ;
        RECT 62.870 105.460 63.160 105.505 ;
        RECT 64.705 105.460 64.995 105.505 ;
        RECT 59.290 105.320 64.995 105.460 ;
        RECT 59.290 105.275 59.580 105.320 ;
        RECT 62.870 105.275 63.160 105.320 ;
        RECT 64.705 105.275 64.995 105.320 ;
        RECT 69.770 105.460 70.060 105.505 ;
        RECT 71.150 105.460 71.440 105.505 ;
        RECT 69.770 105.320 71.440 105.460 ;
        RECT 69.770 105.275 70.060 105.320 ;
        RECT 71.150 105.275 71.440 105.320 ;
        RECT 26.530 104.935 26.820 105.165 ;
        RECT 34.795 105.120 35.115 105.180 ;
        RECT 36.650 105.120 36.940 105.165 ;
        RECT 37.110 105.120 37.400 105.165 ;
        RECT 34.795 104.980 37.400 105.120 ;
        RECT 24.215 104.240 24.535 104.500 ;
        RECT 26.605 104.440 26.745 104.935 ;
        RECT 34.795 104.920 35.115 104.980 ;
        RECT 36.650 104.935 36.940 104.980 ;
        RECT 37.110 104.935 37.400 104.980 ;
        RECT 38.490 105.120 38.780 105.165 ;
        RECT 45.835 105.120 46.155 105.180 ;
        RECT 38.490 104.980 46.155 105.120 ;
        RECT 38.490 104.935 38.780 104.980 ;
        RECT 45.835 104.920 46.155 104.980 ;
        RECT 47.230 105.120 47.520 105.165 ;
        RECT 49.055 105.120 49.375 105.180 ;
        RECT 47.230 104.980 49.375 105.120 ;
        RECT 47.230 104.935 47.520 104.980 ;
        RECT 49.055 104.920 49.375 104.980 ;
        RECT 55.050 105.120 55.340 105.165 ;
        RECT 57.795 105.120 58.115 105.180 ;
        RECT 55.050 104.980 58.115 105.120 ;
        RECT 55.050 104.935 55.340 104.980 ;
        RECT 57.795 104.920 58.115 104.980 ;
        RECT 60.095 105.120 60.415 105.180 ;
        RECT 65.170 105.120 65.460 105.165 ;
        RECT 60.095 104.980 65.460 105.120 ;
        RECT 71.225 105.120 71.365 105.275 ;
        RECT 72.055 105.260 72.375 105.520 ;
        RECT 77.070 105.300 77.360 105.615 ;
        RECT 78.955 105.600 79.275 105.660 ;
        RECT 80.010 105.615 80.660 105.660 ;
        RECT 82.650 105.615 82.940 105.845 ;
        RECT 86.775 105.800 87.095 105.860 ;
        RECT 87.350 105.800 87.640 105.845 ;
        RECT 90.590 105.800 91.240 105.845 ;
        RECT 86.775 105.660 91.240 105.800 ;
        RECT 86.775 105.600 87.095 105.660 ;
        RECT 87.350 105.615 87.940 105.660 ;
        RECT 90.590 105.615 91.240 105.660 ;
        RECT 78.150 105.460 78.440 105.505 ;
        RECT 81.730 105.460 82.020 105.505 ;
        RECT 83.565 105.460 83.855 105.505 ;
        RECT 78.150 105.320 83.855 105.460 ;
        RECT 78.150 105.275 78.440 105.320 ;
        RECT 81.730 105.275 82.020 105.320 ;
        RECT 83.565 105.275 83.855 105.320 ;
        RECT 84.030 105.460 84.320 105.505 ;
        RECT 85.855 105.460 86.175 105.520 ;
        RECT 84.030 105.320 86.175 105.460 ;
        RECT 84.030 105.275 84.320 105.320 ;
        RECT 85.855 105.260 86.175 105.320 ;
        RECT 87.650 105.300 87.940 105.615 ;
        RECT 93.215 105.600 93.535 105.860 ;
        RECT 101.955 105.800 102.275 105.860 ;
        RECT 108.485 105.845 108.625 106.000 ;
        RECT 109.775 105.940 110.095 106.000 ;
        RECT 102.530 105.800 102.820 105.845 ;
        RECT 105.770 105.800 106.420 105.845 ;
        RECT 101.955 105.660 106.420 105.800 ;
        RECT 101.955 105.600 102.275 105.660 ;
        RECT 102.530 105.615 103.120 105.660 ;
        RECT 105.770 105.615 106.420 105.660 ;
        RECT 108.410 105.615 108.700 105.845 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 88.730 105.460 89.020 105.505 ;
        RECT 92.310 105.460 92.600 105.505 ;
        RECT 94.145 105.460 94.435 105.505 ;
        RECT 88.730 105.320 94.435 105.460 ;
        RECT 88.730 105.275 89.020 105.320 ;
        RECT 92.310 105.275 92.600 105.320 ;
        RECT 94.145 105.275 94.435 105.320 ;
        RECT 94.610 105.460 94.900 105.505 ;
        RECT 96.895 105.460 97.215 105.520 ;
        RECT 94.610 105.320 97.215 105.460 ;
        RECT 94.610 105.275 94.900 105.320 ;
        RECT 96.895 105.260 97.215 105.320 ;
        RECT 97.830 105.460 98.120 105.505 ;
        RECT 98.735 105.460 99.055 105.520 ;
        RECT 97.830 105.320 99.055 105.460 ;
        RECT 97.830 105.275 98.120 105.320 ;
        RECT 98.735 105.260 99.055 105.320 ;
        RECT 102.830 105.300 103.120 105.615 ;
        RECT 103.910 105.460 104.200 105.505 ;
        RECT 107.490 105.460 107.780 105.505 ;
        RECT 109.325 105.460 109.615 105.505 ;
        RECT 103.910 105.320 109.615 105.460 ;
        RECT 103.910 105.275 104.200 105.320 ;
        RECT 107.490 105.275 107.780 105.320 ;
        RECT 109.325 105.275 109.615 105.320 ;
        RECT 109.790 105.460 110.080 105.505 ;
        RECT 110.695 105.460 111.015 105.520 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 109.790 105.320 111.015 105.460 ;
        RECT 109.790 105.275 110.080 105.320 ;
        RECT 110.695 105.260 111.015 105.320 ;
        RECT 72.515 105.120 72.835 105.180 ;
        RECT 71.225 104.980 72.835 105.120 ;
        RECT 60.095 104.920 60.415 104.980 ;
        RECT 65.170 104.935 65.460 104.980 ;
        RECT 72.515 104.920 72.835 104.980 ;
        RECT 73.910 105.120 74.200 105.165 ;
        RECT 75.735 105.120 76.055 105.180 ;
        RECT 73.910 104.980 76.055 105.120 ;
        RECT 73.910 104.935 74.200 104.980 ;
        RECT 75.735 104.920 76.055 104.980 ;
        RECT 84.490 104.935 84.780 105.165 ;
        RECT 99.195 105.120 99.515 105.180 ;
        RECT 99.670 105.120 99.960 105.165 ;
        RECT 99.195 104.980 99.960 105.120 ;
        RECT 30.770 104.780 31.060 104.825 ;
        RECT 33.890 104.780 34.180 104.825 ;
        RECT 35.780 104.780 36.070 104.825 ;
        RECT 30.770 104.640 36.070 104.780 ;
        RECT 30.770 104.595 31.060 104.640 ;
        RECT 33.890 104.595 34.180 104.640 ;
        RECT 35.780 104.595 36.070 104.640 ;
        RECT 37.980 104.780 38.270 104.825 ;
        RECT 39.870 104.780 40.160 104.825 ;
        RECT 42.990 104.780 43.280 104.825 ;
        RECT 37.980 104.640 43.280 104.780 ;
        RECT 37.980 104.595 38.270 104.640 ;
        RECT 39.870 104.595 40.160 104.640 ;
        RECT 42.990 104.595 43.280 104.640 ;
        RECT 59.290 104.780 59.580 104.825 ;
        RECT 62.410 104.780 62.700 104.825 ;
        RECT 64.300 104.780 64.590 104.825 ;
        RECT 59.290 104.640 64.590 104.780 ;
        RECT 59.290 104.595 59.580 104.640 ;
        RECT 62.410 104.595 62.700 104.640 ;
        RECT 64.300 104.595 64.590 104.640 ;
        RECT 78.150 104.780 78.440 104.825 ;
        RECT 81.270 104.780 81.560 104.825 ;
        RECT 83.160 104.780 83.450 104.825 ;
        RECT 78.150 104.640 83.450 104.780 ;
        RECT 84.565 104.780 84.705 104.935 ;
        RECT 99.195 104.920 99.515 104.980 ;
        RECT 99.670 104.935 99.960 104.980 ;
        RECT 85.855 104.780 86.175 104.840 ;
        RECT 84.565 104.640 86.175 104.780 ;
        RECT 78.150 104.595 78.440 104.640 ;
        RECT 81.270 104.595 81.560 104.640 ;
        RECT 83.160 104.595 83.450 104.640 ;
        RECT 85.855 104.580 86.175 104.640 ;
        RECT 88.730 104.780 89.020 104.825 ;
        RECT 91.850 104.780 92.140 104.825 ;
        RECT 93.740 104.780 94.030 104.825 ;
        RECT 88.730 104.640 94.030 104.780 ;
        RECT 88.730 104.595 89.020 104.640 ;
        RECT 91.850 104.595 92.140 104.640 ;
        RECT 93.740 104.595 94.030 104.640 ;
        RECT 103.910 104.780 104.200 104.825 ;
        RECT 107.030 104.780 107.320 104.825 ;
        RECT 108.920 104.780 109.210 104.825 ;
        RECT 103.910 104.640 109.210 104.780 ;
        RECT 103.910 104.595 104.200 104.640 ;
        RECT 107.030 104.595 107.320 104.640 ;
        RECT 108.920 104.595 109.210 104.640 ;
        RECT 35.255 104.440 35.575 104.500 ;
        RECT 26.605 104.300 35.575 104.440 ;
        RECT 35.255 104.240 35.575 104.300 ;
        RECT 69.295 104.240 69.615 104.500 ;
        RECT 98.290 104.440 98.580 104.485 ;
        RECT 101.955 104.440 102.275 104.500 ;
        RECT 98.290 104.300 102.275 104.440 ;
        RECT 98.290 104.255 98.580 104.300 ;
        RECT 101.955 104.240 102.275 104.300 ;
        RECT 18.165 103.620 112.465 104.100 ;
        RECT 32.955 103.420 33.275 103.480 ;
        RECT 38.950 103.420 39.240 103.465 ;
        RECT 32.955 103.280 39.240 103.420 ;
        RECT 32.955 103.220 33.275 103.280 ;
        RECT 38.950 103.235 39.240 103.280 ;
        RECT 41.710 103.420 42.000 103.465 ;
        RECT 42.615 103.420 42.935 103.480 ;
        RECT 41.710 103.280 42.935 103.420 ;
        RECT 41.710 103.235 42.000 103.280 ;
        RECT 42.615 103.220 42.935 103.280 ;
        RECT 58.255 103.220 58.575 103.480 ;
        RECT 59.635 103.220 59.955 103.480 ;
        RECT 77.130 103.420 77.420 103.465 ;
        RECT 78.955 103.420 79.275 103.480 ;
        RECT 77.130 103.280 79.275 103.420 ;
        RECT 77.130 103.235 77.420 103.280 ;
        RECT 78.955 103.220 79.275 103.280 ;
        RECT 79.415 103.420 79.735 103.480 ;
        RECT 82.190 103.420 82.480 103.465 ;
        RECT 79.415 103.280 82.480 103.420 ;
        RECT 79.415 103.220 79.735 103.280 ;
        RECT 82.190 103.235 82.480 103.280 ;
        RECT 96.895 103.420 97.215 103.480 ;
        RECT 96.895 103.280 98.505 103.420 ;
        RECT 96.895 103.220 97.215 103.280 ;
        RECT 26.630 103.080 26.920 103.125 ;
        RECT 29.750 103.080 30.040 103.125 ;
        RECT 31.640 103.080 31.930 103.125 ;
        RECT 26.630 102.940 31.930 103.080 ;
        RECT 26.630 102.895 26.920 102.940 ;
        RECT 29.750 102.895 30.040 102.940 ;
        RECT 31.640 102.895 31.930 102.940 ;
        RECT 63.740 103.080 64.030 103.125 ;
        RECT 65.630 103.080 65.920 103.125 ;
        RECT 68.750 103.080 69.040 103.125 ;
        RECT 63.740 102.940 69.040 103.080 ;
        RECT 63.740 102.895 64.030 102.940 ;
        RECT 65.630 102.895 65.920 102.940 ;
        RECT 68.750 102.895 69.040 102.940 ;
        RECT 92.870 103.080 93.160 103.125 ;
        RECT 95.990 103.080 96.280 103.125 ;
        RECT 97.880 103.080 98.170 103.125 ;
        RECT 92.870 102.940 98.170 103.080 ;
        RECT 92.870 102.895 93.160 102.940 ;
        RECT 95.990 102.895 96.280 102.940 ;
        RECT 97.880 102.895 98.170 102.940 ;
        RECT 31.115 102.540 31.435 102.800 ;
        RECT 32.510 102.740 32.800 102.785 ;
        RECT 34.795 102.740 35.115 102.800 ;
        RECT 32.510 102.600 35.115 102.740 ;
        RECT 32.510 102.555 32.800 102.600 ;
        RECT 34.795 102.540 35.115 102.600 ;
        RECT 60.095 102.740 60.415 102.800 ;
        RECT 62.870 102.740 63.160 102.785 ;
        RECT 60.095 102.600 63.160 102.740 ;
        RECT 60.095 102.540 60.415 102.600 ;
        RECT 62.870 102.555 63.160 102.600 ;
        RECT 64.250 102.740 64.540 102.785 ;
        RECT 66.535 102.740 66.855 102.800 ;
        RECT 64.250 102.600 66.855 102.740 ;
        RECT 64.250 102.555 64.540 102.600 ;
        RECT 66.535 102.540 66.855 102.600 ;
        RECT 88.630 102.740 88.920 102.785 ;
        RECT 95.055 102.740 95.375 102.800 ;
        RECT 88.630 102.600 95.375 102.740 ;
        RECT 88.630 102.555 88.920 102.600 ;
        RECT 95.055 102.540 95.375 102.600 ;
        RECT 97.355 102.540 97.675 102.800 ;
        RECT 98.365 102.740 98.505 103.280 ;
        RECT 104.830 103.080 105.120 103.125 ;
        RECT 107.950 103.080 108.240 103.125 ;
        RECT 109.840 103.080 110.130 103.125 ;
        RECT 104.830 102.940 110.130 103.080 ;
        RECT 104.830 102.895 105.120 102.940 ;
        RECT 107.950 102.895 108.240 102.940 ;
        RECT 109.840 102.895 110.130 102.940 ;
        RECT 98.750 102.740 99.040 102.785 ;
        RECT 98.365 102.600 99.040 102.740 ;
        RECT 98.750 102.555 99.040 102.600 ;
        RECT 100.590 102.740 100.880 102.785 ;
        RECT 104.255 102.740 104.575 102.800 ;
        RECT 100.590 102.600 104.575 102.740 ;
        RECT 100.590 102.555 100.880 102.600 ;
        RECT 104.255 102.540 104.575 102.600 ;
        RECT 108.855 102.740 109.175 102.800 ;
        RECT 109.330 102.740 109.620 102.785 ;
        RECT 108.855 102.600 109.620 102.740 ;
        RECT 108.855 102.540 109.175 102.600 ;
        RECT 109.330 102.555 109.620 102.600 ;
        RECT 110.695 102.540 111.015 102.800 ;
        RECT 24.215 102.400 24.535 102.460 ;
        RECT 25.550 102.400 25.840 102.420 ;
        RECT 24.215 102.260 25.840 102.400 ;
        RECT 24.215 102.200 24.535 102.260 ;
        RECT 21.455 102.060 21.775 102.120 ;
        RECT 25.550 102.105 25.840 102.260 ;
        RECT 26.630 102.400 26.920 102.445 ;
        RECT 30.210 102.400 30.500 102.445 ;
        RECT 32.045 102.400 32.335 102.445 ;
        RECT 26.630 102.260 32.335 102.400 ;
        RECT 26.630 102.215 26.920 102.260 ;
        RECT 30.210 102.215 30.500 102.260 ;
        RECT 32.045 102.215 32.335 102.260 ;
        RECT 33.415 102.400 33.735 102.460 ;
        RECT 39.410 102.400 39.700 102.445 ;
        RECT 41.250 102.400 41.540 102.445 ;
        RECT 33.415 102.260 41.540 102.400 ;
        RECT 33.415 102.200 33.735 102.260 ;
        RECT 39.410 102.215 39.700 102.260 ;
        RECT 41.250 102.215 41.540 102.260 ;
        RECT 55.035 102.400 55.355 102.460 ;
        RECT 57.810 102.400 58.100 102.445 ;
        RECT 59.190 102.400 59.480 102.445 ;
        RECT 55.035 102.260 59.480 102.400 ;
        RECT 55.035 102.200 55.355 102.260 ;
        RECT 57.810 102.215 58.100 102.260 ;
        RECT 59.190 102.215 59.480 102.260 ;
        RECT 63.335 102.400 63.625 102.445 ;
        RECT 65.170 102.400 65.460 102.445 ;
        RECT 68.750 102.400 69.040 102.445 ;
        RECT 63.335 102.260 69.040 102.400 ;
        RECT 63.335 102.215 63.625 102.260 ;
        RECT 65.170 102.215 65.460 102.260 ;
        RECT 68.750 102.215 69.040 102.260 ;
        RECT 22.390 102.060 22.680 102.105 ;
        RECT 21.455 101.920 22.680 102.060 ;
        RECT 21.455 101.860 21.775 101.920 ;
        RECT 22.390 101.875 22.680 101.920 ;
        RECT 25.250 102.060 25.840 102.105 ;
        RECT 28.490 102.060 29.140 102.105 ;
        RECT 25.250 101.920 29.140 102.060 ;
        RECT 25.250 101.875 25.540 101.920 ;
        RECT 28.490 101.875 29.140 101.920 ;
        RECT 66.530 102.060 67.180 102.105 ;
        RECT 69.295 102.060 69.615 102.120 ;
        RECT 69.830 102.105 70.120 102.420 ;
        RECT 72.515 102.400 72.835 102.460 ;
        RECT 76.670 102.400 76.960 102.445 ;
        RECT 82.650 102.400 82.940 102.445 ;
        RECT 86.315 102.400 86.635 102.460 ;
        RECT 72.515 102.260 86.635 102.400 ;
        RECT 72.515 102.200 72.835 102.260 ;
        RECT 76.670 102.215 76.960 102.260 ;
        RECT 82.650 102.215 82.940 102.260 ;
        RECT 86.315 102.200 86.635 102.260 ;
        RECT 69.830 102.060 70.420 102.105 ;
        RECT 66.530 101.920 70.420 102.060 ;
        RECT 66.530 101.875 67.180 101.920 ;
        RECT 69.295 101.860 69.615 101.920 ;
        RECT 70.130 101.875 70.420 101.920 ;
        RECT 72.055 102.060 72.375 102.120 ;
        RECT 91.790 102.105 92.080 102.420 ;
        RECT 92.870 102.400 93.160 102.445 ;
        RECT 96.450 102.400 96.740 102.445 ;
        RECT 98.285 102.400 98.575 102.445 ;
        RECT 92.870 102.260 98.575 102.400 ;
        RECT 92.870 102.215 93.160 102.260 ;
        RECT 96.450 102.215 96.740 102.260 ;
        RECT 98.285 102.215 98.575 102.260 ;
        RECT 101.955 102.400 102.275 102.460 ;
        RECT 103.750 102.400 104.040 102.420 ;
        RECT 101.955 102.260 104.040 102.400 ;
        RECT 101.955 102.200 102.275 102.260 ;
        RECT 72.990 102.060 73.280 102.105 ;
        RECT 72.055 101.920 73.280 102.060 ;
        RECT 72.055 101.860 72.375 101.920 ;
        RECT 72.990 101.875 73.280 101.920 ;
        RECT 91.490 102.060 92.080 102.105 ;
        RECT 94.135 102.060 94.455 102.120 ;
        RECT 103.750 102.105 104.040 102.260 ;
        RECT 104.830 102.400 105.120 102.445 ;
        RECT 108.410 102.400 108.700 102.445 ;
        RECT 110.245 102.400 110.535 102.445 ;
        RECT 104.830 102.260 110.535 102.400 ;
        RECT 104.830 102.215 105.120 102.260 ;
        RECT 108.410 102.215 108.700 102.260 ;
        RECT 110.245 102.215 110.535 102.260 ;
        RECT 94.730 102.060 95.380 102.105 ;
        RECT 91.490 101.920 95.380 102.060 ;
        RECT 91.490 101.875 91.780 101.920 ;
        RECT 94.135 101.860 94.455 101.920 ;
        RECT 94.730 101.875 95.380 101.920 ;
        RECT 103.450 102.060 104.040 102.105 ;
        RECT 106.690 102.060 107.340 102.105 ;
        RECT 103.450 101.920 107.340 102.060 ;
        RECT 103.450 101.875 103.740 101.920 ;
        RECT 106.690 101.875 107.340 101.920 ;
        RECT 17.370 100.900 112.465 101.380 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 17.400 193.435 18.940 193.805 ;
        RECT 40.975 193.435 42.515 193.805 ;
        RECT 64.550 193.435 66.090 193.805 ;
        RECT 88.125 193.435 89.665 193.805 ;
        RECT 105.665 192.610 105.925 192.930 ;
        RECT 108.885 192.610 109.145 192.930 ;
        RECT 20.565 192.270 20.825 192.590 ;
        RECT 28.385 192.270 28.645 192.590 ;
        RECT 44.025 192.270 44.285 192.590 ;
        RECT 44.945 192.270 45.205 192.590 ;
        RECT 51.385 192.270 51.645 192.590 ;
        RECT 70.245 192.270 70.505 192.590 ;
        RECT 75.305 192.270 75.565 192.590 ;
        RECT 87.725 192.270 87.985 192.590 ;
        RECT 94.625 192.270 94.885 192.590 ;
        RECT 98.765 192.270 99.025 192.590 ;
        RECT 17.400 187.995 18.940 188.365 ;
        RECT 20.625 187.150 20.765 192.270 ;
        RECT 21.025 191.250 21.285 191.570 ;
        RECT 21.085 189.190 21.225 191.250 ;
        RECT 23.785 189.550 24.045 189.870 ;
        RECT 21.025 188.870 21.285 189.190 ;
        RECT 23.845 187.230 23.985 189.550 ;
        RECT 25.165 189.270 25.425 189.530 ;
        RECT 25.165 189.210 26.285 189.270 ;
        RECT 25.225 189.130 26.285 189.210 ;
        RECT 23.845 187.150 24.445 187.230 ;
        RECT 20.565 186.830 20.825 187.150 ;
        RECT 23.845 187.090 24.505 187.150 ;
        RECT 24.245 186.830 24.505 187.090 ;
        RECT 20.625 184.090 20.765 186.830 ;
        RECT 24.305 184.430 24.445 186.830 ;
        RECT 26.145 186.810 26.285 189.130 ;
        RECT 26.545 188.530 26.805 188.850 ;
        RECT 26.605 187.830 26.745 188.530 ;
        RECT 28.445 187.830 28.585 192.270 ;
        RECT 31.605 191.250 31.865 191.570 ;
        RECT 43.565 191.250 43.825 191.570 ;
        RECT 29.185 190.715 30.725 191.085 ;
        RECT 31.665 189.870 31.805 191.250 ;
        RECT 31.605 189.550 31.865 189.870 ;
        RECT 32.985 189.550 33.245 189.870 ;
        RECT 26.545 187.510 26.805 187.830 ;
        RECT 28.385 187.510 28.645 187.830 ;
        RECT 25.625 186.490 25.885 186.810 ;
        RECT 26.085 186.490 26.345 186.810 ;
        RECT 27.465 186.490 27.725 186.810 ;
        RECT 31.145 186.490 31.405 186.810 ;
        RECT 24.705 185.810 24.965 186.130 ;
        RECT 24.245 184.110 24.505 184.430 ;
        RECT 20.565 183.770 20.825 184.090 ;
        RECT 20.105 183.090 20.365 183.410 ;
        RECT 17.400 182.555 18.940 182.925 ;
        RECT 20.165 178.310 20.305 183.090 ;
        RECT 20.105 177.990 20.365 178.310 ;
        RECT 17.400 177.115 18.940 177.485 ;
        RECT 17.400 171.675 18.940 172.045 ;
        RECT 20.625 170.830 20.765 183.770 ;
        RECT 24.765 183.750 24.905 185.810 ;
        RECT 25.685 185.110 25.825 186.490 ;
        RECT 25.625 184.790 25.885 185.110 ;
        RECT 22.405 183.430 22.665 183.750 ;
        RECT 24.705 183.430 24.965 183.750 ;
        RECT 22.465 182.390 22.605 183.430 ;
        RECT 22.405 182.070 22.665 182.390 ;
        RECT 27.525 181.710 27.665 186.490 ;
        RECT 29.185 185.275 30.725 185.645 ;
        RECT 31.205 185.110 31.345 186.490 ;
        RECT 28.845 184.790 29.105 185.110 ;
        RECT 31.145 184.790 31.405 185.110 ;
        RECT 27.465 181.390 27.725 181.710 ;
        RECT 26.085 180.370 26.345 180.690 ;
        RECT 24.705 178.670 24.965 178.990 ;
        RECT 24.765 176.270 24.905 178.670 ;
        RECT 26.145 176.950 26.285 180.370 ;
        RECT 28.905 178.650 29.045 184.790 ;
        RECT 29.765 184.110 30.025 184.430 ;
        RECT 29.825 181.030 29.965 184.110 ;
        RECT 33.045 183.410 33.185 189.550 ;
        RECT 38.505 188.870 38.765 189.190 ;
        RECT 36.205 187.170 36.465 187.490 ;
        RECT 36.265 185.110 36.405 187.170 ;
        RECT 38.565 185.110 38.705 188.870 ;
        RECT 40.345 188.530 40.605 188.850 ;
        RECT 36.205 184.790 36.465 185.110 ;
        RECT 38.505 184.790 38.765 185.110 ;
        RECT 38.965 184.110 39.225 184.430 ;
        RECT 33.905 183.770 34.165 184.090 ;
        RECT 32.985 183.090 33.245 183.410 ;
        RECT 33.045 182.470 33.185 183.090 ;
        RECT 33.045 182.390 33.645 182.470 ;
        RECT 33.045 182.330 33.705 182.390 ;
        RECT 33.445 182.070 33.705 182.330 ;
        RECT 31.145 181.390 31.405 181.710 ;
        RECT 29.765 180.710 30.025 181.030 ;
        RECT 29.185 179.835 30.725 180.205 ;
        RECT 28.845 178.330 29.105 178.650 ;
        RECT 27.925 177.990 28.185 178.310 ;
        RECT 27.985 176.950 28.125 177.990 ;
        RECT 26.085 176.630 26.345 176.950 ;
        RECT 27.925 176.630 28.185 176.950 ;
        RECT 24.705 175.950 24.965 176.270 ;
        RECT 24.765 172.870 24.905 175.950 ;
        RECT 24.705 172.550 24.965 172.870 ;
        RECT 23.785 170.850 24.045 171.170 ;
        RECT 20.565 170.510 20.825 170.830 ;
        RECT 21.945 170.510 22.205 170.830 ;
        RECT 22.005 167.770 22.145 170.510 ;
        RECT 23.845 168.790 23.985 170.850 ;
        RECT 28.905 170.490 29.045 178.330 ;
        RECT 29.185 174.395 30.725 174.765 ;
        RECT 31.205 173.630 31.345 181.390 ;
        RECT 32.525 181.050 32.785 181.370 ;
        RECT 32.585 178.990 32.725 181.050 ;
        RECT 33.445 180.370 33.705 180.690 ;
        RECT 32.525 178.670 32.785 178.990 ;
        RECT 31.605 177.650 31.865 177.970 ;
        RECT 31.665 174.230 31.805 177.650 ;
        RECT 32.065 176.290 32.325 176.610 ;
        RECT 32.585 176.350 32.725 178.670 ;
        RECT 33.505 178.310 33.645 180.370 ;
        RECT 33.445 177.990 33.705 178.310 ;
        RECT 32.125 174.230 32.265 176.290 ;
        RECT 32.585 176.210 33.185 176.350 ;
        RECT 33.045 175.930 33.185 176.210 ;
        RECT 32.985 175.610 33.245 175.930 ;
        RECT 31.605 173.910 31.865 174.230 ;
        RECT 32.065 173.910 32.325 174.230 ;
        RECT 31.205 173.490 31.805 173.630 ;
        RECT 28.845 170.170 29.105 170.490 ;
        RECT 31.145 170.170 31.405 170.490 ;
        RECT 29.185 168.955 30.725 169.325 ;
        RECT 23.785 168.470 24.045 168.790 ;
        RECT 27.465 167.790 27.725 168.110 ;
        RECT 27.925 167.790 28.185 168.110 ;
        RECT 21.945 167.625 22.205 167.770 ;
        RECT 21.935 167.255 22.215 167.625 ;
        RECT 27.525 167.510 27.665 167.790 ;
        RECT 17.400 166.235 18.940 166.605 ;
        RECT 21.025 162.010 21.285 162.330 ;
        RECT 17.400 160.795 18.940 161.165 ;
        RECT 21.085 157.910 21.225 162.010 ;
        RECT 22.005 161.990 22.145 167.255 ;
        RECT 25.625 167.110 25.885 167.430 ;
        RECT 27.065 167.370 27.665 167.510 ;
        RECT 22.865 166.770 23.125 167.090 ;
        RECT 22.925 165.730 23.065 166.770 ;
        RECT 24.705 165.750 24.965 166.070 ;
        RECT 22.865 165.410 23.125 165.730 ;
        RECT 21.945 161.670 22.205 161.990 ;
        RECT 24.245 159.860 24.505 159.950 ;
        RECT 24.765 159.860 24.905 165.750 ;
        RECT 25.685 159.950 25.825 167.110 ;
        RECT 27.065 163.350 27.205 167.370 ;
        RECT 27.465 166.770 27.725 167.090 ;
        RECT 27.525 164.370 27.665 166.770 ;
        RECT 27.465 164.050 27.725 164.370 ;
        RECT 27.005 163.030 27.265 163.350 ;
        RECT 26.085 161.330 26.345 161.650 ;
        RECT 26.145 159.950 26.285 161.330 ;
        RECT 24.245 159.720 24.905 159.860 ;
        RECT 24.245 159.630 24.505 159.720 ;
        RECT 25.625 159.630 25.885 159.950 ;
        RECT 26.085 159.630 26.345 159.950 ;
        RECT 23.325 158.610 23.585 158.930 ;
        RECT 21.025 157.590 21.285 157.910 ;
        RECT 22.865 157.590 23.125 157.910 ;
        RECT 22.925 156.890 23.065 157.590 ;
        RECT 22.865 156.570 23.125 156.890 ;
        RECT 21.945 156.230 22.205 156.550 ;
        RECT 20.565 155.890 20.825 156.210 ;
        RECT 17.400 155.355 18.940 155.725 ;
        RECT 20.625 151.110 20.765 155.890 ;
        RECT 22.005 154.850 22.145 156.230 ;
        RECT 21.945 154.530 22.205 154.850 ;
        RECT 22.925 154.510 23.065 156.570 ;
        RECT 22.865 154.190 23.125 154.510 ;
        RECT 21.025 153.850 21.285 154.170 ;
        RECT 20.565 150.790 20.825 151.110 ;
        RECT 20.105 150.450 20.365 150.770 ;
        RECT 17.400 149.915 18.940 150.285 ;
        RECT 20.165 149.410 20.305 150.450 ;
        RECT 20.105 149.090 20.365 149.410 ;
        RECT 20.565 145.350 20.825 145.670 ;
        RECT 17.400 144.475 18.940 144.845 ;
        RECT 20.625 141.250 20.765 145.350 ;
        RECT 20.565 140.930 20.825 141.250 ;
        RECT 21.085 140.570 21.225 153.850 ;
        RECT 21.945 145.070 22.205 145.330 ;
        RECT 21.545 145.010 22.205 145.070 ;
        RECT 21.545 144.930 22.145 145.010 ;
        RECT 21.545 144.310 21.685 144.930 ;
        RECT 21.485 143.990 21.745 144.310 ;
        RECT 21.945 143.650 22.205 143.970 ;
        RECT 22.005 141.590 22.145 143.650 ;
        RECT 22.865 143.310 23.125 143.630 ;
        RECT 22.405 142.290 22.665 142.610 ;
        RECT 21.945 141.270 22.205 141.590 ;
        RECT 22.465 140.570 22.605 142.290 ;
        RECT 22.925 141.590 23.065 143.310 ;
        RECT 22.865 141.270 23.125 141.590 ;
        RECT 21.025 140.250 21.285 140.570 ;
        RECT 22.405 140.250 22.665 140.570 ;
        RECT 17.400 139.035 18.940 139.405 ;
        RECT 17.400 133.595 18.940 133.965 ;
        RECT 23.385 133.430 23.525 158.610 ;
        RECT 26.145 156.890 26.285 159.630 ;
        RECT 27.065 159.610 27.205 163.030 ;
        RECT 27.525 159.610 27.665 164.050 ;
        RECT 27.985 160.630 28.125 167.790 ;
        RECT 31.205 167.770 31.345 170.170 ;
        RECT 31.665 167.770 31.805 173.490 ;
        RECT 32.065 172.550 32.325 172.870 ;
        RECT 32.125 172.270 32.265 172.550 ;
        RECT 33.505 172.530 33.645 177.990 ;
        RECT 32.125 172.130 32.725 172.270 ;
        RECT 33.445 172.210 33.705 172.530 ;
        RECT 32.065 171.190 32.325 171.510 ;
        RECT 32.125 168.790 32.265 171.190 ;
        RECT 32.585 170.830 32.725 172.130 ;
        RECT 32.525 170.510 32.785 170.830 ;
        RECT 32.985 170.510 33.245 170.830 ;
        RECT 32.065 168.470 32.325 168.790 ;
        RECT 28.845 167.450 29.105 167.770 ;
        RECT 31.145 167.450 31.405 167.770 ;
        RECT 31.605 167.450 31.865 167.770 ;
        RECT 32.525 167.680 32.785 167.770 ;
        RECT 33.045 167.680 33.185 170.510 ;
        RECT 32.525 167.540 33.185 167.680 ;
        RECT 32.525 167.450 32.785 167.540 ;
        RECT 28.905 160.630 29.045 167.450 ;
        RECT 29.765 166.770 30.025 167.090 ;
        RECT 29.825 165.730 29.965 166.770 ;
        RECT 32.585 166.070 32.725 167.450 ;
        RECT 32.985 166.770 33.245 167.090 ;
        RECT 32.525 165.750 32.785 166.070 ;
        RECT 29.765 165.410 30.025 165.730 ;
        RECT 32.525 165.070 32.785 165.390 ;
        RECT 32.065 164.730 32.325 165.050 ;
        RECT 29.185 163.515 30.725 163.885 ;
        RECT 32.125 163.350 32.265 164.730 ;
        RECT 32.065 163.030 32.325 163.350 ;
        RECT 32.585 162.670 32.725 165.070 ;
        RECT 32.525 162.350 32.785 162.670 ;
        RECT 27.925 160.310 28.185 160.630 ;
        RECT 28.845 160.310 29.105 160.630 ;
        RECT 31.605 159.630 31.865 159.950 ;
        RECT 27.005 159.290 27.265 159.610 ;
        RECT 27.465 159.290 27.725 159.610 ;
        RECT 27.065 157.570 27.205 159.290 ;
        RECT 29.185 158.075 30.725 158.445 ;
        RECT 27.005 157.250 27.265 157.570 ;
        RECT 26.085 156.570 26.345 156.890 ;
        RECT 23.785 155.890 24.045 156.210 ;
        RECT 25.625 155.890 25.885 156.210 ;
        RECT 23.845 149.410 23.985 155.890 ;
        RECT 25.685 154.850 25.825 155.890 ;
        RECT 25.625 154.530 25.885 154.850 ;
        RECT 27.065 154.170 27.205 157.250 ;
        RECT 29.305 156.910 29.565 157.230 ;
        RECT 31.145 156.910 31.405 157.230 ;
        RECT 29.365 155.190 29.505 156.910 ;
        RECT 27.925 154.870 28.185 155.190 ;
        RECT 29.305 154.870 29.565 155.190 ;
        RECT 27.005 153.850 27.265 154.170 ;
        RECT 26.545 152.150 26.805 152.470 ;
        RECT 23.785 149.090 24.045 149.410 ;
        RECT 25.625 148.750 25.885 149.070 ;
        RECT 25.685 147.110 25.825 148.750 ;
        RECT 25.225 147.030 25.825 147.110 ;
        RECT 25.165 146.970 25.825 147.030 ;
        RECT 25.165 146.710 25.425 146.970 ;
        RECT 25.225 140.910 25.365 146.710 ;
        RECT 25.165 140.590 25.425 140.910 ;
        RECT 23.325 133.110 23.585 133.430 ;
        RECT 24.705 132.430 24.965 132.750 ;
        RECT 23.325 131.410 23.585 131.730 ;
        RECT 23.385 129.350 23.525 131.410 ;
        RECT 24.765 130.030 24.905 132.430 ;
        RECT 26.085 132.090 26.345 132.410 ;
        RECT 25.625 131.750 25.885 132.070 ;
        RECT 25.165 131.410 25.425 131.730 ;
        RECT 24.705 129.710 24.965 130.030 ;
        RECT 23.325 129.030 23.585 129.350 ;
        RECT 24.765 129.010 24.905 129.710 ;
        RECT 24.705 128.690 24.965 129.010 ;
        RECT 17.400 128.155 18.940 128.525 ;
        RECT 24.765 127.990 24.905 128.690 ;
        RECT 24.705 127.670 24.965 127.990 ;
        RECT 25.225 127.310 25.365 131.410 ;
        RECT 24.245 126.990 24.505 127.310 ;
        RECT 25.165 126.990 25.425 127.310 ;
        RECT 21.485 125.970 21.745 126.290 ;
        RECT 21.545 124.590 21.685 125.970 ;
        RECT 24.305 125.270 24.445 126.990 ;
        RECT 25.685 126.970 25.825 131.750 ;
        RECT 26.145 130.710 26.285 132.090 ;
        RECT 26.085 130.390 26.345 130.710 ;
        RECT 24.705 126.650 24.965 126.970 ;
        RECT 25.625 126.650 25.885 126.970 ;
        RECT 24.245 124.950 24.505 125.270 ;
        RECT 21.485 124.270 21.745 124.590 ;
        RECT 21.025 123.590 21.285 123.910 ;
        RECT 17.400 122.715 18.940 123.085 ;
        RECT 21.085 122.550 21.225 123.590 ;
        RECT 24.765 123.570 24.905 126.650 ;
        RECT 24.705 123.250 24.965 123.570 ;
        RECT 21.025 122.230 21.285 122.550 ;
        RECT 22.865 122.230 23.125 122.550 ;
        RECT 22.925 118.810 23.065 122.230 ;
        RECT 23.785 121.890 24.045 122.210 ;
        RECT 22.865 118.490 23.125 118.810 ;
        RECT 17.400 117.275 18.940 117.645 ;
        RECT 23.845 117.110 23.985 121.890 ;
        RECT 24.765 119.490 24.905 123.250 ;
        RECT 26.145 121.950 26.285 130.390 ;
        RECT 25.685 121.870 26.285 121.950 ;
        RECT 25.625 121.810 26.285 121.870 ;
        RECT 25.625 121.550 25.885 121.810 ;
        RECT 26.145 119.490 26.285 121.810 ;
        RECT 24.705 119.170 24.965 119.490 ;
        RECT 26.085 119.170 26.345 119.490 ;
        RECT 24.705 117.810 24.965 118.130 ;
        RECT 23.785 116.790 24.045 117.110 ;
        RECT 24.765 116.430 24.905 117.810 ;
        RECT 26.145 116.430 26.285 119.170 ;
        RECT 24.705 116.110 24.965 116.430 ;
        RECT 26.085 116.110 26.345 116.430 ;
        RECT 23.325 112.710 23.585 113.030 ;
        RECT 17.400 111.835 18.940 112.205 ;
        RECT 23.385 108.950 23.525 112.710 ;
        RECT 26.605 111.330 26.745 152.150 ;
        RECT 27.065 148.730 27.205 153.850 ;
        RECT 27.005 148.410 27.265 148.730 ;
        RECT 27.065 140.910 27.205 148.410 ;
        RECT 27.985 145.330 28.125 154.870 ;
        RECT 29.185 152.635 30.725 153.005 ;
        RECT 31.205 152.470 31.345 156.910 ;
        RECT 31.665 154.170 31.805 159.630 ;
        RECT 31.605 153.850 31.865 154.170 ;
        RECT 31.605 153.170 31.865 153.490 ;
        RECT 31.145 152.150 31.405 152.470 ;
        RECT 28.845 151.470 29.105 151.790 ;
        RECT 28.905 146.690 29.045 151.470 ;
        RECT 31.665 151.450 31.805 153.170 ;
        RECT 33.045 151.450 33.185 166.770 ;
        RECT 33.505 160.290 33.645 172.210 ;
        RECT 33.965 168.110 34.105 183.770 ;
        RECT 39.025 182.610 39.165 184.110 ;
        RECT 40.405 183.410 40.545 188.530 ;
        RECT 40.975 187.995 42.515 188.365 ;
        RECT 43.625 187.490 43.765 191.250 ;
        RECT 43.565 187.170 43.825 187.490 ;
        RECT 40.805 185.810 41.065 186.130 ;
        RECT 40.865 184.090 41.005 185.810 ;
        RECT 44.085 184.510 44.225 192.270 ;
        RECT 44.485 191.250 44.745 191.570 ;
        RECT 44.545 189.870 44.685 191.250 ;
        RECT 44.485 189.550 44.745 189.870 ;
        RECT 45.005 185.110 45.145 192.270 ;
        RECT 45.865 189.550 46.125 189.870 ;
        RECT 45.405 188.530 45.665 188.850 ;
        RECT 45.465 187.150 45.605 188.530 ;
        RECT 45.405 186.830 45.665 187.150 ;
        RECT 45.925 186.810 46.065 189.550 ;
        RECT 47.245 189.210 47.505 189.530 ;
        RECT 45.865 186.490 46.125 186.810 ;
        RECT 47.305 185.110 47.445 189.210 ;
        RECT 49.545 188.870 49.805 189.190 ;
        RECT 49.605 187.830 49.745 188.870 ;
        RECT 49.545 187.510 49.805 187.830 ;
        RECT 51.445 187.150 51.585 192.270 ;
        RECT 52.305 191.250 52.565 191.570 ;
        RECT 64.725 191.250 64.985 191.570 ;
        RECT 66.565 191.250 66.825 191.570 ;
        RECT 52.365 189.190 52.505 191.250 ;
        RECT 52.760 190.715 54.300 191.085 ;
        RECT 62.425 189.550 62.685 189.870 ;
        RECT 52.305 188.870 52.565 189.190 ;
        RECT 56.445 188.530 56.705 188.850 ;
        RECT 61.505 188.530 61.765 188.850 ;
        RECT 51.385 186.830 51.645 187.150 ;
        RECT 56.505 186.810 56.645 188.530 ;
        RECT 59.205 186.830 59.465 187.150 ;
        RECT 55.985 186.490 56.245 186.810 ;
        RECT 56.445 186.490 56.705 186.810 ;
        RECT 54.605 186.150 54.865 186.470 ;
        RECT 49.085 185.810 49.345 186.130 ;
        RECT 44.945 184.790 45.205 185.110 ;
        RECT 47.245 184.790 47.505 185.110 ;
        RECT 43.625 184.430 44.225 184.510 ;
        RECT 43.565 184.370 44.225 184.430 ;
        RECT 43.565 184.110 43.825 184.370 ;
        RECT 40.805 183.770 41.065 184.090 ;
        RECT 42.645 183.770 42.905 184.090 ;
        RECT 40.345 183.090 40.605 183.410 ;
        RECT 37.645 182.470 39.165 182.610 ;
        RECT 35.745 181.730 36.005 182.050 ;
        RECT 34.825 181.050 35.085 181.370 ;
        RECT 34.885 172.530 35.025 181.050 ;
        RECT 35.805 179.670 35.945 181.730 ;
        RECT 35.745 179.350 36.005 179.670 ;
        RECT 35.285 178.330 35.545 178.650 ;
        RECT 34.825 172.210 35.085 172.530 ;
        RECT 34.365 170.510 34.625 170.830 ;
        RECT 34.425 168.450 34.565 170.510 ;
        RECT 34.365 168.130 34.625 168.450 ;
        RECT 33.905 167.790 34.165 168.110 ;
        RECT 35.345 167.625 35.485 178.330 ;
        RECT 37.645 178.310 37.785 182.470 ;
        RECT 38.965 181.730 39.225 182.050 ;
        RECT 38.045 181.050 38.305 181.370 ;
        RECT 38.105 179.670 38.245 181.050 ;
        RECT 38.045 179.350 38.305 179.670 ;
        RECT 38.045 178.330 38.305 178.650 ;
        RECT 37.585 177.990 37.845 178.310 ;
        RECT 37.125 176.630 37.385 176.950 ;
        RECT 37.185 173.550 37.325 176.630 ;
        RECT 37.645 175.250 37.785 177.990 ;
        RECT 37.585 174.930 37.845 175.250 ;
        RECT 37.125 173.230 37.385 173.550 ;
        RECT 36.655 170.655 36.935 171.025 ;
        RECT 36.665 170.510 36.925 170.655 ;
        RECT 36.665 169.830 36.925 170.150 ;
        RECT 36.205 169.490 36.465 169.810 ;
        RECT 34.825 167.110 35.085 167.430 ;
        RECT 35.275 167.255 35.555 167.625 ;
        RECT 33.445 159.970 33.705 160.290 ;
        RECT 34.365 156.910 34.625 157.230 ;
        RECT 34.425 155.190 34.565 156.910 ;
        RECT 34.365 154.870 34.625 155.190 ;
        RECT 33.445 151.700 33.705 151.790 ;
        RECT 34.425 151.700 34.565 154.870 ;
        RECT 33.445 151.560 34.565 151.700 ;
        RECT 33.445 151.470 33.705 151.560 ;
        RECT 30.225 151.130 30.485 151.450 ;
        RECT 31.605 151.130 31.865 151.450 ;
        RECT 32.985 151.130 33.245 151.450 ;
        RECT 30.285 149.750 30.425 151.130 ;
        RECT 34.365 150.790 34.625 151.110 ;
        RECT 32.065 150.450 32.325 150.770 ;
        RECT 32.525 150.450 32.785 150.770 ;
        RECT 30.225 149.430 30.485 149.750 ;
        RECT 32.125 149.265 32.265 150.450 ;
        RECT 31.145 148.750 31.405 149.070 ;
        RECT 32.055 148.895 32.335 149.265 ;
        RECT 32.585 149.070 32.725 150.450 ;
        RECT 34.425 149.750 34.565 150.790 ;
        RECT 34.365 149.430 34.625 149.750 ;
        RECT 34.885 149.150 35.025 167.110 ;
        RECT 35.345 167.000 35.485 167.255 ;
        RECT 35.745 167.000 36.005 167.090 ;
        RECT 35.345 166.860 36.005 167.000 ;
        RECT 35.745 166.770 36.005 166.860 ;
        RECT 35.285 165.750 35.545 166.070 ;
        RECT 35.345 156.210 35.485 165.750 ;
        RECT 35.285 155.890 35.545 156.210 ;
        RECT 35.345 154.510 35.485 155.890 ;
        RECT 35.285 154.190 35.545 154.510 ;
        RECT 35.345 153.230 35.485 154.190 ;
        RECT 35.345 153.090 35.945 153.230 ;
        RECT 35.285 152.150 35.545 152.470 ;
        RECT 32.525 148.750 32.785 149.070 ;
        RECT 33.045 149.010 35.025 149.150 ;
        RECT 29.185 147.195 30.725 147.565 ;
        RECT 28.845 146.370 29.105 146.690 ;
        RECT 31.205 146.430 31.345 148.750 ;
        RECT 32.065 148.070 32.325 148.390 ;
        RECT 32.525 148.070 32.785 148.390 ;
        RECT 31.605 146.710 31.865 147.030 ;
        RECT 28.385 145.350 28.645 145.670 ;
        RECT 27.925 145.010 28.185 145.330 ;
        RECT 27.005 140.590 27.265 140.910 ;
        RECT 27.985 140.230 28.125 145.010 ;
        RECT 28.445 141.590 28.585 145.350 ;
        RECT 28.905 143.710 29.045 146.370 ;
        RECT 30.745 146.290 31.345 146.430 ;
        RECT 29.765 145.010 30.025 145.330 ;
        RECT 29.825 143.970 29.965 145.010 ;
        RECT 28.905 143.570 29.505 143.710 ;
        RECT 29.765 143.650 30.025 143.970 ;
        RECT 29.365 143.290 29.505 143.570 ;
        RECT 29.305 142.970 29.565 143.290 ;
        RECT 30.745 143.030 30.885 146.290 ;
        RECT 31.665 146.010 31.805 146.710 ;
        RECT 31.145 145.690 31.405 146.010 ;
        RECT 31.605 145.690 31.865 146.010 ;
        RECT 31.205 143.970 31.345 145.690 ;
        RECT 31.145 143.650 31.405 143.970 ;
        RECT 30.745 142.890 31.345 143.030 ;
        RECT 31.605 142.970 31.865 143.290 ;
        RECT 29.185 141.755 30.725 142.125 ;
        RECT 28.385 141.270 28.645 141.590 ;
        RECT 31.205 141.250 31.345 142.890 ;
        RECT 31.145 140.930 31.405 141.250 ;
        RECT 31.665 140.910 31.805 142.970 ;
        RECT 31.605 140.590 31.865 140.910 ;
        RECT 27.925 139.910 28.185 140.230 ;
        RECT 29.185 136.315 30.725 136.685 ;
        RECT 31.605 135.830 31.865 136.150 ;
        RECT 27.925 133.110 28.185 133.430 ;
        RECT 27.985 132.410 28.125 133.110 ;
        RECT 27.925 132.090 28.185 132.410 ;
        RECT 31.665 132.150 31.805 135.830 ;
        RECT 32.125 132.750 32.265 148.070 ;
        RECT 32.585 146.010 32.725 148.070 ;
        RECT 32.525 145.690 32.785 146.010 ;
        RECT 32.585 144.310 32.725 145.690 ;
        RECT 32.525 143.990 32.785 144.310 ;
        RECT 33.045 140.570 33.185 149.010 ;
        RECT 34.365 146.370 34.625 146.690 ;
        RECT 33.905 145.010 34.165 145.330 ;
        RECT 33.445 141.270 33.705 141.590 ;
        RECT 32.985 140.250 33.245 140.570 ;
        RECT 32.985 136.850 33.245 137.170 ;
        RECT 32.065 132.430 32.325 132.750 ;
        RECT 27.465 129.370 27.725 129.690 ;
        RECT 27.525 127.990 27.665 129.370 ;
        RECT 27.985 127.990 28.125 132.090 ;
        RECT 31.665 132.010 32.265 132.150 ;
        RECT 28.385 131.410 28.645 131.730 ;
        RECT 31.605 131.410 31.865 131.730 ;
        RECT 27.465 127.670 27.725 127.990 ;
        RECT 27.925 127.670 28.185 127.990 ;
        RECT 27.465 123.930 27.725 124.250 ;
        RECT 27.005 120.530 27.265 120.850 ;
        RECT 27.065 117.110 27.205 120.530 ;
        RECT 27.525 119.150 27.665 123.930 ;
        RECT 27.465 118.830 27.725 119.150 ;
        RECT 27.465 118.150 27.725 118.470 ;
        RECT 27.525 117.110 27.665 118.150 ;
        RECT 27.005 116.790 27.265 117.110 ;
        RECT 27.465 116.790 27.725 117.110 ;
        RECT 28.445 113.610 28.585 131.410 ;
        RECT 29.185 130.875 30.725 131.245 ;
        RECT 29.765 130.390 30.025 130.710 ;
        RECT 29.825 129.690 29.965 130.390 ;
        RECT 28.845 129.370 29.105 129.690 ;
        RECT 29.765 129.370 30.025 129.690 ;
        RECT 28.905 124.590 29.045 129.370 ;
        RECT 30.225 128.690 30.485 129.010 ;
        RECT 30.285 127.650 30.425 128.690 ;
        RECT 30.225 127.330 30.485 127.650 ;
        RECT 29.185 125.435 30.725 125.805 ;
        RECT 31.665 125.270 31.805 131.410 ;
        RECT 32.125 125.270 32.265 132.010 ;
        RECT 33.045 130.710 33.185 136.850 ;
        RECT 33.505 133.430 33.645 141.270 ;
        RECT 33.965 140.910 34.105 145.010 ;
        RECT 34.425 143.630 34.565 146.370 ;
        RECT 34.825 145.350 35.085 145.670 ;
        RECT 34.365 143.310 34.625 143.630 ;
        RECT 34.365 142.290 34.625 142.610 ;
        RECT 33.905 140.590 34.165 140.910 ;
        RECT 34.425 140.570 34.565 142.290 ;
        RECT 34.365 140.250 34.625 140.570 ;
        RECT 34.885 135.470 35.025 145.350 ;
        RECT 34.825 135.150 35.085 135.470 ;
        RECT 33.445 133.110 33.705 133.430 ;
        RECT 34.365 132.430 34.625 132.750 ;
        RECT 32.985 130.390 33.245 130.710 ;
        RECT 34.425 129.690 34.565 132.430 ;
        RECT 35.345 130.710 35.485 152.150 ;
        RECT 35.805 151.790 35.945 153.090 ;
        RECT 35.745 151.470 36.005 151.790 ;
        RECT 35.745 142.630 36.005 142.950 ;
        RECT 35.805 137.850 35.945 142.630 ;
        RECT 36.265 138.190 36.405 169.490 ;
        RECT 36.205 137.870 36.465 138.190 ;
        RECT 35.745 137.530 36.005 137.850 ;
        RECT 36.725 135.130 36.865 169.830 ;
        RECT 37.185 168.450 37.325 173.230 ;
        RECT 37.645 173.210 37.785 174.930 ;
        RECT 38.105 174.230 38.245 178.330 ;
        RECT 38.505 177.650 38.765 177.970 ;
        RECT 38.565 176.270 38.705 177.650 ;
        RECT 38.505 175.950 38.765 176.270 ;
        RECT 39.025 175.930 39.165 181.730 ;
        RECT 38.965 175.610 39.225 175.930 ;
        RECT 38.045 173.910 38.305 174.230 ;
        RECT 37.585 172.890 37.845 173.210 ;
        RECT 37.585 172.210 37.845 172.530 ;
        RECT 37.645 170.830 37.785 172.210 ;
        RECT 38.045 170.850 38.305 171.170 ;
        RECT 37.585 170.510 37.845 170.830 ;
        RECT 37.125 168.130 37.385 168.450 ;
        RECT 38.105 168.020 38.245 170.850 ;
        RECT 37.645 167.880 38.245 168.020 ;
        RECT 37.125 167.680 37.385 167.770 ;
        RECT 37.645 167.680 37.785 167.880 ;
        RECT 37.125 167.540 37.785 167.680 ;
        RECT 37.125 167.450 37.385 167.540 ;
        RECT 38.105 161.650 38.245 167.880 ;
        RECT 39.025 165.050 39.165 175.610 ;
        RECT 40.405 171.170 40.545 183.090 ;
        RECT 40.975 182.555 42.515 182.925 ;
        RECT 42.705 182.610 42.845 183.770 ;
        RECT 42.705 182.470 43.305 182.610 ;
        RECT 40.975 177.115 42.515 177.485 ;
        RECT 40.975 171.675 42.515 172.045 ;
        RECT 40.345 170.850 40.605 171.170 ;
        RECT 42.185 170.510 42.445 170.830 ;
        RECT 40.345 170.170 40.605 170.490 ;
        RECT 40.405 167.770 40.545 170.170 ;
        RECT 42.245 167.770 42.385 170.510 ;
        RECT 40.345 167.450 40.605 167.770 ;
        RECT 42.185 167.450 42.445 167.770 ;
        RECT 39.425 166.770 39.685 167.090 ;
        RECT 39.485 165.730 39.625 166.770 ;
        RECT 39.425 165.410 39.685 165.730 ;
        RECT 38.965 164.730 39.225 165.050 ;
        RECT 39.025 162.670 39.165 164.730 ;
        RECT 39.425 164.050 39.685 164.370 ;
        RECT 38.965 162.350 39.225 162.670 ;
        RECT 38.045 161.330 38.305 161.650 ;
        RECT 39.025 159.950 39.165 162.350 ;
        RECT 38.965 159.630 39.225 159.950 ;
        RECT 39.025 157.230 39.165 159.630 ;
        RECT 38.965 156.910 39.225 157.230 ;
        RECT 38.505 153.510 38.765 153.830 ;
        RECT 38.565 151.450 38.705 153.510 ;
        RECT 37.125 151.130 37.385 151.450 ;
        RECT 38.505 151.130 38.765 151.450 ;
        RECT 37.185 150.770 37.325 151.130 ;
        RECT 38.045 150.790 38.305 151.110 ;
        RECT 37.125 150.450 37.385 150.770 ;
        RECT 37.185 148.730 37.325 150.450 ;
        RECT 37.585 148.750 37.845 149.070 ;
        RECT 37.125 148.410 37.385 148.730 ;
        RECT 37.185 146.010 37.325 148.410 ;
        RECT 37.125 145.690 37.385 146.010 ;
        RECT 37.645 143.630 37.785 148.750 ;
        RECT 38.105 146.690 38.245 150.790 ;
        RECT 38.565 149.750 38.705 151.130 ;
        RECT 38.505 149.430 38.765 149.750 ;
        RECT 38.565 147.030 38.705 149.430 ;
        RECT 39.025 149.410 39.165 156.910 ;
        RECT 39.485 154.510 39.625 164.050 ;
        RECT 40.405 163.350 40.545 167.450 ;
        RECT 40.975 166.235 42.515 166.605 ;
        RECT 40.345 163.030 40.605 163.350 ;
        RECT 42.645 162.010 42.905 162.330 ;
        RECT 40.975 160.795 42.515 161.165 ;
        RECT 40.975 155.355 42.515 155.725 ;
        RECT 42.705 154.850 42.845 162.010 ;
        RECT 43.165 160.290 43.305 182.470 ;
        RECT 44.085 178.650 44.225 184.370 ;
        RECT 49.145 183.750 49.285 185.810 ;
        RECT 52.760 185.275 54.300 185.645 ;
        RECT 50.465 183.770 50.725 184.090 ;
        RECT 49.085 183.430 49.345 183.750 ;
        RECT 48.165 183.090 48.425 183.410 ;
        RECT 44.025 178.330 44.285 178.650 ;
        RECT 44.945 178.330 45.205 178.650 ;
        RECT 44.025 177.650 44.285 177.970 ;
        RECT 44.085 176.610 44.225 177.650 ;
        RECT 44.025 176.290 44.285 176.610 ;
        RECT 44.485 175.610 44.745 175.930 ;
        RECT 44.545 174.230 44.685 175.610 ;
        RECT 44.485 173.910 44.745 174.230 ;
        RECT 45.005 173.550 45.145 178.330 ;
        RECT 48.225 176.950 48.365 183.090 ;
        RECT 50.525 178.990 50.665 183.770 ;
        RECT 54.665 183.150 54.805 186.150 ;
        RECT 56.045 185.110 56.185 186.490 ;
        RECT 55.985 184.790 56.245 185.110 ;
        RECT 55.065 183.150 55.325 183.410 ;
        RECT 54.665 183.090 55.325 183.150 ;
        RECT 54.665 183.010 55.265 183.090 ;
        RECT 52.760 179.835 54.300 180.205 ;
        RECT 50.465 178.670 50.725 178.990 ;
        RECT 54.665 178.650 54.805 183.010 ;
        RECT 56.045 180.690 56.185 184.790 ;
        RECT 59.265 183.750 59.405 186.830 ;
        RECT 60.125 186.490 60.385 186.810 ;
        RECT 60.185 184.510 60.325 186.490 ;
        RECT 61.045 185.810 61.305 186.130 ;
        RECT 59.725 184.370 60.325 184.510 ;
        RECT 61.105 184.430 61.245 185.810 ;
        RECT 59.205 183.430 59.465 183.750 ;
        RECT 57.365 183.090 57.625 183.410 ;
        RECT 57.425 182.390 57.565 183.090 ;
        RECT 57.365 182.070 57.625 182.390 ;
        RECT 58.745 181.390 59.005 181.710 ;
        RECT 57.825 181.050 58.085 181.370 ;
        RECT 56.905 180.710 57.165 181.030 ;
        RECT 55.985 180.370 56.245 180.690 ;
        RECT 56.965 178.990 57.105 180.710 ;
        RECT 56.905 178.670 57.165 178.990 ;
        RECT 52.305 178.330 52.565 178.650 ;
        RECT 54.605 178.330 54.865 178.650 ;
        RECT 50.465 177.990 50.725 178.310 ;
        RECT 49.545 177.650 49.805 177.970 ;
        RECT 49.605 176.950 49.745 177.650 ;
        RECT 48.165 176.630 48.425 176.950 ;
        RECT 49.545 176.630 49.805 176.950 ;
        RECT 48.225 173.550 48.365 176.630 ;
        RECT 49.085 175.270 49.345 175.590 ;
        RECT 49.145 173.550 49.285 175.270 ;
        RECT 44.945 173.230 45.205 173.550 ;
        RECT 48.165 173.230 48.425 173.550 ;
        RECT 49.085 173.230 49.345 173.550 ;
        RECT 46.785 172.890 47.045 173.210 ;
        RECT 46.325 172.550 46.585 172.870 ;
        RECT 44.945 170.510 45.205 170.830 ;
        RECT 44.485 169.490 44.745 169.810 ;
        RECT 43.565 166.945 43.825 167.090 ;
        RECT 43.555 166.575 43.835 166.945 ;
        RECT 43.565 162.690 43.825 163.010 ;
        RECT 43.105 159.970 43.365 160.290 ;
        RECT 43.625 159.610 43.765 162.690 ;
        RECT 44.025 162.350 44.285 162.670 ;
        RECT 43.565 159.290 43.825 159.610 ;
        RECT 44.085 157.230 44.225 162.350 ;
        RECT 44.025 156.910 44.285 157.230 ;
        RECT 43.105 156.230 43.365 156.550 ;
        RECT 43.165 155.190 43.305 156.230 ;
        RECT 43.105 154.870 43.365 155.190 ;
        RECT 42.645 154.530 42.905 154.850 ;
        RECT 39.425 154.190 39.685 154.510 ;
        RECT 40.975 149.915 42.515 150.285 ;
        RECT 40.345 149.430 40.605 149.750 ;
        RECT 38.965 149.090 39.225 149.410 ;
        RECT 40.405 149.070 40.545 149.430 ;
        RECT 39.885 148.750 40.145 149.070 ;
        RECT 40.345 148.750 40.605 149.070 ;
        RECT 39.425 148.070 39.685 148.390 ;
        RECT 39.945 148.110 40.085 148.750 ;
        RECT 42.705 148.585 42.845 154.530 ;
        RECT 44.025 154.190 44.285 154.510 ;
        RECT 44.085 153.830 44.225 154.190 ;
        RECT 44.025 153.510 44.285 153.830 ;
        RECT 44.025 152.150 44.285 152.470 ;
        RECT 42.635 148.215 42.915 148.585 ;
        RECT 38.965 147.730 39.225 148.050 ;
        RECT 38.505 146.710 38.765 147.030 ;
        RECT 38.045 146.370 38.305 146.690 ;
        RECT 38.565 146.010 38.705 146.710 ;
        RECT 38.505 145.690 38.765 146.010 ;
        RECT 39.025 145.670 39.165 147.730 ;
        RECT 38.965 145.350 39.225 145.670 ;
        RECT 39.485 143.630 39.625 148.070 ;
        RECT 39.945 147.970 40.545 148.110 ;
        RECT 40.405 143.630 40.545 147.970 ;
        RECT 40.975 144.475 42.515 144.845 ;
        RECT 37.585 143.310 37.845 143.630 ;
        RECT 38.965 143.310 39.225 143.630 ;
        RECT 39.425 143.310 39.685 143.630 ;
        RECT 40.345 143.310 40.605 143.630 ;
        RECT 38.045 140.250 38.305 140.570 ;
        RECT 37.125 137.870 37.385 138.190 ;
        RECT 36.665 134.810 36.925 135.130 ;
        RECT 37.185 134.985 37.325 137.870 ;
        RECT 38.105 135.470 38.245 140.250 ;
        RECT 39.025 138.190 39.165 143.310 ;
        RECT 39.485 138.870 39.625 143.310 ;
        RECT 39.425 138.550 39.685 138.870 ;
        RECT 40.405 138.270 40.545 143.310 ;
        RECT 43.105 142.970 43.365 143.290 ;
        RECT 43.165 140.910 43.305 142.970 ;
        RECT 43.565 142.290 43.825 142.610 ;
        RECT 43.105 140.590 43.365 140.910 ;
        RECT 40.975 139.035 42.515 139.405 ;
        RECT 41.265 138.550 41.525 138.870 ;
        RECT 39.485 138.190 41.005 138.270 ;
        RECT 38.965 137.870 39.225 138.190 ;
        RECT 39.485 138.130 41.065 138.190 ;
        RECT 38.045 135.150 38.305 135.470 ;
        RECT 38.965 135.150 39.225 135.470 ;
        RECT 37.115 134.615 37.395 134.985 ;
        RECT 37.185 132.750 37.325 134.615 ;
        RECT 38.045 134.130 38.305 134.450 ;
        RECT 37.125 132.430 37.385 132.750 ;
        RECT 35.285 130.390 35.545 130.710 ;
        RECT 34.365 129.370 34.625 129.690 ;
        RECT 36.665 129.370 36.925 129.690 ;
        RECT 35.285 126.650 35.545 126.970 ;
        RECT 31.605 124.950 31.865 125.270 ;
        RECT 32.065 124.950 32.325 125.270 ;
        RECT 28.845 124.270 29.105 124.590 ;
        RECT 28.905 121.530 29.045 124.270 ;
        RECT 34.365 123.930 34.625 124.250 ;
        RECT 32.065 123.590 32.325 123.910 ;
        RECT 30.225 123.250 30.485 123.570 ;
        RECT 30.285 121.870 30.425 123.250 ;
        RECT 32.125 122.550 32.265 123.590 ;
        RECT 34.425 122.550 34.565 123.930 ;
        RECT 35.345 122.550 35.485 126.650 ;
        RECT 36.725 124.930 36.865 129.370 ;
        RECT 38.105 129.350 38.245 134.130 ;
        RECT 39.025 133.430 39.165 135.150 ;
        RECT 39.485 134.790 39.625 138.130 ;
        RECT 40.805 137.870 41.065 138.130 ;
        RECT 39.885 135.830 40.145 136.150 ;
        RECT 39.425 134.470 39.685 134.790 ;
        RECT 38.965 133.110 39.225 133.430 ;
        RECT 39.485 132.830 39.625 134.470 ;
        RECT 39.025 132.750 39.625 132.830 ;
        RECT 38.965 132.690 39.625 132.750 ;
        RECT 38.965 132.430 39.225 132.690 ;
        RECT 39.425 132.090 39.685 132.410 ;
        RECT 38.965 129.370 39.225 129.690 ;
        RECT 38.045 129.030 38.305 129.350 ;
        RECT 38.045 126.990 38.305 127.310 ;
        RECT 37.585 126.310 37.845 126.630 ;
        RECT 37.645 125.270 37.785 126.310 ;
        RECT 37.585 124.950 37.845 125.270 ;
        RECT 36.665 124.610 36.925 124.930 ;
        RECT 36.725 123.910 36.865 124.610 ;
        RECT 36.665 123.590 36.925 123.910 ;
        RECT 31.605 122.230 31.865 122.550 ;
        RECT 32.065 122.230 32.325 122.550 ;
        RECT 34.365 122.230 34.625 122.550 ;
        RECT 35.285 122.230 35.545 122.550 ;
        RECT 31.145 121.950 31.405 122.210 ;
        RECT 30.745 121.890 31.405 121.950 ;
        RECT 29.765 121.550 30.025 121.870 ;
        RECT 30.225 121.550 30.485 121.870 ;
        RECT 30.745 121.810 31.345 121.890 ;
        RECT 28.845 121.210 29.105 121.530 ;
        RECT 29.825 120.850 29.965 121.550 ;
        RECT 30.745 121.530 30.885 121.810 ;
        RECT 30.685 121.210 30.945 121.530 ;
        RECT 31.665 120.850 31.805 122.230 ;
        RECT 37.645 122.210 37.785 124.950 ;
        RECT 34.825 121.890 35.085 122.210 ;
        RECT 37.585 121.890 37.845 122.210 ;
        RECT 29.765 120.530 30.025 120.850 ;
        RECT 31.605 120.530 31.865 120.850 ;
        RECT 32.065 120.530 32.325 120.850 ;
        RECT 29.185 119.995 30.725 120.365 ;
        RECT 30.685 116.110 30.945 116.430 ;
        RECT 30.745 115.830 30.885 116.110 ;
        RECT 30.745 115.690 31.345 115.830 ;
        RECT 29.185 114.555 30.725 114.925 ;
        RECT 28.445 113.470 29.045 113.610 ;
        RECT 28.385 112.710 28.645 113.030 ;
        RECT 28.445 111.670 28.585 112.710 ;
        RECT 28.385 111.350 28.645 111.670 ;
        RECT 26.545 111.010 26.805 111.330 ;
        RECT 28.905 110.990 29.045 113.470 ;
        RECT 31.205 113.030 31.345 115.690 ;
        RECT 32.125 113.370 32.265 120.530 ;
        RECT 34.885 119.150 35.025 121.890 ;
        RECT 38.105 121.870 38.245 126.990 ;
        RECT 39.025 126.970 39.165 129.370 ;
        RECT 39.485 127.990 39.625 132.090 ;
        RECT 39.425 127.670 39.685 127.990 ;
        RECT 38.965 126.650 39.225 126.970 ;
        RECT 38.045 121.550 38.305 121.870 ;
        RECT 35.285 121.210 35.545 121.530 ;
        RECT 36.665 121.210 36.925 121.530 ;
        RECT 35.345 119.150 35.485 121.210 ;
        RECT 34.825 118.830 35.085 119.150 ;
        RECT 35.285 118.830 35.545 119.150 ;
        RECT 32.985 118.490 33.245 118.810 ;
        RECT 32.525 115.770 32.785 116.090 ;
        RECT 32.585 113.710 32.725 115.770 ;
        RECT 33.045 114.390 33.185 118.490 ;
        RECT 34.885 116.090 35.025 118.830 ;
        RECT 36.725 118.810 36.865 121.210 ;
        RECT 38.505 120.530 38.765 120.850 ;
        RECT 36.665 118.490 36.925 118.810 ;
        RECT 38.565 118.470 38.705 120.530 ;
        RECT 38.505 118.150 38.765 118.470 ;
        RECT 39.025 118.130 39.165 126.650 ;
        RECT 36.205 117.810 36.465 118.130 ;
        RECT 36.665 117.810 36.925 118.130 ;
        RECT 37.585 117.810 37.845 118.130 ;
        RECT 38.965 117.810 39.225 118.130 ;
        RECT 36.265 116.770 36.405 117.810 ;
        RECT 36.205 116.450 36.465 116.770 ;
        RECT 34.825 115.770 35.085 116.090 ;
        RECT 32.985 114.070 33.245 114.390 ;
        RECT 32.525 113.390 32.785 113.710 ;
        RECT 34.365 113.390 34.625 113.710 ;
        RECT 32.065 113.050 32.325 113.370 ;
        RECT 33.445 113.050 33.705 113.370 ;
        RECT 31.145 112.710 31.405 113.030 ;
        RECT 28.845 110.670 29.105 110.990 ;
        RECT 31.605 110.330 31.865 110.650 ;
        RECT 31.145 109.650 31.405 109.970 ;
        RECT 29.185 109.115 30.725 109.485 ;
        RECT 23.325 108.630 23.585 108.950 ;
        RECT 23.785 107.610 24.045 107.930 ;
        RECT 26.085 107.610 26.345 107.930 ;
        RECT 17.400 106.395 18.940 106.765 ;
        RECT 23.845 105.550 23.985 107.610 ;
        RECT 25.625 107.270 25.885 107.590 ;
        RECT 25.685 106.230 25.825 107.270 ;
        RECT 25.625 105.910 25.885 106.230 ;
        RECT 23.785 105.230 24.045 105.550 ;
        RECT 24.245 104.210 24.505 104.530 ;
        RECT 24.305 102.490 24.445 104.210 ;
        RECT 24.245 102.170 24.505 102.490 ;
        RECT 21.485 101.830 21.745 102.150 ;
        RECT 17.400 100.955 18.940 101.325 ;
        RECT 21.545 98.340 21.685 101.830 ;
        RECT 26.145 98.340 26.285 107.610 ;
        RECT 29.185 103.675 30.725 104.045 ;
        RECT 31.205 102.830 31.345 109.650 ;
        RECT 31.145 102.510 31.405 102.830 ;
        RECT 31.665 102.230 31.805 110.330 ;
        RECT 33.505 106.230 33.645 113.050 ;
        RECT 34.425 110.560 34.565 113.390 ;
        RECT 36.725 113.370 36.865 117.810 ;
        RECT 37.645 117.110 37.785 117.810 ;
        RECT 37.585 116.790 37.845 117.110 ;
        RECT 39.945 113.610 40.085 135.830 ;
        RECT 41.325 135.550 41.465 138.550 ;
        RECT 43.165 138.530 43.305 140.590 ;
        RECT 43.105 138.210 43.365 138.530 ;
        RECT 43.165 137.590 43.305 138.210 ;
        RECT 43.625 138.190 43.765 142.290 ;
        RECT 43.565 137.870 43.825 138.190 ;
        RECT 43.165 137.450 43.765 137.590 ;
        RECT 40.865 135.410 43.305 135.550 ;
        RECT 40.865 135.130 41.005 135.410 ;
        RECT 43.165 135.130 43.305 135.410 ;
        RECT 40.345 134.985 40.605 135.130 ;
        RECT 40.335 134.615 40.615 134.985 ;
        RECT 40.805 134.810 41.065 135.130 ;
        RECT 43.105 134.810 43.365 135.130 ;
        RECT 40.975 133.595 42.515 133.965 ;
        RECT 43.625 133.090 43.765 137.450 ;
        RECT 43.565 132.770 43.825 133.090 ;
        RECT 40.805 132.090 41.065 132.410 ;
        RECT 40.865 130.710 41.005 132.090 ;
        RECT 43.105 131.410 43.365 131.730 ;
        RECT 43.565 131.410 43.825 131.730 ;
        RECT 40.805 130.390 41.065 130.710 ;
        RECT 42.645 129.710 42.905 130.030 ;
        RECT 40.975 128.155 42.515 128.525 ;
        RECT 42.705 127.990 42.845 129.710 ;
        RECT 42.645 127.670 42.905 127.990 ;
        RECT 42.645 127.220 42.905 127.310 ;
        RECT 43.165 127.220 43.305 131.410 ;
        RECT 43.625 130.710 43.765 131.410 ;
        RECT 43.565 130.390 43.825 130.710 ;
        RECT 42.645 127.080 43.305 127.220 ;
        RECT 42.645 126.990 42.905 127.080 ;
        RECT 43.565 126.990 43.825 127.310 ;
        RECT 40.805 126.650 41.065 126.970 ;
        RECT 42.185 126.650 42.445 126.970 ;
        RECT 40.865 124.590 41.005 126.650 ;
        RECT 40.805 124.270 41.065 124.590 ;
        RECT 42.245 123.480 42.385 126.650 ;
        RECT 43.105 124.950 43.365 125.270 ;
        RECT 42.245 123.340 42.845 123.480 ;
        RECT 40.975 122.715 42.515 123.085 ;
        RECT 40.975 117.275 42.515 117.645 ;
        RECT 42.705 117.110 42.845 123.340 ;
        RECT 43.165 122.550 43.305 124.950 ;
        RECT 43.105 122.230 43.365 122.550 ;
        RECT 43.625 121.780 43.765 126.990 ;
        RECT 44.085 126.290 44.225 152.150 ;
        RECT 44.545 138.190 44.685 169.490 ;
        RECT 45.005 168.110 45.145 170.510 ;
        RECT 45.865 169.490 46.125 169.810 ;
        RECT 44.945 167.790 45.205 168.110 ;
        RECT 45.405 166.770 45.665 167.090 ;
        RECT 44.945 164.050 45.205 164.370 ;
        RECT 45.005 159.610 45.145 164.050 ;
        RECT 45.465 160.630 45.605 166.770 ;
        RECT 45.405 160.310 45.665 160.630 ;
        RECT 44.945 159.290 45.205 159.610 ;
        RECT 45.005 157.230 45.145 159.290 ;
        RECT 44.945 156.910 45.205 157.230 ;
        RECT 44.945 155.890 45.205 156.210 ;
        RECT 45.005 151.790 45.145 155.890 ;
        RECT 45.405 152.150 45.665 152.470 ;
        RECT 45.465 151.985 45.605 152.150 ;
        RECT 44.945 151.470 45.205 151.790 ;
        RECT 45.395 151.615 45.675 151.985 ;
        RECT 45.925 151.790 46.065 169.490 ;
        RECT 46.385 154.170 46.525 172.550 ;
        RECT 46.845 171.170 46.985 172.890 ;
        RECT 46.785 170.850 47.045 171.170 ;
        RECT 47.705 170.510 47.965 170.830 ;
        RECT 47.765 167.770 47.905 170.510 ;
        RECT 48.225 167.770 48.365 173.230 ;
        RECT 49.605 173.210 49.745 176.630 ;
        RECT 50.525 174.230 50.665 177.990 ;
        RECT 52.365 176.950 52.505 178.330 ;
        RECT 52.305 176.630 52.565 176.950 ;
        RECT 52.760 174.395 54.300 174.765 ;
        RECT 50.465 173.910 50.725 174.230 ;
        RECT 54.145 173.230 54.405 173.550 ;
        RECT 49.545 172.890 49.805 173.210 ;
        RECT 54.205 171.510 54.345 173.230 ;
        RECT 49.085 171.190 49.345 171.510 ;
        RECT 54.145 171.190 54.405 171.510 ;
        RECT 49.145 170.830 49.285 171.190 ;
        RECT 49.085 170.510 49.345 170.830 ;
        RECT 50.005 170.510 50.265 170.830 ;
        RECT 52.295 170.655 52.575 171.025 ;
        RECT 49.545 169.830 49.805 170.150 ;
        RECT 48.625 168.470 48.885 168.790 ;
        RECT 47.705 167.450 47.965 167.770 ;
        RECT 48.165 167.450 48.425 167.770 ;
        RECT 46.785 167.110 47.045 167.430 ;
        RECT 46.845 165.730 46.985 167.110 ;
        RECT 46.785 165.410 47.045 165.730 ;
        RECT 47.245 164.390 47.505 164.710 ;
        RECT 47.305 163.010 47.445 164.390 ;
        RECT 47.245 162.690 47.505 163.010 ;
        RECT 47.765 162.865 47.905 167.450 ;
        RECT 48.685 166.070 48.825 168.470 ;
        RECT 49.605 167.770 49.745 169.830 ;
        RECT 50.065 168.110 50.205 170.510 ;
        RECT 50.005 167.790 50.265 168.110 ;
        RECT 49.545 167.450 49.805 167.770 ;
        RECT 50.465 166.830 50.725 167.090 ;
        RECT 50.465 166.770 51.125 166.830 ;
        RECT 51.845 166.770 52.105 167.090 ;
        RECT 50.525 166.690 51.125 166.770 ;
        RECT 48.625 165.750 48.885 166.070 ;
        RECT 50.465 165.750 50.725 166.070 ;
        RECT 49.085 165.070 49.345 165.390 ;
        RECT 47.695 162.495 47.975 162.865 ;
        RECT 49.145 160.630 49.285 165.070 ;
        RECT 50.005 164.050 50.265 164.370 ;
        RECT 50.065 162.330 50.205 164.050 ;
        RECT 50.005 162.010 50.265 162.330 ;
        RECT 50.005 161.330 50.265 161.650 ;
        RECT 49.085 160.310 49.345 160.630 ;
        RECT 49.545 160.310 49.805 160.630 ;
        RECT 49.605 159.950 49.745 160.310 ;
        RECT 50.065 159.950 50.205 161.330 ;
        RECT 49.545 159.630 49.805 159.950 ;
        RECT 50.005 159.630 50.265 159.950 ;
        RECT 49.085 158.950 49.345 159.270 ;
        RECT 47.705 158.610 47.965 158.930 ;
        RECT 47.245 157.250 47.505 157.570 ;
        RECT 47.305 156.890 47.445 157.250 ;
        RECT 46.785 156.570 47.045 156.890 ;
        RECT 47.245 156.570 47.505 156.890 ;
        RECT 46.845 154.510 46.985 156.570 ;
        RECT 47.305 154.850 47.445 156.570 ;
        RECT 47.245 154.530 47.505 154.850 ;
        RECT 46.785 154.190 47.045 154.510 ;
        RECT 46.325 153.850 46.585 154.170 ;
        RECT 47.245 153.850 47.505 154.170 ;
        RECT 45.865 151.470 46.125 151.790 ;
        RECT 46.785 151.130 47.045 151.450 ;
        RECT 45.865 150.790 46.125 151.110 ;
        RECT 44.945 148.470 45.205 148.730 ;
        RECT 44.945 148.410 45.605 148.470 ;
        RECT 45.005 148.330 45.605 148.410 ;
        RECT 44.945 147.730 45.205 148.050 ;
        RECT 45.005 143.710 45.145 147.730 ;
        RECT 45.465 146.350 45.605 148.330 ;
        RECT 45.925 147.030 46.065 150.790 ;
        RECT 46.845 149.410 46.985 151.130 ;
        RECT 46.785 149.090 47.045 149.410 ;
        RECT 45.865 146.710 46.125 147.030 ;
        RECT 45.405 146.030 45.665 146.350 ;
        RECT 45.465 144.310 45.605 146.030 ;
        RECT 46.325 145.690 46.585 146.010 ;
        RECT 45.405 143.990 45.665 144.310 ;
        RECT 45.005 143.570 45.605 143.710 ;
        RECT 45.465 142.950 45.605 143.570 ;
        RECT 45.405 142.630 45.665 142.950 ;
        RECT 44.945 142.290 45.205 142.610 ;
        RECT 45.005 140.910 45.145 142.290 ;
        RECT 44.945 140.590 45.205 140.910 ;
        RECT 44.485 137.870 44.745 138.190 ;
        RECT 44.485 136.850 44.745 137.170 ;
        RECT 44.025 125.970 44.285 126.290 ;
        RECT 44.025 121.780 44.285 121.870 ;
        RECT 43.625 121.640 44.285 121.780 ;
        RECT 44.025 121.550 44.285 121.640 ;
        RECT 43.565 120.870 43.825 121.190 ;
        RECT 42.645 116.790 42.905 117.110 ;
        RECT 41.265 116.450 41.525 116.770 ;
        RECT 41.325 114.390 41.465 116.450 ;
        RECT 41.265 114.070 41.525 114.390 ;
        RECT 39.945 113.470 40.545 113.610 ;
        RECT 36.665 113.050 36.925 113.370 ;
        RECT 34.825 112.370 35.085 112.690 ;
        RECT 34.885 111.330 35.025 112.370 ;
        RECT 40.405 111.330 40.545 113.470 ;
        RECT 42.705 113.030 42.845 116.790 ;
        RECT 43.625 113.370 43.765 120.870 ;
        RECT 44.085 118.810 44.225 121.550 ;
        RECT 44.025 118.490 44.285 118.810 ;
        RECT 44.025 113.730 44.285 114.050 ;
        RECT 43.565 113.050 43.825 113.370 ;
        RECT 42.645 112.710 42.905 113.030 ;
        RECT 40.975 111.835 42.515 112.205 ;
        RECT 34.825 111.010 35.085 111.330 ;
        RECT 40.345 111.010 40.605 111.330 ;
        RECT 34.825 110.560 35.085 110.650 ;
        RECT 34.425 110.420 35.085 110.560 ;
        RECT 34.425 108.270 34.565 110.420 ;
        RECT 34.825 110.330 35.085 110.420 ;
        RECT 37.115 110.135 37.395 110.505 ;
        RECT 34.365 108.180 34.625 108.270 ;
        RECT 34.365 108.040 35.025 108.180 ;
        RECT 34.365 107.950 34.625 108.040 ;
        RECT 33.445 105.910 33.705 106.230 ;
        RECT 32.985 105.570 33.245 105.890 ;
        RECT 33.045 103.510 33.185 105.570 ;
        RECT 32.985 103.190 33.245 103.510 ;
        RECT 33.505 102.490 33.645 105.910 ;
        RECT 34.885 105.210 35.025 108.040 ;
        RECT 37.185 107.930 37.325 110.135 ;
        RECT 38.045 109.650 38.305 109.970 ;
        RECT 37.125 107.610 37.385 107.930 ;
        RECT 38.105 105.890 38.245 109.650 ;
        RECT 39.885 107.270 40.145 107.590 ;
        RECT 42.645 107.270 42.905 107.590 ;
        RECT 38.045 105.570 38.305 105.890 ;
        RECT 34.825 104.890 35.085 105.210 ;
        RECT 34.885 102.830 35.025 104.890 ;
        RECT 35.285 104.210 35.545 104.530 ;
        RECT 34.825 102.510 35.085 102.830 ;
        RECT 30.745 102.090 31.805 102.230 ;
        RECT 33.445 102.170 33.705 102.490 ;
        RECT 30.745 98.340 30.885 102.090 ;
        RECT 35.345 98.340 35.485 104.210 ;
        RECT 39.945 98.340 40.085 107.270 ;
        RECT 40.975 106.395 42.515 106.765 ;
        RECT 42.705 103.510 42.845 107.270 ;
        RECT 44.085 105.630 44.225 113.730 ;
        RECT 44.545 110.990 44.685 136.850 ;
        RECT 44.945 135.150 45.205 135.470 ;
        RECT 45.005 133.430 45.145 135.150 ;
        RECT 44.945 133.110 45.205 133.430 ;
        RECT 45.465 132.410 45.605 142.630 ;
        RECT 45.865 140.590 46.125 140.910 ;
        RECT 45.925 136.150 46.065 140.590 ;
        RECT 45.865 135.830 46.125 136.150 ;
        RECT 45.405 132.090 45.665 132.410 ;
        RECT 45.405 130.620 45.665 130.710 ;
        RECT 45.005 130.480 45.665 130.620 ;
        RECT 45.005 125.270 45.145 130.480 ;
        RECT 45.405 130.390 45.665 130.480 ;
        RECT 45.405 128.690 45.665 129.010 ;
        RECT 44.945 124.950 45.205 125.270 ;
        RECT 44.945 123.930 45.205 124.250 ;
        RECT 45.005 122.550 45.145 123.930 ;
        RECT 44.945 122.230 45.205 122.550 ;
        RECT 45.465 118.550 45.605 128.690 ;
        RECT 45.865 126.540 46.125 126.630 ;
        RECT 46.385 126.540 46.525 145.690 ;
        RECT 47.305 142.610 47.445 153.850 ;
        RECT 47.765 151.790 47.905 158.610 ;
        RECT 49.145 156.890 49.285 158.950 ;
        RECT 49.545 157.590 49.805 157.910 ;
        RECT 49.085 156.570 49.345 156.890 ;
        RECT 48.625 153.170 48.885 153.490 ;
        RECT 48.165 152.150 48.425 152.470 ;
        RECT 47.705 151.470 47.965 151.790 ;
        RECT 47.245 142.290 47.505 142.610 ;
        RECT 47.245 136.850 47.505 137.170 ;
        RECT 47.305 127.310 47.445 136.850 ;
        RECT 47.705 135.490 47.965 135.810 ;
        RECT 47.245 126.990 47.505 127.310 ;
        RECT 47.765 126.710 47.905 135.490 ;
        RECT 48.225 127.310 48.365 152.150 ;
        RECT 48.685 147.790 48.825 153.170 ;
        RECT 49.085 150.450 49.345 150.770 ;
        RECT 49.145 149.750 49.285 150.450 ;
        RECT 49.085 149.430 49.345 149.750 ;
        RECT 48.685 147.650 49.285 147.790 ;
        RECT 48.625 140.250 48.885 140.570 ;
        RECT 48.685 138.870 48.825 140.250 ;
        RECT 48.625 138.550 48.885 138.870 ;
        RECT 48.615 133.935 48.895 134.305 ;
        RECT 48.685 129.690 48.825 133.935 ;
        RECT 49.145 130.030 49.285 147.650 ;
        RECT 49.605 146.545 49.745 157.590 ;
        RECT 50.005 156.800 50.265 156.890 ;
        RECT 50.525 156.800 50.665 165.750 ;
        RECT 50.985 165.390 51.125 166.690 ;
        RECT 50.925 165.070 51.185 165.390 ;
        RECT 50.985 163.010 51.125 165.070 ;
        RECT 50.925 162.690 51.185 163.010 ;
        RECT 50.005 156.660 50.665 156.800 ;
        RECT 50.005 156.570 50.265 156.660 ;
        RECT 49.995 155.695 50.275 156.065 ;
        RECT 50.065 152.130 50.205 155.695 ;
        RECT 50.005 151.810 50.265 152.130 ;
        RECT 50.065 151.450 50.205 151.810 ;
        RECT 50.985 151.450 51.125 162.690 ;
        RECT 51.385 158.610 51.645 158.930 ;
        RECT 50.005 151.130 50.265 151.450 ;
        RECT 50.925 151.130 51.185 151.450 ;
        RECT 50.925 149.090 51.185 149.410 ;
        RECT 50.005 147.730 50.265 148.050 ;
        RECT 49.535 146.175 49.815 146.545 ;
        RECT 50.065 146.010 50.205 147.730 ;
        RECT 50.985 147.030 51.125 149.090 ;
        RECT 50.925 146.710 51.185 147.030 ;
        RECT 51.445 146.430 51.585 158.610 ;
        RECT 50.985 146.290 51.585 146.430 ;
        RECT 50.005 145.690 50.265 146.010 ;
        RECT 49.545 145.350 49.805 145.670 ;
        RECT 49.605 142.610 49.745 145.350 ;
        RECT 49.545 142.290 49.805 142.610 ;
        RECT 49.605 138.270 49.745 142.290 ;
        RECT 50.465 140.250 50.725 140.570 ;
        RECT 50.005 139.570 50.265 139.890 ;
        RECT 50.065 138.870 50.205 139.570 ;
        RECT 50.005 138.550 50.265 138.870 ;
        RECT 49.605 138.130 50.205 138.270 ;
        RECT 49.545 134.470 49.805 134.790 ;
        RECT 49.605 133.430 49.745 134.470 ;
        RECT 49.545 133.110 49.805 133.430 ;
        RECT 50.065 132.750 50.205 138.130 ;
        RECT 50.525 135.470 50.665 140.250 ;
        RECT 50.985 137.850 51.125 146.290 ;
        RECT 51.385 141.270 51.645 141.590 ;
        RECT 50.925 137.530 51.185 137.850 ;
        RECT 50.465 135.150 50.725 135.470 ;
        RECT 50.005 132.430 50.265 132.750 ;
        RECT 49.545 131.410 49.805 131.730 ;
        RECT 49.605 130.030 49.745 131.410 ;
        RECT 49.085 129.710 49.345 130.030 ;
        RECT 49.545 129.710 49.805 130.030 ;
        RECT 48.625 129.370 48.885 129.690 ;
        RECT 48.165 126.990 48.425 127.310 ;
        RECT 47.765 126.570 49.285 126.710 ;
        RECT 45.865 126.400 46.525 126.540 ;
        RECT 45.865 126.310 46.125 126.400 ;
        RECT 45.865 123.250 46.125 123.570 ;
        RECT 45.925 119.150 46.065 123.250 ;
        RECT 45.865 118.830 46.125 119.150 ;
        RECT 45.465 118.410 46.065 118.550 ;
        RECT 45.405 115.770 45.665 116.090 ;
        RECT 45.465 114.050 45.605 115.770 ;
        RECT 45.405 113.730 45.665 114.050 ;
        RECT 45.925 110.990 46.065 118.410 ;
        RECT 46.385 116.090 46.525 126.400 ;
        RECT 46.775 124.415 47.055 124.785 ;
        RECT 46.845 124.250 46.985 124.415 ;
        RECT 47.705 124.270 47.965 124.590 ;
        RECT 46.785 123.930 47.045 124.250 ;
        RECT 46.785 123.250 47.045 123.570 ;
        RECT 46.845 121.530 46.985 123.250 ;
        RECT 46.785 121.210 47.045 121.530 ;
        RECT 46.845 119.830 46.985 121.210 ;
        RECT 47.765 121.190 47.905 124.270 ;
        RECT 48.625 121.550 48.885 121.870 ;
        RECT 47.705 120.870 47.965 121.190 ;
        RECT 48.685 119.830 48.825 121.550 ;
        RECT 46.785 119.510 47.045 119.830 ;
        RECT 48.625 119.510 48.885 119.830 ;
        RECT 46.845 116.430 46.985 119.510 ;
        RECT 46.785 116.110 47.045 116.430 ;
        RECT 46.325 115.770 46.585 116.090 ;
        RECT 46.845 113.710 46.985 116.110 ;
        RECT 47.705 115.770 47.965 116.090 ;
        RECT 46.785 113.390 47.045 113.710 ;
        RECT 44.485 110.670 44.745 110.990 ;
        RECT 45.865 110.670 46.125 110.990 ;
        RECT 45.865 109.990 46.125 110.310 ;
        RECT 44.085 105.490 44.685 105.630 ;
        RECT 42.645 103.190 42.905 103.510 ;
        RECT 40.975 100.955 42.515 101.325 ;
        RECT 44.545 98.340 44.685 105.490 ;
        RECT 45.925 105.210 46.065 109.990 ;
        RECT 46.325 109.650 46.585 109.970 ;
        RECT 46.385 108.270 46.525 109.650 ;
        RECT 47.765 108.270 47.905 115.770 ;
        RECT 49.145 110.990 49.285 126.570 ;
        RECT 50.925 125.970 51.185 126.290 ;
        RECT 50.985 121.780 51.125 125.970 ;
        RECT 51.445 122.550 51.585 141.270 ;
        RECT 51.905 140.570 52.045 166.770 ;
        RECT 52.365 164.710 52.505 170.655 ;
        RECT 52.760 168.955 54.300 169.325 ;
        RECT 52.305 164.390 52.565 164.710 ;
        RECT 52.365 160.630 52.505 164.390 ;
        RECT 52.760 163.515 54.300 163.885 ;
        RECT 54.665 162.670 54.805 178.330 ;
        RECT 56.965 176.610 57.105 178.670 ;
        RECT 57.885 176.950 58.025 181.050 ;
        RECT 58.805 180.690 58.945 181.390 ;
        RECT 59.265 181.370 59.405 183.430 ;
        RECT 59.725 181.790 59.865 184.370 ;
        RECT 61.045 184.110 61.305 184.430 ;
        RECT 61.045 183.090 61.305 183.410 ;
        RECT 61.105 182.050 61.245 183.090 ;
        RECT 59.725 181.710 60.325 181.790 ;
        RECT 61.045 181.730 61.305 182.050 ;
        RECT 59.665 181.650 60.325 181.710 ;
        RECT 59.665 181.390 59.925 181.650 ;
        RECT 59.205 181.050 59.465 181.370 ;
        RECT 58.745 180.370 59.005 180.690 ;
        RECT 60.185 179.670 60.325 181.650 ;
        RECT 61.045 180.370 61.305 180.690 ;
        RECT 60.125 179.350 60.385 179.670 ;
        RECT 58.745 177.650 59.005 177.970 ;
        RECT 60.125 177.650 60.385 177.970 ;
        RECT 57.825 176.630 58.085 176.950 ;
        RECT 56.905 176.290 57.165 176.610 ;
        RECT 58.805 176.270 58.945 177.650 ;
        RECT 59.665 176.290 59.925 176.610 ;
        RECT 58.745 175.950 59.005 176.270 ;
        RECT 59.725 173.890 59.865 176.290 ;
        RECT 59.665 173.800 59.925 173.890 ;
        RECT 59.265 173.660 59.925 173.800 ;
        RECT 59.265 171.025 59.405 173.660 ;
        RECT 59.665 173.570 59.925 173.660 ;
        RECT 59.665 172.890 59.925 173.210 ;
        RECT 59.725 171.170 59.865 172.890 ;
        RECT 57.365 170.510 57.625 170.830 ;
        RECT 59.195 170.655 59.475 171.025 ;
        RECT 59.665 170.850 59.925 171.170 ;
        RECT 59.205 170.510 59.465 170.655 ;
        RECT 57.425 166.070 57.565 170.510 ;
        RECT 58.285 169.830 58.545 170.150 ;
        RECT 57.825 169.490 58.085 169.810 ;
        RECT 57.885 167.770 58.025 169.490 ;
        RECT 57.825 167.450 58.085 167.770 ;
        RECT 57.365 165.750 57.625 166.070 ;
        RECT 56.445 165.410 56.705 165.730 ;
        RECT 54.605 162.350 54.865 162.670 ;
        RECT 52.305 160.310 52.565 160.630 ;
        RECT 56.505 160.290 56.645 165.410 ;
        RECT 56.905 165.300 57.165 165.390 ;
        RECT 57.885 165.300 58.025 167.450 ;
        RECT 58.345 166.070 58.485 169.830 ;
        RECT 59.725 168.790 59.865 170.850 ;
        RECT 59.205 168.470 59.465 168.790 ;
        RECT 59.665 168.470 59.925 168.790 ;
        RECT 59.265 168.190 59.405 168.470 ;
        RECT 60.185 168.190 60.325 177.650 ;
        RECT 61.105 176.350 61.245 180.370 ;
        RECT 61.565 178.650 61.705 188.530 ;
        RECT 62.485 187.830 62.625 189.550 ;
        RECT 64.785 189.190 64.925 191.250 ;
        RECT 64.725 188.870 64.985 189.190 ;
        RECT 64.550 187.995 66.090 188.365 ;
        RECT 62.425 187.510 62.685 187.830 ;
        RECT 66.625 187.490 66.765 191.250 ;
        RECT 70.305 189.530 70.445 192.270 ;
        RECT 69.785 189.210 70.045 189.530 ;
        RECT 70.245 189.210 70.505 189.530 ;
        RECT 66.565 187.170 66.825 187.490 ;
        RECT 61.965 186.830 62.225 187.150 ;
        RECT 62.025 182.390 62.165 186.830 ;
        RECT 69.845 186.810 69.985 189.210 ;
        RECT 64.265 186.490 64.525 186.810 ;
        RECT 69.785 186.490 70.045 186.810 ;
        RECT 63.805 186.150 64.065 186.470 ;
        RECT 62.425 185.810 62.685 186.130 ;
        RECT 61.965 182.070 62.225 182.390 ;
        RECT 62.485 181.710 62.625 185.810 ;
        RECT 63.345 184.790 63.605 185.110 ;
        RECT 62.885 183.770 63.145 184.090 ;
        RECT 62.425 181.390 62.685 181.710 ;
        RECT 61.965 179.350 62.225 179.670 ;
        RECT 61.505 178.330 61.765 178.650 ;
        RECT 61.565 176.950 61.705 178.330 ;
        RECT 61.505 176.630 61.765 176.950 ;
        RECT 61.105 176.210 61.705 176.350 ;
        RECT 61.565 175.590 61.705 176.210 ;
        RECT 61.505 175.270 61.765 175.590 ;
        RECT 61.565 173.550 61.705 175.270 ;
        RECT 62.025 173.550 62.165 179.350 ;
        RECT 62.485 178.990 62.625 181.390 ;
        RECT 62.945 181.370 63.085 183.770 ;
        RECT 62.885 181.050 63.145 181.370 ;
        RECT 63.405 180.690 63.545 184.790 ;
        RECT 63.345 180.370 63.605 180.690 ;
        RECT 62.425 178.670 62.685 178.990 ;
        RECT 62.425 174.930 62.685 175.250 ;
        RECT 61.505 173.230 61.765 173.550 ;
        RECT 61.965 173.230 62.225 173.550 ;
        RECT 61.565 171.510 61.705 173.230 ;
        RECT 61.505 171.190 61.765 171.510 ;
        RECT 61.565 168.870 61.705 171.190 ;
        RECT 62.025 171.170 62.165 173.230 ;
        RECT 61.965 170.850 62.225 171.170 ;
        RECT 61.965 170.170 62.225 170.490 ;
        RECT 59.265 168.050 60.325 168.190 ;
        RECT 59.205 167.625 59.465 167.770 ;
        RECT 59.195 167.510 59.475 167.625 ;
        RECT 59.195 167.370 59.865 167.510 ;
        RECT 59.195 167.255 59.475 167.370 ;
        RECT 58.285 165.750 58.545 166.070 ;
        RECT 56.905 165.160 58.025 165.300 ;
        RECT 56.905 165.070 57.165 165.160 ;
        RECT 59.205 164.050 59.465 164.370 ;
        RECT 58.285 161.670 58.545 161.990 ;
        RECT 58.345 160.630 58.485 161.670 ;
        RECT 58.285 160.310 58.545 160.630 ;
        RECT 56.445 159.970 56.705 160.290 ;
        RECT 59.265 159.950 59.405 164.050 ;
        RECT 53.685 159.630 53.945 159.950 ;
        RECT 57.825 159.630 58.085 159.950 ;
        RECT 59.205 159.630 59.465 159.950 ;
        RECT 53.745 159.465 53.885 159.630 ;
        RECT 53.675 159.095 53.955 159.465 ;
        RECT 54.605 159.290 54.865 159.610 ;
        RECT 53.745 158.840 53.885 159.095 ;
        RECT 54.665 158.930 54.805 159.290 ;
        RECT 52.365 158.700 53.885 158.840 ;
        RECT 52.365 157.230 52.505 158.700 ;
        RECT 54.605 158.610 54.865 158.930 ;
        RECT 52.760 158.075 54.300 158.445 ;
        RECT 52.305 156.910 52.565 157.230 ;
        RECT 53.225 157.140 53.485 157.230 ;
        RECT 52.825 157.000 53.485 157.140 ;
        RECT 52.305 155.890 52.565 156.210 ;
        RECT 52.365 140.910 52.505 155.890 ;
        RECT 52.825 154.510 52.965 157.000 ;
        RECT 53.225 156.910 53.485 157.000 ;
        RECT 54.665 156.890 54.805 158.610 ;
        RECT 57.365 157.590 57.625 157.910 ;
        RECT 57.425 156.890 57.565 157.590 ;
        RECT 57.885 157.230 58.025 159.630 ;
        RECT 57.825 156.910 58.085 157.230 ;
        RECT 54.605 156.570 54.865 156.890 ;
        RECT 57.365 156.570 57.625 156.890 ;
        RECT 57.825 155.890 58.085 156.210 ;
        RECT 59.205 156.065 59.465 156.210 ;
        RECT 57.885 154.850 58.025 155.890 ;
        RECT 59.195 155.695 59.475 156.065 ;
        RECT 57.825 154.530 58.085 154.850 ;
        RECT 52.765 154.190 53.025 154.510 ;
        RECT 55.065 153.170 55.325 153.490 ;
        RECT 52.760 152.635 54.300 153.005 ;
        RECT 52.765 151.470 53.025 151.790 ;
        RECT 52.825 148.050 52.965 151.470 ;
        RECT 54.605 151.130 54.865 151.450 ;
        RECT 52.765 147.730 53.025 148.050 ;
        RECT 52.760 147.195 54.300 147.565 ;
        RECT 54.665 147.030 54.805 151.130 ;
        RECT 55.125 150.770 55.265 153.170 ;
        RECT 57.365 152.150 57.625 152.470 ;
        RECT 55.525 151.470 55.785 151.790 ;
        RECT 55.065 150.450 55.325 150.770 ;
        RECT 54.605 146.710 54.865 147.030 ;
        RECT 55.125 146.010 55.265 150.450 ;
        RECT 55.585 149.945 55.725 151.470 ;
        RECT 55.515 149.575 55.795 149.945 ;
        RECT 55.585 146.350 55.725 149.575 ;
        RECT 57.425 148.640 57.565 152.150 ;
        RECT 59.725 151.985 59.865 167.370 ;
        RECT 60.185 165.390 60.325 168.050 ;
        RECT 61.105 168.730 61.705 168.870 ;
        RECT 61.105 167.770 61.245 168.730 ;
        RECT 61.505 168.130 61.765 168.450 ;
        RECT 61.045 167.450 61.305 167.770 ;
        RECT 60.125 165.070 60.385 165.390 ;
        RECT 60.125 164.050 60.385 164.370 ;
        RECT 60.185 161.650 60.325 164.050 ;
        RECT 61.565 162.330 61.705 168.130 ;
        RECT 62.025 168.110 62.165 170.170 ;
        RECT 61.965 167.790 62.225 168.110 ;
        RECT 61.965 162.865 62.225 163.010 ;
        RECT 61.955 162.495 62.235 162.865 ;
        RECT 61.505 162.010 61.765 162.330 ;
        RECT 60.125 161.330 60.385 161.650 ;
        RECT 61.565 159.950 61.705 162.010 ;
        RECT 62.025 160.630 62.165 162.495 ;
        RECT 61.965 160.310 62.225 160.630 ;
        RECT 61.505 159.630 61.765 159.950 ;
        RECT 60.115 159.095 60.395 159.465 ;
        RECT 60.185 156.210 60.325 159.095 ;
        RECT 61.505 158.610 61.765 158.930 ;
        RECT 61.045 157.590 61.305 157.910 ;
        RECT 60.125 155.890 60.385 156.210 ;
        RECT 59.655 151.615 59.935 151.985 ;
        RECT 58.745 150.450 59.005 150.770 ;
        RECT 58.805 149.070 58.945 150.450 ;
        RECT 58.745 148.750 59.005 149.070 ;
        RECT 60.575 148.895 60.855 149.265 ;
        RECT 57.825 148.640 58.085 148.730 ;
        RECT 57.425 148.500 58.085 148.640 ;
        RECT 55.985 146.710 56.245 147.030 ;
        RECT 55.525 146.030 55.785 146.350 ;
        RECT 55.065 145.690 55.325 146.010 ;
        RECT 54.595 142.775 54.875 143.145 ;
        RECT 54.605 142.630 54.865 142.775 ;
        RECT 52.760 141.755 54.300 142.125 ;
        RECT 52.305 140.590 52.565 140.910 ;
        RECT 51.845 140.250 52.105 140.570 ;
        RECT 55.585 137.850 55.725 146.030 ;
        RECT 56.045 146.010 56.185 146.710 ;
        RECT 55.985 145.690 56.245 146.010 ;
        RECT 56.045 140.910 56.185 145.690 ;
        RECT 57.425 145.670 57.565 148.500 ;
        RECT 57.825 148.410 58.085 148.500 ;
        RECT 58.285 148.070 58.545 148.390 ;
        RECT 58.345 146.690 58.485 148.070 ;
        RECT 58.285 146.370 58.545 146.690 ;
        RECT 57.365 145.350 57.625 145.670 ;
        RECT 55.985 140.590 56.245 140.910 ;
        RECT 57.425 140.480 57.565 145.350 ;
        RECT 58.345 140.570 58.485 146.370 ;
        RECT 58.745 145.010 59.005 145.330 ;
        RECT 58.805 140.570 58.945 145.010 ;
        RECT 57.825 140.480 58.085 140.570 ;
        RECT 57.425 140.340 58.085 140.480 ;
        RECT 57.825 140.250 58.085 140.340 ;
        RECT 58.285 140.250 58.545 140.570 ;
        RECT 58.745 140.250 59.005 140.570 ;
        RECT 59.665 140.250 59.925 140.570 ;
        RECT 57.885 138.190 58.025 140.250 ;
        RECT 58.345 138.190 58.485 140.250 ;
        RECT 59.725 138.190 59.865 140.250 ;
        RECT 60.125 138.550 60.385 138.870 ;
        RECT 57.825 137.870 58.085 138.190 ;
        RECT 58.285 137.870 58.545 138.190 ;
        RECT 58.745 137.870 59.005 138.190 ;
        RECT 59.665 137.870 59.925 138.190 ;
        RECT 55.525 137.530 55.785 137.850 ;
        RECT 55.065 137.190 55.325 137.510 ;
        RECT 52.760 136.315 54.300 136.685 ;
        RECT 53.685 135.830 53.945 136.150 ;
        RECT 52.305 135.150 52.565 135.470 ;
        RECT 53.225 135.380 53.485 135.470 ;
        RECT 52.825 135.240 53.485 135.380 ;
        RECT 51.845 131.410 52.105 131.730 ;
        RECT 51.905 129.690 52.045 131.410 ;
        RECT 51.845 129.370 52.105 129.690 ;
        RECT 52.365 129.350 52.505 135.150 ;
        RECT 52.825 132.070 52.965 135.240 ;
        RECT 53.225 135.150 53.485 135.240 ;
        RECT 53.745 132.750 53.885 135.830 ;
        RECT 54.605 134.130 54.865 134.450 ;
        RECT 54.665 132.750 54.805 134.130 ;
        RECT 53.685 132.430 53.945 132.750 ;
        RECT 54.145 132.430 54.405 132.750 ;
        RECT 54.605 132.430 54.865 132.750 ;
        RECT 53.745 132.070 53.885 132.430 ;
        RECT 52.765 131.750 53.025 132.070 ;
        RECT 53.685 131.750 53.945 132.070 ;
        RECT 54.205 131.730 54.345 132.430 ;
        RECT 54.145 131.410 54.405 131.730 ;
        RECT 52.760 130.875 54.300 131.245 ;
        RECT 52.305 129.030 52.565 129.350 ;
        RECT 52.365 127.310 52.505 129.030 ;
        RECT 52.305 126.990 52.565 127.310 ;
        RECT 51.845 126.650 52.105 126.970 ;
        RECT 51.385 122.230 51.645 122.550 ;
        RECT 51.905 121.870 52.045 126.650 ;
        RECT 52.365 125.270 52.505 126.990 ;
        RECT 52.760 125.435 54.300 125.805 ;
        RECT 52.305 124.950 52.565 125.270 ;
        RECT 51.385 121.780 51.645 121.870 ;
        RECT 50.985 121.640 51.645 121.780 ;
        RECT 51.385 121.550 51.645 121.640 ;
        RECT 51.845 121.550 52.105 121.870 ;
        RECT 51.905 119.830 52.045 121.550 ;
        RECT 52.365 120.850 52.505 124.950 ;
        RECT 53.225 123.590 53.485 123.910 ;
        RECT 52.765 122.230 53.025 122.550 ;
        RECT 52.825 121.870 52.965 122.230 ;
        RECT 52.765 121.550 53.025 121.870 ;
        RECT 53.285 121.530 53.425 123.590 ;
        RECT 53.685 123.250 53.945 123.570 ;
        RECT 55.125 123.310 55.265 137.190 ;
        RECT 55.585 135.470 55.725 137.530 ;
        RECT 58.805 135.470 58.945 137.870 ;
        RECT 60.185 136.150 60.325 138.550 ;
        RECT 60.125 135.830 60.385 136.150 ;
        RECT 55.525 135.150 55.785 135.470 ;
        RECT 58.745 135.150 59.005 135.470 ;
        RECT 55.585 130.030 55.725 135.150 ;
        RECT 55.985 134.985 56.245 135.130 ;
        RECT 55.975 134.615 56.255 134.985 ;
        RECT 56.045 133.090 56.185 134.615 ;
        RECT 57.365 134.130 57.625 134.450 ;
        RECT 60.125 134.310 60.385 134.450 ;
        RECT 59.725 134.170 60.385 134.310 ;
        RECT 60.645 134.305 60.785 148.895 ;
        RECT 61.105 146.010 61.245 157.590 ;
        RECT 61.565 151.110 61.705 158.610 ;
        RECT 61.505 150.790 61.765 151.110 ;
        RECT 62.025 149.070 62.165 160.310 ;
        RECT 62.485 154.510 62.625 174.930 ;
        RECT 63.865 173.550 64.005 186.150 ;
        RECT 64.325 184.430 64.465 186.490 ;
        RECT 65.645 184.790 65.905 185.110 ;
        RECT 64.265 184.110 64.525 184.430 ;
        RECT 65.705 183.750 65.845 184.790 ;
        RECT 69.325 184.110 69.585 184.430 ;
        RECT 66.565 183.770 66.825 184.090 ;
        RECT 68.405 183.770 68.665 184.090 ;
        RECT 65.645 183.430 65.905 183.750 ;
        RECT 64.550 182.555 66.090 182.925 ;
        RECT 66.625 180.690 66.765 183.770 ;
        RECT 68.465 183.410 68.605 183.770 ;
        RECT 68.405 183.090 68.665 183.410 ;
        RECT 66.565 180.370 66.825 180.690 ;
        RECT 68.465 178.650 68.605 183.090 ;
        RECT 69.385 182.050 69.525 184.110 ;
        RECT 69.325 181.730 69.585 182.050 ;
        RECT 70.305 178.990 70.445 189.210 ;
        RECT 74.845 188.870 75.105 189.190 ;
        RECT 74.385 186.830 74.645 187.150 ;
        RECT 71.165 185.810 71.425 186.130 ;
        RECT 71.225 185.110 71.365 185.810 ;
        RECT 71.165 184.790 71.425 185.110 ;
        RECT 71.625 184.790 71.885 185.110 ;
        RECT 71.685 184.430 71.825 184.790 ;
        RECT 71.625 184.110 71.885 184.430 ;
        RECT 74.445 184.090 74.585 186.830 ;
        RECT 74.905 185.110 75.045 188.870 ;
        RECT 75.365 186.130 75.505 192.270 ;
        RECT 75.765 191.930 76.025 192.250 ;
        RECT 78.525 191.930 78.785 192.250 ;
        RECT 75.825 186.130 75.965 191.930 ;
        RECT 76.335 190.715 77.875 191.085 ;
        RECT 78.585 188.850 78.725 191.930 ;
        RECT 82.665 191.250 82.925 191.570 ;
        RECT 81.745 189.210 82.005 189.530 ;
        RECT 78.525 188.530 78.785 188.850 ;
        RECT 78.585 187.830 78.725 188.530 ;
        RECT 78.525 187.510 78.785 187.830 ;
        RECT 75.305 185.810 75.565 186.130 ;
        RECT 75.765 185.810 76.025 186.130 ;
        RECT 74.845 184.790 75.105 185.110 ;
        RECT 74.385 183.770 74.645 184.090 ;
        RECT 71.625 183.090 71.885 183.410 ;
        RECT 71.685 182.610 71.825 183.090 ;
        RECT 70.765 182.470 71.825 182.610 ;
        RECT 70.245 178.670 70.505 178.990 ;
        RECT 68.405 178.330 68.665 178.650 ;
        RECT 67.485 177.650 67.745 177.970 ;
        RECT 64.550 177.115 66.090 177.485 ;
        RECT 67.545 176.610 67.685 177.650 ;
        RECT 67.485 176.290 67.745 176.610 ;
        RECT 63.805 173.230 64.065 173.550 ;
        RECT 63.345 172.550 63.605 172.870 ;
        RECT 62.885 170.850 63.145 171.170 ;
        RECT 62.945 168.110 63.085 170.850 ;
        RECT 62.885 167.790 63.145 168.110 ;
        RECT 62.885 166.770 63.145 167.090 ;
        RECT 62.945 165.730 63.085 166.770 ;
        RECT 62.885 165.410 63.145 165.730 ;
        RECT 62.425 154.190 62.685 154.510 ;
        RECT 62.485 151.450 62.625 154.190 ;
        RECT 62.885 153.850 63.145 154.170 ;
        RECT 62.425 151.130 62.685 151.450 ;
        RECT 61.505 148.750 61.765 149.070 ;
        RECT 61.965 148.750 62.225 149.070 ;
        RECT 61.045 145.690 61.305 146.010 ;
        RECT 61.565 145.670 61.705 148.750 ;
        RECT 62.485 146.010 62.625 151.130 ;
        RECT 62.945 149.750 63.085 153.850 ;
        RECT 62.885 149.430 63.145 149.750 ;
        RECT 62.875 146.175 63.155 146.545 ;
        RECT 62.425 145.690 62.685 146.010 ;
        RECT 61.505 145.350 61.765 145.670 ;
        RECT 61.565 144.310 61.705 145.350 ;
        RECT 61.505 143.990 61.765 144.310 ;
        RECT 61.045 143.310 61.305 143.630 ;
        RECT 61.105 134.985 61.245 143.310 ;
        RECT 62.425 139.570 62.685 139.890 ;
        RECT 62.485 138.870 62.625 139.570 ;
        RECT 62.425 138.550 62.685 138.870 ;
        RECT 62.945 137.590 63.085 146.175 ;
        RECT 63.405 138.190 63.545 172.550 ;
        RECT 63.865 168.020 64.005 173.230 ;
        RECT 66.565 172.550 66.825 172.870 ;
        RECT 64.550 171.675 66.090 172.045 ;
        RECT 64.265 171.025 64.525 171.170 ;
        RECT 64.255 170.655 64.535 171.025 ;
        RECT 64.325 170.060 64.465 170.655 ;
        RECT 64.725 170.060 64.985 170.150 ;
        RECT 64.325 169.920 64.985 170.060 ;
        RECT 64.725 169.830 64.985 169.920 ;
        RECT 64.785 168.450 64.925 169.830 ;
        RECT 64.725 168.130 64.985 168.450 ;
        RECT 64.265 168.020 64.525 168.110 ;
        RECT 63.865 167.880 64.525 168.020 ;
        RECT 64.265 167.790 64.525 167.880 ;
        RECT 66.105 167.790 66.365 168.110 ;
        RECT 64.725 167.450 64.985 167.770 ;
        RECT 66.165 167.625 66.305 167.790 ;
        RECT 64.785 167.000 64.925 167.450 ;
        RECT 66.095 167.255 66.375 167.625 ;
        RECT 66.625 167.090 66.765 172.550 ;
        RECT 67.485 170.510 67.745 170.830 ;
        RECT 67.545 170.150 67.685 170.510 ;
        RECT 68.465 170.490 68.605 178.330 ;
        RECT 70.245 172.210 70.505 172.530 ;
        RECT 68.405 170.170 68.665 170.490 ;
        RECT 67.485 169.830 67.745 170.150 ;
        RECT 67.945 169.830 68.205 170.150 ;
        RECT 67.025 169.490 67.285 169.810 ;
        RECT 67.085 168.790 67.225 169.490 ;
        RECT 67.025 168.470 67.285 168.790 ;
        RECT 63.865 166.860 64.925 167.000 ;
        RECT 63.865 165.390 64.005 166.860 ;
        RECT 66.565 166.770 66.825 167.090 ;
        RECT 64.550 166.235 66.090 166.605 ;
        RECT 63.805 165.070 64.065 165.390 ;
        RECT 65.645 165.070 65.905 165.390 ;
        RECT 63.805 164.050 64.065 164.370 ;
        RECT 64.265 164.050 64.525 164.370 ;
        RECT 63.865 159.950 64.005 164.050 ;
        RECT 64.325 163.010 64.465 164.050 ;
        RECT 65.705 163.350 65.845 165.070 ;
        RECT 66.105 164.730 66.365 165.050 ;
        RECT 65.645 163.030 65.905 163.350 ;
        RECT 64.265 162.690 64.525 163.010 ;
        RECT 66.165 161.650 66.305 164.730 ;
        RECT 67.085 162.330 67.225 168.470 ;
        RECT 66.565 162.010 66.825 162.330 ;
        RECT 67.025 162.010 67.285 162.330 ;
        RECT 68.005 162.070 68.145 169.830 ;
        RECT 68.395 167.255 68.675 167.625 ;
        RECT 68.465 164.370 68.605 167.255 ;
        RECT 70.305 165.050 70.445 172.210 ;
        RECT 69.785 164.730 70.045 165.050 ;
        RECT 70.245 164.730 70.505 165.050 ;
        RECT 68.405 164.050 68.665 164.370 ;
        RECT 68.865 164.050 69.125 164.370 ;
        RECT 66.105 161.330 66.365 161.650 ;
        RECT 64.550 160.795 66.090 161.165 ;
        RECT 66.625 159.950 66.765 162.010 ;
        RECT 68.005 161.930 68.605 162.070 ;
        RECT 67.945 161.330 68.205 161.650 ;
        RECT 68.005 160.290 68.145 161.330 ;
        RECT 67.945 159.970 68.205 160.290 ;
        RECT 63.805 159.630 64.065 159.950 ;
        RECT 66.565 159.630 66.825 159.950 ;
        RECT 63.865 157.230 64.005 159.630 ;
        RECT 63.805 156.910 64.065 157.230 ;
        RECT 63.795 155.695 64.075 156.065 ;
        RECT 63.865 152.130 64.005 155.695 ;
        RECT 64.550 155.355 66.090 155.725 ;
        RECT 66.625 155.190 66.765 159.630 ;
        RECT 68.005 156.890 68.145 159.970 ;
        RECT 67.945 156.570 68.205 156.890 ;
        RECT 66.565 155.100 66.825 155.190 ;
        RECT 65.245 154.960 66.825 155.100 ;
        RECT 64.715 154.335 64.995 154.705 ;
        RECT 64.785 154.170 64.925 154.335 ;
        RECT 64.725 153.850 64.985 154.170 ;
        RECT 63.805 151.810 64.065 152.130 ;
        RECT 63.805 151.305 64.065 151.450 ;
        RECT 63.795 150.935 64.075 151.305 ;
        RECT 63.805 150.450 64.065 150.770 ;
        RECT 65.245 150.680 65.385 154.960 ;
        RECT 66.565 154.870 66.825 154.960 ;
        RECT 68.465 154.850 68.605 161.930 ;
        RECT 66.095 154.335 66.375 154.705 ;
        RECT 68.405 154.530 68.665 154.850 ;
        RECT 66.165 154.170 66.305 154.335 ;
        RECT 67.485 154.190 67.745 154.510 ;
        RECT 66.105 153.850 66.365 154.170 ;
        RECT 66.105 153.400 66.365 153.490 ;
        RECT 65.705 153.260 66.365 153.400 ;
        RECT 65.705 151.450 65.845 153.260 ;
        RECT 66.105 153.170 66.365 153.260 ;
        RECT 67.545 151.985 67.685 154.190 ;
        RECT 67.935 153.655 68.215 154.025 ;
        RECT 68.005 153.490 68.145 153.655 ;
        RECT 67.945 153.170 68.205 153.490 ;
        RECT 67.025 151.470 67.285 151.790 ;
        RECT 67.475 151.615 67.755 151.985 ;
        RECT 65.645 151.130 65.905 151.450 ;
        RECT 66.565 151.130 66.825 151.450 ;
        RECT 66.625 150.680 66.765 151.130 ;
        RECT 65.245 150.540 66.765 150.680 ;
        RECT 63.865 149.750 64.005 150.450 ;
        RECT 64.550 149.915 66.090 150.285 ;
        RECT 63.805 149.430 64.065 149.750 ;
        RECT 64.725 149.265 64.985 149.410 ;
        RECT 64.715 148.895 64.995 149.265 ;
        RECT 66.625 149.070 66.765 150.540 ;
        RECT 67.085 149.410 67.225 151.470 ;
        RECT 68.465 151.450 68.605 154.530 ;
        RECT 68.405 151.190 68.665 151.450 ;
        RECT 67.545 151.130 68.665 151.190 ;
        RECT 67.545 151.050 68.605 151.130 ;
        RECT 67.025 149.090 67.285 149.410 ;
        RECT 67.545 149.070 67.685 151.050 ;
        RECT 67.945 150.450 68.205 150.770 ;
        RECT 68.405 150.450 68.665 150.770 ;
        RECT 66.565 148.750 66.825 149.070 ;
        RECT 67.485 148.750 67.745 149.070 ;
        RECT 66.555 148.215 66.835 148.585 ;
        RECT 67.475 148.215 67.755 148.585 ;
        RECT 66.565 148.070 66.825 148.215 ;
        RECT 67.485 148.070 67.745 148.215 ;
        RECT 66.625 147.790 66.765 148.070 ;
        RECT 66.625 147.650 67.685 147.790 ;
        RECT 63.805 145.010 64.065 145.330 ;
        RECT 66.565 145.010 66.825 145.330 ;
        RECT 63.865 143.970 64.005 145.010 ;
        RECT 64.550 144.475 66.090 144.845 ;
        RECT 63.805 143.650 64.065 143.970 ;
        RECT 66.625 140.820 66.765 145.010 ;
        RECT 66.625 140.680 67.225 140.820 ;
        RECT 66.565 139.910 66.825 140.230 ;
        RECT 64.550 139.035 66.090 139.405 ;
        RECT 66.625 138.870 66.765 139.910 ;
        RECT 66.565 138.550 66.825 138.870 ;
        RECT 67.085 138.270 67.225 140.680 ;
        RECT 66.625 138.190 67.225 138.270 ;
        RECT 63.345 137.870 63.605 138.190 ;
        RECT 66.625 138.130 67.285 138.190 ;
        RECT 62.945 137.450 64.005 137.590 ;
        RECT 61.505 136.850 61.765 137.170 ;
        RECT 61.035 134.615 61.315 134.985 ;
        RECT 55.985 132.770 56.245 133.090 ;
        RECT 57.425 131.730 57.565 134.130 ;
        RECT 59.725 133.510 59.865 134.170 ;
        RECT 60.125 134.130 60.385 134.170 ;
        RECT 60.575 133.935 60.855 134.305 ;
        RECT 61.565 133.510 61.705 136.850 ;
        RECT 61.965 135.830 62.225 136.150 ;
        RECT 63.345 135.830 63.605 136.150 ;
        RECT 59.725 133.430 60.325 133.510 ;
        RECT 59.725 133.370 60.385 133.430 ;
        RECT 60.125 133.110 60.385 133.370 ;
        RECT 60.645 133.370 61.705 133.510 ;
        RECT 58.285 132.430 58.545 132.750 ;
        RECT 57.365 131.410 57.625 131.730 ;
        RECT 57.425 130.030 57.565 131.410 ;
        RECT 58.345 130.030 58.485 132.430 ;
        RECT 55.525 129.710 55.785 130.030 ;
        RECT 57.365 129.710 57.625 130.030 ;
        RECT 58.285 129.710 58.545 130.030 ;
        RECT 60.645 127.650 60.785 133.370 ;
        RECT 61.045 132.770 61.305 133.090 ;
        RECT 62.025 132.830 62.165 135.830 ;
        RECT 62.415 133.935 62.695 134.305 ;
        RECT 61.105 130.370 61.245 132.770 ;
        RECT 61.565 132.690 62.165 132.830 ;
        RECT 61.045 130.050 61.305 130.370 ;
        RECT 60.585 127.330 60.845 127.650 ;
        RECT 59.665 125.970 59.925 126.290 ;
        RECT 61.045 125.970 61.305 126.290 ;
        RECT 59.725 125.270 59.865 125.970 ;
        RECT 59.665 124.950 59.925 125.270 ;
        RECT 61.105 124.590 61.245 125.970 ;
        RECT 61.045 124.270 61.305 124.590 ;
        RECT 57.825 123.590 58.085 123.910 ;
        RECT 53.745 121.530 53.885 123.250 ;
        RECT 55.125 123.170 55.725 123.310 ;
        RECT 55.065 122.230 55.325 122.550 ;
        RECT 53.225 121.210 53.485 121.530 ;
        RECT 53.685 121.210 53.945 121.530 ;
        RECT 54.605 121.210 54.865 121.530 ;
        RECT 52.305 120.530 52.565 120.850 ;
        RECT 51.845 119.510 52.105 119.830 ;
        RECT 52.365 119.150 52.505 120.530 ;
        RECT 52.760 119.995 54.300 120.365 ;
        RECT 52.305 118.830 52.565 119.150 ;
        RECT 54.665 118.470 54.805 121.210 ;
        RECT 55.125 121.190 55.265 122.230 ;
        RECT 55.065 120.870 55.325 121.190 ;
        RECT 54.605 118.150 54.865 118.470 ;
        RECT 55.125 117.870 55.265 120.870 ;
        RECT 54.665 117.730 55.265 117.870 ;
        RECT 54.665 117.110 54.805 117.730 ;
        RECT 54.605 116.790 54.865 117.110 ;
        RECT 52.305 115.090 52.565 115.410 ;
        RECT 52.365 113.030 52.505 115.090 ;
        RECT 52.760 114.555 54.300 114.925 ;
        RECT 52.305 112.710 52.565 113.030 ;
        RECT 49.085 110.670 49.345 110.990 ;
        RECT 55.065 110.330 55.325 110.650 ;
        RECT 52.760 109.115 54.300 109.485 ;
        RECT 46.325 107.950 46.585 108.270 ;
        RECT 47.705 107.950 47.965 108.270 ;
        RECT 54.605 107.950 54.865 108.270 ;
        RECT 52.765 107.270 53.025 107.590 ;
        RECT 52.825 106.230 52.965 107.270 ;
        RECT 52.765 105.910 53.025 106.230 ;
        RECT 45.865 104.890 46.125 105.210 ;
        RECT 49.085 104.890 49.345 105.210 ;
        RECT 49.145 98.340 49.285 104.890 ;
        RECT 52.760 103.675 54.300 104.045 ;
        RECT 54.665 102.910 54.805 107.950 ;
        RECT 55.125 105.890 55.265 110.330 ;
        RECT 55.065 105.570 55.325 105.890 ;
        RECT 53.745 102.770 54.805 102.910 ;
        RECT 53.745 98.340 53.885 102.770 ;
        RECT 55.125 102.490 55.265 105.570 ;
        RECT 55.585 105.550 55.725 123.170 ;
        RECT 57.885 122.210 58.025 123.590 ;
        RECT 57.825 121.890 58.085 122.210 ;
        RECT 56.905 116.450 57.165 116.770 ;
        RECT 56.965 114.390 57.105 116.450 ;
        RECT 56.905 114.070 57.165 114.390 ;
        RECT 57.885 113.370 58.025 121.890 ;
        RECT 61.045 121.550 61.305 121.870 ;
        RECT 59.665 120.870 59.925 121.190 ;
        RECT 59.725 118.470 59.865 120.870 ;
        RECT 59.665 118.150 59.925 118.470 ;
        RECT 60.125 116.110 60.385 116.430 ;
        RECT 59.205 115.770 59.465 116.090 ;
        RECT 59.265 114.390 59.405 115.770 ;
        RECT 59.205 114.070 59.465 114.390 ;
        RECT 57.825 113.050 58.085 113.370 ;
        RECT 59.665 111.010 59.925 111.330 ;
        RECT 57.365 107.270 57.625 107.590 ;
        RECT 57.425 106.230 57.565 107.270 ;
        RECT 57.365 105.910 57.625 106.230 ;
        RECT 55.525 105.230 55.785 105.550 ;
        RECT 58.285 105.230 58.545 105.550 ;
        RECT 57.825 104.890 58.085 105.210 ;
        RECT 57.885 102.910 58.025 104.890 ;
        RECT 58.345 103.510 58.485 105.230 ;
        RECT 59.725 103.510 59.865 111.010 ;
        RECT 60.185 108.270 60.325 116.110 ;
        RECT 61.105 111.670 61.245 121.550 ;
        RECT 61.045 111.350 61.305 111.670 ;
        RECT 60.125 107.950 60.385 108.270 ;
        RECT 60.185 105.210 60.325 107.950 ;
        RECT 61.565 107.930 61.705 132.690 ;
        RECT 61.965 132.090 62.225 132.410 ;
        RECT 62.025 130.710 62.165 132.090 ;
        RECT 61.965 130.390 62.225 130.710 ;
        RECT 62.485 130.110 62.625 133.935 ;
        RECT 63.405 132.750 63.545 135.830 ;
        RECT 63.865 132.830 64.005 137.450 ;
        RECT 66.625 136.150 66.765 138.130 ;
        RECT 67.025 137.870 67.285 138.130 ;
        RECT 66.565 135.830 66.825 136.150 ;
        RECT 66.565 134.470 66.825 134.790 ;
        RECT 64.550 133.595 66.090 133.965 ;
        RECT 66.625 133.430 66.765 134.470 ;
        RECT 66.565 133.110 66.825 133.430 ;
        RECT 63.345 132.430 63.605 132.750 ;
        RECT 63.865 132.690 66.765 132.830 ;
        RECT 62.025 129.970 62.625 130.110 ;
        RECT 62.025 107.930 62.165 129.970 ;
        RECT 63.405 129.690 63.545 132.430 ;
        RECT 63.805 132.090 64.065 132.410 ;
        RECT 63.345 129.370 63.605 129.690 ;
        RECT 62.425 125.970 62.685 126.290 ;
        RECT 62.485 124.250 62.625 125.970 ;
        RECT 62.425 123.930 62.685 124.250 ;
        RECT 63.405 121.870 63.545 129.370 ;
        RECT 63.865 121.870 64.005 132.090 ;
        RECT 64.550 128.155 66.090 128.525 ;
        RECT 66.625 124.670 66.765 132.690 ;
        RECT 67.545 126.290 67.685 147.650 ;
        RECT 68.005 147.030 68.145 150.450 ;
        RECT 68.465 148.585 68.605 150.450 ;
        RECT 68.395 148.215 68.675 148.585 ;
        RECT 67.945 146.710 68.205 147.030 ;
        RECT 68.005 146.545 68.145 146.710 ;
        RECT 67.935 146.175 68.215 146.545 ;
        RECT 68.925 146.010 69.065 164.050 ;
        RECT 69.325 162.350 69.585 162.670 ;
        RECT 68.865 145.690 69.125 146.010 ;
        RECT 68.865 145.010 69.125 145.330 ;
        RECT 68.925 143.630 69.065 145.010 ;
        RECT 68.865 143.310 69.125 143.630 ;
        RECT 68.405 140.250 68.665 140.570 ;
        RECT 68.465 138.870 68.605 140.250 ;
        RECT 68.405 138.550 68.665 138.870 ;
        RECT 68.865 137.190 69.125 137.510 ;
        RECT 68.405 134.810 68.665 135.130 ;
        RECT 68.465 133.430 68.605 134.810 ;
        RECT 68.405 133.110 68.665 133.430 ;
        RECT 68.925 126.970 69.065 137.190 ;
        RECT 69.385 132.750 69.525 162.350 ;
        RECT 69.845 162.330 69.985 164.730 ;
        RECT 70.305 163.350 70.445 164.730 ;
        RECT 70.245 163.030 70.505 163.350 ;
        RECT 69.785 162.010 70.045 162.330 ;
        RECT 69.845 159.950 69.985 162.010 ;
        RECT 69.785 159.630 70.045 159.950 ;
        RECT 69.845 156.890 69.985 159.630 ;
        RECT 69.785 156.570 70.045 156.890 ;
        RECT 69.785 155.890 70.045 156.210 ;
        RECT 69.325 132.430 69.585 132.750 ;
        RECT 69.325 129.370 69.585 129.690 ;
        RECT 69.385 127.310 69.525 129.370 ;
        RECT 69.845 127.310 69.985 155.890 ;
        RECT 70.245 153.170 70.505 153.490 ;
        RECT 70.305 151.110 70.445 153.170 ;
        RECT 70.245 150.790 70.505 151.110 ;
        RECT 70.305 149.070 70.445 150.790 ;
        RECT 70.765 149.070 70.905 182.470 ;
        RECT 73.925 181.050 74.185 181.370 ;
        RECT 72.545 178.330 72.805 178.650 ;
        RECT 71.165 177.650 71.425 177.970 ;
        RECT 71.225 176.610 71.365 177.650 ;
        RECT 71.165 176.290 71.425 176.610 ;
        RECT 72.605 173.210 72.745 178.330 ;
        RECT 72.545 172.890 72.805 173.210 ;
        RECT 72.085 170.510 72.345 170.830 ;
        RECT 72.145 166.070 72.285 170.510 ;
        RECT 71.625 165.750 71.885 166.070 ;
        RECT 72.085 165.750 72.345 166.070 ;
        RECT 71.685 164.710 71.825 165.750 ;
        RECT 71.625 164.390 71.885 164.710 ;
        RECT 72.605 162.750 72.745 172.890 ;
        RECT 73.985 172.870 74.125 181.050 ;
        RECT 74.445 178.650 74.585 183.770 ;
        RECT 75.365 183.410 75.505 185.810 ;
        RECT 75.825 184.430 75.965 185.810 ;
        RECT 76.335 185.275 77.875 185.645 ;
        RECT 75.765 184.110 76.025 184.430 ;
        RECT 75.305 183.090 75.565 183.410 ;
        RECT 74.845 181.390 75.105 181.710 ;
        RECT 74.385 178.330 74.645 178.650 ;
        RECT 74.445 173.550 74.585 178.330 ;
        RECT 74.905 177.970 75.045 181.390 ;
        RECT 75.825 181.370 75.965 184.110 ;
        RECT 77.605 183.090 77.865 183.410 ;
        RECT 77.665 181.710 77.805 183.090 ;
        RECT 77.605 181.390 77.865 181.710 ;
        RECT 75.765 181.050 76.025 181.370 ;
        RECT 76.335 179.835 77.875 180.205 ;
        RECT 74.845 177.650 75.105 177.970 ;
        RECT 74.385 173.230 74.645 173.550 ;
        RECT 73.925 172.550 74.185 172.870 ;
        RECT 73.985 171.510 74.125 172.550 ;
        RECT 73.925 171.190 74.185 171.510 ;
        RECT 74.385 165.410 74.645 165.730 ;
        RECT 73.925 165.070 74.185 165.390 ;
        RECT 72.145 162.610 72.745 162.750 ;
        RECT 73.005 162.690 73.265 163.010 ;
        RECT 71.625 161.670 71.885 161.990 ;
        RECT 71.685 159.950 71.825 161.670 ;
        RECT 71.625 159.630 71.885 159.950 ;
        RECT 71.165 158.610 71.425 158.930 ;
        RECT 71.225 149.150 71.365 158.610 ;
        RECT 71.685 156.890 71.825 159.630 ;
        RECT 72.145 157.910 72.285 162.610 ;
        RECT 73.065 159.950 73.205 162.690 ;
        RECT 73.985 162.185 74.125 165.070 ;
        RECT 74.445 162.670 74.585 165.410 ;
        RECT 74.385 162.350 74.645 162.670 ;
        RECT 73.915 161.815 74.195 162.185 ;
        RECT 73.005 159.630 73.265 159.950 ;
        RECT 72.085 157.590 72.345 157.910 ;
        RECT 73.065 156.890 73.205 159.630 ;
        RECT 74.445 159.610 74.585 162.350 ;
        RECT 74.385 159.290 74.645 159.610 ;
        RECT 74.445 157.910 74.585 159.290 ;
        RECT 74.385 157.590 74.645 157.910 ;
        RECT 71.625 156.570 71.885 156.890 ;
        RECT 73.005 156.570 73.265 156.890 ;
        RECT 74.385 151.810 74.645 152.130 ;
        RECT 74.445 151.450 74.585 151.810 ;
        RECT 74.905 151.450 75.045 177.650 ;
        RECT 76.335 174.395 77.875 174.765 ;
        RECT 76.335 168.955 77.875 169.325 ;
        RECT 76.335 163.515 77.875 163.885 ;
        RECT 77.145 161.670 77.405 161.990 ;
        RECT 75.305 161.330 75.565 161.650 ;
        RECT 75.765 161.330 76.025 161.650 ;
        RECT 75.365 159.950 75.505 161.330 ;
        RECT 75.305 159.630 75.565 159.950 ;
        RECT 75.825 157.230 75.965 161.330 ;
        RECT 77.205 159.950 77.345 161.670 ;
        RECT 77.145 159.630 77.405 159.950 ;
        RECT 78.065 158.610 78.325 158.930 ;
        RECT 76.335 158.075 77.875 158.445 ;
        RECT 78.125 157.230 78.265 158.610 ;
        RECT 75.765 156.910 76.025 157.230 ;
        RECT 78.065 156.910 78.325 157.230 ;
        RECT 78.065 156.230 78.325 156.550 ;
        RECT 78.125 154.850 78.265 156.230 ;
        RECT 78.065 154.530 78.325 154.850 ;
        RECT 75.305 154.190 75.565 154.510 ;
        RECT 75.365 154.025 75.505 154.190 ;
        RECT 75.295 153.655 75.575 154.025 ;
        RECT 76.335 152.635 77.875 153.005 ;
        RECT 72.085 151.130 72.345 151.450 ;
        RECT 74.385 151.130 74.645 151.450 ;
        RECT 74.845 151.130 75.105 151.450 ;
        RECT 70.245 148.750 70.505 149.070 ;
        RECT 70.705 148.750 70.965 149.070 ;
        RECT 71.225 149.010 71.825 149.150 ;
        RECT 72.145 149.070 72.285 151.130 ;
        RECT 72.545 150.450 72.805 150.770 ;
        RECT 73.005 150.450 73.265 150.770 ;
        RECT 70.705 146.710 70.965 147.030 ;
        RECT 70.245 145.185 70.505 145.330 ;
        RECT 70.235 144.815 70.515 145.185 ;
        RECT 70.245 136.850 70.505 137.170 ;
        RECT 69.325 126.990 69.585 127.310 ;
        RECT 69.785 126.990 70.045 127.310 ;
        RECT 68.865 126.650 69.125 126.970 ;
        RECT 67.945 126.310 68.205 126.630 ;
        RECT 67.485 125.970 67.745 126.290 ;
        RECT 66.625 124.530 67.225 124.670 ;
        RECT 67.085 124.250 67.225 124.530 ;
        RECT 67.025 123.930 67.285 124.250 ;
        RECT 64.550 122.715 66.090 123.085 ;
        RECT 63.345 121.550 63.605 121.870 ;
        RECT 63.805 121.550 64.065 121.870 ;
        RECT 63.865 120.850 64.005 121.550 ;
        RECT 63.805 120.530 64.065 120.850 ;
        RECT 63.865 119.150 64.005 120.530 ;
        RECT 63.805 118.830 64.065 119.150 ;
        RECT 63.865 116.430 64.005 118.830 ;
        RECT 66.565 118.150 66.825 118.470 ;
        RECT 64.550 117.275 66.090 117.645 ;
        RECT 66.625 117.110 66.765 118.150 ;
        RECT 66.565 116.790 66.825 117.110 ;
        RECT 67.085 116.430 67.225 123.930 ;
        RECT 67.485 123.250 67.745 123.570 ;
        RECT 63.805 116.110 64.065 116.430 ;
        RECT 67.025 116.110 67.285 116.430 ;
        RECT 67.085 113.030 67.225 116.110 ;
        RECT 67.545 116.090 67.685 123.250 ;
        RECT 68.005 119.830 68.145 126.310 ;
        RECT 68.865 125.970 69.125 126.290 ;
        RECT 68.405 123.250 68.665 123.570 ;
        RECT 68.465 122.210 68.605 123.250 ;
        RECT 68.405 121.890 68.665 122.210 ;
        RECT 67.945 119.510 68.205 119.830 ;
        RECT 68.005 117.110 68.145 119.510 ;
        RECT 67.945 116.790 68.205 117.110 ;
        RECT 67.485 115.770 67.745 116.090 ;
        RECT 68.925 114.390 69.065 125.970 ;
        RECT 69.385 124.930 69.525 126.990 ;
        RECT 69.325 124.610 69.585 124.930 ;
        RECT 68.865 114.070 69.125 114.390 ;
        RECT 67.025 112.710 67.285 113.030 ;
        RECT 64.550 111.835 66.090 112.205 ;
        RECT 70.305 110.990 70.445 136.850 ;
        RECT 70.765 130.710 70.905 146.710 ;
        RECT 71.165 142.970 71.425 143.290 ;
        RECT 71.225 140.570 71.365 142.970 ;
        RECT 71.165 140.250 71.425 140.570 ;
        RECT 71.225 135.130 71.365 140.250 ;
        RECT 71.685 138.190 71.825 149.010 ;
        RECT 72.085 148.750 72.345 149.070 ;
        RECT 72.085 148.070 72.345 148.390 ;
        RECT 72.145 146.350 72.285 148.070 ;
        RECT 72.085 146.030 72.345 146.350 ;
        RECT 72.605 145.580 72.745 150.450 ;
        RECT 72.145 145.440 72.745 145.580 ;
        RECT 72.145 144.390 72.285 145.440 ;
        RECT 72.145 144.250 72.745 144.390 ;
        RECT 72.085 140.250 72.345 140.570 ;
        RECT 71.625 137.870 71.885 138.190 ;
        RECT 71.165 134.810 71.425 135.130 ;
        RECT 70.705 130.390 70.965 130.710 ;
        RECT 71.225 130.030 71.365 134.810 ;
        RECT 71.165 129.710 71.425 130.030 ;
        RECT 71.225 127.990 71.365 129.710 ;
        RECT 71.165 127.670 71.425 127.990 ;
        RECT 70.705 123.930 70.965 124.250 ;
        RECT 70.765 120.850 70.905 123.930 ;
        RECT 70.705 120.530 70.965 120.850 ;
        RECT 70.765 118.130 70.905 120.530 ;
        RECT 71.225 119.150 71.365 127.670 ;
        RECT 72.145 127.310 72.285 140.250 ;
        RECT 72.605 132.410 72.745 144.250 ;
        RECT 73.065 140.570 73.205 150.450 ;
        RECT 74.445 149.750 74.585 151.130 ;
        RECT 77.145 150.790 77.405 151.110 ;
        RECT 74.385 149.430 74.645 149.750 ;
        RECT 77.205 149.070 77.345 150.790 ;
        RECT 78.585 149.410 78.725 187.510 ;
        RECT 81.285 186.830 81.545 187.150 ;
        RECT 81.345 185.110 81.485 186.830 ;
        RECT 81.805 185.110 81.945 189.210 ;
        RECT 81.285 184.790 81.545 185.110 ;
        RECT 81.745 184.790 82.005 185.110 ;
        RECT 82.725 184.090 82.865 191.250 ;
        RECT 83.585 189.550 83.845 189.870 ;
        RECT 83.645 186.810 83.785 189.550 ;
        RECT 87.785 187.830 87.925 192.270 ;
        RECT 88.645 191.250 88.905 191.570 ;
        RECT 88.705 189.870 88.845 191.250 ;
        RECT 88.645 189.550 88.905 189.870 ;
        RECT 94.685 189.530 94.825 192.270 ;
        RECT 97.845 191.250 98.105 191.570 ;
        RECT 97.905 189.530 98.045 191.250 ;
        RECT 94.625 189.270 94.885 189.530 ;
        RECT 94.225 189.210 94.885 189.270 ;
        RECT 95.545 189.210 95.805 189.530 ;
        RECT 96.005 189.210 96.265 189.530 ;
        RECT 97.845 189.210 98.105 189.530 ;
        RECT 94.225 189.130 94.825 189.210 ;
        RECT 93.245 188.760 93.505 188.850 ;
        RECT 94.225 188.760 94.365 189.130 ;
        RECT 95.085 188.760 95.345 188.850 ;
        RECT 93.245 188.620 94.365 188.760 ;
        RECT 94.685 188.620 95.345 188.760 ;
        RECT 93.245 188.530 93.505 188.620 ;
        RECT 88.125 187.995 89.665 188.365 ;
        RECT 87.725 187.510 87.985 187.830 ;
        RECT 94.685 187.150 94.825 188.620 ;
        RECT 95.085 188.530 95.345 188.620 ;
        RECT 95.605 187.490 95.745 189.210 ;
        RECT 95.545 187.170 95.805 187.490 ;
        RECT 90.025 186.830 90.285 187.150 ;
        RECT 93.245 186.830 93.505 187.150 ;
        RECT 94.625 186.830 94.885 187.150 ;
        RECT 83.585 186.490 83.845 186.810 ;
        RECT 82.665 183.770 82.925 184.090 ;
        RECT 81.745 181.390 82.005 181.710 ;
        RECT 79.905 180.370 80.165 180.690 ;
        RECT 79.965 176.270 80.105 180.370 ;
        RECT 81.285 177.990 81.545 178.310 ;
        RECT 81.345 176.950 81.485 177.990 ;
        RECT 81.285 176.630 81.545 176.950 ;
        RECT 79.905 175.950 80.165 176.270 ;
        RECT 81.805 175.250 81.945 181.390 ;
        RECT 82.665 178.560 82.925 178.650 ;
        RECT 83.645 178.560 83.785 186.490 ;
        RECT 85.885 183.090 86.145 183.410 ;
        RECT 82.665 178.420 83.785 178.560 ;
        RECT 82.665 178.330 82.925 178.420 ;
        RECT 82.725 175.590 82.865 178.330 ;
        RECT 85.945 178.310 86.085 183.090 ;
        RECT 88.125 182.555 89.665 182.925 ;
        RECT 90.085 178.990 90.225 186.830 ;
        RECT 90.485 185.810 90.745 186.130 ;
        RECT 90.545 183.750 90.685 185.810 ;
        RECT 90.485 183.430 90.745 183.750 ;
        RECT 92.325 183.090 92.585 183.410 ;
        RECT 92.385 180.690 92.525 183.090 ;
        RECT 92.325 180.370 92.585 180.690 ;
        RECT 90.025 178.670 90.285 178.990 ;
        RECT 87.265 178.330 87.525 178.650 ;
        RECT 90.085 178.390 90.225 178.670 ;
        RECT 85.885 177.990 86.145 178.310 ;
        RECT 85.425 177.650 85.685 177.970 ;
        RECT 85.485 176.610 85.625 177.650 ;
        RECT 85.425 176.290 85.685 176.610 ;
        RECT 82.665 175.270 82.925 175.590 ;
        RECT 81.745 174.930 82.005 175.250 ;
        RECT 81.285 172.210 81.545 172.530 ;
        RECT 81.345 170.150 81.485 172.210 ;
        RECT 81.805 170.830 81.945 174.930 ;
        RECT 82.725 172.530 82.865 175.270 ;
        RECT 82.665 172.210 82.925 172.530 ;
        RECT 81.745 170.510 82.005 170.830 ;
        RECT 81.285 169.830 81.545 170.150 ;
        RECT 81.345 168.450 81.485 169.830 ;
        RECT 81.285 168.130 81.545 168.450 ;
        RECT 80.825 167.790 81.085 168.110 ;
        RECT 80.365 164.050 80.625 164.370 ;
        RECT 80.425 163.350 80.565 164.050 ;
        RECT 80.365 163.030 80.625 163.350 ;
        RECT 78.985 162.010 79.245 162.330 ;
        RECT 79.045 159.610 79.185 162.010 ;
        RECT 80.425 161.650 80.565 163.030 ;
        RECT 80.885 162.865 81.025 167.790 ;
        RECT 80.815 162.495 81.095 162.865 ;
        RECT 80.825 162.350 81.085 162.495 ;
        RECT 80.365 161.330 80.625 161.650 ;
        RECT 78.985 159.290 79.245 159.610 ;
        RECT 79.045 154.510 79.185 159.290 ;
        RECT 78.985 154.420 79.245 154.510 ;
        RECT 78.985 154.280 80.105 154.420 ;
        RECT 78.985 154.190 79.245 154.280 ;
        RECT 79.965 151.450 80.105 154.280 ;
        RECT 81.805 151.790 81.945 170.510 ;
        RECT 82.725 170.490 82.865 172.210 ;
        RECT 84.045 171.190 84.305 171.510 ;
        RECT 84.105 170.490 84.245 171.190 ;
        RECT 85.425 170.740 85.685 170.830 ;
        RECT 85.945 170.740 86.085 177.990 ;
        RECT 86.805 172.210 87.065 172.530 ;
        RECT 86.865 171.170 87.005 172.210 ;
        RECT 87.325 171.510 87.465 178.330 ;
        RECT 90.085 178.250 90.685 178.390 ;
        RECT 87.725 177.650 87.985 177.970 ;
        RECT 90.025 177.650 90.285 177.970 ;
        RECT 87.785 176.860 87.925 177.650 ;
        RECT 88.125 177.115 89.665 177.485 ;
        RECT 90.085 176.950 90.225 177.650 ;
        RECT 87.785 176.720 88.385 176.860 ;
        RECT 87.725 172.890 87.985 173.210 ;
        RECT 87.265 171.190 87.525 171.510 ;
        RECT 86.805 170.850 87.065 171.170 ;
        RECT 85.425 170.600 86.085 170.740 ;
        RECT 85.425 170.510 85.685 170.600 ;
        RECT 82.665 170.170 82.925 170.490 ;
        RECT 84.045 170.170 84.305 170.490 ;
        RECT 82.205 169.490 82.465 169.810 ;
        RECT 82.265 167.090 82.405 169.490 ;
        RECT 82.725 167.430 82.865 170.170 ;
        RECT 82.665 167.110 82.925 167.430 ;
        RECT 82.205 166.770 82.465 167.090 ;
        RECT 82.265 165.050 82.405 166.770 ;
        RECT 82.725 165.050 82.865 167.110 ;
        RECT 82.205 164.730 82.465 165.050 ;
        RECT 82.665 164.730 82.925 165.050 ;
        RECT 82.725 159.610 82.865 164.730 ;
        RECT 84.045 161.330 84.305 161.650 ;
        RECT 84.105 159.950 84.245 161.330 ;
        RECT 84.045 159.630 84.305 159.950 ;
        RECT 82.665 159.290 82.925 159.610 ;
        RECT 82.725 156.890 82.865 159.290 ;
        RECT 82.665 156.570 82.925 156.890 ;
        RECT 82.725 154.170 82.865 156.570 ;
        RECT 84.505 155.890 84.765 156.210 ;
        RECT 84.965 155.890 85.225 156.210 ;
        RECT 84.565 154.170 84.705 155.890 ;
        RECT 82.665 153.850 82.925 154.170 ;
        RECT 84.505 153.850 84.765 154.170 ;
        RECT 82.665 153.170 82.925 153.490 ;
        RECT 82.725 151.790 82.865 153.170 ;
        RECT 81.745 151.470 82.005 151.790 ;
        RECT 82.665 151.470 82.925 151.790 ;
        RECT 79.905 151.130 80.165 151.450 ;
        RECT 81.745 150.790 82.005 151.110 ;
        RECT 81.285 150.450 81.545 150.770 ;
        RECT 81.345 149.410 81.485 150.450 ;
        RECT 78.525 149.090 78.785 149.410 ;
        RECT 81.285 149.090 81.545 149.410 ;
        RECT 73.925 148.750 74.185 149.070 ;
        RECT 77.145 148.750 77.405 149.070 ;
        RECT 73.465 148.410 73.725 148.730 ;
        RECT 73.005 140.250 73.265 140.570 ;
        RECT 73.005 139.570 73.265 139.890 ;
        RECT 73.065 138.530 73.205 139.570 ;
        RECT 73.005 138.210 73.265 138.530 ;
        RECT 73.525 137.850 73.665 148.410 ;
        RECT 73.985 145.670 74.125 148.750 ;
        RECT 74.845 147.730 75.105 148.050 ;
        RECT 74.905 146.010 75.045 147.730 ;
        RECT 76.335 147.195 77.875 147.565 ;
        RECT 81.805 147.030 81.945 150.790 ;
        RECT 81.745 146.710 82.005 147.030 ;
        RECT 74.385 145.690 74.645 146.010 ;
        RECT 74.845 145.690 75.105 146.010 ;
        RECT 73.925 145.350 74.185 145.670 ;
        RECT 74.445 140.570 74.585 145.690 ;
        RECT 74.905 140.570 75.045 145.690 ;
        RECT 75.765 145.350 76.025 145.670 ;
        RECT 75.825 140.570 75.965 145.350 ;
        RECT 81.805 144.310 81.945 146.710 ;
        RECT 81.745 143.990 82.005 144.310 ;
        RECT 79.905 143.310 80.165 143.630 ;
        RECT 76.335 141.755 77.875 142.125 ;
        RECT 79.965 141.250 80.105 143.310 ;
        RECT 82.725 143.290 82.865 151.470 ;
        RECT 83.585 150.450 83.845 150.770 ;
        RECT 83.645 149.265 83.785 150.450 ;
        RECT 83.575 148.895 83.855 149.265 ;
        RECT 83.645 148.730 83.785 148.895 ;
        RECT 83.585 148.410 83.845 148.730 ;
        RECT 84.045 145.690 84.305 146.010 ;
        RECT 84.105 144.310 84.245 145.690 ;
        RECT 84.045 143.990 84.305 144.310 ;
        RECT 82.665 142.970 82.925 143.290 ;
        RECT 82.725 141.590 82.865 142.970 ;
        RECT 82.665 141.270 82.925 141.590 ;
        RECT 79.905 140.930 80.165 141.250 ;
        RECT 74.385 140.250 74.645 140.570 ;
        RECT 74.845 140.250 75.105 140.570 ;
        RECT 75.765 140.250 76.025 140.570 ;
        RECT 73.465 137.530 73.725 137.850 ;
        RECT 74.445 135.470 74.585 140.250 ;
        RECT 74.385 135.150 74.645 135.470 ;
        RECT 73.005 134.130 73.265 134.450 ;
        RECT 73.065 133.090 73.205 134.130 ;
        RECT 73.005 132.770 73.265 133.090 ;
        RECT 74.445 132.750 74.585 135.150 ;
        RECT 74.905 134.790 75.045 140.250 ;
        RECT 75.825 135.810 75.965 140.250 ;
        RECT 79.965 138.870 80.105 140.930 ;
        RECT 79.905 138.550 80.165 138.870 ;
        RECT 80.365 137.870 80.625 138.190 ;
        RECT 76.335 136.315 77.875 136.685 ;
        RECT 75.765 135.490 76.025 135.810 ;
        RECT 77.145 134.810 77.405 135.130 ;
        RECT 74.845 134.470 75.105 134.790 ;
        RECT 74.905 133.090 75.045 134.470 ;
        RECT 74.845 132.770 75.105 133.090 ;
        RECT 77.205 132.750 77.345 134.810 ;
        RECT 80.425 134.790 80.565 137.870 ;
        RECT 82.205 137.760 82.465 137.850 ;
        RECT 82.725 137.760 82.865 141.270 ;
        RECT 84.045 140.250 84.305 140.570 ;
        RECT 84.105 138.870 84.245 140.250 ;
        RECT 84.045 138.550 84.305 138.870 ;
        RECT 85.025 138.190 85.165 155.890 ;
        RECT 85.485 154.850 85.625 170.510 ;
        RECT 87.265 169.490 87.525 169.810 ;
        RECT 87.325 167.770 87.465 169.490 ;
        RECT 86.805 167.625 87.065 167.770 ;
        RECT 86.795 167.255 87.075 167.625 ;
        RECT 87.265 167.450 87.525 167.770 ;
        RECT 87.265 166.770 87.525 167.090 ;
        RECT 85.885 165.410 86.145 165.730 ;
        RECT 85.945 163.350 86.085 165.410 ;
        RECT 87.325 164.370 87.465 166.770 ;
        RECT 87.265 164.050 87.525 164.370 ;
        RECT 87.785 163.350 87.925 172.890 ;
        RECT 88.245 172.870 88.385 176.720 ;
        RECT 90.025 176.630 90.285 176.950 ;
        RECT 90.545 176.610 90.685 178.250 ;
        RECT 92.385 177.970 92.525 180.370 ;
        RECT 93.305 179.670 93.445 186.830 ;
        RECT 93.705 186.490 93.965 186.810 ;
        RECT 93.765 185.110 93.905 186.490 ;
        RECT 94.165 185.810 94.425 186.130 ;
        RECT 93.705 184.790 93.965 185.110 ;
        RECT 93.245 179.350 93.505 179.670 ;
        RECT 93.765 179.330 93.905 184.790 ;
        RECT 94.225 184.430 94.365 185.810 ;
        RECT 94.165 184.110 94.425 184.430 ;
        RECT 94.685 183.830 94.825 186.830 ;
        RECT 94.225 183.690 94.825 183.830 ;
        RECT 93.705 179.010 93.965 179.330 ;
        RECT 92.325 177.650 92.585 177.970 ;
        RECT 93.705 177.650 93.965 177.970 ;
        RECT 90.485 176.290 90.745 176.610 ;
        RECT 90.485 175.610 90.745 175.930 ;
        RECT 88.185 172.550 88.445 172.870 ;
        RECT 88.125 171.675 89.665 172.045 ;
        RECT 89.565 170.510 89.825 170.830 ;
        RECT 89.625 168.790 89.765 170.510 ;
        RECT 90.025 170.170 90.285 170.490 ;
        RECT 89.565 168.470 89.825 168.790 ;
        RECT 89.105 168.130 89.365 168.450 ;
        RECT 89.165 167.340 89.305 168.130 ;
        RECT 89.565 167.340 89.825 167.430 ;
        RECT 89.165 167.200 89.825 167.340 ;
        RECT 89.565 167.110 89.825 167.200 ;
        RECT 88.125 166.235 89.665 166.605 ;
        RECT 88.185 164.050 88.445 164.370 ;
        RECT 85.885 163.030 86.145 163.350 ;
        RECT 87.725 163.030 87.985 163.350 ;
        RECT 87.255 162.495 87.535 162.865 ;
        RECT 87.265 162.350 87.525 162.495 ;
        RECT 87.785 162.330 87.925 163.030 ;
        RECT 87.725 162.010 87.985 162.330 ;
        RECT 88.245 161.560 88.385 164.050 ;
        RECT 90.085 162.330 90.225 170.170 ;
        RECT 90.025 162.010 90.285 162.330 ;
        RECT 87.785 161.420 88.385 161.560 ;
        RECT 87.785 159.350 87.925 161.420 ;
        RECT 90.025 161.330 90.285 161.650 ;
        RECT 88.125 160.795 89.665 161.165 ;
        RECT 90.085 160.630 90.225 161.330 ;
        RECT 90.025 160.310 90.285 160.630 ;
        RECT 86.345 158.950 86.605 159.270 ;
        RECT 87.785 159.210 88.385 159.350 ;
        RECT 86.405 157.910 86.545 158.950 ;
        RECT 87.725 158.610 87.985 158.930 ;
        RECT 86.345 157.590 86.605 157.910 ;
        RECT 87.785 157.140 87.925 158.610 ;
        RECT 88.245 157.230 88.385 159.210 ;
        RECT 90.025 158.840 90.285 158.930 ;
        RECT 90.545 158.840 90.685 175.610 ;
        RECT 91.405 169.830 91.665 170.150 ;
        RECT 91.465 167.770 91.605 169.830 ;
        RECT 90.945 167.625 91.205 167.770 ;
        RECT 90.935 167.255 91.215 167.625 ;
        RECT 91.405 167.450 91.665 167.770 ;
        RECT 92.325 167.510 92.585 167.770 ;
        RECT 92.785 167.625 93.045 167.770 ;
        RECT 91.925 167.450 92.585 167.510 ;
        RECT 91.925 167.370 92.525 167.450 ;
        RECT 91.925 167.000 92.065 167.370 ;
        RECT 92.775 167.255 93.055 167.625 ;
        RECT 91.465 166.860 92.065 167.000 ;
        RECT 91.465 165.390 91.605 166.860 ;
        RECT 92.325 166.770 92.585 167.090 ;
        RECT 92.785 166.770 93.045 167.090 ;
        RECT 90.945 165.070 91.205 165.390 ;
        RECT 91.405 165.070 91.665 165.390 ;
        RECT 91.005 163.350 91.145 165.070 ;
        RECT 91.465 164.370 91.605 165.070 ;
        RECT 91.405 164.050 91.665 164.370 ;
        RECT 91.865 164.050 92.125 164.370 ;
        RECT 90.945 163.030 91.205 163.350 ;
        RECT 90.945 161.670 91.205 161.990 ;
        RECT 90.025 158.700 90.685 158.840 ;
        RECT 90.025 158.610 90.285 158.700 ;
        RECT 87.325 157.000 87.925 157.140 ;
        RECT 87.325 155.190 87.465 157.000 ;
        RECT 88.185 156.910 88.445 157.230 ;
        RECT 90.085 156.890 90.225 158.610 ;
        RECT 91.005 156.890 91.145 161.670 ;
        RECT 91.405 160.310 91.665 160.630 ;
        RECT 91.465 156.890 91.605 160.310 ;
        RECT 90.025 156.570 90.285 156.890 ;
        RECT 90.945 156.570 91.205 156.890 ;
        RECT 91.405 156.570 91.665 156.890 ;
        RECT 88.125 155.355 89.665 155.725 ;
        RECT 87.265 154.870 87.525 155.190 ;
        RECT 85.425 154.530 85.685 154.850 ;
        RECT 87.325 154.510 87.465 154.870 ;
        RECT 87.265 154.190 87.525 154.510 ;
        RECT 87.725 150.450 87.985 150.770 ;
        RECT 87.785 149.750 87.925 150.450 ;
        RECT 88.125 149.915 89.665 150.285 ;
        RECT 87.725 149.430 87.985 149.750 ;
        RECT 90.085 149.410 90.225 156.570 ;
        RECT 91.405 155.890 91.665 156.210 ;
        RECT 90.485 153.510 90.745 153.830 ;
        RECT 90.025 149.090 90.285 149.410 ;
        RECT 87.255 148.215 87.535 148.585 ;
        RECT 86.805 147.730 87.065 148.050 ;
        RECT 87.325 147.905 87.465 148.215 ;
        RECT 86.865 146.545 87.005 147.730 ;
        RECT 87.255 147.535 87.535 147.905 ;
        RECT 86.795 146.175 87.075 146.545 ;
        RECT 85.885 145.690 86.145 146.010 ;
        RECT 85.945 140.910 86.085 145.690 ;
        RECT 85.885 140.590 86.145 140.910 ;
        RECT 86.865 138.190 87.005 146.175 ;
        RECT 90.545 146.010 90.685 153.510 ;
        RECT 90.945 153.170 91.205 153.490 ;
        RECT 87.725 145.690 87.985 146.010 ;
        RECT 90.485 145.690 90.745 146.010 ;
        RECT 87.785 140.570 87.925 145.690 ;
        RECT 88.125 144.475 89.665 144.845 ;
        RECT 90.025 141.270 90.285 141.590 ;
        RECT 87.725 140.250 87.985 140.570 ;
        RECT 88.125 139.035 89.665 139.405 ;
        RECT 90.085 138.870 90.225 141.270 ;
        RECT 90.485 139.570 90.745 139.890 ;
        RECT 90.025 138.550 90.285 138.870 ;
        RECT 84.965 137.870 85.225 138.190 ;
        RECT 86.805 137.870 87.065 138.190 ;
        RECT 87.725 137.870 87.985 138.190 ;
        RECT 88.175 138.015 88.455 138.385 ;
        RECT 88.185 137.870 88.445 138.015 ;
        RECT 82.205 137.620 82.865 137.760 ;
        RECT 82.205 137.530 82.465 137.620 ;
        RECT 82.725 135.470 82.865 137.620 ;
        RECT 87.785 137.510 87.925 137.870 ;
        RECT 87.725 137.190 87.985 137.510 ;
        RECT 84.045 136.850 84.305 137.170 ;
        RECT 87.265 136.850 87.525 137.170 ;
        RECT 82.665 135.150 82.925 135.470 ;
        RECT 77.605 134.470 77.865 134.790 ;
        RECT 80.365 134.470 80.625 134.790 ;
        RECT 77.665 133.430 77.805 134.470 ;
        RECT 81.285 134.130 81.545 134.450 ;
        RECT 81.345 133.430 81.485 134.130 ;
        RECT 77.605 133.110 77.865 133.430 ;
        RECT 81.285 133.110 81.545 133.430 ;
        RECT 82.205 132.770 82.465 133.090 ;
        RECT 74.385 132.430 74.645 132.750 ;
        RECT 77.145 132.430 77.405 132.750 ;
        RECT 72.545 132.090 72.805 132.410 ;
        RECT 73.925 132.090 74.185 132.410 ;
        RECT 73.005 131.410 73.265 131.730 ;
        RECT 73.465 131.410 73.725 131.730 ;
        RECT 72.085 126.990 72.345 127.310 ;
        RECT 72.545 126.990 72.805 127.310 ;
        RECT 71.625 125.970 71.885 126.290 ;
        RECT 72.085 125.970 72.345 126.290 ;
        RECT 71.685 121.190 71.825 125.970 ;
        RECT 72.145 125.270 72.285 125.970 ;
        RECT 72.085 124.950 72.345 125.270 ;
        RECT 72.605 123.570 72.745 126.990 ;
        RECT 73.065 125.270 73.205 131.410 ;
        RECT 73.525 127.650 73.665 131.410 ;
        RECT 73.985 130.370 74.125 132.090 ;
        RECT 74.385 131.750 74.645 132.070 ;
        RECT 73.925 130.050 74.185 130.370 ;
        RECT 73.465 127.330 73.725 127.650 ;
        RECT 73.005 124.950 73.265 125.270 ;
        RECT 73.465 123.590 73.725 123.910 ;
        RECT 72.545 123.250 72.805 123.570 ;
        RECT 73.005 121.550 73.265 121.870 ;
        RECT 71.625 120.870 71.885 121.190 ;
        RECT 73.065 119.830 73.205 121.550 ;
        RECT 73.005 119.510 73.265 119.830 ;
        RECT 73.525 119.150 73.665 123.590 ;
        RECT 71.165 118.830 71.425 119.150 ;
        RECT 73.465 118.830 73.725 119.150 ;
        RECT 72.085 118.490 72.345 118.810 ;
        RECT 70.705 117.810 70.965 118.130 ;
        RECT 70.765 116.770 70.905 117.810 ;
        RECT 72.145 117.110 72.285 118.490 ;
        RECT 73.525 117.110 73.665 118.830 ;
        RECT 72.085 116.790 72.345 117.110 ;
        RECT 73.465 116.790 73.725 117.110 ;
        RECT 70.705 116.450 70.965 116.770 ;
        RECT 74.445 110.990 74.585 131.750 ;
        RECT 76.335 130.875 77.875 131.245 ;
        RECT 82.265 130.710 82.405 132.770 ;
        RECT 83.125 132.090 83.385 132.410 ;
        RECT 82.205 130.390 82.465 130.710 ;
        RECT 79.435 129.855 79.715 130.225 ;
        RECT 79.505 129.690 79.645 129.855 ;
        RECT 79.445 129.370 79.705 129.690 ;
        RECT 74.845 129.030 75.105 129.350 ;
        RECT 74.905 127.390 75.045 129.030 ;
        RECT 75.765 127.670 76.025 127.990 ;
        RECT 75.825 127.390 75.965 127.670 ;
        RECT 74.905 127.250 75.965 127.390 ;
        RECT 83.185 127.310 83.325 132.090 ;
        RECT 74.905 123.570 75.045 127.250 ;
        RECT 83.125 126.990 83.385 127.310 ;
        RECT 75.305 126.880 75.565 126.970 ;
        RECT 75.305 126.740 75.965 126.880 ;
        RECT 75.305 126.650 75.565 126.740 ;
        RECT 74.845 123.250 75.105 123.570 ;
        RECT 74.905 122.210 75.045 123.250 ;
        RECT 74.845 121.890 75.105 122.210 ;
        RECT 75.825 121.530 75.965 126.740 ;
        RECT 78.065 125.970 78.325 126.290 ;
        RECT 79.445 125.970 79.705 126.290 ;
        RECT 76.335 125.435 77.875 125.805 ;
        RECT 78.125 121.870 78.265 125.970 ;
        RECT 79.505 123.910 79.645 125.970 ;
        RECT 83.185 124.590 83.325 126.990 ;
        RECT 83.125 124.270 83.385 124.590 ;
        RECT 81.285 123.930 81.545 124.250 ;
        RECT 79.445 123.590 79.705 123.910 ;
        RECT 81.345 122.550 81.485 123.930 ;
        RECT 81.285 122.230 81.545 122.550 ;
        RECT 78.065 121.550 78.325 121.870 ;
        RECT 75.765 121.210 76.025 121.530 ;
        RECT 75.825 119.150 75.965 121.210 ;
        RECT 81.285 120.530 81.545 120.850 ;
        RECT 76.335 119.995 77.875 120.365 ;
        RECT 75.765 118.830 76.025 119.150 ;
        RECT 75.825 116.090 75.965 118.830 ;
        RECT 79.905 117.810 80.165 118.130 ;
        RECT 80.825 117.810 81.085 118.130 ;
        RECT 78.525 116.450 78.785 116.770 ;
        RECT 75.765 115.770 76.025 116.090 ;
        RECT 76.335 114.555 77.875 114.925 ;
        RECT 78.585 114.390 78.725 116.450 ;
        RECT 78.525 114.070 78.785 114.390 ;
        RECT 79.965 113.370 80.105 117.810 ;
        RECT 80.885 117.110 81.025 117.810 ;
        RECT 80.825 116.790 81.085 117.110 ;
        RECT 80.825 115.770 81.085 116.090 ;
        RECT 80.885 114.390 81.025 115.770 ;
        RECT 80.825 114.070 81.085 114.390 ;
        RECT 77.145 113.050 77.405 113.370 ;
        RECT 79.905 113.050 80.165 113.370 ;
        RECT 77.205 111.330 77.345 113.050 ;
        RECT 77.145 111.010 77.405 111.330 ;
        RECT 81.345 110.990 81.485 120.530 ;
        RECT 83.185 116.090 83.325 124.270 ;
        RECT 83.125 115.770 83.385 116.090 ;
        RECT 70.245 110.670 70.505 110.990 ;
        RECT 74.385 110.670 74.645 110.990 ;
        RECT 81.285 110.670 81.545 110.990 ;
        RECT 84.105 110.650 84.245 136.850 ;
        RECT 84.965 134.130 85.225 134.450 ;
        RECT 85.025 132.750 85.165 134.130 ;
        RECT 84.965 132.430 85.225 132.750 ;
        RECT 86.805 127.390 87.065 127.650 ;
        RECT 86.405 127.330 87.065 127.390 ;
        RECT 86.405 127.250 87.005 127.330 ;
        RECT 85.885 125.970 86.145 126.290 ;
        RECT 85.945 122.550 86.085 125.970 ;
        RECT 86.405 125.270 86.545 127.250 ;
        RECT 86.805 126.650 87.065 126.970 ;
        RECT 86.865 125.270 87.005 126.650 ;
        RECT 87.325 125.270 87.465 136.850 ;
        RECT 90.085 135.470 90.225 138.550 ;
        RECT 90.025 135.150 90.285 135.470 ;
        RECT 88.125 133.595 89.665 133.965 ;
        RECT 89.565 132.770 89.825 133.090 ;
        RECT 89.625 130.710 89.765 132.770 ;
        RECT 89.565 130.390 89.825 130.710 ;
        RECT 87.725 129.370 87.985 129.690 ;
        RECT 86.345 124.950 86.605 125.270 ;
        RECT 86.805 124.950 87.065 125.270 ;
        RECT 87.265 124.950 87.525 125.270 ;
        RECT 87.785 124.930 87.925 129.370 ;
        RECT 88.125 128.155 89.665 128.525 ;
        RECT 87.725 124.610 87.985 124.930 ;
        RECT 87.265 123.930 87.525 124.250 ;
        RECT 86.805 123.590 87.065 123.910 ;
        RECT 85.885 122.230 86.145 122.550 ;
        RECT 86.865 121.780 87.005 123.590 ;
        RECT 87.325 122.550 87.465 123.930 ;
        RECT 88.125 122.715 89.665 123.085 ;
        RECT 87.265 122.230 87.525 122.550 ;
        RECT 87.265 121.780 87.525 121.870 ;
        RECT 86.865 121.640 87.525 121.780 ;
        RECT 87.265 121.550 87.525 121.640 ;
        RECT 87.325 117.110 87.465 121.550 ;
        RECT 90.025 121.210 90.285 121.530 ;
        RECT 87.725 120.530 87.985 120.850 ;
        RECT 87.265 116.790 87.525 117.110 ;
        RECT 86.805 116.450 87.065 116.770 ;
        RECT 85.885 115.770 86.145 116.090 ;
        RECT 62.885 110.330 63.145 110.650 ;
        RECT 66.105 110.330 66.365 110.650 ;
        RECT 67.485 110.330 67.745 110.650 ;
        RECT 72.545 110.330 72.805 110.650 ;
        RECT 84.045 110.330 84.305 110.650 ;
        RECT 61.505 107.610 61.765 107.930 ;
        RECT 61.965 107.610 62.225 107.930 ;
        RECT 60.125 104.890 60.385 105.210 ;
        RECT 58.285 103.190 58.545 103.510 ;
        RECT 59.665 103.190 59.925 103.510 ;
        RECT 57.885 102.770 58.485 102.910 ;
        RECT 60.185 102.830 60.325 104.890 ;
        RECT 55.065 102.170 55.325 102.490 ;
        RECT 58.345 98.340 58.485 102.770 ;
        RECT 60.125 102.510 60.385 102.830 ;
        RECT 62.945 98.340 63.085 110.330 ;
        RECT 66.165 108.950 66.305 110.330 ;
        RECT 67.025 109.880 67.285 109.970 ;
        RECT 66.625 109.740 67.285 109.880 ;
        RECT 66.105 108.630 66.365 108.950 ;
        RECT 63.805 106.930 64.065 107.250 ;
        RECT 63.865 105.890 64.005 106.930 ;
        RECT 64.550 106.395 66.090 106.765 ;
        RECT 63.805 105.570 64.065 105.890 ;
        RECT 66.625 102.830 66.765 109.740 ;
        RECT 67.025 109.650 67.285 109.740 ;
        RECT 67.545 108.950 67.685 110.330 ;
        RECT 67.485 108.630 67.745 108.950 ;
        RECT 67.485 107.950 67.745 108.270 ;
        RECT 66.565 102.510 66.825 102.830 ;
        RECT 64.550 100.955 66.090 101.325 ;
        RECT 67.545 98.340 67.685 107.950 ;
        RECT 70.705 107.270 70.965 107.590 ;
        RECT 70.765 106.230 70.905 107.270 ;
        RECT 70.705 105.910 70.965 106.230 ;
        RECT 72.075 106.055 72.355 106.425 ;
        RECT 72.145 105.550 72.285 106.055 ;
        RECT 72.085 105.230 72.345 105.550 ;
        RECT 72.605 105.210 72.745 110.330 ;
        RECT 78.525 109.650 78.785 109.970 ;
        RECT 84.045 109.650 84.305 109.970 ;
        RECT 76.335 109.115 77.875 109.485 ;
        RECT 73.005 107.270 73.265 107.590 ;
        RECT 73.065 106.230 73.205 107.270 ;
        RECT 78.585 106.230 78.725 109.650 ;
        RECT 84.105 108.270 84.245 109.650 ;
        RECT 85.945 108.950 86.085 115.770 ;
        RECT 86.865 114.390 87.005 116.450 ;
        RECT 86.805 114.070 87.065 114.390 ;
        RECT 87.785 113.370 87.925 120.530 ;
        RECT 90.085 119.830 90.225 121.210 ;
        RECT 90.025 119.510 90.285 119.830 ;
        RECT 88.125 117.275 89.665 117.645 ;
        RECT 89.565 115.770 89.825 116.090 ;
        RECT 89.625 114.390 89.765 115.770 ;
        RECT 89.565 114.070 89.825 114.390 ;
        RECT 87.725 113.050 87.985 113.370 ;
        RECT 88.125 111.835 89.665 112.205 ;
        RECT 86.345 110.670 86.605 110.990 ;
        RECT 86.405 110.310 86.545 110.670 ;
        RECT 86.345 109.990 86.605 110.310 ;
        RECT 85.885 108.630 86.145 108.950 ;
        RECT 85.945 108.270 86.085 108.630 ;
        RECT 81.285 107.950 81.545 108.270 ;
        RECT 84.045 107.950 84.305 108.270 ;
        RECT 85.885 107.950 86.145 108.270 ;
        RECT 79.445 107.270 79.705 107.590 ;
        RECT 73.005 105.910 73.265 106.230 ;
        RECT 78.525 105.910 78.785 106.230 ;
        RECT 78.985 105.570 79.245 105.890 ;
        RECT 72.545 104.890 72.805 105.210 ;
        RECT 75.765 104.890 76.025 105.210 ;
        RECT 69.325 104.210 69.585 104.530 ;
        RECT 69.385 102.150 69.525 104.210 ;
        RECT 72.605 102.490 72.745 104.890 ;
        RECT 75.825 102.910 75.965 104.890 ;
        RECT 76.335 103.675 77.875 104.045 ;
        RECT 79.045 103.510 79.185 105.570 ;
        RECT 79.505 103.510 79.645 107.270 ;
        RECT 78.985 103.190 79.245 103.510 ;
        RECT 79.445 103.190 79.705 103.510 ;
        RECT 75.825 102.770 76.885 102.910 ;
        RECT 72.545 102.170 72.805 102.490 ;
        RECT 69.325 101.830 69.585 102.150 ;
        RECT 72.085 101.830 72.345 102.150 ;
        RECT 72.145 98.340 72.285 101.830 ;
        RECT 76.745 98.340 76.885 102.770 ;
        RECT 81.345 98.340 81.485 107.950 ;
        RECT 85.945 105.550 86.085 107.950 ;
        RECT 85.885 105.230 86.145 105.550 ;
        RECT 85.885 104.550 86.145 104.870 ;
        RECT 85.945 98.340 86.085 104.550 ;
        RECT 86.405 102.490 86.545 109.990 ;
        RECT 86.805 109.650 87.065 109.970 ;
        RECT 86.865 105.890 87.005 109.650 ;
        RECT 90.545 108.950 90.685 139.570 ;
        RECT 91.005 137.850 91.145 153.170 ;
        RECT 91.465 141.250 91.605 155.890 ;
        RECT 91.405 140.930 91.665 141.250 ;
        RECT 91.925 140.570 92.065 164.050 ;
        RECT 92.385 143.630 92.525 166.770 ;
        RECT 92.845 146.010 92.985 166.770 ;
        RECT 93.245 159.970 93.505 160.290 ;
        RECT 93.305 156.890 93.445 159.970 ;
        RECT 93.765 156.890 93.905 177.650 ;
        RECT 93.245 156.570 93.505 156.890 ;
        RECT 93.705 156.570 93.965 156.890 ;
        RECT 93.305 156.210 93.445 156.570 ;
        RECT 93.245 155.890 93.505 156.210 ;
        RECT 93.305 154.850 93.445 155.890 ;
        RECT 93.695 155.695 93.975 156.065 ;
        RECT 93.245 154.530 93.505 154.850 ;
        RECT 93.245 153.910 93.505 154.170 ;
        RECT 93.765 153.910 93.905 155.695 ;
        RECT 93.245 153.850 93.905 153.910 ;
        RECT 93.305 153.770 93.905 153.850 ;
        RECT 93.245 153.170 93.505 153.490 ;
        RECT 93.305 146.350 93.445 153.170 ;
        RECT 93.765 150.770 93.905 153.770 ;
        RECT 94.225 151.790 94.365 183.690 ;
        RECT 95.085 181.730 95.345 182.050 ;
        RECT 95.145 179.670 95.285 181.730 ;
        RECT 95.085 179.350 95.345 179.670 ;
        RECT 95.605 174.310 95.745 187.170 ;
        RECT 96.065 178.650 96.205 189.210 ;
        RECT 98.825 187.830 98.965 192.270 ;
        RECT 101.985 191.590 102.245 191.910 ;
        RECT 99.910 190.715 101.450 191.085 ;
        RECT 98.765 187.510 99.025 187.830 ;
        RECT 102.045 186.810 102.185 191.590 ;
        RECT 103.365 191.250 103.625 191.570 ;
        RECT 103.425 189.870 103.565 191.250 ;
        RECT 103.365 189.550 103.625 189.870 ;
        RECT 105.725 189.530 105.865 192.610 ;
        RECT 108.425 191.930 108.685 192.250 ;
        RECT 108.485 189.870 108.625 191.930 ;
        RECT 108.425 189.550 108.685 189.870 ;
        RECT 105.665 189.210 105.925 189.530 ;
        RECT 105.205 188.530 105.465 188.850 ;
        RECT 101.985 186.490 102.245 186.810 ;
        RECT 99.910 185.275 101.450 185.645 ;
        RECT 102.045 184.090 102.185 186.490 ;
        RECT 105.265 184.090 105.405 188.530 ;
        RECT 108.485 187.230 108.625 189.550 ;
        RECT 108.945 187.830 109.085 192.610 ;
        RECT 108.885 187.510 109.145 187.830 ;
        RECT 108.485 187.090 109.085 187.230 ;
        RECT 96.925 183.770 97.185 184.090 ;
        RECT 98.305 183.830 98.565 184.090 ;
        RECT 97.905 183.770 98.565 183.830 ;
        RECT 101.985 183.770 102.245 184.090 ;
        RECT 105.205 183.770 105.465 184.090 ;
        RECT 96.985 181.370 97.125 183.770 ;
        RECT 97.905 183.690 98.505 183.770 ;
        RECT 96.925 181.050 97.185 181.370 ;
        RECT 96.005 178.330 96.265 178.650 ;
        RECT 96.465 178.330 96.725 178.650 ;
        RECT 96.525 176.270 96.665 178.330 ;
        RECT 96.465 175.950 96.725 176.270 ;
        RECT 94.625 173.910 94.885 174.230 ;
        RECT 95.605 174.170 96.205 174.310 ;
        RECT 94.685 171.510 94.825 173.910 ;
        RECT 95.545 173.230 95.805 173.550 ;
        RECT 95.605 171.510 95.745 173.230 ;
        RECT 94.625 171.190 94.885 171.510 ;
        RECT 95.545 171.190 95.805 171.510 ;
        RECT 94.685 170.490 94.825 171.190 ;
        RECT 94.625 170.170 94.885 170.490 ;
        RECT 94.685 167.770 94.825 170.170 ;
        RECT 94.625 167.450 94.885 167.770 ;
        RECT 95.085 166.770 95.345 167.090 ;
        RECT 95.545 166.770 95.805 167.090 ;
        RECT 95.145 165.730 95.285 166.770 ;
        RECT 95.085 165.410 95.345 165.730 ;
        RECT 95.605 165.390 95.745 166.770 ;
        RECT 95.545 165.070 95.805 165.390 ;
        RECT 94.625 162.350 94.885 162.670 ;
        RECT 94.685 162.185 94.825 162.350 ;
        RECT 94.615 161.815 94.895 162.185 ;
        RECT 95.605 161.990 95.745 165.070 ;
        RECT 95.545 161.670 95.805 161.990 ;
        RECT 95.075 159.775 95.355 160.145 ;
        RECT 95.085 159.630 95.345 159.775 ;
        RECT 95.545 159.630 95.805 159.950 ;
        RECT 95.605 159.350 95.745 159.630 ;
        RECT 95.145 159.210 95.745 159.350 ;
        RECT 94.625 158.610 94.885 158.930 ;
        RECT 94.165 151.470 94.425 151.790 ;
        RECT 94.165 150.790 94.425 151.110 ;
        RECT 93.705 150.450 93.965 150.770 ;
        RECT 93.705 149.430 93.965 149.750 ;
        RECT 93.765 149.265 93.905 149.430 ;
        RECT 93.695 148.895 93.975 149.265 ;
        RECT 94.225 149.070 94.365 150.790 ;
        RECT 94.165 148.750 94.425 149.070 ;
        RECT 94.165 148.070 94.425 148.390 ;
        RECT 93.705 146.710 93.965 147.030 ;
        RECT 93.245 146.030 93.505 146.350 ;
        RECT 92.785 145.690 93.045 146.010 ;
        RECT 92.325 143.310 92.585 143.630 ;
        RECT 92.785 141.270 93.045 141.590 ;
        RECT 92.325 140.590 92.585 140.910 ;
        RECT 91.405 140.250 91.665 140.570 ;
        RECT 91.865 140.250 92.125 140.570 ;
        RECT 91.465 139.630 91.605 140.250 ;
        RECT 91.465 139.490 92.065 139.630 ;
        RECT 91.395 138.015 91.675 138.385 ;
        RECT 91.465 137.850 91.605 138.015 ;
        RECT 90.945 137.530 91.205 137.850 ;
        RECT 91.405 137.530 91.665 137.850 ;
        RECT 91.405 134.130 91.665 134.450 ;
        RECT 91.465 133.430 91.605 134.130 ;
        RECT 91.925 133.430 92.065 139.490 ;
        RECT 92.385 134.450 92.525 140.590 ;
        RECT 92.325 134.130 92.585 134.450 ;
        RECT 91.405 133.110 91.665 133.430 ;
        RECT 91.865 133.110 92.125 133.430 ;
        RECT 91.925 129.690 92.065 133.110 ;
        RECT 92.385 132.410 92.525 134.130 ;
        RECT 92.325 132.090 92.585 132.410 ;
        RECT 92.385 130.710 92.525 132.090 ;
        RECT 92.325 130.390 92.585 130.710 ;
        RECT 91.865 129.370 92.125 129.690 ;
        RECT 91.925 127.650 92.065 129.370 ;
        RECT 91.865 127.330 92.125 127.650 ;
        RECT 92.845 125.270 92.985 141.270 ;
        RECT 93.245 135.490 93.505 135.810 ;
        RECT 93.305 129.690 93.445 135.490 ;
        RECT 93.245 129.370 93.505 129.690 ;
        RECT 93.765 127.310 93.905 146.710 ;
        RECT 94.225 146.010 94.365 148.070 ;
        RECT 94.165 145.690 94.425 146.010 ;
        RECT 94.685 143.290 94.825 158.610 ;
        RECT 95.145 156.890 95.285 159.210 ;
        RECT 95.545 156.910 95.805 157.230 ;
        RECT 95.085 156.570 95.345 156.890 ;
        RECT 95.605 156.745 95.745 156.910 ;
        RECT 95.145 155.190 95.285 156.570 ;
        RECT 95.535 156.375 95.815 156.745 ;
        RECT 95.545 155.890 95.805 156.210 ;
        RECT 95.085 154.870 95.345 155.190 ;
        RECT 95.145 151.450 95.285 154.870 ;
        RECT 95.605 154.510 95.745 155.890 ;
        RECT 96.065 154.850 96.205 174.170 ;
        RECT 96.525 172.530 96.665 175.950 ;
        RECT 96.985 175.930 97.125 181.050 ;
        RECT 96.925 175.610 97.185 175.930 ;
        RECT 96.985 174.230 97.125 175.610 ;
        RECT 96.925 173.910 97.185 174.230 ;
        RECT 96.985 173.550 97.125 173.910 ;
        RECT 96.925 173.230 97.185 173.550 ;
        RECT 96.925 172.550 97.185 172.870 ;
        RECT 96.465 172.210 96.725 172.530 ;
        RECT 96.985 171.510 97.125 172.550 ;
        RECT 96.925 171.190 97.185 171.510 ;
        RECT 97.375 167.255 97.655 167.625 ;
        RECT 96.925 166.770 97.185 167.090 ;
        RECT 96.465 165.070 96.725 165.390 ;
        RECT 96.525 162.330 96.665 165.070 ;
        RECT 96.465 162.010 96.725 162.330 ;
        RECT 96.465 161.330 96.725 161.650 ;
        RECT 96.525 157.570 96.665 161.330 ;
        RECT 96.465 157.250 96.725 157.570 ;
        RECT 96.005 154.530 96.265 154.850 ;
        RECT 95.545 154.190 95.805 154.510 ;
        RECT 95.605 152.130 95.745 154.190 ;
        RECT 95.545 151.810 95.805 152.130 ;
        RECT 95.085 151.130 95.345 151.450 ;
        RECT 96.465 151.130 96.725 151.450 ;
        RECT 95.085 150.450 95.345 150.770 ;
        RECT 95.545 150.450 95.805 150.770 ;
        RECT 95.145 146.350 95.285 150.450 ;
        RECT 95.085 146.030 95.345 146.350 ;
        RECT 95.605 146.010 95.745 150.450 ;
        RECT 96.005 146.710 96.265 147.030 ;
        RECT 95.545 145.690 95.805 146.010 ;
        RECT 94.155 142.775 94.435 143.145 ;
        RECT 94.625 142.970 94.885 143.290 ;
        RECT 95.545 142.970 95.805 143.290 ;
        RECT 94.225 138.190 94.365 142.775 ;
        RECT 95.075 140.735 95.355 141.105 ;
        RECT 94.625 140.250 94.885 140.570 ;
        RECT 94.685 138.530 94.825 140.250 ;
        RECT 94.625 138.210 94.885 138.530 ;
        RECT 94.165 137.870 94.425 138.190 ;
        RECT 94.625 137.530 94.885 137.850 ;
        RECT 94.685 135.810 94.825 137.530 ;
        RECT 94.165 135.490 94.425 135.810 ;
        RECT 94.625 135.490 94.885 135.810 ;
        RECT 93.705 126.990 93.965 127.310 ;
        RECT 92.785 124.950 93.045 125.270 ;
        RECT 92.785 124.270 93.045 124.590 ;
        RECT 92.845 121.870 92.985 124.270 ;
        RECT 92.785 121.550 93.045 121.870 ;
        RECT 94.225 110.990 94.365 135.490 ;
        RECT 95.145 135.130 95.285 140.735 ;
        RECT 95.605 140.570 95.745 142.970 ;
        RECT 95.545 140.250 95.805 140.570 ;
        RECT 95.605 138.385 95.745 140.250 ;
        RECT 95.535 138.015 95.815 138.385 ;
        RECT 95.545 136.850 95.805 137.170 ;
        RECT 95.605 135.130 95.745 136.850 ;
        RECT 95.085 134.810 95.345 135.130 ;
        RECT 95.545 134.810 95.805 135.130 ;
        RECT 96.065 134.310 96.205 146.710 ;
        RECT 96.525 143.630 96.665 151.130 ;
        RECT 96.985 146.010 97.125 166.770 ;
        RECT 97.445 165.390 97.585 167.255 ;
        RECT 97.385 165.070 97.645 165.390 ;
        RECT 97.445 162.330 97.585 165.070 ;
        RECT 97.385 162.010 97.645 162.330 ;
        RECT 97.905 159.950 98.045 183.690 ;
        RECT 100.605 183.090 100.865 183.410 ;
        RECT 101.065 183.090 101.325 183.410 ;
        RECT 104.745 183.090 105.005 183.410 ;
        RECT 108.425 183.090 108.685 183.410 ;
        RECT 100.665 181.710 100.805 183.090 ;
        RECT 100.605 181.390 100.865 181.710 ;
        RECT 101.125 180.690 101.265 183.090 ;
        RECT 104.805 182.050 104.945 183.090 ;
        RECT 108.485 182.050 108.625 183.090 ;
        RECT 108.945 182.050 109.085 187.090 ;
        RECT 104.745 181.730 105.005 182.050 ;
        RECT 108.425 181.730 108.685 182.050 ;
        RECT 108.885 181.730 109.145 182.050 ;
        RECT 99.225 180.370 99.485 180.690 ;
        RECT 101.065 180.370 101.325 180.690 ;
        RECT 98.305 175.610 98.565 175.930 ;
        RECT 98.365 172.870 98.505 175.610 ;
        RECT 98.765 173.570 99.025 173.890 ;
        RECT 98.305 172.550 98.565 172.870 ;
        RECT 98.825 165.730 98.965 173.570 ;
        RECT 98.765 165.410 99.025 165.730 ;
        RECT 97.385 159.630 97.645 159.950 ;
        RECT 97.845 159.630 98.105 159.950 ;
        RECT 98.765 159.630 99.025 159.950 ;
        RECT 97.445 157.230 97.585 159.630 ;
        RECT 98.825 157.570 98.965 159.630 ;
        RECT 98.765 157.250 99.025 157.570 ;
        RECT 97.385 156.910 97.645 157.230 ;
        RECT 99.285 156.890 99.425 180.370 ;
        RECT 99.910 179.835 101.450 180.205 ;
        RECT 105.665 178.330 105.925 178.650 ;
        RECT 102.445 177.650 102.705 177.970 ;
        RECT 102.505 176.610 102.645 177.650 ;
        RECT 102.445 176.290 102.705 176.610 ;
        RECT 101.985 174.930 102.245 175.250 ;
        RECT 99.910 174.395 101.450 174.765 ;
        RECT 101.525 171.080 101.785 171.170 ;
        RECT 102.045 171.080 102.185 174.930 ;
        RECT 102.905 172.210 103.165 172.530 ;
        RECT 103.825 172.210 104.085 172.530 ;
        RECT 101.525 170.940 102.185 171.080 ;
        RECT 101.525 170.850 101.785 170.940 ;
        RECT 101.585 169.810 101.725 170.850 ;
        RECT 102.965 170.490 103.105 172.210 ;
        RECT 103.885 171.510 104.025 172.210 ;
        RECT 105.725 171.510 105.865 178.330 ;
        RECT 107.045 177.650 107.305 177.970 ;
        RECT 107.105 173.550 107.245 177.650 ;
        RECT 108.945 175.930 109.085 181.730 ;
        RECT 108.885 175.610 109.145 175.930 ;
        RECT 108.425 174.930 108.685 175.250 ;
        RECT 108.485 174.230 108.625 174.930 ;
        RECT 108.425 173.910 108.685 174.230 ;
        RECT 108.945 173.550 109.085 175.610 ;
        RECT 107.045 173.230 107.305 173.550 ;
        RECT 108.885 173.230 109.145 173.550 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 103.825 171.190 104.085 171.510 ;
        RECT 105.665 171.190 105.925 171.510 ;
        RECT 102.905 170.170 103.165 170.490 ;
        RECT 101.985 169.830 102.245 170.150 ;
        RECT 101.525 169.490 101.785 169.810 ;
        RECT 99.910 168.955 101.450 169.325 ;
        RECT 102.045 168.110 102.185 169.830 ;
        RECT 101.985 168.020 102.245 168.110 ;
        RECT 101.985 167.880 102.645 168.020 ;
        RECT 101.985 167.790 102.245 167.880 ;
        RECT 101.985 166.770 102.245 167.090 ;
        RECT 102.045 164.370 102.185 166.770 ;
        RECT 101.985 164.050 102.245 164.370 ;
        RECT 99.910 163.515 101.450 163.885 ;
        RECT 102.045 162.330 102.185 164.050 ;
        RECT 102.505 162.580 102.645 167.880 ;
        RECT 102.965 167.090 103.105 170.170 ;
        RECT 102.905 166.770 103.165 167.090 ;
        RECT 107.505 166.770 107.765 167.090 ;
        RECT 102.965 166.070 103.105 166.770 ;
        RECT 102.905 165.750 103.165 166.070 ;
        RECT 107.565 165.730 107.705 166.770 ;
        RECT 107.505 165.410 107.765 165.730 ;
        RECT 108.945 165.390 109.085 173.230 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 108.885 165.070 109.145 165.390 ;
        RECT 103.825 162.690 104.085 163.010 ;
        RECT 102.905 162.580 103.165 162.670 ;
        RECT 102.505 162.440 103.165 162.580 ;
        RECT 102.905 162.350 103.165 162.440 ;
        RECT 103.885 162.330 104.025 162.690 ;
        RECT 101.985 162.010 102.245 162.330 ;
        RECT 103.825 162.010 104.085 162.330 ;
        RECT 105.205 162.010 105.465 162.330 ;
        RECT 107.965 162.010 108.225 162.330 ;
        RECT 101.985 161.330 102.245 161.650 ;
        RECT 102.445 161.330 102.705 161.650 ;
        RECT 102.045 160.630 102.185 161.330 ;
        RECT 101.985 160.310 102.245 160.630 ;
        RECT 102.505 159.270 102.645 161.330 ;
        RECT 102.445 158.950 102.705 159.270 ;
        RECT 99.910 158.075 101.450 158.445 ;
        RECT 102.505 156.890 102.645 158.950 ;
        RECT 103.885 157.230 104.025 162.010 ;
        RECT 105.265 160.290 105.405 162.010 ;
        RECT 105.205 159.970 105.465 160.290 ;
        RECT 108.025 159.465 108.165 162.010 ;
        RECT 108.945 159.860 109.085 165.070 ;
        RECT 109.805 161.330 110.065 161.650 ;
        RECT 109.345 159.860 109.605 159.950 ;
        RECT 108.945 159.720 109.605 159.860 ;
        RECT 107.955 159.095 108.235 159.465 ;
        RECT 103.825 156.910 104.085 157.230 ;
        RECT 99.225 156.570 99.485 156.890 ;
        RECT 102.445 156.570 102.705 156.890 ;
        RECT 97.385 155.890 97.645 156.210 ;
        RECT 96.925 145.690 97.185 146.010 ;
        RECT 96.465 143.310 96.725 143.630 ;
        RECT 96.525 141.590 96.665 143.310 ;
        RECT 96.465 141.270 96.725 141.590 ;
        RECT 96.925 140.930 97.185 141.250 ;
        RECT 96.985 139.890 97.125 140.930 ;
        RECT 96.925 139.570 97.185 139.890 ;
        RECT 96.985 138.870 97.125 139.570 ;
        RECT 96.925 138.550 97.185 138.870 ;
        RECT 96.465 135.830 96.725 136.150 ;
        RECT 96.525 135.380 96.665 135.830 ;
        RECT 97.445 135.470 97.585 155.890 ;
        RECT 102.505 154.510 102.645 156.570 ;
        RECT 102.445 154.190 102.705 154.510 ;
        RECT 98.765 153.850 99.025 154.170 ;
        RECT 98.305 151.130 98.565 151.450 ;
        RECT 97.845 150.450 98.105 150.770 ;
        RECT 97.905 149.070 98.045 150.450 ;
        RECT 97.845 148.750 98.105 149.070 ;
        RECT 97.905 147.905 98.045 148.750 ;
        RECT 98.365 148.050 98.505 151.130 ;
        RECT 98.825 149.750 98.965 153.850 ;
        RECT 99.910 152.635 101.450 153.005 ;
        RECT 103.885 151.870 104.025 156.910 ;
        RECT 106.585 153.170 106.845 153.490 ;
        RECT 103.425 151.790 104.025 151.870 ;
        RECT 106.645 151.790 106.785 153.170 ;
        RECT 103.365 151.730 104.025 151.790 ;
        RECT 103.365 151.470 103.625 151.730 ;
        RECT 99.225 150.450 99.485 150.770 ;
        RECT 98.765 149.430 99.025 149.750 ;
        RECT 99.285 149.410 99.425 150.450 ;
        RECT 99.225 149.090 99.485 149.410 ;
        RECT 97.835 147.535 98.115 147.905 ;
        RECT 98.305 147.730 98.565 148.050 ;
        RECT 97.905 144.310 98.045 147.535 ;
        RECT 97.845 143.990 98.105 144.310 ;
        RECT 98.365 143.630 98.505 147.730 ;
        RECT 99.285 146.010 99.425 149.090 ;
        RECT 101.985 147.730 102.245 148.050 ;
        RECT 102.445 147.730 102.705 148.050 ;
        RECT 99.910 147.195 101.450 147.565 ;
        RECT 102.045 146.350 102.185 147.730 ;
        RECT 102.505 146.690 102.645 147.730 ;
        RECT 102.445 146.370 102.705 146.690 ;
        RECT 101.985 146.030 102.245 146.350 ;
        RECT 99.225 145.690 99.485 146.010 ;
        RECT 99.225 143.650 99.485 143.970 ;
        RECT 98.305 143.310 98.565 143.630 ;
        RECT 98.365 143.145 98.505 143.310 ;
        RECT 98.295 142.775 98.575 143.145 ;
        RECT 97.845 142.290 98.105 142.610 ;
        RECT 96.525 135.240 97.125 135.380 ;
        RECT 96.065 134.170 96.665 134.310 ;
        RECT 94.625 132.430 94.885 132.750 ;
        RECT 94.685 130.710 94.825 132.430 ;
        RECT 94.625 130.390 94.885 130.710 ;
        RECT 96.525 127.310 96.665 134.170 ;
        RECT 94.625 126.990 94.885 127.310 ;
        RECT 96.465 126.990 96.725 127.310 ;
        RECT 94.685 124.590 94.825 126.990 ;
        RECT 95.545 125.970 95.805 126.290 ;
        RECT 95.605 124.930 95.745 125.970 ;
        RECT 95.545 124.610 95.805 124.930 ;
        RECT 94.625 124.270 94.885 124.590 ;
        RECT 96.005 123.930 96.265 124.250 ;
        RECT 96.065 121.530 96.205 123.930 ;
        RECT 96.985 122.550 97.125 135.240 ;
        RECT 97.385 135.150 97.645 135.470 ;
        RECT 97.905 134.310 98.045 142.290 ;
        RECT 98.365 140.570 98.505 142.775 ;
        RECT 98.765 142.630 99.025 142.950 ;
        RECT 98.305 140.250 98.565 140.570 ;
        RECT 98.305 134.470 98.565 134.790 ;
        RECT 97.445 134.170 98.045 134.310 ;
        RECT 97.445 125.270 97.585 134.170 ;
        RECT 98.365 133.430 98.505 134.470 ;
        RECT 98.305 133.110 98.565 133.430 ;
        RECT 97.385 124.950 97.645 125.270 ;
        RECT 98.305 124.270 98.565 124.590 ;
        RECT 96.925 122.230 97.185 122.550 ;
        RECT 94.625 121.210 94.885 121.530 ;
        RECT 96.005 121.210 96.265 121.530 ;
        RECT 94.685 116.090 94.825 121.210 ;
        RECT 96.065 117.110 96.205 121.210 ;
        RECT 97.385 120.530 97.645 120.850 ;
        RECT 96.925 119.060 97.185 119.150 ;
        RECT 96.525 118.920 97.185 119.060 ;
        RECT 96.005 116.790 96.265 117.110 ;
        RECT 94.625 115.770 94.885 116.090 ;
        RECT 96.525 114.390 96.665 118.920 ;
        RECT 96.925 118.830 97.185 118.920 ;
        RECT 96.925 116.110 97.185 116.430 ;
        RECT 96.465 114.070 96.725 114.390 ;
        RECT 94.165 110.670 94.425 110.990 ;
        RECT 93.245 109.990 93.505 110.310 ;
        RECT 91.865 109.650 92.125 109.970 ;
        RECT 90.485 108.630 90.745 108.950 ;
        RECT 90.485 107.950 90.745 108.270 ;
        RECT 88.125 106.395 89.665 106.765 ;
        RECT 86.805 105.570 87.065 105.890 ;
        RECT 86.345 102.170 86.605 102.490 ;
        RECT 88.125 100.955 89.665 101.325 ;
        RECT 90.545 98.340 90.685 107.950 ;
        RECT 91.925 107.590 92.065 109.650 ;
        RECT 91.865 107.270 92.125 107.590 ;
        RECT 93.305 105.890 93.445 109.990 ;
        RECT 95.545 109.650 95.805 109.970 ;
        RECT 95.605 108.270 95.745 109.650 ;
        RECT 96.985 108.270 97.125 116.110 ;
        RECT 97.445 113.370 97.585 120.530 ;
        RECT 98.365 117.110 98.505 124.270 ;
        RECT 98.825 121.950 98.965 142.630 ;
        RECT 99.285 140.570 99.425 143.650 ;
        RECT 102.045 143.630 102.185 146.030 ;
        RECT 101.985 143.310 102.245 143.630 ;
        RECT 99.910 141.755 101.450 142.125 ;
        RECT 102.505 140.910 102.645 146.370 ;
        RECT 103.885 146.010 104.025 151.730 ;
        RECT 106.585 151.470 106.845 151.790 ;
        RECT 108.945 151.110 109.085 159.720 ;
        RECT 109.345 159.630 109.605 159.720 ;
        RECT 109.865 159.610 110.005 161.330 ;
        RECT 109.805 159.290 110.065 159.610 ;
        RECT 108.885 150.790 109.145 151.110 ;
        RECT 110.725 150.790 110.985 151.110 ;
        RECT 105.205 149.090 105.465 149.410 ;
        RECT 105.265 147.030 105.405 149.090 ;
        RECT 110.785 149.070 110.925 150.790 ;
        RECT 110.725 148.750 110.985 149.070 ;
        RECT 108.885 148.410 109.145 148.730 ;
        RECT 108.945 147.030 109.085 148.410 ;
        RECT 105.205 146.710 105.465 147.030 ;
        RECT 108.885 146.710 109.145 147.030 ;
        RECT 103.825 145.690 104.085 146.010 ;
        RECT 103.885 143.630 104.025 145.690 ;
        RECT 107.505 145.350 107.765 145.670 ;
        RECT 105.665 145.010 105.925 145.330 ;
        RECT 103.825 143.310 104.085 143.630 ;
        RECT 99.685 140.590 99.945 140.910 ;
        RECT 102.445 140.590 102.705 140.910 ;
        RECT 99.225 140.250 99.485 140.570 ;
        RECT 99.745 138.190 99.885 140.590 ;
        RECT 99.685 137.870 99.945 138.190 ;
        RECT 101.985 137.190 102.245 137.510 ;
        RECT 99.910 136.315 101.450 136.685 ;
        RECT 99.225 135.830 99.485 136.150 ;
        RECT 99.285 133.430 99.425 135.830 ;
        RECT 102.045 133.430 102.185 137.190 ;
        RECT 99.225 133.110 99.485 133.430 ;
        RECT 101.985 133.110 102.245 133.430 ;
        RECT 102.505 132.410 102.645 140.590 ;
        RECT 103.885 137.850 104.025 143.310 ;
        RECT 103.825 137.530 104.085 137.850 ;
        RECT 104.745 134.810 105.005 135.130 ;
        RECT 104.805 133.430 104.945 134.810 ;
        RECT 104.745 133.110 105.005 133.430 ;
        RECT 102.445 132.090 102.705 132.410 ;
        RECT 99.910 130.875 101.450 131.245 ;
        RECT 104.745 126.990 105.005 127.310 ;
        RECT 99.225 126.650 99.485 126.970 ;
        RECT 99.285 123.570 99.425 126.650 ;
        RECT 99.910 125.435 101.450 125.805 ;
        RECT 100.145 124.270 100.405 124.590 ;
        RECT 99.225 123.250 99.485 123.570 ;
        RECT 99.285 122.550 99.425 123.250 ;
        RECT 99.225 122.230 99.485 122.550 ;
        RECT 98.825 121.810 99.425 121.950 ;
        RECT 98.765 118.830 99.025 119.150 ;
        RECT 98.305 116.790 98.565 117.110 ;
        RECT 98.825 116.430 98.965 118.830 ;
        RECT 98.765 116.110 99.025 116.430 ;
        RECT 97.385 113.050 97.645 113.370 ;
        RECT 99.285 110.990 99.425 121.810 ;
        RECT 100.205 121.190 100.345 124.270 ;
        RECT 102.445 123.590 102.705 123.910 ;
        RECT 102.505 121.870 102.645 123.590 ;
        RECT 104.805 121.870 104.945 126.990 ;
        RECT 102.445 121.550 102.705 121.870 ;
        RECT 104.745 121.550 105.005 121.870 ;
        RECT 100.145 120.870 100.405 121.190 ;
        RECT 99.910 119.995 101.450 120.365 ;
        RECT 102.505 119.830 102.645 121.550 ;
        RECT 102.445 119.510 102.705 119.830 ;
        RECT 100.605 117.810 100.865 118.130 ;
        RECT 100.665 116.770 100.805 117.810 ;
        RECT 100.605 116.450 100.865 116.770 ;
        RECT 102.505 116.090 102.645 119.510 ;
        RECT 104.805 118.810 104.945 121.550 ;
        RECT 105.205 120.530 105.465 120.850 ;
        RECT 104.745 118.490 105.005 118.810 ;
        RECT 105.265 118.470 105.405 120.530 ;
        RECT 105.205 118.150 105.465 118.470 ;
        RECT 102.445 115.770 102.705 116.090 ;
        RECT 99.910 114.555 101.450 114.925 ;
        RECT 105.725 110.990 105.865 145.010 ;
        RECT 106.585 143.310 106.845 143.630 ;
        RECT 106.125 142.290 106.385 142.610 ;
        RECT 106.185 140.230 106.325 142.290 ;
        RECT 106.645 141.590 106.785 143.310 ;
        RECT 106.585 141.270 106.845 141.590 ;
        RECT 106.125 139.910 106.385 140.230 ;
        RECT 106.125 137.530 106.385 137.850 ;
        RECT 106.185 135.130 106.325 137.530 ;
        RECT 106.585 136.850 106.845 137.170 ;
        RECT 106.645 135.130 106.785 136.850 ;
        RECT 106.125 134.810 106.385 135.130 ;
        RECT 106.585 134.810 106.845 135.130 ;
        RECT 107.045 123.250 107.305 123.570 ;
        RECT 107.105 116.430 107.245 123.250 ;
        RECT 107.045 116.110 107.305 116.430 ;
        RECT 107.565 110.990 107.705 145.350 ;
        RECT 108.885 142.290 109.145 142.610 ;
        RECT 108.945 140.910 109.085 142.290 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 108.885 140.590 109.145 140.910 ;
        RECT 110.725 140.250 110.985 140.570 ;
        RECT 108.885 137.870 109.145 138.190 ;
        RECT 108.945 136.150 109.085 137.870 ;
        RECT 110.785 137.850 110.925 140.250 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 110.725 137.530 110.985 137.850 ;
        RECT 108.885 135.830 109.145 136.150 ;
        RECT 110.785 127.310 110.925 137.530 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 110.725 126.990 110.985 127.310 ;
        RECT 108.885 126.650 109.145 126.970 ;
        RECT 108.945 125.270 109.085 126.650 ;
        RECT 108.885 124.950 109.145 125.270 ;
        RECT 108.885 120.530 109.145 120.850 ;
        RECT 108.945 119.150 109.085 120.530 ;
        RECT 110.785 119.150 110.925 126.990 ;
        RECT 108.885 118.830 109.145 119.150 ;
        RECT 110.725 118.830 110.985 119.150 ;
        RECT 110.785 116.430 110.925 118.830 ;
        RECT 110.725 116.110 110.985 116.430 ;
        RECT 99.225 110.670 99.485 110.990 ;
        RECT 105.665 110.670 105.925 110.990 ;
        RECT 107.505 110.670 107.765 110.990 ;
        RECT 98.765 110.330 99.025 110.650 ;
        RECT 109.805 110.330 110.065 110.650 ;
        RECT 95.545 107.950 95.805 108.270 ;
        RECT 96.925 107.950 97.185 108.270 ;
        RECT 94.165 107.270 94.425 107.590 ;
        RECT 93.245 105.570 93.505 105.890 ;
        RECT 94.225 102.150 94.365 107.270 ;
        RECT 96.985 105.550 97.125 107.950 ;
        RECT 98.825 107.930 98.965 110.330 ;
        RECT 108.885 109.990 109.145 110.310 ;
        RECT 101.985 109.650 102.245 109.970 ;
        RECT 105.665 109.650 105.925 109.970 ;
        RECT 99.910 109.115 101.450 109.485 ;
        RECT 98.765 107.610 99.025 107.930 ;
        RECT 97.385 106.930 97.645 107.250 ;
        RECT 96.925 105.230 97.185 105.550 ;
        RECT 96.985 103.510 97.125 105.230 ;
        RECT 96.925 103.190 97.185 103.510 ;
        RECT 97.445 102.830 97.585 106.930 ;
        RECT 98.825 105.550 98.965 107.610 ;
        RECT 102.045 105.890 102.185 109.650 ;
        RECT 105.725 107.590 105.865 109.650 ;
        RECT 105.665 107.270 105.925 107.590 ;
        RECT 108.425 106.930 108.685 107.250 ;
        RECT 101.985 105.570 102.245 105.890 ;
        RECT 98.765 105.230 99.025 105.550 ;
        RECT 99.225 104.890 99.485 105.210 ;
        RECT 95.085 102.510 95.345 102.830 ;
        RECT 97.385 102.510 97.645 102.830 ;
        RECT 94.165 101.830 94.425 102.150 ;
        RECT 95.145 98.340 95.285 102.510 ;
        RECT 99.285 102.400 99.425 104.890 ;
        RECT 101.985 104.210 102.245 104.530 ;
        RECT 99.910 103.675 101.450 104.045 ;
        RECT 102.045 102.490 102.185 104.210 ;
        RECT 104.285 102.510 104.545 102.830 ;
        RECT 99.285 102.260 99.885 102.400 ;
        RECT 99.745 98.340 99.885 102.260 ;
        RECT 101.985 102.170 102.245 102.490 ;
        RECT 104.345 98.340 104.485 102.510 ;
        RECT 108.485 102.230 108.625 106.930 ;
        RECT 108.945 102.830 109.085 109.990 ;
        RECT 109.345 109.650 109.605 109.970 ;
        RECT 109.405 108.270 109.545 109.650 ;
        RECT 109.345 107.950 109.605 108.270 ;
        RECT 109.865 106.230 110.005 110.330 ;
        RECT 110.785 108.270 110.925 116.110 ;
        RECT 112.565 110.670 112.825 110.990 ;
        RECT 112.625 110.505 112.765 110.670 ;
        RECT 112.555 110.135 112.835 110.505 ;
        RECT 110.725 107.950 110.985 108.270 ;
        RECT 109.805 105.910 110.065 106.230 ;
        RECT 110.785 105.550 110.925 107.950 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 110.725 105.230 110.985 105.550 ;
        RECT 110.785 102.830 110.925 105.230 ;
        RECT 108.885 102.510 109.145 102.830 ;
        RECT 110.725 102.510 110.985 102.830 ;
        RECT 108.485 102.090 109.085 102.230 ;
        RECT 108.945 98.340 109.085 102.090 ;
        RECT 21.475 96.340 21.755 98.340 ;
        RECT 26.075 96.340 26.355 98.340 ;
        RECT 30.675 96.340 30.955 98.340 ;
        RECT 35.275 96.340 35.555 98.340 ;
        RECT 39.875 96.340 40.155 98.340 ;
        RECT 44.475 96.340 44.755 98.340 ;
        RECT 49.075 96.340 49.355 98.340 ;
        RECT 53.675 96.340 53.955 98.340 ;
        RECT 58.275 96.340 58.555 98.340 ;
        RECT 62.875 96.340 63.155 98.340 ;
        RECT 67.475 96.340 67.755 98.340 ;
        RECT 72.075 96.340 72.355 98.340 ;
        RECT 76.675 96.340 76.955 98.340 ;
        RECT 81.275 96.340 81.555 98.340 ;
        RECT 85.875 96.340 86.155 98.340 ;
        RECT 90.475 96.340 90.755 98.340 ;
        RECT 95.075 96.340 95.355 98.340 ;
        RECT 99.675 96.340 99.955 98.340 ;
        RECT 104.275 96.340 104.555 98.340 ;
        RECT 108.875 96.340 109.155 98.340 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 17.380 193.455 18.960 193.785 ;
        RECT 40.955 193.455 42.535 193.785 ;
        RECT 64.530 193.455 66.110 193.785 ;
        RECT 88.105 193.455 89.685 193.785 ;
        RECT 29.165 190.735 30.745 191.065 ;
        RECT 52.740 190.735 54.320 191.065 ;
        RECT 76.315 190.735 77.895 191.065 ;
        RECT 99.890 190.735 101.470 191.065 ;
        RECT 17.380 188.015 18.960 188.345 ;
        RECT 40.955 188.015 42.535 188.345 ;
        RECT 64.530 188.015 66.110 188.345 ;
        RECT 88.105 188.015 89.685 188.345 ;
        RECT 29.165 185.295 30.745 185.625 ;
        RECT 52.740 185.295 54.320 185.625 ;
        RECT 76.315 185.295 77.895 185.625 ;
        RECT 99.890 185.295 101.470 185.625 ;
        RECT 17.380 182.575 18.960 182.905 ;
        RECT 40.955 182.575 42.535 182.905 ;
        RECT 64.530 182.575 66.110 182.905 ;
        RECT 88.105 182.575 89.685 182.905 ;
        RECT 29.165 179.855 30.745 180.185 ;
        RECT 52.740 179.855 54.320 180.185 ;
        RECT 76.315 179.855 77.895 180.185 ;
        RECT 99.890 179.855 101.470 180.185 ;
        RECT 17.380 177.135 18.960 177.465 ;
        RECT 40.955 177.135 42.535 177.465 ;
        RECT 64.530 177.135 66.110 177.465 ;
        RECT 88.105 177.135 89.685 177.465 ;
        RECT 29.165 174.415 30.745 174.745 ;
        RECT 52.740 174.415 54.320 174.745 ;
        RECT 76.315 174.415 77.895 174.745 ;
        RECT 99.890 174.415 101.470 174.745 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 17.380 171.695 18.960 172.025 ;
        RECT 40.955 171.695 42.535 172.025 ;
        RECT 64.530 171.695 66.110 172.025 ;
        RECT 88.105 171.695 89.685 172.025 ;
        RECT 36.630 170.990 36.960 171.005 ;
        RECT 52.270 170.990 52.600 171.005 ;
        RECT 36.630 170.690 52.600 170.990 ;
        RECT 36.630 170.675 36.960 170.690 ;
        RECT 52.270 170.675 52.600 170.690 ;
        RECT 59.170 170.990 59.500 171.005 ;
        RECT 64.230 170.990 64.560 171.005 ;
        RECT 59.170 170.690 64.560 170.990 ;
        RECT 59.170 170.675 59.500 170.690 ;
        RECT 64.230 170.675 64.560 170.690 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 29.165 168.975 30.745 169.305 ;
        RECT 52.740 168.975 54.320 169.305 ;
        RECT 76.315 168.975 77.895 169.305 ;
        RECT 99.890 168.975 101.470 169.305 ;
        RECT 21.910 167.590 22.240 167.605 ;
        RECT 35.250 167.590 35.580 167.605 ;
        RECT 21.910 167.290 35.580 167.590 ;
        RECT 21.910 167.275 22.240 167.290 ;
        RECT 35.250 167.275 35.580 167.290 ;
        RECT 59.170 167.590 59.500 167.605 ;
        RECT 66.070 167.590 66.400 167.605 ;
        RECT 59.170 167.290 66.400 167.590 ;
        RECT 59.170 167.275 59.500 167.290 ;
        RECT 66.070 167.275 66.400 167.290 ;
        RECT 68.370 167.590 68.700 167.605 ;
        RECT 86.770 167.590 87.100 167.605 ;
        RECT 90.910 167.590 91.240 167.605 ;
        RECT 92.750 167.590 93.080 167.605 ;
        RECT 97.350 167.590 97.680 167.605 ;
        RECT 68.370 167.290 97.680 167.590 ;
        RECT 68.370 167.275 68.700 167.290 ;
        RECT 86.770 167.275 87.100 167.290 ;
        RECT 90.910 167.275 91.240 167.290 ;
        RECT 92.750 167.275 93.080 167.290 ;
        RECT 97.350 167.275 97.680 167.290 ;
        RECT 43.530 166.910 43.860 166.925 ;
        RECT 48.335 166.910 48.715 166.920 ;
        RECT 43.530 166.610 48.715 166.910 ;
        RECT 43.530 166.595 43.860 166.610 ;
        RECT 48.335 166.600 48.715 166.610 ;
        RECT 17.380 166.255 18.960 166.585 ;
        RECT 40.955 166.255 42.535 166.585 ;
        RECT 64.530 166.255 66.110 166.585 ;
        RECT 88.105 166.255 89.685 166.585 ;
        RECT 29.165 163.535 30.745 163.865 ;
        RECT 52.740 163.535 54.320 163.865 ;
        RECT 76.315 163.535 77.895 163.865 ;
        RECT 99.890 163.535 101.470 163.865 ;
        RECT 47.670 162.830 48.000 162.845 ;
        RECT 61.930 162.830 62.260 162.845 ;
        RECT 47.670 162.530 62.260 162.830 ;
        RECT 47.670 162.515 48.000 162.530 ;
        RECT 61.930 162.515 62.260 162.530 ;
        RECT 80.790 162.830 81.120 162.845 ;
        RECT 87.230 162.830 87.560 162.845 ;
        RECT 80.790 162.530 87.560 162.830 ;
        RECT 80.790 162.515 81.120 162.530 ;
        RECT 87.230 162.515 87.560 162.530 ;
        RECT 73.890 162.150 74.220 162.165 ;
        RECT 94.590 162.160 94.920 162.165 ;
        RECT 94.335 162.150 94.920 162.160 ;
        RECT 73.890 161.835 74.435 162.150 ;
        RECT 94.335 161.850 95.145 162.150 ;
        RECT 94.335 161.840 94.920 161.850 ;
        RECT 94.590 161.835 94.920 161.840 ;
        RECT 17.380 160.815 18.960 161.145 ;
        RECT 40.955 160.815 42.535 161.145 ;
        RECT 64.530 160.815 66.110 161.145 ;
        RECT 74.135 160.110 74.435 161.835 ;
        RECT 88.105 160.815 89.685 161.145 ;
        RECT 75.015 160.110 75.395 160.120 ;
        RECT 95.050 160.110 95.380 160.125 ;
        RECT 74.135 159.810 95.380 160.110 ;
        RECT 75.015 159.800 75.395 159.810 ;
        RECT 95.050 159.795 95.380 159.810 ;
        RECT 53.650 159.430 53.980 159.445 ;
        RECT 60.090 159.430 60.420 159.445 ;
        RECT 53.650 159.130 60.420 159.430 ;
        RECT 53.650 159.115 53.980 159.130 ;
        RECT 60.090 159.115 60.420 159.130 ;
        RECT 107.930 159.430 108.260 159.445 ;
        RECT 113.225 159.430 115.225 159.580 ;
        RECT 107.930 159.130 115.225 159.430 ;
        RECT 107.930 159.115 108.260 159.130 ;
        RECT 113.225 158.980 115.225 159.130 ;
        RECT 29.165 158.095 30.745 158.425 ;
        RECT 52.740 158.095 54.320 158.425 ;
        RECT 76.315 158.095 77.895 158.425 ;
        RECT 99.890 158.095 101.470 158.425 ;
        RECT 95.510 156.710 95.840 156.725 ;
        RECT 94.375 156.410 95.840 156.710 ;
        RECT 49.970 156.030 50.300 156.045 ;
        RECT 59.170 156.030 59.500 156.045 ;
        RECT 63.770 156.030 64.100 156.045 ;
        RECT 49.970 155.730 64.100 156.030 ;
        RECT 49.970 155.715 50.300 155.730 ;
        RECT 59.170 155.715 59.500 155.730 ;
        RECT 63.770 155.715 64.100 155.730 ;
        RECT 93.670 156.030 94.000 156.045 ;
        RECT 94.375 156.030 94.675 156.410 ;
        RECT 95.510 156.395 95.840 156.410 ;
        RECT 93.670 155.730 94.675 156.030 ;
        RECT 93.670 155.715 94.000 155.730 ;
        RECT 17.380 155.375 18.960 155.705 ;
        RECT 40.955 155.375 42.535 155.705 ;
        RECT 64.530 155.375 66.110 155.705 ;
        RECT 88.105 155.375 89.685 155.705 ;
        RECT 64.690 154.670 65.020 154.685 ;
        RECT 66.070 154.670 66.400 154.685 ;
        RECT 64.690 154.370 66.400 154.670 ;
        RECT 64.690 154.355 65.020 154.370 ;
        RECT 66.070 154.355 66.400 154.370 ;
        RECT 67.910 153.990 68.240 154.005 ;
        RECT 75.270 153.990 75.600 154.005 ;
        RECT 67.910 153.690 75.600 153.990 ;
        RECT 67.910 153.675 68.240 153.690 ;
        RECT 75.270 153.675 75.600 153.690 ;
        RECT 29.165 152.655 30.745 152.985 ;
        RECT 52.740 152.655 54.320 152.985 ;
        RECT 76.315 152.655 77.895 152.985 ;
        RECT 99.890 152.655 101.470 152.985 ;
        RECT 36.375 151.950 36.755 151.960 ;
        RECT 45.370 151.950 45.700 151.965 ;
        RECT 36.375 151.650 45.700 151.950 ;
        RECT 36.375 151.640 36.755 151.650 ;
        RECT 45.370 151.635 45.700 151.650 ;
        RECT 59.630 151.950 59.960 151.965 ;
        RECT 67.450 151.950 67.780 151.965 ;
        RECT 59.630 151.650 67.780 151.950 ;
        RECT 59.630 151.635 59.960 151.650 ;
        RECT 63.770 151.270 64.100 151.285 ;
        RECT 63.095 150.970 64.100 151.270 ;
        RECT 17.380 149.935 18.960 150.265 ;
        RECT 40.955 149.935 42.535 150.265 ;
        RECT 55.490 149.910 55.820 149.925 ;
        RECT 63.095 149.910 63.395 150.970 ;
        RECT 63.770 150.955 64.100 150.970 ;
        RECT 64.530 149.935 66.110 150.265 ;
        RECT 55.490 149.610 63.395 149.910 ;
        RECT 55.490 149.595 55.820 149.610 ;
        RECT 32.030 149.230 32.360 149.245 ;
        RECT 60.550 149.230 60.880 149.245 ;
        RECT 32.030 148.930 60.880 149.230 ;
        RECT 63.095 149.230 63.395 149.610 ;
        RECT 64.690 149.230 65.020 149.245 ;
        RECT 63.095 148.930 65.020 149.230 ;
        RECT 32.030 148.915 32.360 148.930 ;
        RECT 60.550 148.915 60.880 148.930 ;
        RECT 64.690 148.915 65.020 148.930 ;
        RECT 66.545 148.565 66.845 151.650 ;
        RECT 67.450 151.635 67.780 151.650 ;
        RECT 88.105 149.935 89.685 150.265 ;
        RECT 83.550 149.230 83.880 149.245 ;
        RECT 93.670 149.230 94.000 149.245 ;
        RECT 83.550 148.930 94.000 149.230 ;
        RECT 83.550 148.915 83.880 148.930 ;
        RECT 93.670 148.915 94.000 148.930 ;
        RECT 42.610 148.550 42.940 148.565 ;
        RECT 42.610 148.235 43.155 148.550 ;
        RECT 66.530 148.235 66.860 148.565 ;
        RECT 67.450 148.550 67.780 148.565 ;
        RECT 68.370 148.550 68.700 148.565 ;
        RECT 87.230 148.550 87.560 148.565 ;
        RECT 67.450 148.250 87.560 148.550 ;
        RECT 67.450 148.235 67.780 148.250 ;
        RECT 68.370 148.235 68.700 148.250 ;
        RECT 87.230 148.235 87.560 148.250 ;
        RECT 42.855 147.870 43.155 148.235 ;
        RECT 46.495 147.870 46.875 147.880 ;
        RECT 42.855 147.570 46.875 147.870 ;
        RECT 46.495 147.560 46.875 147.570 ;
        RECT 87.230 147.870 87.560 147.885 ;
        RECT 97.810 147.870 98.140 147.885 ;
        RECT 87.230 147.570 98.140 147.870 ;
        RECT 87.230 147.555 87.560 147.570 ;
        RECT 97.810 147.555 98.140 147.570 ;
        RECT 29.165 147.215 30.745 147.545 ;
        RECT 52.740 147.215 54.320 147.545 ;
        RECT 76.315 147.215 77.895 147.545 ;
        RECT 99.890 147.215 101.470 147.545 ;
        RECT 49.510 146.510 49.840 146.525 ;
        RECT 62.850 146.510 63.180 146.525 ;
        RECT 49.510 146.210 63.180 146.510 ;
        RECT 49.510 146.195 49.840 146.210 ;
        RECT 62.850 146.195 63.180 146.210 ;
        RECT 67.910 146.510 68.240 146.525 ;
        RECT 86.770 146.510 87.100 146.525 ;
        RECT 67.910 146.210 87.100 146.510 ;
        RECT 67.910 146.195 68.240 146.210 ;
        RECT 86.770 146.195 87.100 146.210 ;
        RECT 70.210 145.160 70.540 145.165 ;
        RECT 70.210 145.150 70.795 145.160 ;
        RECT 69.985 144.850 70.795 145.150 ;
        RECT 70.210 144.840 70.795 144.850 ;
        RECT 70.210 144.835 70.540 144.840 ;
        RECT 17.380 144.495 18.960 144.825 ;
        RECT 40.955 144.495 42.535 144.825 ;
        RECT 64.530 144.495 66.110 144.825 ;
        RECT 88.105 144.495 89.685 144.825 ;
        RECT 46.495 144.470 46.875 144.480 ;
        RECT 46.495 144.170 53.275 144.470 ;
        RECT 46.495 144.160 46.875 144.170 ;
        RECT 52.975 143.110 53.275 144.170 ;
        RECT 54.570 143.110 54.900 143.125 ;
        RECT 75.015 143.110 75.395 143.120 ;
        RECT 52.975 142.810 75.395 143.110 ;
        RECT 54.570 142.795 54.900 142.810 ;
        RECT 75.015 142.800 75.395 142.810 ;
        RECT 94.130 143.110 94.460 143.125 ;
        RECT 98.270 143.110 98.600 143.125 ;
        RECT 94.130 142.810 98.600 143.110 ;
        RECT 94.130 142.795 94.460 142.810 ;
        RECT 98.270 142.795 98.600 142.810 ;
        RECT 29.165 141.775 30.745 142.105 ;
        RECT 52.740 141.775 54.320 142.105 ;
        RECT 76.315 141.775 77.895 142.105 ;
        RECT 99.890 141.775 101.470 142.105 ;
        RECT 94.335 141.070 94.715 141.080 ;
        RECT 95.050 141.070 95.380 141.085 ;
        RECT 94.335 140.770 95.380 141.070 ;
        RECT 94.335 140.760 94.715 140.770 ;
        RECT 95.050 140.755 95.380 140.770 ;
        RECT 17.380 139.055 18.960 139.385 ;
        RECT 40.955 139.055 42.535 139.385 ;
        RECT 64.530 139.055 66.110 139.385 ;
        RECT 88.105 139.055 89.685 139.385 ;
        RECT 88.150 138.350 88.480 138.365 ;
        RECT 91.370 138.350 91.700 138.365 ;
        RECT 95.510 138.350 95.840 138.365 ;
        RECT 88.150 138.050 95.840 138.350 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 88.150 138.035 88.480 138.050 ;
        RECT 91.370 138.035 91.700 138.050 ;
        RECT 95.510 138.035 95.840 138.050 ;
        RECT 29.165 136.335 30.745 136.665 ;
        RECT 52.740 136.335 54.320 136.665 ;
        RECT 76.315 136.335 77.895 136.665 ;
        RECT 99.890 136.335 101.470 136.665 ;
        RECT 37.090 134.950 37.420 134.965 ;
        RECT 40.310 134.950 40.640 134.965 ;
        RECT 55.950 134.950 56.280 134.965 ;
        RECT 37.090 134.650 56.280 134.950 ;
        RECT 37.090 134.635 37.420 134.650 ;
        RECT 40.310 134.635 40.640 134.650 ;
        RECT 55.950 134.635 56.280 134.650 ;
        RECT 61.010 134.950 61.340 134.965 ;
        RECT 113.225 134.950 115.225 135.100 ;
        RECT 61.010 134.650 115.225 134.950 ;
        RECT 61.010 134.635 61.340 134.650 ;
        RECT 113.225 134.500 115.225 134.650 ;
        RECT 48.590 134.280 48.920 134.285 ;
        RECT 48.335 134.270 48.920 134.280 ;
        RECT 48.135 133.970 48.920 134.270 ;
        RECT 48.335 133.960 48.920 133.970 ;
        RECT 48.590 133.955 48.920 133.960 ;
        RECT 60.550 134.270 60.880 134.285 ;
        RECT 62.390 134.270 62.720 134.285 ;
        RECT 60.550 133.970 62.720 134.270 ;
        RECT 60.550 133.955 60.880 133.970 ;
        RECT 62.390 133.955 62.720 133.970 ;
        RECT 17.380 133.615 18.960 133.945 ;
        RECT 40.955 133.615 42.535 133.945 ;
        RECT 64.530 133.615 66.110 133.945 ;
        RECT 88.105 133.615 89.685 133.945 ;
        RECT 29.165 130.895 30.745 131.225 ;
        RECT 52.740 130.895 54.320 131.225 ;
        RECT 76.315 130.895 77.895 131.225 ;
        RECT 99.890 130.895 101.470 131.225 ;
        RECT 75.015 130.190 75.395 130.200 ;
        RECT 79.410 130.190 79.740 130.205 ;
        RECT 75.015 129.890 79.740 130.190 ;
        RECT 75.015 129.880 75.395 129.890 ;
        RECT 79.410 129.875 79.740 129.890 ;
        RECT 17.380 128.175 18.960 128.505 ;
        RECT 40.955 128.175 42.535 128.505 ;
        RECT 64.530 128.175 66.110 128.505 ;
        RECT 88.105 128.175 89.685 128.505 ;
        RECT 29.165 125.455 30.745 125.785 ;
        RECT 52.740 125.455 54.320 125.785 ;
        RECT 76.315 125.455 77.895 125.785 ;
        RECT 99.890 125.455 101.470 125.785 ;
        RECT 46.750 124.760 47.080 124.765 ;
        RECT 46.495 124.750 47.080 124.760 ;
        RECT 46.495 124.450 47.305 124.750 ;
        RECT 46.495 124.440 47.080 124.450 ;
        RECT 46.750 124.435 47.080 124.440 ;
        RECT 17.380 122.735 18.960 123.065 ;
        RECT 40.955 122.735 42.535 123.065 ;
        RECT 64.530 122.735 66.110 123.065 ;
        RECT 88.105 122.735 89.685 123.065 ;
        RECT 29.165 120.015 30.745 120.345 ;
        RECT 52.740 120.015 54.320 120.345 ;
        RECT 76.315 120.015 77.895 120.345 ;
        RECT 99.890 120.015 101.470 120.345 ;
        RECT 17.380 117.295 18.960 117.625 ;
        RECT 40.955 117.295 42.535 117.625 ;
        RECT 64.530 117.295 66.110 117.625 ;
        RECT 88.105 117.295 89.685 117.625 ;
        RECT 29.165 114.575 30.745 114.905 ;
        RECT 52.740 114.575 54.320 114.905 ;
        RECT 76.315 114.575 77.895 114.905 ;
        RECT 99.890 114.575 101.470 114.905 ;
        RECT 17.380 111.855 18.960 112.185 ;
        RECT 40.955 111.855 42.535 112.185 ;
        RECT 64.530 111.855 66.110 112.185 ;
        RECT 88.105 111.855 89.685 112.185 ;
        RECT 36.375 110.470 36.755 110.480 ;
        RECT 37.090 110.470 37.420 110.485 ;
        RECT 36.375 110.170 37.420 110.470 ;
        RECT 36.375 110.160 36.755 110.170 ;
        RECT 37.090 110.155 37.420 110.170 ;
        RECT 112.530 110.470 112.860 110.485 ;
        RECT 113.225 110.470 115.225 110.620 ;
        RECT 112.530 110.170 115.225 110.470 ;
        RECT 112.530 110.155 112.860 110.170 ;
        RECT 113.225 110.020 115.225 110.170 ;
        RECT 29.165 109.135 30.745 109.465 ;
        RECT 52.740 109.135 54.320 109.465 ;
        RECT 76.315 109.135 77.895 109.465 ;
        RECT 99.890 109.135 101.470 109.465 ;
        RECT 17.380 106.415 18.960 106.745 ;
        RECT 40.955 106.415 42.535 106.745 ;
        RECT 64.530 106.415 66.110 106.745 ;
        RECT 88.105 106.415 89.685 106.745 ;
        RECT 70.415 106.390 70.795 106.400 ;
        RECT 72.050 106.390 72.380 106.405 ;
        RECT 70.415 106.090 72.380 106.390 ;
        RECT 70.415 106.080 70.795 106.090 ;
        RECT 72.050 106.075 72.380 106.090 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 29.165 103.695 30.745 104.025 ;
        RECT 52.740 103.695 54.320 104.025 ;
        RECT 76.315 103.695 77.895 104.025 ;
        RECT 99.890 103.695 101.470 104.025 ;
        RECT 17.380 100.975 18.960 101.305 ;
        RECT 40.955 100.975 42.535 101.305 ;
        RECT 64.530 100.975 66.110 101.305 ;
        RECT 88.105 100.975 89.685 101.305 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 17.370 100.900 18.970 193.860 ;
        RECT 29.155 100.900 30.755 193.860 ;
        RECT 36.400 151.635 36.730 151.965 ;
        RECT 36.415 110.485 36.715 151.635 ;
        RECT 36.400 110.155 36.730 110.485 ;
        RECT 40.945 100.900 42.545 193.860 ;
        RECT 48.360 166.595 48.690 166.925 ;
        RECT 46.520 147.555 46.850 147.885 ;
        RECT 46.535 144.485 46.835 147.555 ;
        RECT 46.520 144.155 46.850 144.485 ;
        RECT 46.535 124.765 46.835 144.155 ;
        RECT 48.375 134.285 48.675 166.595 ;
        RECT 48.360 133.955 48.690 134.285 ;
        RECT 46.520 124.435 46.850 124.765 ;
        RECT 52.730 100.900 54.330 193.860 ;
        RECT 64.520 100.900 66.120 193.860 ;
        RECT 75.040 159.795 75.370 160.125 ;
        RECT 70.440 144.835 70.770 145.165 ;
        RECT 70.455 106.405 70.755 144.835 ;
        RECT 75.055 143.125 75.355 159.795 ;
        RECT 75.040 142.795 75.370 143.125 ;
        RECT 75.055 130.205 75.355 142.795 ;
        RECT 75.040 129.875 75.370 130.205 ;
        RECT 70.440 106.075 70.770 106.405 ;
        RECT 76.305 100.900 77.905 193.860 ;
        RECT 88.095 100.900 89.695 193.860 ;
        RECT 94.360 161.835 94.690 162.165 ;
        RECT 94.375 141.085 94.675 161.835 ;
        RECT 94.360 140.755 94.690 141.085 ;
        RECT 99.880 100.900 101.480 193.860 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

