VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 11.955 215.865 12.125 216.055 ;
        RECT 16.555 215.865 16.725 216.055 ;
        RECT 22.075 215.865 22.245 216.055 ;
        RECT 23.915 215.865 24.085 216.055 ;
        RECT 29.435 215.865 29.605 216.055 ;
        RECT 34.955 215.865 35.125 216.055 ;
        RECT 36.795 215.865 36.965 216.055 ;
        RECT 42.315 215.865 42.485 216.055 ;
        RECT 47.835 215.865 48.005 216.055 ;
        RECT 49.675 215.865 49.845 216.055 ;
        RECT 55.195 215.865 55.365 216.055 ;
        RECT 60.715 215.865 60.885 216.055 ;
        RECT 62.555 215.865 62.725 216.055 ;
        RECT 68.075 215.865 68.245 216.055 ;
        RECT 73.595 215.865 73.765 216.055 ;
        RECT 75.435 215.865 75.605 216.055 ;
        RECT 80.955 215.865 81.125 216.055 ;
        RECT 86.475 215.865 86.645 216.055 ;
        RECT 88.315 215.865 88.485 216.055 ;
        RECT 93.835 215.865 94.005 216.055 ;
        RECT 99.355 215.865 99.525 216.055 ;
        RECT 101.195 215.865 101.365 216.055 ;
        RECT 106.715 215.865 106.885 216.055 ;
        RECT 112.235 215.865 112.405 216.055 ;
        RECT 113.210 215.915 113.330 216.025 ;
        RECT 118.675 215.865 118.845 216.055 ;
        RECT 124.195 215.865 124.365 216.055 ;
        RECT 125.575 215.865 125.745 216.055 ;
        RECT 11.815 215.055 13.185 215.865 ;
        RECT 13.195 215.055 16.865 215.865 ;
        RECT 16.875 215.055 22.385 215.865 ;
        RECT 22.405 214.995 22.835 215.780 ;
        RECT 22.855 215.055 24.225 215.865 ;
        RECT 24.235 215.055 29.745 215.865 ;
        RECT 29.755 215.055 35.265 215.865 ;
        RECT 35.285 214.995 35.715 215.780 ;
        RECT 35.735 215.055 37.105 215.865 ;
        RECT 37.115 215.055 42.625 215.865 ;
        RECT 42.635 215.055 48.145 215.865 ;
        RECT 48.165 214.995 48.595 215.780 ;
        RECT 48.615 215.055 49.985 215.865 ;
        RECT 49.995 215.055 55.505 215.865 ;
        RECT 55.515 215.055 61.025 215.865 ;
        RECT 61.045 214.995 61.475 215.780 ;
        RECT 61.495 215.055 62.865 215.865 ;
        RECT 62.875 215.055 68.385 215.865 ;
        RECT 68.395 215.055 73.905 215.865 ;
        RECT 73.925 214.995 74.355 215.780 ;
        RECT 74.375 215.055 75.745 215.865 ;
        RECT 75.755 215.055 81.265 215.865 ;
        RECT 81.275 215.055 86.785 215.865 ;
        RECT 86.805 214.995 87.235 215.780 ;
        RECT 87.255 215.055 88.625 215.865 ;
        RECT 88.635 215.055 94.145 215.865 ;
        RECT 94.155 215.055 99.665 215.865 ;
        RECT 99.685 214.995 100.115 215.780 ;
        RECT 100.135 215.055 101.505 215.865 ;
        RECT 101.515 215.055 107.025 215.865 ;
        RECT 107.035 215.055 112.545 215.865 ;
        RECT 112.565 214.995 112.995 215.780 ;
        RECT 113.475 215.055 118.985 215.865 ;
        RECT 118.995 215.055 124.505 215.865 ;
        RECT 124.515 215.055 125.885 215.865 ;
      LAYER nwell ;
        RECT 11.620 211.835 126.080 214.665 ;
      LAYER pwell ;
        RECT 11.815 210.635 13.185 211.445 ;
        RECT 13.195 210.635 16.865 211.445 ;
        RECT 16.875 210.635 22.385 211.445 ;
        RECT 22.405 210.720 22.835 211.505 ;
        RECT 23.315 210.635 26.065 211.445 ;
        RECT 26.075 210.635 31.585 211.445 ;
        RECT 31.595 210.635 37.105 211.445 ;
        RECT 37.115 210.635 42.625 211.445 ;
        RECT 42.635 210.635 48.145 211.445 ;
        RECT 48.165 210.720 48.595 211.505 ;
        RECT 49.075 210.635 51.825 211.445 ;
        RECT 51.835 210.635 57.345 211.445 ;
        RECT 57.355 210.635 62.865 211.445 ;
        RECT 62.875 210.635 68.385 211.445 ;
        RECT 68.395 210.635 73.905 211.445 ;
        RECT 73.925 210.720 74.355 211.505 ;
        RECT 74.835 210.635 77.585 211.445 ;
        RECT 77.595 210.635 83.105 211.445 ;
        RECT 83.115 210.635 88.625 211.445 ;
        RECT 88.635 210.635 94.145 211.445 ;
        RECT 94.155 210.635 99.665 211.445 ;
        RECT 99.685 210.720 100.115 211.505 ;
        RECT 100.595 210.635 102.425 211.445 ;
        RECT 102.435 210.635 107.945 211.445 ;
        RECT 107.955 210.635 113.465 211.445 ;
        RECT 113.475 210.635 118.985 211.445 ;
        RECT 118.995 210.635 124.505 211.445 ;
        RECT 124.515 210.635 125.885 211.445 ;
        RECT 11.955 210.425 12.125 210.635 ;
        RECT 16.555 210.445 16.725 210.635 ;
        RECT 18.395 210.425 18.565 210.615 ;
        RECT 22.075 210.445 22.245 210.635 ;
        RECT 23.050 210.475 23.170 210.585 ;
        RECT 23.915 210.425 24.085 210.615 ;
        RECT 25.755 210.445 25.925 210.635 ;
        RECT 29.435 210.425 29.605 210.615 ;
        RECT 31.275 210.445 31.445 210.635 ;
        RECT 34.955 210.425 35.125 210.615 ;
        RECT 35.930 210.475 36.050 210.585 ;
        RECT 36.795 210.445 36.965 210.635 ;
        RECT 38.635 210.425 38.805 210.615 ;
        RECT 42.315 210.445 42.485 210.635 ;
        RECT 44.155 210.425 44.325 210.615 ;
        RECT 47.835 210.445 48.005 210.635 ;
        RECT 48.810 210.475 48.930 210.585 ;
        RECT 49.675 210.425 49.845 210.615 ;
        RECT 51.515 210.445 51.685 210.635 ;
        RECT 55.195 210.425 55.365 210.615 ;
        RECT 57.035 210.445 57.205 210.635 ;
        RECT 60.715 210.425 60.885 210.615 ;
        RECT 61.690 210.475 61.810 210.585 ;
        RECT 62.555 210.445 62.725 210.635 ;
        RECT 64.395 210.425 64.565 210.615 ;
        RECT 68.075 210.445 68.245 210.635 ;
        RECT 69.915 210.425 70.085 210.615 ;
        RECT 73.595 210.445 73.765 210.635 ;
        RECT 74.570 210.475 74.690 210.585 ;
        RECT 75.435 210.425 75.605 210.615 ;
        RECT 77.275 210.445 77.445 210.635 ;
        RECT 80.955 210.425 81.125 210.615 ;
        RECT 82.795 210.445 82.965 210.635 ;
        RECT 86.475 210.425 86.645 210.615 ;
        RECT 87.450 210.475 87.570 210.585 ;
        RECT 88.315 210.445 88.485 210.635 ;
        RECT 90.155 210.425 90.325 210.615 ;
        RECT 93.835 210.445 94.005 210.635 ;
        RECT 95.675 210.425 95.845 210.615 ;
        RECT 99.355 210.445 99.525 210.635 ;
        RECT 100.330 210.475 100.450 210.585 ;
        RECT 101.195 210.425 101.365 210.615 ;
        RECT 102.115 210.445 102.285 210.635 ;
        RECT 106.715 210.425 106.885 210.615 ;
        RECT 107.635 210.445 107.805 210.635 ;
        RECT 112.235 210.425 112.405 210.615 ;
        RECT 113.155 210.585 113.325 210.635 ;
        RECT 113.155 210.475 113.330 210.585 ;
        RECT 113.155 210.445 113.325 210.475 ;
        RECT 118.675 210.425 118.845 210.635 ;
        RECT 124.195 210.425 124.365 210.635 ;
        RECT 125.575 210.425 125.745 210.635 ;
        RECT 11.815 209.615 13.185 210.425 ;
        RECT 13.195 209.615 18.705 210.425 ;
        RECT 18.715 209.615 24.225 210.425 ;
        RECT 24.235 209.615 29.745 210.425 ;
        RECT 29.755 209.615 35.265 210.425 ;
        RECT 35.285 209.555 35.715 210.340 ;
        RECT 36.195 209.615 38.945 210.425 ;
        RECT 38.955 209.615 44.465 210.425 ;
        RECT 44.475 209.615 49.985 210.425 ;
        RECT 49.995 209.615 55.505 210.425 ;
        RECT 55.515 209.615 61.025 210.425 ;
        RECT 61.045 209.555 61.475 210.340 ;
        RECT 61.955 209.615 64.705 210.425 ;
        RECT 64.715 209.615 70.225 210.425 ;
        RECT 70.235 209.615 75.745 210.425 ;
        RECT 75.755 209.615 81.265 210.425 ;
        RECT 81.275 209.615 86.785 210.425 ;
        RECT 86.805 209.555 87.235 210.340 ;
        RECT 87.715 209.615 90.465 210.425 ;
        RECT 90.475 209.615 95.985 210.425 ;
        RECT 95.995 209.615 101.505 210.425 ;
        RECT 101.515 209.615 107.025 210.425 ;
        RECT 107.035 209.615 112.545 210.425 ;
        RECT 112.565 209.555 112.995 210.340 ;
        RECT 113.475 209.615 118.985 210.425 ;
        RECT 118.995 209.615 124.505 210.425 ;
        RECT 124.515 209.615 125.885 210.425 ;
      LAYER nwell ;
        RECT 11.620 206.395 126.080 209.225 ;
      LAYER pwell ;
        RECT 11.815 205.195 13.185 206.005 ;
        RECT 13.195 205.195 16.865 206.005 ;
        RECT 16.875 205.195 22.385 206.005 ;
        RECT 22.405 205.280 22.835 206.065 ;
        RECT 23.315 205.195 26.065 206.005 ;
        RECT 26.075 205.195 31.585 206.005 ;
        RECT 31.595 205.195 37.105 206.005 ;
        RECT 37.115 205.195 42.625 206.005 ;
        RECT 42.635 205.195 48.145 206.005 ;
        RECT 48.165 205.280 48.595 206.065 ;
        RECT 49.075 205.195 51.825 206.005 ;
        RECT 51.835 205.195 57.345 206.005 ;
        RECT 57.355 205.195 62.865 206.005 ;
        RECT 62.875 205.195 68.385 206.005 ;
        RECT 68.395 205.195 73.905 206.005 ;
        RECT 73.925 205.280 74.355 206.065 ;
        RECT 74.835 205.195 77.585 206.005 ;
        RECT 77.595 205.195 83.105 206.005 ;
        RECT 83.115 205.195 88.625 206.005 ;
        RECT 88.635 205.195 94.145 206.005 ;
        RECT 94.155 205.195 99.665 206.005 ;
        RECT 99.685 205.280 100.115 206.065 ;
        RECT 100.595 205.195 102.425 206.005 ;
        RECT 102.435 205.195 107.945 206.005 ;
        RECT 107.955 205.195 113.465 206.005 ;
        RECT 113.475 205.195 118.985 206.005 ;
        RECT 118.995 205.195 124.505 206.005 ;
        RECT 124.515 205.195 125.885 206.005 ;
        RECT 11.955 204.985 12.125 205.195 ;
        RECT 16.555 205.005 16.725 205.195 ;
        RECT 18.395 204.985 18.565 205.175 ;
        RECT 22.075 205.005 22.245 205.195 ;
        RECT 23.050 205.035 23.170 205.145 ;
        RECT 23.915 204.985 24.085 205.175 ;
        RECT 25.755 205.005 25.925 205.195 ;
        RECT 29.435 204.985 29.605 205.175 ;
        RECT 31.275 205.005 31.445 205.195 ;
        RECT 34.955 204.985 35.125 205.175 ;
        RECT 35.930 205.035 36.050 205.145 ;
        RECT 36.795 205.005 36.965 205.195 ;
        RECT 38.635 204.985 38.805 205.175 ;
        RECT 42.315 205.005 42.485 205.195 ;
        RECT 44.155 204.985 44.325 205.175 ;
        RECT 47.835 205.005 48.005 205.195 ;
        RECT 48.810 205.035 48.930 205.145 ;
        RECT 49.675 204.985 49.845 205.175 ;
        RECT 51.515 205.005 51.685 205.195 ;
        RECT 55.195 204.985 55.365 205.175 ;
        RECT 57.035 205.005 57.205 205.195 ;
        RECT 60.715 204.985 60.885 205.175 ;
        RECT 61.690 205.035 61.810 205.145 ;
        RECT 62.555 205.005 62.725 205.195 ;
        RECT 64.395 204.985 64.565 205.175 ;
        RECT 68.075 205.005 68.245 205.195 ;
        RECT 69.915 204.985 70.085 205.175 ;
        RECT 73.595 205.005 73.765 205.195 ;
        RECT 74.570 205.035 74.690 205.145 ;
        RECT 75.435 204.985 75.605 205.175 ;
        RECT 77.275 205.005 77.445 205.195 ;
        RECT 80.955 204.985 81.125 205.175 ;
        RECT 82.795 205.005 82.965 205.195 ;
        RECT 86.475 204.985 86.645 205.175 ;
        RECT 87.450 205.035 87.570 205.145 ;
        RECT 88.315 205.005 88.485 205.195 ;
        RECT 90.155 204.985 90.325 205.175 ;
        RECT 93.835 205.005 94.005 205.195 ;
        RECT 95.675 204.985 95.845 205.175 ;
        RECT 99.355 205.005 99.525 205.195 ;
        RECT 100.330 205.035 100.450 205.145 ;
        RECT 101.195 204.985 101.365 205.175 ;
        RECT 102.115 205.005 102.285 205.195 ;
        RECT 106.715 204.985 106.885 205.175 ;
        RECT 107.635 205.005 107.805 205.195 ;
        RECT 112.235 204.985 112.405 205.175 ;
        RECT 113.155 205.145 113.325 205.195 ;
        RECT 113.155 205.035 113.330 205.145 ;
        RECT 113.155 205.005 113.325 205.035 ;
        RECT 118.675 204.985 118.845 205.195 ;
        RECT 124.195 204.985 124.365 205.195 ;
        RECT 125.575 204.985 125.745 205.195 ;
        RECT 11.815 204.175 13.185 204.985 ;
        RECT 13.195 204.175 18.705 204.985 ;
        RECT 18.715 204.175 24.225 204.985 ;
        RECT 24.235 204.175 29.745 204.985 ;
        RECT 29.755 204.175 35.265 204.985 ;
        RECT 35.285 204.115 35.715 204.900 ;
        RECT 36.195 204.175 38.945 204.985 ;
        RECT 38.955 204.175 44.465 204.985 ;
        RECT 44.475 204.175 49.985 204.985 ;
        RECT 49.995 204.175 55.505 204.985 ;
        RECT 55.515 204.175 61.025 204.985 ;
        RECT 61.045 204.115 61.475 204.900 ;
        RECT 61.955 204.175 64.705 204.985 ;
        RECT 64.715 204.175 70.225 204.985 ;
        RECT 70.235 204.175 75.745 204.985 ;
        RECT 75.755 204.175 81.265 204.985 ;
        RECT 81.275 204.175 86.785 204.985 ;
        RECT 86.805 204.115 87.235 204.900 ;
        RECT 87.715 204.175 90.465 204.985 ;
        RECT 90.475 204.175 95.985 204.985 ;
        RECT 95.995 204.175 101.505 204.985 ;
        RECT 101.515 204.175 107.025 204.985 ;
        RECT 107.035 204.175 112.545 204.985 ;
        RECT 112.565 204.115 112.995 204.900 ;
        RECT 113.475 204.175 118.985 204.985 ;
        RECT 118.995 204.175 124.505 204.985 ;
        RECT 124.515 204.175 125.885 204.985 ;
      LAYER nwell ;
        RECT 11.620 200.955 126.080 203.785 ;
      LAYER pwell ;
        RECT 11.815 199.755 13.185 200.565 ;
        RECT 13.195 199.755 16.865 200.565 ;
        RECT 16.875 199.755 22.385 200.565 ;
        RECT 22.405 199.840 22.835 200.625 ;
        RECT 23.315 199.755 26.065 200.565 ;
        RECT 26.075 199.755 31.585 200.565 ;
        RECT 31.595 199.755 37.105 200.565 ;
        RECT 37.115 199.755 42.625 200.565 ;
        RECT 42.635 199.755 48.145 200.565 ;
        RECT 48.165 199.840 48.595 200.625 ;
        RECT 49.075 199.755 51.825 200.565 ;
        RECT 51.835 199.755 57.345 200.565 ;
        RECT 57.355 199.755 62.865 200.565 ;
        RECT 62.875 199.755 68.385 200.565 ;
        RECT 68.395 199.755 73.905 200.565 ;
        RECT 73.925 199.840 74.355 200.625 ;
        RECT 74.835 199.755 77.585 200.565 ;
        RECT 77.595 199.755 83.105 200.565 ;
        RECT 83.115 199.755 88.625 200.565 ;
        RECT 88.635 199.755 94.145 200.565 ;
        RECT 94.155 199.755 99.665 200.565 ;
        RECT 99.685 199.840 100.115 200.625 ;
        RECT 100.595 199.755 102.425 200.565 ;
        RECT 102.435 199.755 107.945 200.565 ;
        RECT 107.955 199.755 113.465 200.565 ;
        RECT 113.475 199.755 118.985 200.565 ;
        RECT 118.995 199.755 124.505 200.565 ;
        RECT 124.515 199.755 125.885 200.565 ;
        RECT 11.955 199.545 12.125 199.755 ;
        RECT 16.555 199.565 16.725 199.755 ;
        RECT 18.395 199.545 18.565 199.735 ;
        RECT 22.075 199.565 22.245 199.755 ;
        RECT 23.050 199.595 23.170 199.705 ;
        RECT 23.915 199.545 24.085 199.735 ;
        RECT 25.755 199.565 25.925 199.755 ;
        RECT 29.435 199.545 29.605 199.735 ;
        RECT 31.275 199.565 31.445 199.755 ;
        RECT 34.955 199.545 35.125 199.735 ;
        RECT 35.930 199.595 36.050 199.705 ;
        RECT 36.795 199.565 36.965 199.755 ;
        RECT 38.635 199.545 38.805 199.735 ;
        RECT 42.315 199.565 42.485 199.755 ;
        RECT 44.155 199.545 44.325 199.735 ;
        RECT 47.835 199.565 48.005 199.755 ;
        RECT 48.810 199.595 48.930 199.705 ;
        RECT 49.675 199.545 49.845 199.735 ;
        RECT 51.515 199.565 51.685 199.755 ;
        RECT 55.195 199.545 55.365 199.735 ;
        RECT 57.035 199.565 57.205 199.755 ;
        RECT 60.715 199.545 60.885 199.735 ;
        RECT 62.555 199.545 62.725 199.755 ;
        RECT 68.075 199.565 68.245 199.755 ;
        RECT 71.755 199.545 71.925 199.735 ;
        RECT 73.595 199.565 73.765 199.755 ;
        RECT 74.570 199.595 74.690 199.705 ;
        RECT 75.435 199.545 75.605 199.735 ;
        RECT 77.275 199.565 77.445 199.755 ;
        RECT 80.955 199.545 81.125 199.735 ;
        RECT 82.795 199.565 82.965 199.755 ;
        RECT 86.475 199.545 86.645 199.735 ;
        RECT 87.450 199.595 87.570 199.705 ;
        RECT 88.315 199.565 88.485 199.755 ;
        RECT 90.155 199.545 90.325 199.735 ;
        RECT 93.835 199.565 94.005 199.755 ;
        RECT 95.675 199.545 95.845 199.735 ;
        RECT 99.355 199.565 99.525 199.755 ;
        RECT 100.330 199.595 100.450 199.705 ;
        RECT 101.195 199.545 101.365 199.735 ;
        RECT 102.115 199.565 102.285 199.755 ;
        RECT 106.715 199.545 106.885 199.735 ;
        RECT 107.635 199.565 107.805 199.755 ;
        RECT 112.235 199.545 112.405 199.735 ;
        RECT 113.155 199.705 113.325 199.755 ;
        RECT 113.155 199.595 113.330 199.705 ;
        RECT 113.155 199.565 113.325 199.595 ;
        RECT 118.675 199.545 118.845 199.755 ;
        RECT 124.195 199.545 124.365 199.755 ;
        RECT 125.575 199.545 125.745 199.755 ;
        RECT 11.815 198.735 13.185 199.545 ;
        RECT 13.195 198.735 18.705 199.545 ;
        RECT 18.715 198.735 24.225 199.545 ;
        RECT 24.235 198.735 29.745 199.545 ;
        RECT 29.755 198.735 35.265 199.545 ;
        RECT 35.285 198.675 35.715 199.460 ;
        RECT 36.195 198.735 38.945 199.545 ;
        RECT 38.955 198.735 44.465 199.545 ;
        RECT 44.475 198.735 49.985 199.545 ;
        RECT 49.995 198.735 55.505 199.545 ;
        RECT 55.515 198.735 61.025 199.545 ;
        RECT 61.045 198.675 61.475 199.460 ;
        RECT 61.495 198.735 62.865 199.545 ;
        RECT 62.875 198.865 72.065 199.545 ;
        RECT 62.875 198.635 63.795 198.865 ;
        RECT 66.625 198.645 67.555 198.865 ;
        RECT 72.075 198.735 75.745 199.545 ;
        RECT 75.755 198.735 81.265 199.545 ;
        RECT 81.275 198.735 86.785 199.545 ;
        RECT 86.805 198.675 87.235 199.460 ;
        RECT 87.715 198.735 90.465 199.545 ;
        RECT 90.475 198.735 95.985 199.545 ;
        RECT 95.995 198.735 101.505 199.545 ;
        RECT 101.515 198.735 107.025 199.545 ;
        RECT 107.035 198.735 112.545 199.545 ;
        RECT 112.565 198.675 112.995 199.460 ;
        RECT 113.475 198.735 118.985 199.545 ;
        RECT 118.995 198.735 124.505 199.545 ;
        RECT 124.515 198.735 125.885 199.545 ;
      LAYER nwell ;
        RECT 11.620 195.515 126.080 198.345 ;
      LAYER pwell ;
        RECT 11.815 194.315 13.185 195.125 ;
        RECT 13.195 194.315 16.865 195.125 ;
        RECT 16.875 194.315 22.385 195.125 ;
        RECT 22.405 194.400 22.835 195.185 ;
        RECT 23.315 194.315 26.065 195.125 ;
        RECT 26.075 194.315 31.585 195.125 ;
        RECT 31.595 194.315 37.105 195.125 ;
        RECT 37.115 194.315 42.625 195.125 ;
        RECT 42.635 194.315 48.145 195.125 ;
        RECT 48.165 194.400 48.595 195.185 ;
        RECT 49.075 194.315 52.745 195.125 ;
        RECT 52.755 194.315 58.265 195.125 ;
        RECT 62.785 194.995 63.715 195.215 ;
        RECT 66.435 194.995 68.645 195.225 ;
        RECT 58.275 194.315 68.645 194.995 ;
        RECT 68.865 194.315 70.215 195.225 ;
        RECT 70.235 194.315 73.905 195.125 ;
        RECT 73.925 194.400 74.355 195.185 ;
        RECT 74.385 194.315 75.735 195.225 ;
        RECT 75.755 194.995 76.675 195.225 ;
        RECT 79.505 194.995 80.435 195.215 ;
        RECT 75.755 194.315 84.945 194.995 ;
        RECT 84.955 194.315 88.625 195.125 ;
        RECT 88.635 194.315 94.145 195.125 ;
        RECT 94.155 194.315 99.665 195.125 ;
        RECT 99.685 194.400 100.115 195.185 ;
        RECT 100.595 194.315 102.425 195.125 ;
        RECT 102.435 194.315 107.945 195.125 ;
        RECT 107.955 194.315 113.465 195.125 ;
        RECT 113.475 194.315 118.985 195.125 ;
        RECT 118.995 194.315 124.505 195.125 ;
        RECT 124.515 194.315 125.885 195.125 ;
        RECT 11.955 194.105 12.125 194.315 ;
        RECT 16.555 194.125 16.725 194.315 ;
        RECT 18.395 194.105 18.565 194.295 ;
        RECT 22.075 194.125 22.245 194.315 ;
        RECT 23.050 194.155 23.170 194.265 ;
        RECT 23.915 194.105 24.085 194.295 ;
        RECT 25.755 194.125 25.925 194.315 ;
        RECT 29.435 194.105 29.605 194.295 ;
        RECT 31.275 194.125 31.445 194.315 ;
        RECT 34.955 194.105 35.125 194.295 ;
        RECT 35.930 194.155 36.050 194.265 ;
        RECT 36.795 194.125 36.965 194.315 ;
        RECT 38.635 194.105 38.805 194.295 ;
        RECT 42.315 194.125 42.485 194.315 ;
        RECT 44.155 194.105 44.325 194.295 ;
        RECT 47.835 194.125 48.005 194.315 ;
        RECT 48.810 194.155 48.930 194.265 ;
        RECT 49.675 194.105 49.845 194.295 ;
        RECT 52.435 194.125 52.605 194.315 ;
        RECT 55.195 194.105 55.365 194.295 ;
        RECT 57.955 194.125 58.125 194.315 ;
        RECT 58.415 194.125 58.585 194.315 ;
        RECT 60.715 194.105 60.885 194.295 ;
        RECT 63.015 194.105 63.185 194.295 ;
        RECT 63.475 194.105 63.645 194.295 ;
        RECT 65.315 194.150 65.475 194.260 ;
        RECT 65.775 194.105 65.945 194.295 ;
        RECT 67.620 194.105 67.790 194.295 ;
        RECT 69.915 194.125 70.085 194.315 ;
        RECT 71.295 194.150 71.455 194.260 ;
        RECT 73.595 194.125 73.765 194.315 ;
        RECT 74.515 194.105 74.685 194.315 ;
        RECT 83.715 194.105 83.885 194.295 ;
        RECT 84.635 194.125 84.805 194.315 ;
        RECT 85.095 194.105 85.265 194.295 ;
        RECT 86.475 194.105 86.645 194.295 ;
        RECT 88.315 194.125 88.485 194.315 ;
        RECT 90.615 194.105 90.785 194.295 ;
        RECT 93.835 194.125 94.005 194.315 ;
        RECT 96.135 194.105 96.305 194.295 ;
        RECT 99.355 194.125 99.525 194.315 ;
        RECT 100.330 194.155 100.450 194.265 ;
        RECT 102.115 194.125 102.285 194.315 ;
        RECT 105.335 194.105 105.505 194.295 ;
        RECT 105.795 194.105 105.965 194.295 ;
        RECT 107.230 194.155 107.350 194.265 ;
        RECT 107.635 194.105 107.805 194.315 ;
        RECT 112.235 194.105 112.405 194.295 ;
        RECT 113.155 194.265 113.325 194.315 ;
        RECT 113.155 194.155 113.330 194.265 ;
        RECT 113.155 194.125 113.325 194.155 ;
        RECT 118.675 194.105 118.845 194.315 ;
        RECT 124.195 194.105 124.365 194.315 ;
        RECT 125.575 194.105 125.745 194.315 ;
        RECT 11.815 193.295 13.185 194.105 ;
        RECT 13.195 193.295 18.705 194.105 ;
        RECT 18.715 193.295 24.225 194.105 ;
        RECT 24.235 193.295 29.745 194.105 ;
        RECT 29.755 193.295 35.265 194.105 ;
        RECT 35.285 193.235 35.715 194.020 ;
        RECT 36.195 193.295 38.945 194.105 ;
        RECT 38.955 193.295 44.465 194.105 ;
        RECT 44.475 193.295 49.985 194.105 ;
        RECT 49.995 193.295 55.505 194.105 ;
        RECT 55.515 193.295 61.025 194.105 ;
        RECT 61.045 193.235 61.475 194.020 ;
        RECT 61.495 193.295 63.325 194.105 ;
        RECT 63.345 193.195 64.695 194.105 ;
        RECT 65.635 193.425 67.465 194.105 ;
        RECT 66.120 193.195 67.465 193.425 ;
        RECT 67.475 193.195 70.395 194.105 ;
        RECT 71.615 193.195 74.725 194.105 ;
        RECT 74.835 193.425 84.025 194.105 ;
        RECT 74.835 193.195 75.755 193.425 ;
        RECT 78.585 193.205 79.515 193.425 ;
        RECT 84.045 193.195 85.395 194.105 ;
        RECT 85.415 193.295 86.785 194.105 ;
        RECT 86.805 193.235 87.235 194.020 ;
        RECT 87.255 193.295 90.925 194.105 ;
        RECT 90.935 193.295 96.445 194.105 ;
        RECT 96.455 193.425 105.645 194.105 ;
        RECT 96.455 193.195 97.375 193.425 ;
        RECT 100.205 193.205 101.135 193.425 ;
        RECT 105.665 193.195 107.015 194.105 ;
        RECT 107.495 193.325 108.865 194.105 ;
        RECT 108.875 193.295 112.545 194.105 ;
        RECT 112.565 193.235 112.995 194.020 ;
        RECT 113.475 193.295 118.985 194.105 ;
        RECT 118.995 193.295 124.505 194.105 ;
        RECT 124.515 193.295 125.885 194.105 ;
      LAYER nwell ;
        RECT 11.620 190.075 126.080 192.905 ;
      LAYER pwell ;
        RECT 11.815 188.875 13.185 189.685 ;
        RECT 13.195 188.875 16.865 189.685 ;
        RECT 16.875 188.875 22.385 189.685 ;
        RECT 22.405 188.960 22.835 189.745 ;
        RECT 23.315 188.875 26.065 189.685 ;
        RECT 26.075 188.875 31.585 189.685 ;
        RECT 31.595 188.875 37.105 189.685 ;
        RECT 37.115 188.875 42.625 189.685 ;
        RECT 42.635 188.875 48.145 189.685 ;
        RECT 48.165 188.960 48.595 189.745 ;
        RECT 49.075 188.875 52.745 189.685 ;
        RECT 52.755 188.875 58.265 189.685 ;
        RECT 58.275 188.875 63.785 189.685 ;
        RECT 68.375 189.555 69.305 189.785 ;
        RECT 70.895 189.555 73.895 189.785 ;
        RECT 63.795 188.875 65.625 189.555 ;
        RECT 65.635 188.875 69.305 189.555 ;
        RECT 69.315 189.465 73.895 189.555 ;
        RECT 69.315 189.105 73.905 189.465 ;
        RECT 69.315 188.875 70.885 189.105 ;
        RECT 72.975 188.915 73.905 189.105 ;
        RECT 73.925 188.960 74.355 189.745 ;
        RECT 74.685 189.555 75.615 189.785 ;
        RECT 72.975 188.875 73.895 188.915 ;
        RECT 74.685 188.875 76.520 189.555 ;
        RECT 76.675 188.875 78.505 189.555 ;
        RECT 78.985 188.875 80.335 189.785 ;
        RECT 80.355 188.875 81.725 189.655 ;
        RECT 81.735 188.875 84.485 189.685 ;
        RECT 84.495 188.875 90.005 189.685 ;
        RECT 90.025 188.875 91.375 189.785 ;
        RECT 92.315 188.875 93.685 189.655 ;
        RECT 94.615 188.875 98.285 189.685 ;
        RECT 98.305 188.875 99.655 189.785 ;
        RECT 99.685 188.960 100.115 189.745 ;
        RECT 100.595 188.875 102.425 189.685 ;
        RECT 102.435 189.555 103.355 189.785 ;
        RECT 106.185 189.555 107.115 189.775 ;
        RECT 102.435 188.875 111.625 189.555 ;
        RECT 111.635 188.875 113.465 189.685 ;
        RECT 113.475 188.875 118.985 189.685 ;
        RECT 118.995 188.875 124.505 189.685 ;
        RECT 124.515 188.875 125.885 189.685 ;
        RECT 11.955 188.665 12.125 188.875 ;
        RECT 16.555 188.685 16.725 188.875 ;
        RECT 18.395 188.665 18.565 188.855 ;
        RECT 22.075 188.685 22.245 188.875 ;
        RECT 23.050 188.715 23.170 188.825 ;
        RECT 23.915 188.665 24.085 188.855 ;
        RECT 25.755 188.685 25.925 188.875 ;
        RECT 29.435 188.665 29.605 188.855 ;
        RECT 31.275 188.685 31.445 188.875 ;
        RECT 34.955 188.665 35.125 188.855 ;
        RECT 36.795 188.685 36.965 188.875 ;
        RECT 38.175 188.665 38.345 188.855 ;
        RECT 38.635 188.665 38.805 188.855 ;
        RECT 42.315 188.685 42.485 188.875 ;
        RECT 47.835 188.685 48.005 188.875 ;
        RECT 48.755 188.825 48.925 188.855 ;
        RECT 48.755 188.715 48.930 188.825 ;
        RECT 48.755 188.665 48.925 188.715 ;
        RECT 50.135 188.665 50.305 188.855 ;
        RECT 50.595 188.665 50.765 188.855 ;
        RECT 52.030 188.715 52.150 188.825 ;
        RECT 52.435 188.665 52.605 188.875 ;
        RECT 54.735 188.665 54.905 188.855 ;
        RECT 55.250 188.715 55.370 188.825 ;
        RECT 57.955 188.685 58.125 188.875 ;
        RECT 60.715 188.665 60.885 188.855 ;
        RECT 63.475 188.685 63.645 188.875 ;
        RECT 63.935 188.685 64.105 188.875 ;
        RECT 64.855 188.665 65.025 188.855 ;
        RECT 65.775 188.685 65.945 188.875 ;
        RECT 66.235 188.665 66.405 188.855 ;
        RECT 68.535 188.665 68.705 188.855 ;
        RECT 11.815 187.855 13.185 188.665 ;
        RECT 13.195 187.855 18.705 188.665 ;
        RECT 18.715 187.855 24.225 188.665 ;
        RECT 24.235 187.855 29.745 188.665 ;
        RECT 29.755 187.855 35.265 188.665 ;
        RECT 35.285 187.795 35.715 188.580 ;
        RECT 35.735 187.855 38.485 188.665 ;
        RECT 38.505 187.755 39.855 188.665 ;
        RECT 39.875 187.985 49.065 188.665 ;
        RECT 39.875 187.755 40.795 187.985 ;
        RECT 43.625 187.765 44.555 187.985 ;
        RECT 49.075 187.855 50.445 188.665 ;
        RECT 50.465 187.755 51.815 188.665 ;
        RECT 52.295 187.885 53.665 188.665 ;
        RECT 53.685 187.755 55.035 188.665 ;
        RECT 55.515 187.855 61.025 188.665 ;
        RECT 61.045 187.795 61.475 188.580 ;
        RECT 61.495 187.855 65.165 188.665 ;
        RECT 65.175 187.885 66.545 188.665 ;
        RECT 66.555 187.985 68.845 188.665 ;
        RECT 68.995 188.635 69.165 188.855 ;
        RECT 69.455 188.685 69.625 188.875 ;
        RECT 76.355 188.855 76.520 188.875 ;
        RECT 72.675 188.710 72.835 188.820 ;
        RECT 73.135 188.665 73.305 188.855 ;
        RECT 76.355 188.685 76.530 188.855 ;
        RECT 76.815 188.685 76.985 188.875 ;
        RECT 77.275 188.710 77.435 188.820 ;
        RECT 78.710 188.715 78.830 188.825 ;
        RECT 79.115 188.685 79.285 188.875 ;
        RECT 80.495 188.685 80.665 188.875 ;
        RECT 76.360 188.665 76.530 188.685 ;
        RECT 80.955 188.665 81.125 188.855 ;
        RECT 84.175 188.685 84.345 188.875 ;
        RECT 86.475 188.665 86.645 188.855 ;
        RECT 89.695 188.685 89.865 188.875 ;
        RECT 91.075 188.685 91.245 188.875 ;
        RECT 91.995 188.720 92.155 188.830 ;
        RECT 92.455 188.685 92.625 188.875 ;
        RECT 94.295 188.720 94.455 188.830 ;
        RECT 96.135 188.665 96.305 188.855 ;
        RECT 97.975 188.665 98.145 188.875 ;
        RECT 98.435 188.685 98.605 188.875 ;
        RECT 100.330 188.715 100.450 188.825 ;
        RECT 101.840 188.665 102.010 188.855 ;
        RECT 102.115 188.685 102.285 188.875 ;
        RECT 105.980 188.665 106.150 188.855 ;
        RECT 106.770 188.715 106.890 188.825 ;
        RECT 109.475 188.665 109.645 188.855 ;
        RECT 109.935 188.665 110.105 188.855 ;
        RECT 111.315 188.685 111.485 188.875 ;
        RECT 112.235 188.665 112.405 188.855 ;
        RECT 113.155 188.825 113.325 188.875 ;
        RECT 113.155 188.715 113.330 188.825 ;
        RECT 113.155 188.685 113.325 188.715 ;
        RECT 118.675 188.665 118.845 188.875 ;
        RECT 124.195 188.665 124.365 188.875 ;
        RECT 125.575 188.665 125.745 188.875 ;
        RECT 71.120 188.635 72.065 188.665 ;
        RECT 68.995 188.435 72.065 188.635 ;
        RECT 66.555 187.755 67.475 187.985 ;
        RECT 68.855 187.955 72.065 188.435 ;
        RECT 72.995 187.985 75.285 188.665 ;
        RECT 68.855 187.755 69.785 187.955 ;
        RECT 71.120 187.755 72.065 187.955 ;
        RECT 74.365 187.755 75.285 187.985 ;
        RECT 75.295 187.755 76.645 188.665 ;
        RECT 77.595 187.855 81.265 188.665 ;
        RECT 81.275 187.855 86.785 188.665 ;
        RECT 86.805 187.795 87.235 188.580 ;
        RECT 87.255 187.985 96.445 188.665 ;
        RECT 87.255 187.755 88.175 187.985 ;
        RECT 91.005 187.765 91.935 187.985 ;
        RECT 96.455 187.855 98.285 188.665 ;
        RECT 98.525 187.985 102.425 188.665 ;
        RECT 102.665 187.985 106.565 188.665 ;
        RECT 101.495 187.755 102.425 187.985 ;
        RECT 105.635 187.755 106.565 187.985 ;
        RECT 107.035 187.855 109.785 188.665 ;
        RECT 109.795 187.885 111.165 188.665 ;
        RECT 111.175 187.855 112.545 188.665 ;
        RECT 112.565 187.795 112.995 188.580 ;
        RECT 113.475 187.855 118.985 188.665 ;
        RECT 118.995 187.855 124.505 188.665 ;
        RECT 124.515 187.855 125.885 188.665 ;
      LAYER nwell ;
        RECT 11.620 184.635 126.080 187.465 ;
      LAYER pwell ;
        RECT 11.815 183.435 13.185 184.245 ;
        RECT 13.195 183.435 16.865 184.245 ;
        RECT 16.875 183.435 22.385 184.245 ;
        RECT 22.405 183.520 22.835 184.305 ;
        RECT 23.315 183.435 26.985 184.245 ;
        RECT 26.995 183.435 32.505 184.245 ;
        RECT 32.525 183.435 33.875 184.345 ;
        RECT 38.405 184.115 39.335 184.335 ;
        RECT 42.165 184.115 43.085 184.345 ;
        RECT 33.895 183.435 43.085 184.115 ;
        RECT 44.015 184.115 44.945 184.345 ;
        RECT 44.015 183.435 47.915 184.115 ;
        RECT 48.165 183.520 48.595 184.305 ;
        RECT 48.615 184.115 49.535 184.345 ;
        RECT 52.365 184.115 53.295 184.335 ;
        RECT 48.615 183.435 57.805 184.115 ;
        RECT 58.275 183.435 61.945 184.245 ;
        RECT 61.965 183.435 63.315 184.345 ;
        RECT 65.990 184.115 66.910 184.345 ;
        RECT 63.445 183.435 66.910 184.115 ;
        RECT 67.935 184.145 68.865 184.345 ;
        RECT 70.200 184.145 71.145 184.345 ;
        RECT 67.935 183.665 71.145 184.145 ;
        RECT 68.075 183.465 71.145 183.665 ;
        RECT 11.955 183.225 12.125 183.435 ;
        RECT 16.555 183.245 16.725 183.435 ;
        RECT 18.395 183.225 18.565 183.415 ;
        RECT 22.075 183.245 22.245 183.435 ;
        RECT 23.050 183.275 23.170 183.385 ;
        RECT 23.915 183.225 24.085 183.415 ;
        RECT 26.675 183.245 26.845 183.435 ;
        RECT 29.435 183.225 29.605 183.415 ;
        RECT 32.195 183.245 32.365 183.435 ;
        RECT 32.655 183.245 32.825 183.435 ;
        RECT 34.035 183.245 34.205 183.435 ;
        RECT 34.955 183.225 35.125 183.415 ;
        RECT 39.095 183.225 39.265 183.415 ;
        RECT 40.475 183.225 40.645 183.415 ;
        RECT 41.210 183.225 41.380 183.415 ;
        RECT 43.695 183.280 43.855 183.390 ;
        RECT 44.430 183.245 44.600 183.435 ;
        RECT 45.130 183.275 45.250 183.385 ;
        RECT 45.535 183.225 45.705 183.415 ;
        RECT 50.320 183.225 50.490 183.415 ;
        RECT 57.495 183.245 57.665 183.435 ;
        RECT 58.010 183.275 58.130 183.385 ;
        RECT 59.795 183.225 59.965 183.415 ;
        RECT 60.715 183.270 60.875 183.380 ;
        RECT 61.635 183.245 61.805 183.435 ;
        RECT 63.015 183.245 63.185 183.435 ;
        RECT 63.475 183.245 63.645 183.435 ;
        RECT 67.615 183.280 67.775 183.390 ;
        RECT 68.075 183.245 68.245 183.465 ;
        RECT 70.200 183.435 71.145 183.465 ;
        RECT 71.155 183.435 73.445 184.345 ;
        RECT 73.925 183.520 74.355 184.305 ;
        RECT 74.835 183.435 76.665 184.245 ;
        RECT 76.675 183.435 82.185 184.245 ;
        RECT 82.205 183.435 83.555 184.345 ;
        RECT 84.045 183.435 85.395 184.345 ;
        RECT 85.415 183.435 88.165 184.245 ;
        RECT 91.375 184.115 92.305 184.345 ;
        RECT 88.405 183.435 92.305 184.115 ;
        RECT 92.315 183.435 94.145 184.245 ;
        RECT 94.155 183.435 99.665 184.245 ;
        RECT 99.685 183.520 100.115 184.305 ;
        RECT 100.595 183.435 102.425 184.245 ;
        RECT 102.435 183.435 103.805 184.215 ;
        RECT 103.825 183.435 105.175 184.345 ;
        RECT 105.195 184.115 106.115 184.345 ;
        RECT 108.945 184.115 109.875 184.335 ;
        RECT 105.195 183.435 114.385 184.115 ;
        RECT 115.315 183.435 118.985 184.245 ;
        RECT 118.995 183.435 124.505 184.245 ;
        RECT 124.515 183.435 125.885 184.245 ;
        RECT 70.375 183.225 70.545 183.415 ;
        RECT 73.130 183.245 73.300 183.435 ;
        RECT 73.595 183.385 73.765 183.415 ;
        RECT 73.595 183.275 73.770 183.385 ;
        RECT 74.110 183.275 74.230 183.385 ;
        RECT 74.570 183.275 74.690 183.385 ;
        RECT 73.595 183.225 73.765 183.275 ;
        RECT 76.355 183.245 76.525 183.435 ;
        RECT 76.815 183.225 76.985 183.415 ;
        RECT 81.875 183.245 82.045 183.435 ;
        RECT 83.255 183.245 83.425 183.435 ;
        RECT 83.770 183.275 83.890 183.385 ;
        RECT 85.095 183.245 85.265 183.435 ;
        RECT 86.475 183.225 86.645 183.415 ;
        RECT 87.855 183.245 88.025 183.435 ;
        RECT 88.315 183.225 88.485 183.415 ;
        RECT 88.830 183.275 88.950 183.385 ;
        RECT 91.535 183.225 91.705 183.415 ;
        RECT 91.720 183.245 91.890 183.435 ;
        RECT 93.835 183.245 94.005 183.435 ;
        RECT 97.055 183.225 97.225 183.415 ;
        RECT 98.435 183.225 98.605 183.415 ;
        RECT 98.950 183.275 99.070 183.385 ;
        RECT 99.355 183.245 99.525 183.435 ;
        RECT 100.330 183.275 100.450 183.385 ;
        RECT 101.655 183.225 101.825 183.415 ;
        RECT 102.115 183.225 102.285 183.435 ;
        RECT 102.575 183.245 102.745 183.435 ;
        RECT 103.955 183.245 104.125 183.435 ;
        RECT 106.900 183.225 107.070 183.415 ;
        RECT 111.040 183.225 111.210 183.415 ;
        RECT 112.235 183.270 112.395 183.380 ;
        RECT 113.210 183.275 113.330 183.385 ;
        RECT 114.075 183.245 114.245 183.435 ;
        RECT 114.995 183.280 115.155 183.390 ;
        RECT 118.675 183.225 118.845 183.435 ;
        RECT 124.195 183.225 124.365 183.435 ;
        RECT 125.575 183.225 125.745 183.435 ;
        RECT 11.815 182.415 13.185 183.225 ;
        RECT 13.195 182.415 18.705 183.225 ;
        RECT 18.715 182.415 24.225 183.225 ;
        RECT 24.235 182.415 29.745 183.225 ;
        RECT 29.755 182.415 35.265 183.225 ;
        RECT 35.285 182.355 35.715 183.140 ;
        RECT 35.735 182.415 39.405 183.225 ;
        RECT 39.415 182.445 40.785 183.225 ;
        RECT 40.795 182.545 44.695 183.225 ;
        RECT 40.795 182.315 41.725 182.545 ;
        RECT 45.395 182.445 46.765 183.225 ;
        RECT 47.005 182.545 50.905 183.225 ;
        RECT 49.975 182.315 50.905 182.545 ;
        RECT 50.915 182.545 60.105 183.225 ;
        RECT 50.915 182.315 51.835 182.545 ;
        RECT 54.665 182.325 55.595 182.545 ;
        RECT 61.045 182.355 61.475 183.140 ;
        RECT 61.495 182.545 70.685 183.225 ;
        RECT 61.495 182.315 62.415 182.545 ;
        RECT 65.245 182.325 66.175 182.545 ;
        RECT 70.695 182.315 73.805 183.225 ;
        RECT 74.375 182.415 77.125 183.225 ;
        RECT 77.505 182.545 86.785 183.225 ;
        RECT 77.505 182.425 79.840 182.545 ;
        RECT 77.505 182.315 78.425 182.425 ;
        RECT 84.505 182.325 85.425 182.545 ;
        RECT 86.805 182.355 87.235 183.140 ;
        RECT 87.255 182.445 88.625 183.225 ;
        RECT 89.095 182.415 91.845 183.225 ;
        RECT 91.855 182.415 97.365 183.225 ;
        RECT 97.385 182.315 98.735 183.225 ;
        RECT 99.215 182.415 101.965 183.225 ;
        RECT 101.985 182.315 103.335 183.225 ;
        RECT 103.585 182.545 107.485 183.225 ;
        RECT 107.725 182.545 111.625 183.225 ;
        RECT 106.555 182.315 107.485 182.545 ;
        RECT 110.695 182.315 111.625 182.545 ;
        RECT 112.565 182.355 112.995 183.140 ;
        RECT 113.475 182.415 118.985 183.225 ;
        RECT 118.995 182.415 124.505 183.225 ;
        RECT 124.515 182.415 125.885 183.225 ;
      LAYER nwell ;
        RECT 11.620 179.195 126.080 182.025 ;
      LAYER pwell ;
        RECT 11.815 177.995 13.185 178.805 ;
        RECT 13.195 177.995 16.865 178.805 ;
        RECT 16.875 177.995 22.385 178.805 ;
        RECT 22.405 178.080 22.835 178.865 ;
        RECT 22.855 177.995 24.225 178.805 ;
        RECT 24.235 177.995 27.905 178.805 ;
        RECT 27.915 177.995 33.425 178.805 ;
        RECT 33.435 177.995 38.945 178.805 ;
        RECT 41.610 178.675 42.530 178.905 ;
        RECT 45.835 178.675 46.765 178.905 ;
        RECT 39.065 177.995 42.530 178.675 ;
        RECT 42.865 177.995 46.765 178.675 ;
        RECT 46.775 177.995 48.145 178.805 ;
        RECT 48.165 178.080 48.595 178.865 ;
        RECT 49.075 177.995 51.825 178.805 ;
        RECT 55.035 178.675 55.965 178.905 ;
        RECT 52.065 177.995 55.965 178.675 ;
        RECT 56.435 177.995 57.805 178.775 ;
        RECT 57.815 177.995 60.565 178.805 ;
        RECT 60.575 177.995 66.085 178.805 ;
        RECT 66.095 177.995 68.705 178.905 ;
        RECT 68.855 177.995 70.225 178.805 ;
        RECT 70.235 177.995 73.905 178.805 ;
        RECT 73.925 178.080 74.355 178.865 ;
        RECT 77.575 178.675 78.505 178.905 ;
        RECT 74.605 177.995 78.505 178.675 ;
        RECT 78.885 178.795 79.805 178.905 ;
        RECT 78.885 178.675 81.220 178.795 ;
        RECT 85.885 178.675 86.805 178.895 ;
        RECT 78.885 177.995 88.165 178.675 ;
        RECT 88.635 177.995 90.465 178.805 ;
        RECT 94.985 178.675 95.915 178.895 ;
        RECT 98.745 178.675 99.665 178.905 ;
        RECT 90.475 177.995 99.665 178.675 ;
        RECT 99.685 178.080 100.115 178.865 ;
        RECT 100.595 177.995 103.345 178.805 ;
        RECT 103.355 178.675 104.275 178.905 ;
        RECT 107.105 178.675 108.035 178.895 ;
        RECT 103.355 177.995 112.545 178.675 ;
        RECT 113.475 177.995 118.985 178.805 ;
        RECT 118.995 177.995 124.505 178.805 ;
        RECT 124.515 177.995 125.885 178.805 ;
        RECT 11.955 177.785 12.125 177.995 ;
        RECT 13.390 177.835 13.510 177.945 ;
        RECT 16.555 177.805 16.725 177.995 ;
        RECT 18.855 177.785 19.025 177.975 ;
        RECT 22.075 177.805 22.245 177.995 ;
        RECT 23.915 177.805 24.085 177.995 ;
        RECT 24.375 177.785 24.545 177.975 ;
        RECT 27.595 177.805 27.765 177.995 ;
        RECT 29.895 177.785 30.065 177.975 ;
        RECT 30.355 177.785 30.525 177.975 ;
        RECT 33.115 177.805 33.285 177.995 ;
        RECT 34.955 177.785 35.125 177.975 ;
        RECT 35.930 177.835 36.050 177.945 ;
        RECT 37.715 177.785 37.885 177.975 ;
        RECT 38.175 177.785 38.345 177.975 ;
        RECT 38.635 177.805 38.805 177.995 ;
        RECT 39.095 177.805 39.265 177.995 ;
        RECT 46.180 177.805 46.350 177.995 ;
        RECT 47.835 177.805 48.005 177.995 ;
        RECT 48.295 177.785 48.465 177.975 ;
        RECT 48.810 177.835 48.930 177.945 ;
        RECT 49.675 177.785 49.845 177.975 ;
        RECT 51.515 177.805 51.685 177.995 ;
        RECT 55.195 177.785 55.365 177.975 ;
        RECT 55.380 177.805 55.550 177.995 ;
        RECT 56.170 177.835 56.290 177.945 ;
        RECT 56.575 177.785 56.745 177.995 ;
        RECT 57.090 177.835 57.210 177.945 ;
        RECT 60.255 177.805 60.425 177.995 ;
        RECT 60.715 177.785 60.885 177.975 ;
        RECT 63.935 177.785 64.105 177.975 ;
        RECT 65.775 177.805 65.945 177.995 ;
        RECT 66.240 177.805 66.410 177.995 ;
        RECT 69.455 177.785 69.625 177.975 ;
        RECT 69.915 177.805 70.085 177.995 ;
        RECT 73.595 177.805 73.765 177.995 ;
        RECT 70.015 177.785 70.085 177.805 ;
        RECT 74.055 177.785 74.225 177.975 ;
        RECT 74.520 177.785 74.690 177.975 ;
        RECT 77.920 177.805 78.090 177.995 ;
        RECT 80.680 177.785 80.850 177.975 ;
        RECT 84.820 177.785 84.990 177.975 ;
        RECT 85.555 177.785 85.725 177.975 ;
        RECT 87.855 177.805 88.025 177.995 ;
        RECT 88.315 177.945 88.485 177.975 ;
        RECT 88.315 177.835 88.490 177.945 ;
        RECT 88.315 177.785 88.485 177.835 ;
        RECT 88.775 177.785 88.945 177.975 ;
        RECT 90.155 177.805 90.325 177.995 ;
        RECT 90.615 177.805 90.785 177.995 ;
        RECT 98.895 177.785 99.065 177.975 ;
        RECT 100.330 177.835 100.450 177.945 ;
        RECT 102.760 177.785 102.930 177.975 ;
        RECT 103.035 177.805 103.205 177.995 ;
        RECT 106.715 177.785 106.885 177.975 ;
        RECT 108.095 177.785 108.265 177.975 ;
        RECT 108.555 177.785 108.725 177.975 ;
        RECT 110.855 177.785 111.025 177.975 ;
        RECT 111.315 177.785 111.485 177.975 ;
        RECT 112.235 177.805 112.405 177.995 ;
        RECT 113.155 177.840 113.315 177.950 ;
        RECT 113.615 177.830 113.775 177.940 ;
        RECT 118.675 177.805 118.845 177.995 ;
        RECT 122.815 177.785 122.985 177.975 ;
        RECT 124.195 177.785 124.365 177.995 ;
        RECT 125.575 177.785 125.745 177.995 ;
        RECT 11.815 176.975 13.185 177.785 ;
        RECT 13.655 176.975 19.165 177.785 ;
        RECT 19.175 176.975 24.685 177.785 ;
        RECT 24.695 176.975 30.205 177.785 ;
        RECT 30.225 176.875 31.575 177.785 ;
        RECT 31.595 176.975 35.265 177.785 ;
        RECT 35.285 176.915 35.715 177.700 ;
        RECT 36.195 176.975 38.025 177.785 ;
        RECT 38.045 176.875 39.395 177.785 ;
        RECT 39.415 177.105 48.605 177.785 ;
        RECT 39.415 176.875 40.335 177.105 ;
        RECT 43.165 176.885 44.095 177.105 ;
        RECT 48.615 176.975 49.985 177.785 ;
        RECT 49.995 176.975 55.505 177.785 ;
        RECT 55.525 176.875 56.875 177.785 ;
        RECT 57.355 176.975 61.025 177.785 ;
        RECT 61.045 176.915 61.475 177.700 ;
        RECT 61.495 176.975 64.245 177.785 ;
        RECT 64.255 176.975 69.765 177.785 ;
        RECT 70.015 177.555 72.285 177.785 ;
        RECT 70.015 176.875 72.770 177.555 ;
        RECT 72.995 176.975 74.365 177.785 ;
        RECT 74.375 176.875 76.985 177.785 ;
        RECT 77.365 177.105 81.265 177.785 ;
        RECT 81.505 177.105 85.405 177.785 ;
        RECT 80.335 176.875 81.265 177.105 ;
        RECT 84.475 176.875 85.405 177.105 ;
        RECT 85.415 177.005 86.785 177.785 ;
        RECT 86.805 176.915 87.235 177.700 ;
        RECT 87.255 176.975 88.625 177.785 ;
        RECT 88.645 176.875 89.995 177.785 ;
        RECT 90.015 177.105 99.205 177.785 ;
        RECT 99.445 177.105 103.345 177.785 ;
        RECT 90.015 176.875 90.935 177.105 ;
        RECT 93.765 176.885 94.695 177.105 ;
        RECT 102.415 176.875 103.345 177.105 ;
        RECT 103.450 177.105 106.915 177.785 ;
        RECT 103.450 176.875 104.370 177.105 ;
        RECT 107.035 176.975 108.405 177.785 ;
        RECT 108.415 177.005 109.785 177.785 ;
        RECT 109.795 176.975 111.165 177.785 ;
        RECT 111.185 176.875 112.535 177.785 ;
        RECT 112.565 176.915 112.995 177.700 ;
        RECT 113.935 177.105 123.125 177.785 ;
        RECT 113.935 176.875 114.855 177.105 ;
        RECT 117.685 176.885 118.615 177.105 ;
        RECT 123.135 176.975 124.505 177.785 ;
        RECT 124.515 176.975 125.885 177.785 ;
      LAYER nwell ;
        RECT 11.620 173.755 126.080 176.585 ;
      LAYER pwell ;
        RECT 11.815 172.555 13.185 173.365 ;
        RECT 13.195 172.555 16.865 173.365 ;
        RECT 16.875 172.555 22.385 173.365 ;
        RECT 22.405 172.640 22.835 173.425 ;
        RECT 23.785 172.555 25.135 173.465 ;
        RECT 25.165 172.555 26.515 173.465 ;
        RECT 26.535 172.555 27.905 173.335 ;
        RECT 27.915 173.235 28.835 173.465 ;
        RECT 31.665 173.235 32.595 173.455 ;
        RECT 27.915 172.555 37.105 173.235 ;
        RECT 37.115 172.555 38.485 173.335 ;
        RECT 38.495 172.555 40.325 173.365 ;
        RECT 40.335 172.555 45.845 173.365 ;
        RECT 45.855 172.555 47.225 173.335 ;
        RECT 48.165 172.640 48.595 173.425 ;
        RECT 48.615 172.555 50.445 173.365 ;
        RECT 50.465 172.555 51.815 173.465 ;
        RECT 52.205 173.355 53.125 173.465 ;
        RECT 52.205 173.235 54.540 173.355 ;
        RECT 59.205 173.235 60.125 173.455 ;
        RECT 52.205 172.555 61.485 173.235 ;
        RECT 62.415 172.555 66.085 173.365 ;
        RECT 66.335 172.785 69.090 173.465 ;
        RECT 70.895 173.235 73.895 173.465 ;
        RECT 69.315 173.145 73.895 173.235 ;
        RECT 69.315 172.785 73.905 173.145 ;
        RECT 66.335 172.555 68.605 172.785 ;
        RECT 69.315 172.555 70.885 172.785 ;
        RECT 72.975 172.595 73.905 172.785 ;
        RECT 73.925 172.640 74.355 173.425 ;
        RECT 74.615 172.785 77.370 173.465 ;
        RECT 72.975 172.555 73.895 172.595 ;
        RECT 74.615 172.555 76.885 172.785 ;
        RECT 78.065 172.555 79.415 173.465 ;
        RECT 79.435 173.235 80.355 173.465 ;
        RECT 83.185 173.235 84.115 173.455 ;
        RECT 79.435 172.555 88.625 173.235 ;
        RECT 89.095 172.555 92.765 173.365 ;
        RECT 95.975 173.235 96.905 173.465 ;
        RECT 93.005 172.555 96.905 173.235 ;
        RECT 96.915 172.555 98.285 173.335 ;
        RECT 98.295 172.555 99.665 173.365 ;
        RECT 99.685 172.640 100.115 173.425 ;
        RECT 100.595 172.555 103.345 173.365 ;
        RECT 103.355 172.555 104.725 173.335 ;
        RECT 105.655 172.555 111.165 173.365 ;
        RECT 111.185 172.555 112.535 173.465 ;
        RECT 112.555 173.235 113.475 173.465 ;
        RECT 116.305 173.235 117.235 173.455 ;
        RECT 112.555 172.555 121.745 173.235 ;
        RECT 121.755 172.555 123.585 173.235 ;
        RECT 124.515 172.555 125.885 173.365 ;
        RECT 11.955 172.345 12.125 172.555 ;
        RECT 13.390 172.395 13.510 172.505 ;
        RECT 16.555 172.365 16.725 172.555 ;
        RECT 17.015 172.345 17.185 172.535 ;
        RECT 22.075 172.365 22.245 172.555 ;
        RECT 23.455 172.400 23.615 172.510 ;
        RECT 23.915 172.365 24.085 172.555 ;
        RECT 25.295 172.365 25.465 172.555 ;
        RECT 26.675 172.345 26.845 172.555 ;
        RECT 27.190 172.395 27.310 172.505 ;
        RECT 27.595 172.345 27.765 172.535 ;
        RECT 34.680 172.345 34.850 172.535 ;
        RECT 36.795 172.365 36.965 172.555 ;
        RECT 38.175 172.365 38.345 172.555 ;
        RECT 40.015 172.365 40.185 172.555 ;
        RECT 44.615 172.345 44.785 172.535 ;
        RECT 45.535 172.365 45.705 172.555 ;
        RECT 45.995 172.365 46.165 172.555 ;
        RECT 47.835 172.400 47.995 172.510 ;
        RECT 50.135 172.365 50.305 172.555 ;
        RECT 51.515 172.365 51.685 172.555 ;
        RECT 55.195 172.345 55.365 172.535 ;
        RECT 59.060 172.345 59.230 172.535 ;
        RECT 60.715 172.345 60.885 172.535 ;
        RECT 61.175 172.365 61.345 172.555 ;
        RECT 62.095 172.400 62.255 172.510 ;
        RECT 63.935 172.345 64.105 172.535 ;
        RECT 64.855 172.390 65.015 172.500 ;
        RECT 65.775 172.365 65.945 172.555 ;
        RECT 66.335 172.535 66.405 172.555 ;
        RECT 66.235 172.365 66.405 172.535 ;
        RECT 68.535 172.345 68.705 172.535 ;
        RECT 68.995 172.345 69.165 172.535 ;
        RECT 69.455 172.365 69.625 172.555 ;
        RECT 74.615 172.535 74.685 172.555 ;
        RECT 73.135 172.365 73.305 172.535 ;
        RECT 73.135 172.345 73.205 172.365 ;
        RECT 73.595 172.345 73.765 172.535 ;
        RECT 74.515 172.365 74.685 172.535 ;
        RECT 76.410 172.395 76.530 172.505 ;
        RECT 77.790 172.395 77.910 172.505 ;
        RECT 78.195 172.365 78.365 172.555 ;
        RECT 79.115 172.345 79.285 172.535 ;
        RECT 84.635 172.345 84.805 172.535 ;
        RECT 85.095 172.345 85.265 172.535 ;
        RECT 86.530 172.395 86.650 172.505 ;
        RECT 88.315 172.345 88.485 172.555 ;
        RECT 88.830 172.395 88.950 172.505 ;
        RECT 90.615 172.345 90.785 172.535 ;
        RECT 92.455 172.365 92.625 172.555 ;
        RECT 94.290 172.345 94.460 172.535 ;
        RECT 95.675 172.345 95.845 172.535 ;
        RECT 96.320 172.365 96.490 172.555 ;
        RECT 97.055 172.365 97.225 172.555 ;
        RECT 99.355 172.345 99.525 172.555 ;
        RECT 100.330 172.395 100.450 172.505 ;
        RECT 100.735 172.345 100.905 172.535 ;
        RECT 103.035 172.365 103.205 172.555 ;
        RECT 103.495 172.345 103.665 172.535 ;
        RECT 103.960 172.345 104.130 172.535 ;
        RECT 104.415 172.365 104.585 172.555 ;
        RECT 105.335 172.400 105.495 172.510 ;
        RECT 108.095 172.390 108.255 172.500 ;
        RECT 110.855 172.365 111.025 172.555 ;
        RECT 111.315 172.365 111.485 172.555 ;
        RECT 111.960 172.345 112.130 172.535 ;
        RECT 116.560 172.345 116.730 172.535 ;
        RECT 117.295 172.345 117.465 172.535 ;
        RECT 118.730 172.395 118.850 172.505 ;
        RECT 119.135 172.345 119.305 172.535 ;
        RECT 120.570 172.395 120.690 172.505 ;
        RECT 121.435 172.365 121.605 172.555 ;
        RECT 123.275 172.365 123.445 172.555 ;
        RECT 124.195 172.345 124.365 172.535 ;
        RECT 125.575 172.345 125.745 172.555 ;
        RECT 11.815 171.535 13.185 172.345 ;
        RECT 13.655 171.535 17.325 172.345 ;
        RECT 17.705 171.665 26.985 172.345 ;
        RECT 27.565 171.665 31.030 172.345 ;
        RECT 31.365 171.665 35.265 172.345 ;
        RECT 17.705 171.545 20.040 171.665 ;
        RECT 17.705 171.435 18.625 171.545 ;
        RECT 24.705 171.445 25.625 171.665 ;
        RECT 30.110 171.435 31.030 171.665 ;
        RECT 34.335 171.435 35.265 171.665 ;
        RECT 35.285 171.475 35.715 172.260 ;
        RECT 35.735 171.665 44.925 172.345 ;
        RECT 46.225 171.665 55.505 172.345 ;
        RECT 55.745 171.665 59.645 172.345 ;
        RECT 35.735 171.435 36.655 171.665 ;
        RECT 39.485 171.445 40.415 171.665 ;
        RECT 46.225 171.545 48.560 171.665 ;
        RECT 46.225 171.435 47.145 171.545 ;
        RECT 53.225 171.445 54.145 171.665 ;
        RECT 58.715 171.435 59.645 171.665 ;
        RECT 59.655 171.565 61.025 172.345 ;
        RECT 61.045 171.475 61.475 172.260 ;
        RECT 61.505 171.665 64.245 172.345 ;
        RECT 65.175 171.535 68.845 172.345 ;
        RECT 68.865 171.435 70.215 172.345 ;
        RECT 70.935 172.115 73.205 172.345 ;
        RECT 70.450 171.435 73.205 172.115 ;
        RECT 73.455 171.665 76.195 172.345 ;
        RECT 76.675 171.535 79.425 172.345 ;
        RECT 79.435 171.535 84.945 172.345 ;
        RECT 84.955 171.565 86.325 172.345 ;
        RECT 86.805 171.475 87.235 172.260 ;
        RECT 87.265 171.435 88.615 172.345 ;
        RECT 89.095 171.535 90.925 172.345 ;
        RECT 91.130 171.435 94.605 172.345 ;
        RECT 94.615 171.535 95.985 172.345 ;
        RECT 95.995 171.535 99.665 172.345 ;
        RECT 99.675 171.565 101.045 172.345 ;
        RECT 101.055 171.535 103.805 172.345 ;
        RECT 103.815 171.435 107.290 172.345 ;
        RECT 108.645 171.665 112.545 172.345 ;
        RECT 111.615 171.435 112.545 171.665 ;
        RECT 112.565 171.475 112.995 172.260 ;
        RECT 113.245 171.665 117.145 172.345 ;
        RECT 116.215 171.435 117.145 171.665 ;
        RECT 117.155 171.565 118.525 172.345 ;
        RECT 118.995 171.565 120.365 172.345 ;
        RECT 120.835 171.535 124.505 172.345 ;
        RECT 124.515 171.535 125.885 172.345 ;
      LAYER nwell ;
        RECT 11.620 168.315 126.080 171.145 ;
      LAYER pwell ;
        RECT 11.815 167.115 13.185 167.925 ;
        RECT 13.195 167.115 16.865 167.925 ;
        RECT 16.885 167.115 18.235 168.025 ;
        RECT 21.455 167.795 22.385 168.025 ;
        RECT 18.485 167.115 22.385 167.795 ;
        RECT 22.405 167.200 22.835 167.985 ;
        RECT 22.855 167.795 23.775 168.025 ;
        RECT 26.605 167.795 27.535 168.015 ;
        RECT 22.855 167.115 32.045 167.795 ;
        RECT 32.055 167.115 35.725 167.925 ;
        RECT 35.745 167.115 37.095 168.025 ;
        RECT 40.315 167.795 41.245 168.025 ;
        RECT 37.345 167.115 41.245 167.795 ;
        RECT 41.255 167.115 42.625 167.895 ;
        RECT 42.635 167.115 44.005 167.925 ;
        RECT 47.215 167.795 48.145 168.025 ;
        RECT 44.245 167.115 48.145 167.795 ;
        RECT 48.165 167.200 48.595 167.985 ;
        RECT 49.075 167.115 50.905 167.925 ;
        RECT 50.915 167.115 52.285 167.895 ;
        RECT 52.755 167.115 54.585 167.925 ;
        RECT 54.605 167.115 55.955 168.025 ;
        RECT 56.115 167.115 58.725 168.025 ;
        RECT 58.875 167.115 61.485 168.025 ;
        RECT 61.495 167.115 67.005 167.925 ;
        RECT 67.025 167.115 69.765 167.795 ;
        RECT 69.775 167.115 71.145 167.895 ;
        RECT 71.155 167.795 72.500 168.025 ;
        RECT 71.155 167.115 72.985 167.795 ;
        RECT 73.925 167.200 74.355 167.985 ;
        RECT 74.375 167.115 78.045 167.925 ;
        RECT 78.055 167.115 83.565 167.925 ;
        RECT 83.575 167.115 92.680 167.795 ;
        RECT 93.705 167.115 95.055 168.025 ;
        RECT 98.275 167.795 99.205 168.025 ;
        RECT 95.305 167.115 99.205 167.795 ;
        RECT 99.685 167.200 100.115 167.985 ;
        RECT 101.250 167.115 104.725 168.025 ;
        RECT 104.735 167.115 106.565 167.925 ;
        RECT 106.585 167.115 107.935 168.025 ;
        RECT 107.955 167.795 108.875 168.025 ;
        RECT 111.705 167.795 112.635 168.015 ;
        RECT 107.955 167.115 117.145 167.795 ;
        RECT 117.155 167.115 118.525 167.895 ;
        RECT 118.995 167.115 124.505 167.925 ;
        RECT 124.515 167.115 125.885 167.925 ;
        RECT 11.955 166.905 12.125 167.115 ;
        RECT 14.255 166.905 14.425 167.095 ;
        RECT 16.555 166.925 16.725 167.115 ;
        RECT 17.935 166.925 18.105 167.115 ;
        RECT 21.800 167.095 21.970 167.115 ;
        RECT 19.775 166.905 19.945 167.095 ;
        RECT 20.235 166.905 20.405 167.095 ;
        RECT 21.800 166.925 22.060 167.095 ;
        RECT 31.735 166.925 31.905 167.115 ;
        RECT 21.890 166.905 22.060 166.925 ;
        RECT 34.495 166.905 34.665 167.095 ;
        RECT 35.010 166.955 35.130 167.065 ;
        RECT 35.415 166.925 35.585 167.115 ;
        RECT 35.875 166.925 36.045 167.115 ;
        RECT 37.255 166.905 37.425 167.095 ;
        RECT 37.720 166.905 37.890 167.095 ;
        RECT 40.660 166.925 40.830 167.115 ;
        RECT 41.395 166.925 41.565 167.115 ;
        RECT 41.855 166.950 42.015 167.060 ;
        RECT 42.320 166.905 42.490 167.095 ;
        RECT 43.695 166.925 43.865 167.115 ;
        RECT 46.000 166.905 46.170 167.095 ;
        RECT 47.560 166.925 47.730 167.115 ;
        RECT 48.810 166.955 48.930 167.065 ;
        RECT 50.595 166.925 50.765 167.115 ;
        RECT 51.055 166.905 51.225 167.115 ;
        RECT 52.490 166.955 52.610 167.065 ;
        RECT 54.275 166.925 54.445 167.115 ;
        RECT 54.735 166.925 54.905 167.115 ;
        RECT 58.410 166.925 58.580 167.115 ;
        RECT 60.715 166.905 60.885 167.095 ;
        RECT 61.170 166.925 61.340 167.115 ;
        RECT 62.555 166.905 62.725 167.095 ;
        RECT 65.315 166.905 65.485 167.095 ;
        RECT 65.830 166.955 65.950 167.065 ;
        RECT 66.695 166.925 66.865 167.115 ;
        RECT 67.615 166.905 67.785 167.095 ;
        RECT 69.455 166.905 69.625 167.115 ;
        RECT 69.915 166.905 70.085 167.095 ;
        RECT 70.835 166.925 71.005 167.115 ;
        RECT 72.675 166.925 72.845 167.115 ;
        RECT 73.595 166.960 73.755 167.070 ;
        RECT 74.055 166.905 74.225 167.095 ;
        RECT 75.435 166.905 75.605 167.095 ;
        RECT 76.815 166.905 76.985 167.095 ;
        RECT 77.735 166.925 77.905 167.115 ;
        RECT 83.255 166.925 83.425 167.115 ;
        RECT 83.715 166.925 83.885 167.115 ;
        RECT 86.475 166.905 86.645 167.095 ;
        RECT 87.450 166.955 87.570 167.065 ;
        RECT 92.455 166.905 92.625 167.095 ;
        RECT 93.375 166.960 93.535 167.070 ;
        RECT 93.835 166.905 94.005 167.095 ;
        RECT 94.755 166.925 94.925 167.115 ;
        RECT 95.215 166.905 95.385 167.095 ;
        RECT 95.675 166.905 95.845 167.095 ;
        RECT 98.620 166.925 98.790 167.115 ;
        RECT 99.410 166.955 99.530 167.065 ;
        RECT 100.735 166.960 100.895 167.070 ;
        RECT 104.410 166.925 104.580 167.115 ;
        RECT 106.255 166.925 106.425 167.115 ;
        RECT 106.715 166.925 106.885 167.115 ;
        RECT 107.175 166.905 107.345 167.095 ;
        RECT 111.040 166.905 111.210 167.095 ;
        RECT 112.235 166.950 112.395 167.060 ;
        RECT 115.455 166.905 115.625 167.095 ;
        RECT 115.915 166.905 116.085 167.095 ;
        RECT 116.835 166.925 117.005 167.115 ;
        RECT 118.215 166.905 118.385 167.115 ;
        RECT 118.675 167.065 118.845 167.095 ;
        RECT 118.675 166.955 118.850 167.065 ;
        RECT 118.675 166.905 118.845 166.955 ;
        RECT 120.515 166.950 120.675 167.060 ;
        RECT 124.195 166.905 124.365 167.115 ;
        RECT 125.575 166.905 125.745 167.115 ;
        RECT 11.815 166.095 13.185 166.905 ;
        RECT 13.195 166.095 14.565 166.905 ;
        RECT 14.575 166.095 20.085 166.905 ;
        RECT 20.095 166.125 21.465 166.905 ;
        RECT 21.475 166.225 25.375 166.905 ;
        RECT 25.615 166.225 34.805 166.905 ;
        RECT 21.475 165.995 22.405 166.225 ;
        RECT 25.615 165.995 26.535 166.225 ;
        RECT 29.365 166.005 30.295 166.225 ;
        RECT 35.285 166.035 35.715 166.820 ;
        RECT 35.735 166.095 37.565 166.905 ;
        RECT 37.575 165.995 41.050 166.905 ;
        RECT 42.175 165.995 45.650 166.905 ;
        RECT 45.855 165.995 49.330 166.905 ;
        RECT 49.535 166.095 51.365 166.905 ;
        RECT 51.745 166.225 61.025 166.905 ;
        RECT 51.745 166.105 54.080 166.225 ;
        RECT 51.745 165.995 52.665 166.105 ;
        RECT 58.745 166.005 59.665 166.225 ;
        RECT 61.045 166.035 61.475 166.820 ;
        RECT 61.495 166.125 62.865 166.905 ;
        RECT 62.885 166.225 65.625 166.905 ;
        RECT 66.095 166.095 67.925 166.905 ;
        RECT 67.935 166.225 69.765 166.905 ;
        RECT 69.775 166.225 71.605 166.905 ;
        RECT 67.935 165.995 69.280 166.225 ;
        RECT 70.260 165.995 71.605 166.225 ;
        RECT 71.645 165.995 74.365 166.905 ;
        RECT 74.375 166.125 75.745 166.905 ;
        RECT 75.755 166.095 77.125 166.905 ;
        RECT 77.505 166.225 86.785 166.905 ;
        RECT 77.505 166.105 79.840 166.225 ;
        RECT 77.505 165.995 78.425 166.105 ;
        RECT 84.505 166.005 85.425 166.225 ;
        RECT 86.805 166.035 87.235 166.820 ;
        RECT 87.950 166.225 92.765 166.905 ;
        RECT 92.775 166.125 94.145 166.905 ;
        RECT 94.155 166.095 95.525 166.905 ;
        RECT 95.535 166.225 104.640 166.905 ;
        RECT 104.735 166.095 107.485 166.905 ;
        RECT 107.725 166.225 111.625 166.905 ;
        RECT 110.695 165.995 111.625 166.225 ;
        RECT 112.565 166.035 112.995 166.820 ;
        RECT 113.015 166.095 115.765 166.905 ;
        RECT 115.785 165.995 117.135 166.905 ;
        RECT 117.155 166.095 118.525 166.905 ;
        RECT 118.535 166.125 119.905 166.905 ;
        RECT 120.835 166.095 124.505 166.905 ;
        RECT 124.515 166.095 125.885 166.905 ;
      LAYER nwell ;
        RECT 11.620 162.875 126.080 165.705 ;
      LAYER pwell ;
        RECT 11.815 161.675 13.185 162.485 ;
        RECT 13.195 161.675 16.865 162.485 ;
        RECT 16.875 161.675 22.385 162.485 ;
        RECT 22.405 161.760 22.835 162.545 ;
        RECT 23.315 161.675 28.825 162.485 ;
        RECT 31.490 162.355 32.410 162.585 ;
        RECT 28.945 161.675 32.410 162.355 ;
        RECT 32.515 161.675 33.885 162.485 ;
        RECT 33.895 161.675 35.265 162.455 ;
        RECT 35.470 161.675 38.945 162.585 ;
        RECT 38.955 161.675 48.060 162.355 ;
        RECT 48.165 161.760 48.595 162.545 ;
        RECT 49.075 161.675 51.825 162.485 ;
        RECT 55.035 162.355 55.965 162.585 ;
        RECT 52.065 161.675 55.965 162.355 ;
        RECT 56.345 162.475 57.265 162.585 ;
        RECT 56.345 162.355 58.680 162.475 ;
        RECT 63.345 162.355 64.265 162.575 ;
        RECT 56.345 161.675 65.625 162.355 ;
        RECT 66.095 161.675 67.925 162.485 ;
        RECT 67.935 161.675 69.305 162.455 ;
        RECT 69.800 162.355 71.145 162.585 ;
        RECT 69.315 161.675 71.145 162.355 ;
        RECT 71.155 161.675 73.875 162.585 ;
        RECT 73.925 161.760 74.355 162.545 ;
        RECT 74.835 161.675 76.665 162.485 ;
        RECT 79.875 162.355 80.805 162.585 ;
        RECT 76.905 161.675 80.805 162.355 ;
        RECT 81.185 162.475 82.105 162.585 ;
        RECT 81.185 162.355 83.520 162.475 ;
        RECT 88.185 162.355 89.105 162.575 ;
        RECT 90.475 162.355 91.395 162.585 ;
        RECT 94.225 162.355 95.155 162.575 ;
        RECT 81.185 161.675 90.465 162.355 ;
        RECT 90.475 161.675 99.665 162.355 ;
        RECT 99.685 161.760 100.115 162.545 ;
        RECT 100.135 161.675 103.610 162.585 ;
        RECT 103.815 161.675 107.290 162.585 ;
        RECT 107.955 161.675 113.465 162.485 ;
        RECT 113.475 162.355 114.395 162.585 ;
        RECT 117.225 162.355 118.155 162.575 ;
        RECT 113.475 161.675 122.665 162.355 ;
        RECT 122.675 161.675 124.505 162.485 ;
        RECT 124.515 161.675 125.885 162.485 ;
        RECT 11.955 161.465 12.125 161.675 ;
        RECT 13.795 161.510 13.955 161.620 ;
        RECT 16.555 161.485 16.725 161.675 ;
        RECT 19.315 161.465 19.485 161.655 ;
        RECT 22.075 161.485 22.245 161.675 ;
        RECT 23.050 161.515 23.170 161.625 ;
        RECT 23.180 161.465 23.350 161.655 ;
        RECT 28.515 161.485 28.685 161.675 ;
        RECT 28.975 161.465 29.145 161.675 ;
        RECT 32.840 161.465 33.010 161.655 ;
        RECT 33.575 161.485 33.745 161.675 ;
        RECT 34.955 161.465 35.125 161.675 ;
        RECT 36.335 161.510 36.495 161.620 ;
        RECT 38.630 161.485 38.800 161.675 ;
        RECT 39.095 161.485 39.265 161.675 ;
        RECT 51.515 161.655 51.685 161.675 ;
        RECT 40.010 161.465 40.180 161.655 ;
        RECT 48.810 161.515 48.930 161.625 ;
        RECT 51.050 161.465 51.220 161.655 ;
        RECT 51.515 161.485 51.690 161.655 ;
        RECT 55.380 161.485 55.550 161.675 ;
        RECT 51.520 161.465 51.690 161.485 ;
        RECT 56.115 161.465 56.285 161.655 ;
        RECT 59.980 161.465 60.150 161.655 ;
        RECT 60.770 161.515 60.890 161.625 ;
        RECT 61.635 161.465 61.805 161.655 ;
        RECT 64.395 161.465 64.565 161.655 ;
        RECT 65.315 161.485 65.485 161.675 ;
        RECT 65.830 161.515 65.950 161.625 ;
        RECT 66.235 161.465 66.405 161.655 ;
        RECT 67.615 161.485 67.785 161.675 ;
        RECT 68.075 161.465 68.245 161.655 ;
        RECT 68.995 161.485 69.165 161.675 ;
        RECT 69.455 161.485 69.625 161.675 ;
        RECT 69.915 161.465 70.085 161.655 ;
        RECT 70.430 161.515 70.550 161.625 ;
        RECT 71.295 161.485 71.465 161.675 ;
        RECT 72.215 161.465 72.385 161.655 ;
        RECT 73.595 161.465 73.765 161.655 ;
        RECT 74.055 161.465 74.225 161.655 ;
        RECT 74.570 161.515 74.690 161.625 ;
        RECT 76.355 161.485 76.525 161.675 ;
        RECT 80.030 161.465 80.200 161.655 ;
        RECT 80.220 161.485 80.390 161.675 ;
        RECT 81.875 161.465 82.045 161.655 ;
        RECT 85.740 161.465 85.910 161.655 ;
        RECT 86.530 161.515 86.650 161.625 ;
        RECT 87.395 161.465 87.565 161.655 ;
        RECT 89.695 161.465 89.865 161.655 ;
        RECT 90.155 161.625 90.325 161.675 ;
        RECT 90.155 161.515 90.330 161.625 ;
        RECT 90.155 161.485 90.325 161.515 ;
        RECT 90.615 161.465 90.785 161.655 ;
        RECT 92.915 161.465 93.085 161.655 ;
        RECT 99.355 161.485 99.525 161.675 ;
        RECT 100.280 161.485 100.450 161.675 ;
        RECT 102.575 161.465 102.745 161.655 ;
        RECT 103.960 161.485 104.130 161.675 ;
        RECT 104.415 161.465 104.585 161.655 ;
        RECT 104.880 161.465 105.050 161.655 ;
        RECT 107.690 161.515 107.810 161.625 ;
        RECT 108.610 161.515 108.730 161.625 ;
        RECT 112.235 161.465 112.405 161.655 ;
        RECT 113.155 161.485 113.325 161.675 ;
        RECT 116.560 161.465 116.730 161.655 ;
        RECT 117.350 161.515 117.470 161.625 ;
        RECT 117.755 161.465 117.925 161.655 ;
        RECT 119.190 161.515 119.310 161.625 ;
        RECT 119.595 161.465 119.765 161.655 ;
        RECT 122.355 161.485 122.525 161.675 ;
        RECT 124.195 161.465 124.365 161.675 ;
        RECT 125.575 161.465 125.745 161.675 ;
        RECT 11.815 160.655 13.185 161.465 ;
        RECT 14.115 160.655 19.625 161.465 ;
        RECT 19.865 160.785 23.765 161.465 ;
        RECT 22.835 160.555 23.765 160.785 ;
        RECT 23.775 160.655 29.285 161.465 ;
        RECT 29.525 160.785 33.425 161.465 ;
        RECT 32.495 160.555 33.425 160.785 ;
        RECT 33.435 160.655 35.265 161.465 ;
        RECT 35.285 160.595 35.715 161.380 ;
        RECT 36.850 160.555 40.325 161.465 ;
        RECT 40.355 160.555 51.365 161.465 ;
        RECT 51.375 160.555 54.850 161.465 ;
        RECT 55.055 160.655 56.425 161.465 ;
        RECT 56.665 160.785 60.565 161.465 ;
        RECT 59.635 160.555 60.565 160.785 ;
        RECT 61.045 160.595 61.475 161.380 ;
        RECT 61.495 160.685 62.865 161.465 ;
        RECT 62.875 160.655 64.705 161.465 ;
        RECT 64.715 160.785 66.545 161.465 ;
        RECT 66.555 160.785 68.385 161.465 ;
        RECT 68.395 160.785 70.225 161.465 ;
        RECT 70.695 160.785 72.525 161.465 ;
        RECT 64.715 160.555 66.060 160.785 ;
        RECT 66.555 160.555 67.900 160.785 ;
        RECT 68.395 160.555 69.740 160.785 ;
        RECT 70.695 160.555 72.040 160.785 ;
        RECT 72.535 160.655 73.905 161.465 ;
        RECT 73.915 160.785 76.655 161.465 ;
        RECT 76.870 160.555 80.345 161.465 ;
        RECT 80.355 160.655 82.185 161.465 ;
        RECT 82.425 160.785 86.325 161.465 ;
        RECT 85.395 160.555 86.325 160.785 ;
        RECT 86.805 160.595 87.235 161.380 ;
        RECT 87.255 160.685 88.625 161.465 ;
        RECT 88.645 160.555 89.995 161.465 ;
        RECT 90.475 160.685 91.845 161.465 ;
        RECT 91.865 160.555 93.215 161.465 ;
        RECT 93.605 160.785 102.885 161.465 ;
        RECT 93.605 160.665 95.940 160.785 ;
        RECT 93.605 160.555 94.525 160.665 ;
        RECT 100.605 160.565 101.525 160.785 ;
        RECT 102.895 160.655 104.725 161.465 ;
        RECT 104.735 160.555 108.210 161.465 ;
        RECT 108.875 160.655 112.545 161.465 ;
        RECT 112.565 160.595 112.995 161.380 ;
        RECT 113.245 160.785 117.145 161.465 ;
        RECT 116.215 160.555 117.145 160.785 ;
        RECT 117.625 160.555 118.975 161.465 ;
        RECT 119.455 160.685 120.825 161.465 ;
        RECT 120.835 160.655 124.505 161.465 ;
        RECT 124.515 160.655 125.885 161.465 ;
      LAYER nwell ;
        RECT 11.620 157.435 126.080 160.265 ;
      LAYER pwell ;
        RECT 11.815 156.235 13.185 157.045 ;
        RECT 13.195 156.915 14.115 157.145 ;
        RECT 16.945 156.915 17.875 157.135 ;
        RECT 13.195 156.235 22.385 156.915 ;
        RECT 22.405 156.320 22.835 157.105 ;
        RECT 22.855 156.235 24.225 157.015 ;
        RECT 24.235 156.235 26.065 157.045 ;
        RECT 26.085 156.235 27.435 157.145 ;
        RECT 27.540 156.235 36.645 156.915 ;
        RECT 37.310 156.235 40.785 157.145 ;
        RECT 40.795 156.235 44.270 157.145 ;
        RECT 44.475 156.235 47.950 157.145 ;
        RECT 48.165 156.320 48.595 157.105 ;
        RECT 49.075 156.235 51.825 157.045 ;
        RECT 55.035 156.915 55.965 157.145 ;
        RECT 52.065 156.235 55.965 156.915 ;
        RECT 56.345 157.035 57.265 157.145 ;
        RECT 56.345 156.915 58.680 157.035 ;
        RECT 63.345 156.915 64.265 157.135 ;
        RECT 67.040 156.915 68.385 157.145 ;
        RECT 68.880 156.915 70.225 157.145 ;
        RECT 56.345 156.235 65.625 156.915 ;
        RECT 66.555 156.235 68.385 156.915 ;
        RECT 68.395 156.235 70.225 156.915 ;
        RECT 71.155 156.915 72.500 157.145 ;
        RECT 71.155 156.235 72.985 156.915 ;
        RECT 73.925 156.320 74.355 157.105 ;
        RECT 74.375 156.235 76.205 157.045 ;
        RECT 76.215 156.235 79.690 157.145 ;
        RECT 83.555 156.915 84.485 157.145 ;
        RECT 80.585 156.235 84.485 156.915 ;
        RECT 84.865 157.035 85.785 157.145 ;
        RECT 84.865 156.915 87.200 157.035 ;
        RECT 91.865 156.915 92.785 157.135 ;
        RECT 84.865 156.235 94.145 156.915 ;
        RECT 94.165 156.235 95.515 157.145 ;
        RECT 98.735 156.915 99.665 157.145 ;
        RECT 95.765 156.235 99.665 156.915 ;
        RECT 99.685 156.320 100.115 157.105 ;
        RECT 100.135 156.235 101.505 157.015 ;
        RECT 102.635 156.235 104.725 157.045 ;
        RECT 105.655 156.235 109.130 157.145 ;
        RECT 113.455 156.915 114.385 157.145 ;
        RECT 110.485 156.235 114.385 156.915 ;
        RECT 114.765 157.035 115.685 157.145 ;
        RECT 114.765 156.915 117.100 157.035 ;
        RECT 121.765 156.915 122.685 157.135 ;
        RECT 114.765 156.235 124.045 156.915 ;
        RECT 124.515 156.235 125.885 157.045 ;
        RECT 11.955 156.025 12.125 156.235 ;
        RECT 14.255 156.025 14.425 156.215 ;
        RECT 22.075 156.045 22.245 156.235 ;
        RECT 23.455 156.025 23.625 156.215 ;
        RECT 23.915 156.045 24.085 156.235 ;
        RECT 24.375 156.070 24.535 156.180 ;
        RECT 25.755 156.025 25.925 156.235 ;
        RECT 26.215 156.045 26.385 156.235 ;
        RECT 34.955 156.025 35.125 156.215 ;
        RECT 36.335 156.045 36.505 156.235 ;
        RECT 36.850 156.075 36.970 156.185 ;
        RECT 38.175 156.025 38.345 156.215 ;
        RECT 39.555 156.025 39.725 156.215 ;
        RECT 40.470 156.045 40.640 156.235 ;
        RECT 40.940 156.045 41.110 156.235 ;
        RECT 43.235 156.025 43.405 156.215 ;
        RECT 43.700 156.025 43.870 156.215 ;
        RECT 44.620 156.045 44.790 156.235 ;
        RECT 47.380 156.025 47.550 156.215 ;
        RECT 48.810 156.075 48.930 156.185 ;
        RECT 51.060 156.025 51.230 156.215 ;
        RECT 51.515 156.045 51.685 156.235 ;
        RECT 54.790 156.075 54.910 156.185 ;
        RECT 55.380 156.045 55.550 156.235 ;
        RECT 56.575 156.025 56.745 156.215 ;
        RECT 57.035 156.025 57.205 156.215 ;
        RECT 58.415 156.025 58.585 156.215 ;
        RECT 59.795 156.025 59.965 156.215 ;
        RECT 62.555 156.025 62.725 156.215 ;
        RECT 65.315 156.045 65.485 156.235 ;
        RECT 66.235 156.025 66.405 156.215 ;
        RECT 66.695 156.045 66.865 156.235 ;
        RECT 68.535 156.045 68.705 156.235 ;
        RECT 68.990 156.025 69.160 156.215 ;
        RECT 70.835 156.080 70.995 156.190 ;
        RECT 72.675 156.025 72.845 156.235 ;
        RECT 73.595 156.080 73.755 156.190 ;
        RECT 75.895 156.045 76.065 156.235 ;
        RECT 76.360 156.215 76.530 156.235 ;
        RECT 76.350 156.045 76.530 156.215 ;
        RECT 76.350 156.025 76.520 156.045 ;
        RECT 76.820 156.025 76.990 156.215 ;
        RECT 80.090 156.075 80.210 156.185 ;
        RECT 80.955 156.070 81.115 156.180 ;
        RECT 83.900 156.045 84.070 156.235 ;
        RECT 86.475 156.025 86.645 156.215 ;
        RECT 87.450 156.075 87.570 156.185 ;
        RECT 90.155 156.025 90.325 156.215 ;
        RECT 93.835 156.045 94.005 156.235 ;
        RECT 94.295 156.045 94.465 156.235 ;
        RECT 95.675 156.025 95.845 156.215 ;
        RECT 99.080 156.045 99.250 156.235 ;
        RECT 100.275 156.045 100.445 156.235 ;
        RECT 101.195 156.025 101.365 156.215 ;
        RECT 101.710 156.075 101.830 156.185 ;
        RECT 104.415 156.045 104.585 156.235 ;
        RECT 104.870 156.025 105.040 156.215 ;
        RECT 105.340 156.190 105.510 156.215 ;
        RECT 105.335 156.080 105.510 156.190 ;
        RECT 105.340 156.025 105.510 156.080 ;
        RECT 105.800 156.045 105.970 156.235 ;
        RECT 109.935 156.080 110.095 156.190 ;
        RECT 112.235 156.025 112.405 156.215 ;
        RECT 113.800 156.045 113.970 156.235 ;
        RECT 114.075 156.025 114.245 156.215 ;
        RECT 116.830 156.025 117.000 156.215 ;
        RECT 118.675 156.025 118.845 156.215 ;
        RECT 123.735 156.045 123.905 156.235 ;
        RECT 124.195 156.185 124.365 156.215 ;
        RECT 124.195 156.075 124.370 156.185 ;
        RECT 124.195 156.025 124.365 156.075 ;
        RECT 125.575 156.025 125.745 156.235 ;
        RECT 11.815 155.215 13.185 156.025 ;
        RECT 13.205 155.115 14.555 156.025 ;
        RECT 14.575 155.345 23.765 156.025 ;
        RECT 14.575 155.115 15.495 155.345 ;
        RECT 18.325 155.125 19.255 155.345 ;
        RECT 24.695 155.245 26.065 156.025 ;
        RECT 26.075 155.345 35.265 156.025 ;
        RECT 26.075 155.115 26.995 155.345 ;
        RECT 29.825 155.125 30.755 155.345 ;
        RECT 35.285 155.155 35.715 155.940 ;
        RECT 36.395 155.215 38.485 156.025 ;
        RECT 38.495 155.215 39.865 156.025 ;
        RECT 39.875 155.215 43.545 156.025 ;
        RECT 43.555 155.115 47.030 156.025 ;
        RECT 47.235 155.115 50.710 156.025 ;
        RECT 50.915 155.115 54.390 156.025 ;
        RECT 55.055 155.215 56.885 156.025 ;
        RECT 56.905 155.115 58.255 156.025 ;
        RECT 58.285 155.115 59.635 156.025 ;
        RECT 59.655 155.245 61.025 156.025 ;
        RECT 61.045 155.155 61.475 155.940 ;
        RECT 61.495 155.215 62.865 156.025 ;
        RECT 62.875 155.215 66.545 156.025 ;
        RECT 66.695 155.115 69.305 156.025 ;
        RECT 69.315 155.215 72.985 156.025 ;
        RECT 73.190 155.115 76.665 156.025 ;
        RECT 76.675 155.115 80.150 156.025 ;
        RECT 81.275 155.215 86.785 156.025 ;
        RECT 86.805 155.155 87.235 155.940 ;
        RECT 87.715 155.215 90.465 156.025 ;
        RECT 90.475 155.215 95.985 156.025 ;
        RECT 95.995 155.215 101.505 156.025 ;
        RECT 101.710 155.115 105.185 156.025 ;
        RECT 105.195 155.115 108.670 156.025 ;
        RECT 108.875 155.215 112.545 156.025 ;
        RECT 112.565 155.155 112.995 155.940 ;
        RECT 113.015 155.215 114.385 156.025 ;
        RECT 114.535 155.115 117.145 156.025 ;
        RECT 117.155 155.215 118.985 156.025 ;
        RECT 118.995 155.215 124.505 156.025 ;
        RECT 124.515 155.215 125.885 156.025 ;
      LAYER nwell ;
        RECT 11.620 151.995 126.080 154.825 ;
      LAYER pwell ;
        RECT 11.815 150.795 13.185 151.605 ;
        RECT 13.195 151.475 14.115 151.705 ;
        RECT 16.945 151.475 17.875 151.695 ;
        RECT 13.195 150.795 22.385 151.475 ;
        RECT 22.405 150.880 22.835 151.665 ;
        RECT 22.855 151.475 23.785 151.705 ;
        RECT 27.915 151.475 28.835 151.705 ;
        RECT 31.665 151.475 32.595 151.695 ;
        RECT 22.855 150.795 26.755 151.475 ;
        RECT 27.915 150.795 37.105 151.475 ;
        RECT 37.115 150.795 38.485 151.575 ;
        RECT 38.955 150.795 41.705 151.605 ;
        RECT 41.910 150.795 45.385 151.705 ;
        RECT 45.395 150.795 48.145 151.605 ;
        RECT 48.165 150.880 48.595 151.665 ;
        RECT 49.075 150.795 50.905 151.605 ;
        RECT 50.915 150.795 54.390 151.705 ;
        RECT 55.515 150.795 59.185 151.605 ;
        RECT 59.195 150.795 64.705 151.605 ;
        RECT 64.715 150.795 70.225 151.605 ;
        RECT 70.430 150.795 73.905 151.705 ;
        RECT 73.925 150.880 74.355 151.665 ;
        RECT 74.375 150.795 76.205 151.605 ;
        RECT 76.215 150.795 79.690 151.705 ;
        RECT 79.895 150.795 83.370 151.705 ;
        RECT 83.575 150.795 84.945 151.605 ;
        RECT 84.955 150.795 90.465 151.605 ;
        RECT 90.475 150.795 95.985 151.605 ;
        RECT 95.995 150.795 99.470 151.705 ;
        RECT 99.685 150.880 100.115 151.665 ;
        RECT 100.135 150.795 101.505 151.605 ;
        RECT 101.515 150.795 104.990 151.705 ;
        RECT 106.115 150.795 109.590 151.705 ;
        RECT 110.255 150.795 112.865 151.705 ;
        RECT 113.015 151.475 113.935 151.705 ;
        RECT 116.765 151.475 117.695 151.695 ;
        RECT 113.015 150.795 122.205 151.475 ;
        RECT 122.675 150.795 124.505 151.605 ;
        RECT 124.515 150.795 125.885 151.605 ;
        RECT 11.955 150.585 12.125 150.795 ;
        RECT 13.390 150.635 13.510 150.745 ;
        RECT 15.175 150.585 15.345 150.775 ;
        RECT 15.635 150.585 15.805 150.775 ;
        RECT 17.935 150.585 18.105 150.775 ;
        RECT 18.395 150.585 18.565 150.775 ;
        RECT 20.050 150.585 20.220 150.775 ;
        RECT 22.075 150.605 22.245 150.795 ;
        RECT 23.270 150.605 23.440 150.795 ;
        RECT 25.295 150.585 25.465 150.775 ;
        RECT 25.755 150.585 25.925 150.775 ;
        RECT 27.595 150.640 27.755 150.750 ;
        RECT 30.540 150.585 30.710 150.775 ;
        RECT 34.680 150.585 34.850 150.775 ;
        RECT 36.795 150.585 36.965 150.795 ;
        RECT 38.175 150.605 38.345 150.795 ;
        RECT 38.635 150.745 38.805 150.775 ;
        RECT 38.635 150.635 38.810 150.745 ;
        RECT 38.635 150.585 38.805 150.635 ;
        RECT 39.100 150.585 39.270 150.775 ;
        RECT 41.395 150.605 41.565 150.795 ;
        RECT 45.070 150.605 45.240 150.795 ;
        RECT 45.990 150.585 46.160 150.775 ;
        RECT 46.510 150.635 46.630 150.745 ;
        RECT 47.835 150.605 48.005 150.795 ;
        RECT 48.810 150.635 48.930 150.745 ;
        RECT 49.215 150.585 49.385 150.775 ;
        RECT 49.680 150.585 49.850 150.775 ;
        RECT 50.595 150.605 50.765 150.795 ;
        RECT 51.060 150.605 51.230 150.795 ;
        RECT 53.410 150.635 53.530 150.745 ;
        RECT 55.195 150.585 55.365 150.775 ;
        RECT 58.875 150.605 59.045 150.795 ;
        RECT 60.715 150.585 60.885 150.775 ;
        RECT 63.015 150.585 63.185 150.775 ;
        RECT 63.475 150.585 63.645 150.775 ;
        RECT 64.395 150.605 64.565 150.795 ;
        RECT 64.910 150.635 65.030 150.745 ;
        RECT 65.315 150.585 65.485 150.775 ;
        RECT 68.995 150.585 69.165 150.775 ;
        RECT 69.455 150.585 69.625 150.775 ;
        RECT 69.915 150.605 70.085 150.795 ;
        RECT 72.675 150.585 72.845 150.775 ;
        RECT 73.190 150.635 73.310 150.745 ;
        RECT 73.590 150.605 73.760 150.795 ;
        RECT 75.895 150.585 76.065 150.795 ;
        RECT 76.360 150.585 76.530 150.795 ;
        RECT 80.040 150.605 80.210 150.795 ;
        RECT 80.955 150.585 81.125 150.775 ;
        RECT 84.635 150.605 84.805 150.795 ;
        RECT 86.475 150.585 86.645 150.775 ;
        RECT 88.315 150.585 88.485 150.775 ;
        RECT 88.830 150.635 88.950 150.745 ;
        RECT 90.155 150.605 90.325 150.795 ;
        RECT 95.675 150.605 95.845 150.795 ;
        RECT 96.140 150.605 96.310 150.795 ;
        RECT 97.975 150.585 98.145 150.775 ;
        RECT 98.895 150.630 99.055 150.740 ;
        RECT 101.195 150.605 101.365 150.795 ;
        RECT 101.660 150.605 101.830 150.795 ;
        RECT 104.415 150.585 104.585 150.775 ;
        RECT 105.795 150.640 105.955 150.750 ;
        RECT 106.260 150.605 106.430 150.795 ;
        RECT 11.815 149.775 13.185 150.585 ;
        RECT 13.655 149.775 15.485 150.585 ;
        RECT 15.505 149.675 16.855 150.585 ;
        RECT 16.885 149.675 18.235 150.585 ;
        RECT 18.255 149.805 19.625 150.585 ;
        RECT 19.635 149.905 23.535 150.585 ;
        RECT 19.635 149.675 20.565 149.905 ;
        RECT 23.775 149.775 25.605 150.585 ;
        RECT 25.625 149.675 26.975 150.585 ;
        RECT 27.225 149.905 31.125 150.585 ;
        RECT 31.365 149.905 35.265 150.585 ;
        RECT 30.195 149.675 31.125 149.905 ;
        RECT 34.335 149.675 35.265 149.905 ;
        RECT 35.285 149.715 35.715 150.500 ;
        RECT 35.735 149.805 37.105 150.585 ;
        RECT 37.115 149.775 38.945 150.585 ;
        RECT 38.955 149.675 42.430 150.585 ;
        RECT 42.830 149.675 46.305 150.585 ;
        RECT 46.775 149.775 49.525 150.585 ;
        RECT 49.535 149.675 53.010 150.585 ;
        RECT 53.675 149.775 55.505 150.585 ;
        RECT 55.515 149.775 61.025 150.585 ;
        RECT 61.045 149.715 61.475 150.500 ;
        RECT 61.495 149.775 63.325 150.585 ;
        RECT 63.345 149.675 64.695 150.585 ;
        RECT 65.175 149.805 66.545 150.585 ;
        RECT 66.555 149.775 69.305 150.585 ;
        RECT 69.315 149.905 71.145 150.585 ;
        RECT 69.800 149.675 71.145 149.905 ;
        RECT 71.155 149.905 72.985 150.585 ;
        RECT 71.155 149.675 72.500 149.905 ;
        RECT 73.455 149.775 76.205 150.585 ;
        RECT 76.215 149.675 79.690 150.585 ;
        RECT 79.895 149.775 81.265 150.585 ;
        RECT 81.275 149.775 86.785 150.585 ;
        RECT 86.805 149.715 87.235 150.500 ;
        RECT 87.265 149.675 88.615 150.585 ;
        RECT 89.095 149.905 98.285 150.585 ;
        RECT 89.095 149.675 90.015 149.905 ;
        RECT 92.845 149.685 93.775 149.905 ;
        RECT 99.215 149.775 104.725 150.585 ;
        RECT 104.735 150.555 105.680 150.585 ;
        RECT 107.170 150.555 107.340 150.775 ;
        RECT 108.555 150.585 108.725 150.775 ;
        RECT 109.990 150.635 110.110 150.745 ;
        RECT 110.400 150.605 110.570 150.795 ;
        RECT 112.235 150.585 112.405 150.775 ;
        RECT 113.210 150.635 113.330 150.745 ;
        RECT 115.915 150.585 116.085 150.775 ;
        RECT 117.295 150.585 117.465 150.775 ;
        RECT 117.755 150.585 117.925 150.775 ;
        RECT 121.895 150.605 122.065 150.795 ;
        RECT 122.410 150.635 122.530 150.745 ;
        RECT 124.195 150.585 124.365 150.795 ;
        RECT 125.575 150.585 125.745 150.795 ;
        RECT 104.735 149.875 107.485 150.555 ;
        RECT 104.735 149.675 105.680 149.875 ;
        RECT 107.495 149.775 108.865 150.585 ;
        RECT 108.875 149.775 112.545 150.585 ;
        RECT 112.565 149.715 112.995 150.500 ;
        RECT 113.475 149.775 116.225 150.585 ;
        RECT 116.245 149.675 117.595 150.585 ;
        RECT 117.615 149.805 118.985 150.585 ;
        RECT 118.995 149.775 124.505 150.585 ;
        RECT 124.515 149.775 125.885 150.585 ;
      LAYER nwell ;
        RECT 11.620 146.555 126.080 149.385 ;
      LAYER pwell ;
        RECT 11.815 145.355 13.185 146.165 ;
        RECT 13.195 145.355 16.865 146.165 ;
        RECT 16.875 145.355 22.385 146.165 ;
        RECT 22.405 145.440 22.835 146.225 ;
        RECT 23.775 145.355 27.445 146.165 ;
        RECT 27.455 145.355 32.965 146.165 ;
        RECT 32.975 145.355 38.485 146.165 ;
        RECT 38.690 145.355 42.165 146.265 ;
        RECT 42.370 145.355 45.845 146.265 ;
        RECT 46.315 145.355 48.145 146.165 ;
        RECT 48.165 145.440 48.595 146.225 ;
        RECT 48.615 145.355 52.285 146.165 ;
        RECT 52.295 145.355 55.770 146.265 ;
        RECT 55.975 145.355 59.450 146.265 ;
        RECT 68.855 146.035 70.200 146.265 ;
        RECT 59.740 145.355 68.845 146.035 ;
        RECT 68.855 145.355 70.685 146.035 ;
        RECT 71.155 145.355 73.875 146.265 ;
        RECT 73.925 145.440 74.355 146.225 ;
        RECT 74.860 146.035 76.205 146.265 ;
        RECT 76.700 146.035 78.045 146.265 ;
        RECT 74.375 145.355 76.205 146.035 ;
        RECT 76.215 145.355 78.045 146.035 ;
        RECT 78.975 145.355 82.645 146.165 ;
        RECT 83.025 146.155 83.945 146.265 ;
        RECT 83.025 146.035 85.360 146.155 ;
        RECT 90.025 146.035 90.945 146.255 ;
        RECT 83.025 145.355 92.305 146.035 ;
        RECT 92.325 145.355 93.675 146.265 ;
        RECT 94.155 145.355 95.525 146.135 ;
        RECT 95.535 145.355 96.905 146.165 ;
        RECT 98.720 146.065 99.665 146.265 ;
        RECT 96.915 145.385 99.665 146.065 ;
        RECT 99.685 145.440 100.115 146.225 ;
        RECT 11.955 145.145 12.125 145.355 ;
        RECT 13.390 145.195 13.510 145.305 ;
        RECT 16.555 145.165 16.725 145.355 ;
        RECT 22.075 145.165 22.245 145.355 ;
        RECT 22.995 145.145 23.165 145.335 ;
        RECT 23.455 145.200 23.615 145.310 ;
        RECT 23.915 145.190 24.075 145.300 ;
        RECT 27.135 145.165 27.305 145.355 ;
        RECT 29.435 145.145 29.605 145.335 ;
        RECT 32.655 145.165 32.825 145.355 ;
        RECT 34.955 145.145 35.125 145.335 ;
        RECT 36.335 145.190 36.495 145.300 ;
        RECT 38.175 145.165 38.345 145.355 ;
        RECT 11.815 144.335 13.185 145.145 ;
        RECT 14.025 144.465 23.305 145.145 ;
        RECT 14.025 144.345 16.360 144.465 ;
        RECT 14.025 144.235 14.945 144.345 ;
        RECT 21.025 144.245 21.945 144.465 ;
        RECT 24.235 144.335 29.745 145.145 ;
        RECT 29.755 144.335 35.265 145.145 ;
        RECT 36.655 145.115 37.600 145.145 ;
        RECT 39.090 145.115 39.260 145.335 ;
        RECT 39.610 145.195 39.730 145.305 ;
        RECT 41.850 145.165 42.020 145.355 ;
        RECT 39.875 145.115 40.820 145.145 ;
        RECT 42.310 145.115 42.480 145.335 ;
        RECT 42.780 145.145 42.950 145.335 ;
        RECT 45.530 145.165 45.700 145.355 ;
        RECT 46.050 145.195 46.170 145.305 ;
        RECT 47.835 145.165 48.005 145.355 ;
        RECT 51.515 145.145 51.685 145.335 ;
        RECT 51.975 145.145 52.145 145.355 ;
        RECT 52.440 145.165 52.610 145.355 ;
        RECT 53.360 145.145 53.530 145.335 ;
        RECT 56.120 145.165 56.290 145.355 ;
        RECT 60.440 145.145 60.610 145.335 ;
        RECT 68.535 145.165 68.705 145.355 ;
        RECT 70.375 145.165 70.545 145.355 ;
        RECT 70.835 145.305 71.005 145.335 ;
        RECT 70.835 145.195 71.010 145.305 ;
        RECT 70.835 145.145 71.005 145.195 ;
        RECT 71.295 145.165 71.465 145.355 ;
        RECT 73.595 145.145 73.765 145.335 ;
        RECT 74.055 145.145 74.225 145.335 ;
        RECT 74.515 145.165 74.685 145.355 ;
        RECT 75.950 145.195 76.070 145.305 ;
        RECT 76.355 145.145 76.525 145.355 ;
        RECT 78.655 145.200 78.815 145.310 ;
        RECT 82.335 145.145 82.505 145.355 ;
        RECT 86.200 145.145 86.370 145.335 ;
        RECT 87.450 145.195 87.570 145.305 ;
        RECT 87.855 145.145 88.025 145.335 ;
        RECT 91.995 145.165 92.165 145.355 ;
        RECT 92.640 145.145 92.810 145.335 ;
        RECT 93.375 145.165 93.545 145.355 ;
        RECT 93.890 145.195 94.010 145.305 ;
        RECT 94.295 145.165 94.465 145.355 ;
        RECT 94.755 145.145 94.925 145.335 ;
        RECT 96.595 145.165 96.765 145.355 ;
        RECT 97.060 145.165 97.230 145.385 ;
        RECT 98.720 145.355 99.665 145.385 ;
        RECT 100.595 145.355 102.425 146.165 ;
        RECT 102.435 145.355 105.910 146.265 ;
        RECT 106.575 145.355 110.050 146.265 ;
        RECT 114.375 146.035 115.305 146.265 ;
        RECT 111.405 145.355 115.305 146.035 ;
        RECT 115.775 145.355 117.605 146.165 ;
        RECT 117.625 145.355 118.975 146.265 ;
        RECT 119.455 145.355 120.825 146.135 ;
        RECT 120.835 145.355 124.505 146.165 ;
        RECT 124.515 145.355 125.885 146.165 ;
        RECT 100.275 145.305 100.445 145.335 ;
        RECT 100.275 145.195 100.450 145.305 ;
        RECT 100.275 145.145 100.445 145.195 ;
        RECT 102.115 145.165 102.285 145.355 ;
        RECT 102.580 145.165 102.750 145.355 ;
        RECT 35.285 144.275 35.715 145.060 ;
        RECT 36.655 144.435 39.405 145.115 ;
        RECT 39.875 144.435 42.625 145.115 ;
        RECT 36.655 144.235 37.600 144.435 ;
        RECT 39.875 144.235 40.820 144.435 ;
        RECT 42.635 144.235 46.110 145.145 ;
        RECT 46.315 144.335 51.825 145.145 ;
        RECT 51.835 144.365 53.205 145.145 ;
        RECT 53.215 144.235 56.690 145.145 ;
        RECT 57.125 144.465 61.025 145.145 ;
        RECT 60.095 144.235 61.025 144.465 ;
        RECT 61.045 144.275 61.475 145.060 ;
        RECT 61.865 144.465 71.145 145.145 ;
        RECT 71.165 144.465 73.905 145.145 ;
        RECT 73.915 144.465 75.745 145.145 ;
        RECT 76.215 144.465 78.955 145.145 ;
        RECT 61.865 144.345 64.200 144.465 ;
        RECT 61.865 144.235 62.785 144.345 ;
        RECT 68.865 144.245 69.785 144.465 ;
        RECT 74.400 144.235 75.745 144.465 ;
        RECT 78.975 144.335 82.645 145.145 ;
        RECT 82.885 144.465 86.785 145.145 ;
        RECT 85.855 144.235 86.785 144.465 ;
        RECT 86.805 144.275 87.235 145.060 ;
        RECT 87.715 144.365 89.085 145.145 ;
        RECT 89.325 144.465 93.225 145.145 ;
        RECT 92.295 144.235 93.225 144.465 ;
        RECT 93.235 144.335 95.065 145.145 ;
        RECT 95.075 144.335 100.585 145.145 ;
        RECT 100.595 145.115 101.540 145.145 ;
        RECT 103.030 145.115 103.200 145.335 ;
        RECT 103.495 145.145 103.665 145.335 ;
        RECT 106.310 145.195 106.430 145.305 ;
        RECT 106.720 145.165 106.890 145.355 ;
        RECT 107.180 145.145 107.350 145.335 ;
        RECT 110.855 145.200 111.015 145.310 ;
        RECT 112.235 145.145 112.405 145.335 ;
        RECT 114.075 145.145 114.245 145.335 ;
        RECT 114.720 145.165 114.890 145.355 ;
        RECT 115.510 145.195 115.630 145.305 ;
        RECT 117.295 145.165 117.465 145.355 ;
        RECT 117.755 145.165 117.925 145.355 ;
        RECT 119.190 145.195 119.310 145.305 ;
        RECT 119.595 145.165 119.765 145.355 ;
        RECT 123.735 145.145 123.905 145.335 ;
        RECT 124.195 145.305 124.365 145.355 ;
        RECT 124.195 145.195 124.370 145.305 ;
        RECT 124.195 145.165 124.365 145.195 ;
        RECT 125.575 145.145 125.745 145.355 ;
        RECT 100.595 144.435 103.345 145.115 ;
        RECT 103.465 144.465 106.930 145.145 ;
        RECT 100.595 144.235 101.540 144.435 ;
        RECT 106.010 144.235 106.930 144.465 ;
        RECT 107.035 144.235 110.510 145.145 ;
        RECT 110.715 144.335 112.545 145.145 ;
        RECT 112.565 144.275 112.995 145.060 ;
        RECT 113.015 144.335 114.385 145.145 ;
        RECT 114.765 144.465 124.045 145.145 ;
        RECT 114.765 144.345 117.100 144.465 ;
        RECT 114.765 144.235 115.685 144.345 ;
        RECT 121.765 144.245 122.685 144.465 ;
        RECT 124.515 144.335 125.885 145.145 ;
      LAYER nwell ;
        RECT 11.620 141.115 126.080 143.945 ;
      LAYER pwell ;
        RECT 11.815 139.915 13.185 140.725 ;
        RECT 13.655 139.915 15.485 140.725 ;
        RECT 15.495 139.915 21.005 140.725 ;
        RECT 21.015 139.915 22.385 140.695 ;
        RECT 22.405 140.000 22.835 140.785 ;
        RECT 22.865 139.915 24.215 140.825 ;
        RECT 24.235 139.915 26.065 140.725 ;
        RECT 29.275 140.595 30.205 140.825 ;
        RECT 33.195 140.735 34.145 140.825 ;
        RECT 26.305 139.915 30.205 140.595 ;
        RECT 30.215 139.915 32.045 140.725 ;
        RECT 32.215 139.915 34.145 140.735 ;
        RECT 34.355 140.625 35.300 140.825 ;
        RECT 37.115 140.625 38.060 140.825 ;
        RECT 41.015 140.735 41.965 140.825 ;
        RECT 34.355 139.945 37.105 140.625 ;
        RECT 37.115 139.945 39.865 140.625 ;
        RECT 34.355 139.915 35.300 139.945 ;
        RECT 11.955 139.705 12.125 139.915 ;
        RECT 13.390 139.755 13.510 139.865 ;
        RECT 13.795 139.750 13.955 139.860 ;
        RECT 15.175 139.705 15.345 139.915 ;
        RECT 19.040 139.705 19.210 139.895 ;
        RECT 20.695 139.725 20.865 139.915 ;
        RECT 21.155 139.725 21.325 139.915 ;
        RECT 22.995 139.725 23.165 139.915 ;
        RECT 25.755 139.725 25.925 139.915 ;
        RECT 28.975 139.705 29.145 139.895 ;
        RECT 29.620 139.725 29.790 139.915 ;
        RECT 30.355 139.705 30.525 139.895 ;
        RECT 30.870 139.755 30.990 139.865 ;
        RECT 31.735 139.725 31.905 139.915 ;
        RECT 32.215 139.895 32.365 139.915 ;
        RECT 32.195 139.725 32.365 139.895 ;
        RECT 34.680 139.705 34.850 139.895 ;
        RECT 35.875 139.725 36.045 139.895 ;
        RECT 36.790 139.725 36.960 139.945 ;
        RECT 37.115 139.915 38.060 139.945 ;
        RECT 39.550 139.725 39.720 139.945 ;
        RECT 40.035 139.915 41.965 140.735 ;
        RECT 42.635 139.915 48.145 140.725 ;
        RECT 48.165 140.000 48.595 140.785 ;
        RECT 48.615 140.595 49.535 140.825 ;
        RECT 52.365 140.595 53.295 140.815 ;
        RECT 48.615 139.915 57.805 140.595 ;
        RECT 57.815 139.915 61.290 140.825 ;
        RECT 61.955 139.915 63.785 140.725 ;
        RECT 64.165 140.715 65.085 140.825 ;
        RECT 64.165 140.595 66.500 140.715 ;
        RECT 71.165 140.595 72.085 140.815 ;
        RECT 64.165 139.915 73.445 140.595 ;
        RECT 73.925 140.000 74.355 140.785 ;
        RECT 75.295 140.625 76.240 140.825 ;
        RECT 75.295 139.945 78.045 140.625 ;
        RECT 75.295 139.915 76.240 139.945 ;
        RECT 40.035 139.895 40.185 139.915 ;
        RECT 40.015 139.725 40.185 139.895 ;
        RECT 42.370 139.755 42.490 139.865 ;
        RECT 35.895 139.705 36.045 139.725 ;
        RECT 40.015 139.705 40.165 139.725 ;
        RECT 43.695 139.705 43.865 139.895 ;
        RECT 11.815 138.895 13.185 139.705 ;
        RECT 14.125 138.795 15.475 139.705 ;
        RECT 15.725 139.025 19.625 139.705 ;
        RECT 18.695 138.795 19.625 139.025 ;
        RECT 20.005 139.025 29.285 139.705 ;
        RECT 20.005 138.905 22.340 139.025 ;
        RECT 20.005 138.795 20.925 138.905 ;
        RECT 27.005 138.805 27.925 139.025 ;
        RECT 29.295 138.925 30.665 139.705 ;
        RECT 31.365 139.025 35.265 139.705 ;
        RECT 34.335 138.795 35.265 139.025 ;
        RECT 35.285 138.835 35.715 139.620 ;
        RECT 35.895 138.885 37.825 139.705 ;
        RECT 36.875 138.795 37.825 138.885 ;
        RECT 38.235 138.885 40.165 139.705 ;
        RECT 40.335 138.895 44.005 139.705 ;
        RECT 44.160 139.675 44.330 139.895 ;
        RECT 46.970 139.755 47.090 139.865 ;
        RECT 47.380 139.705 47.550 139.895 ;
        RECT 47.835 139.725 48.005 139.915 ;
        RECT 51.110 139.755 51.230 139.865 ;
        RECT 52.435 139.705 52.605 139.895 ;
        RECT 52.950 139.755 53.070 139.865 ;
        RECT 53.630 139.705 53.800 139.895 ;
        RECT 57.495 139.725 57.665 139.915 ;
        RECT 57.960 139.725 58.130 139.915 ;
        RECT 60.715 139.705 60.885 139.895 ;
        RECT 61.645 139.705 61.815 139.895 ;
        RECT 63.015 139.705 63.185 139.895 ;
        RECT 63.475 139.725 63.645 139.915 ;
        RECT 66.750 139.755 66.870 139.865 ;
        RECT 67.155 139.705 67.325 139.895 ;
        RECT 68.535 139.705 68.705 139.895 ;
        RECT 71.755 139.705 71.925 139.895 ;
        RECT 73.135 139.725 73.305 139.915 ;
        RECT 77.730 139.895 77.900 139.945 ;
        RECT 78.055 139.915 81.530 140.825 ;
        RECT 82.105 140.715 83.025 140.825 ;
        RECT 82.105 140.595 84.440 140.715 ;
        RECT 89.105 140.595 90.025 140.815 ;
        RECT 82.105 139.915 91.385 140.595 ;
        RECT 91.395 139.915 93.225 140.725 ;
        RECT 95.040 140.625 95.985 140.825 ;
        RECT 93.235 139.945 95.985 140.625 ;
        RECT 73.650 139.755 73.770 139.865 ;
        RECT 74.975 139.760 75.135 139.870 ;
        RECT 77.275 139.705 77.445 139.895 ;
        RECT 77.730 139.725 77.910 139.895 ;
        RECT 78.200 139.725 78.370 139.915 ;
        RECT 81.470 139.755 81.590 139.865 ;
        RECT 77.740 139.705 77.910 139.725 ;
        RECT 85.095 139.705 85.265 139.895 ;
        RECT 86.475 139.705 86.645 139.895 ;
        RECT 87.395 139.705 87.565 139.895 ;
        RECT 89.695 139.705 89.865 139.895 ;
        RECT 91.075 139.725 91.245 139.915 ;
        RECT 92.915 139.725 93.085 139.915 ;
        RECT 93.380 139.895 93.550 139.945 ;
        RECT 95.040 139.915 95.985 139.945 ;
        RECT 95.995 139.915 99.470 140.825 ;
        RECT 99.685 140.000 100.115 140.785 ;
        RECT 100.135 139.915 103.805 140.725 ;
        RECT 103.815 139.915 107.290 140.825 ;
        RECT 107.495 139.915 109.325 140.725 ;
        RECT 112.535 140.595 113.465 140.825 ;
        RECT 116.675 140.595 117.605 140.825 ;
        RECT 109.565 139.915 113.465 140.595 ;
        RECT 113.705 139.915 117.605 140.595 ;
        RECT 117.625 139.915 118.975 140.825 ;
        RECT 119.455 139.915 120.825 140.695 ;
        RECT 120.835 139.915 124.505 140.725 ;
        RECT 124.515 139.915 125.885 140.725 ;
        RECT 93.375 139.725 93.550 139.895 ;
        RECT 96.140 139.725 96.310 139.915 ;
        RECT 93.375 139.705 93.545 139.725 ;
        RECT 98.895 139.705 99.065 139.895 ;
        RECT 45.820 139.675 46.765 139.705 ;
        RECT 44.015 138.995 46.765 139.675 ;
        RECT 38.235 138.795 39.185 138.885 ;
        RECT 45.820 138.795 46.765 138.995 ;
        RECT 47.235 138.795 50.710 139.705 ;
        RECT 51.385 138.795 52.735 139.705 ;
        RECT 53.215 139.025 57.115 139.705 ;
        RECT 53.215 138.795 54.145 139.025 ;
        RECT 57.355 138.895 61.025 139.705 ;
        RECT 61.045 138.835 61.475 139.620 ;
        RECT 61.495 138.925 62.865 139.705 ;
        RECT 62.985 139.025 66.450 139.705 ;
        RECT 65.530 138.795 66.450 139.025 ;
        RECT 67.025 138.795 68.375 139.705 ;
        RECT 68.395 138.795 71.605 139.705 ;
        RECT 71.615 139.025 73.445 139.705 ;
        RECT 72.100 138.795 73.445 139.025 ;
        RECT 73.915 138.895 77.585 139.705 ;
        RECT 77.595 138.795 81.070 139.705 ;
        RECT 81.735 138.895 85.405 139.705 ;
        RECT 85.425 138.795 86.775 139.705 ;
        RECT 86.805 138.835 87.235 139.620 ;
        RECT 87.255 138.925 88.625 139.705 ;
        RECT 88.635 138.895 90.005 139.705 ;
        RECT 90.015 138.895 93.685 139.705 ;
        RECT 93.695 138.895 99.205 139.705 ;
        RECT 99.215 139.675 100.160 139.705 ;
        RECT 101.650 139.675 101.820 139.895 ;
        RECT 103.495 139.725 103.665 139.915 ;
        RECT 103.960 139.725 104.130 139.915 ;
        RECT 101.975 139.675 102.920 139.705 ;
        RECT 104.410 139.675 104.580 139.895 ;
        RECT 104.880 139.705 105.050 139.895 ;
        RECT 109.015 139.725 109.185 139.915 ;
        RECT 111.960 139.705 112.130 139.895 ;
        RECT 112.880 139.725 113.050 139.915 ;
        RECT 113.155 139.705 113.325 139.895 ;
        RECT 117.020 139.725 117.190 139.915 ;
        RECT 117.755 139.725 117.925 139.915 ;
        RECT 119.190 139.755 119.310 139.865 ;
        RECT 119.595 139.725 119.765 139.915 ;
        RECT 123.735 139.705 123.905 139.895 ;
        RECT 124.195 139.865 124.365 139.915 ;
        RECT 124.195 139.755 124.370 139.865 ;
        RECT 124.195 139.725 124.365 139.755 ;
        RECT 125.575 139.705 125.745 139.915 ;
        RECT 99.215 138.995 101.965 139.675 ;
        RECT 101.975 138.995 104.725 139.675 ;
        RECT 99.215 138.795 100.160 138.995 ;
        RECT 101.975 138.795 102.920 138.995 ;
        RECT 104.735 138.795 108.210 139.705 ;
        RECT 108.645 139.025 112.545 139.705 ;
        RECT 111.615 138.795 112.545 139.025 ;
        RECT 112.565 138.835 112.995 139.620 ;
        RECT 113.025 138.795 114.375 139.705 ;
        RECT 114.765 139.025 124.045 139.705 ;
        RECT 114.765 138.905 117.100 139.025 ;
        RECT 114.765 138.795 115.685 138.905 ;
        RECT 121.765 138.805 122.685 139.025 ;
        RECT 124.515 138.895 125.885 139.705 ;
      LAYER nwell ;
        RECT 11.620 135.675 126.080 138.505 ;
      LAYER pwell ;
        RECT 11.815 134.475 13.185 135.285 ;
        RECT 14.115 134.475 17.785 135.285 ;
        RECT 20.995 135.155 21.925 135.385 ;
        RECT 18.025 134.475 21.925 135.155 ;
        RECT 22.405 134.560 22.835 135.345 ;
        RECT 23.775 134.475 27.445 135.285 ;
        RECT 27.825 135.275 28.745 135.385 ;
        RECT 27.825 135.155 30.160 135.275 ;
        RECT 34.825 135.155 35.745 135.375 ;
        RECT 27.825 134.475 37.105 135.155 ;
        RECT 37.115 134.475 38.485 135.255 ;
        RECT 38.955 134.475 42.625 135.285 ;
        RECT 42.635 134.475 48.145 135.285 ;
        RECT 48.165 134.560 48.595 135.345 ;
        RECT 48.615 134.475 49.985 135.285 ;
        RECT 49.995 134.475 55.505 135.285 ;
        RECT 55.515 134.475 61.025 135.285 ;
        RECT 64.235 135.155 65.165 135.385 ;
        RECT 61.265 134.475 65.165 135.155 ;
        RECT 65.635 134.475 67.005 135.255 ;
        RECT 67.015 134.475 68.385 135.285 ;
        RECT 68.395 134.475 73.905 135.285 ;
        RECT 73.925 134.560 74.355 135.345 ;
        RECT 74.375 134.475 75.745 135.285 ;
        RECT 75.755 135.185 76.700 135.385 ;
        RECT 75.755 134.505 78.505 135.185 ;
        RECT 75.755 134.475 76.700 134.505 ;
        RECT 11.955 134.265 12.125 134.475 ;
        RECT 13.390 134.315 13.510 134.425 ;
        RECT 13.795 134.320 13.955 134.430 ;
        RECT 17.475 134.285 17.645 134.475 ;
        RECT 21.340 134.285 21.510 134.475 ;
        RECT 22.130 134.315 22.250 134.425 ;
        RECT 22.995 134.265 23.165 134.455 ;
        RECT 23.455 134.320 23.615 134.430 ;
        RECT 24.375 134.265 24.545 134.455 ;
        RECT 25.295 134.310 25.455 134.420 ;
        RECT 27.135 134.285 27.305 134.475 ;
        RECT 28.975 134.265 29.145 134.455 ;
        RECT 29.435 134.265 29.605 134.455 ;
        RECT 30.815 134.265 30.985 134.455 ;
        RECT 32.250 134.315 32.370 134.425 ;
        RECT 34.955 134.265 35.125 134.455 ;
        RECT 36.795 134.285 36.965 134.475 ;
        RECT 38.175 134.285 38.345 134.475 ;
        RECT 38.690 134.315 38.810 134.425 ;
        RECT 40.935 134.265 41.105 134.455 ;
        RECT 41.395 134.285 41.565 134.455 ;
        RECT 42.315 134.285 42.485 134.475 ;
        RECT 41.415 134.265 41.565 134.285 ;
        RECT 11.815 133.455 13.185 134.265 ;
        RECT 14.025 133.585 23.305 134.265 ;
        RECT 14.025 133.465 16.360 133.585 ;
        RECT 14.025 133.355 14.945 133.465 ;
        RECT 21.025 133.365 21.945 133.585 ;
        RECT 23.315 133.485 24.685 134.265 ;
        RECT 25.615 133.455 29.285 134.265 ;
        RECT 29.305 133.355 30.655 134.265 ;
        RECT 30.685 133.355 32.035 134.265 ;
        RECT 32.515 133.455 35.265 134.265 ;
        RECT 35.285 133.395 35.715 134.180 ;
        RECT 35.735 133.455 41.245 134.265 ;
        RECT 41.415 133.445 43.345 134.265 ;
        RECT 42.395 133.355 43.345 133.445 ;
        RECT 43.555 134.235 44.500 134.265 ;
        RECT 45.990 134.235 46.160 134.455 ;
        RECT 47.835 134.265 48.005 134.475 ;
        RECT 48.300 134.265 48.470 134.455 ;
        RECT 49.675 134.285 49.845 134.475 ;
        RECT 52.895 134.265 53.065 134.455 ;
        RECT 55.195 134.285 55.365 134.475 ;
        RECT 56.760 134.265 56.930 134.455 ;
        RECT 57.550 134.315 57.670 134.425 ;
        RECT 57.955 134.265 58.125 134.455 ;
        RECT 60.715 134.265 60.885 134.475 ;
        RECT 64.580 134.285 64.750 134.475 ;
        RECT 65.370 134.315 65.490 134.425 ;
        RECT 65.775 134.285 65.945 134.475 ;
        RECT 68.075 134.285 68.245 134.475 ;
        RECT 70.835 134.265 71.005 134.455 ;
        RECT 71.755 134.310 71.915 134.420 ;
        RECT 73.595 134.285 73.765 134.475 ;
        RECT 75.435 134.285 75.605 134.475 ;
        RECT 77.275 134.265 77.445 134.455 ;
        RECT 77.740 134.265 77.910 134.455 ;
        RECT 78.190 134.285 78.360 134.505 ;
        RECT 78.975 134.475 82.645 135.285 ;
        RECT 85.855 135.155 86.785 135.385 ;
        RECT 82.885 134.475 86.785 135.155 ;
        RECT 87.255 134.475 92.765 135.285 ;
        RECT 95.975 135.155 96.905 135.385 ;
        RECT 93.005 134.475 96.905 135.155 ;
        RECT 96.915 134.475 99.665 135.285 ;
        RECT 99.685 134.560 100.115 135.345 ;
        RECT 100.605 134.475 101.955 135.385 ;
        RECT 105.175 135.155 106.105 135.385 ;
        RECT 102.205 134.475 106.105 135.155 ;
        RECT 106.115 134.475 107.485 135.255 ;
        RECT 107.955 134.475 111.625 135.285 ;
        RECT 112.005 135.275 112.925 135.385 ;
        RECT 112.005 135.155 114.340 135.275 ;
        RECT 119.005 135.155 119.925 135.375 ;
        RECT 112.005 134.475 121.285 135.155 ;
        RECT 121.755 134.475 124.505 135.285 ;
        RECT 124.515 134.475 125.885 135.285 ;
        RECT 78.710 134.315 78.830 134.425 ;
        RECT 82.335 134.265 82.505 134.475 ;
        RECT 86.200 134.265 86.370 134.475 ;
        RECT 86.990 134.315 87.110 134.425 ;
        RECT 87.395 134.265 87.565 134.455 ;
        RECT 92.455 134.285 92.625 134.475 ;
        RECT 96.320 134.285 96.490 134.475 ;
        RECT 97.975 134.265 98.145 134.455 ;
        RECT 99.355 134.285 99.525 134.475 ;
        RECT 100.330 134.315 100.450 134.425 ;
        RECT 100.735 134.285 100.905 134.475 ;
        RECT 105.520 134.285 105.690 134.475 ;
        RECT 107.175 134.285 107.345 134.475 ;
        RECT 107.635 134.425 107.805 134.455 ;
        RECT 107.635 134.315 107.810 134.425 ;
        RECT 107.635 134.265 107.805 134.315 ;
        RECT 109.935 134.285 110.105 134.455 ;
        RECT 110.450 134.315 110.570 134.425 ;
        RECT 111.315 134.285 111.485 134.475 ;
        RECT 109.935 134.265 110.085 134.285 ;
        RECT 112.235 134.265 112.405 134.455 ;
        RECT 113.210 134.315 113.330 134.425 ;
        RECT 116.835 134.265 117.005 134.455 ;
        RECT 117.295 134.265 117.465 134.455 ;
        RECT 118.730 134.315 118.850 134.425 ;
        RECT 120.975 134.285 121.145 134.475 ;
        RECT 121.490 134.315 121.610 134.425 ;
        RECT 124.195 134.265 124.365 134.475 ;
        RECT 125.575 134.265 125.745 134.475 ;
        RECT 43.555 133.555 46.305 134.235 ;
        RECT 43.555 133.355 44.500 133.555 ;
        RECT 46.315 133.455 48.145 134.265 ;
        RECT 48.155 133.355 51.630 134.265 ;
        RECT 51.835 133.455 53.205 134.265 ;
        RECT 53.445 133.585 57.345 134.265 ;
        RECT 56.415 133.355 57.345 133.585 ;
        RECT 57.815 133.485 59.185 134.265 ;
        RECT 59.195 133.455 61.025 134.265 ;
        RECT 61.045 133.395 61.475 134.180 ;
        RECT 61.865 133.585 71.145 134.265 ;
        RECT 61.865 133.465 64.200 133.585 ;
        RECT 61.865 133.355 62.785 133.465 ;
        RECT 68.865 133.365 69.785 133.585 ;
        RECT 72.075 133.455 77.585 134.265 ;
        RECT 77.595 133.355 81.070 134.265 ;
        RECT 81.275 133.455 82.645 134.265 ;
        RECT 82.885 133.585 86.785 134.265 ;
        RECT 85.855 133.355 86.785 133.585 ;
        RECT 86.805 133.395 87.235 134.180 ;
        RECT 87.255 133.485 88.625 134.265 ;
        RECT 89.005 133.585 98.285 134.265 ;
        RECT 98.665 133.585 107.945 134.265 ;
        RECT 89.005 133.465 91.340 133.585 ;
        RECT 89.005 133.355 89.925 133.465 ;
        RECT 96.005 133.365 96.925 133.585 ;
        RECT 98.665 133.465 101.000 133.585 ;
        RECT 98.665 133.355 99.585 133.465 ;
        RECT 105.665 133.365 106.585 133.585 ;
        RECT 108.155 133.445 110.085 134.265 ;
        RECT 110.715 133.455 112.545 134.265 ;
        RECT 108.155 133.355 109.105 133.445 ;
        RECT 112.565 133.395 112.995 134.180 ;
        RECT 113.475 133.455 117.145 134.265 ;
        RECT 117.155 133.485 118.525 134.265 ;
        RECT 118.995 133.455 124.505 134.265 ;
        RECT 124.515 133.455 125.885 134.265 ;
      LAYER nwell ;
        RECT 11.620 130.235 126.080 133.065 ;
      LAYER pwell ;
        RECT 11.815 129.035 13.185 129.845 ;
        RECT 13.195 129.035 16.865 129.845 ;
        RECT 16.885 129.035 18.235 129.945 ;
        RECT 21.455 129.715 22.385 129.945 ;
        RECT 18.485 129.035 22.385 129.715 ;
        RECT 22.405 129.120 22.835 129.905 ;
        RECT 22.855 129.035 26.525 129.845 ;
        RECT 27.895 129.715 28.815 129.935 ;
        RECT 34.895 129.835 35.815 129.945 ;
        RECT 40.555 129.855 41.505 129.945 ;
        RECT 33.480 129.715 35.815 129.835 ;
        RECT 26.535 129.035 35.815 129.715 ;
        RECT 36.665 129.035 39.405 129.715 ;
        RECT 39.575 129.035 41.505 129.855 ;
        RECT 43.520 129.745 44.465 129.945 ;
        RECT 41.715 129.065 44.465 129.745 ;
        RECT 11.955 128.825 12.125 129.035 ;
        RECT 13.795 128.870 13.955 128.980 ;
        RECT 16.555 128.845 16.725 129.035 ;
        RECT 17.015 128.845 17.185 129.035 ;
        RECT 21.800 128.845 21.970 129.035 ;
        RECT 23.455 128.825 23.625 129.015 ;
        RECT 24.835 128.825 25.005 129.015 ;
        RECT 25.755 128.870 25.915 128.980 ;
        RECT 26.215 128.825 26.385 129.035 ;
        RECT 26.675 128.845 26.845 129.035 ;
        RECT 27.595 128.845 27.765 129.015 ;
        RECT 27.615 128.825 27.765 128.845 ;
        RECT 30.170 128.825 30.340 129.015 ;
        RECT 34.955 128.825 35.125 129.015 ;
        RECT 36.390 128.875 36.510 128.985 ;
        RECT 36.795 128.825 36.965 129.015 ;
        RECT 39.095 128.845 39.265 129.035 ;
        RECT 39.575 129.015 39.725 129.035 ;
        RECT 39.550 128.845 39.725 129.015 ;
        RECT 11.815 128.015 13.185 128.825 ;
        RECT 14.485 128.145 23.765 128.825 ;
        RECT 14.485 128.025 16.820 128.145 ;
        RECT 14.485 127.915 15.405 128.025 ;
        RECT 21.485 127.925 22.405 128.145 ;
        RECT 23.775 128.045 25.145 128.825 ;
        RECT 26.075 128.045 27.445 128.825 ;
        RECT 27.615 128.005 29.545 128.825 ;
        RECT 28.595 127.915 29.545 128.005 ;
        RECT 29.755 128.145 33.655 128.825 ;
        RECT 29.755 127.915 30.685 128.145 ;
        RECT 33.895 128.015 35.265 128.825 ;
        RECT 35.285 127.955 35.715 128.740 ;
        RECT 35.735 128.015 37.105 128.825 ;
        RECT 37.115 128.795 38.060 128.825 ;
        RECT 39.550 128.795 39.720 128.845 ;
        RECT 40.020 128.825 40.190 129.015 ;
        RECT 41.860 128.845 42.030 129.065 ;
        RECT 43.520 129.035 44.465 129.065 ;
        RECT 44.475 129.035 47.950 129.945 ;
        RECT 48.165 129.120 48.595 129.905 ;
        RECT 49.075 129.035 51.825 129.845 ;
        RECT 52.205 129.835 53.125 129.945 ;
        RECT 52.205 129.715 54.540 129.835 ;
        RECT 59.205 129.715 60.125 129.935 ;
        RECT 52.205 129.035 61.485 129.715 ;
        RECT 61.495 129.035 64.245 129.845 ;
        RECT 64.265 129.035 65.615 129.945 ;
        RECT 72.755 129.855 73.705 129.945 ;
        RECT 66.555 129.035 67.925 129.815 ;
        RECT 67.935 129.035 69.765 129.715 ;
        RECT 69.775 129.035 71.605 129.715 ;
        RECT 71.775 129.035 73.705 129.855 ;
        RECT 73.925 129.120 74.355 129.905 ;
        RECT 74.375 129.035 75.745 129.845 ;
        RECT 77.560 129.745 78.505 129.945 ;
        RECT 75.755 129.065 78.505 129.745 ;
        RECT 44.620 128.845 44.790 129.035 ;
        RECT 48.810 128.875 48.930 128.985 ;
        RECT 51.515 128.845 51.685 129.035 ;
        RECT 54.270 128.825 54.440 129.015 ;
        RECT 54.735 128.825 54.905 129.015 ;
        RECT 59.520 128.825 59.690 129.015 ;
        RECT 60.715 128.870 60.875 128.980 ;
        RECT 61.175 128.845 61.345 129.035 ;
        RECT 62.095 128.870 62.255 128.980 ;
        RECT 62.555 128.825 62.725 129.015 ;
        RECT 63.935 128.825 64.105 129.035 ;
        RECT 64.395 128.845 64.565 129.035 ;
        RECT 66.235 128.825 66.405 129.015 ;
        RECT 66.695 128.845 66.865 129.035 ;
        RECT 69.455 128.845 69.625 129.035 ;
        RECT 69.915 128.825 70.085 129.035 ;
        RECT 71.775 129.015 71.925 129.035 ;
        RECT 71.755 128.845 71.925 129.015 ;
        RECT 72.215 128.845 72.385 129.015 ;
        RECT 72.215 128.825 72.365 128.845 ;
        RECT 74.055 128.825 74.225 129.015 ;
        RECT 74.515 128.845 74.685 129.015 ;
        RECT 75.435 128.845 75.605 129.035 ;
        RECT 75.900 128.845 76.070 129.065 ;
        RECT 77.560 129.035 78.505 129.065 ;
        RECT 78.515 129.035 81.990 129.945 ;
        RECT 83.485 129.835 84.405 129.945 ;
        RECT 83.485 129.715 85.820 129.835 ;
        RECT 90.485 129.715 91.405 129.935 ;
        RECT 83.485 129.035 92.765 129.715 ;
        RECT 92.785 129.035 94.135 129.945 ;
        RECT 94.155 129.035 95.525 129.845 ;
        RECT 95.535 129.035 96.905 129.815 ;
        RECT 96.915 129.035 99.665 129.845 ;
        RECT 99.685 129.120 100.115 129.905 ;
        RECT 100.795 129.855 101.745 129.945 ;
        RECT 106.775 129.855 107.725 129.945 ;
        RECT 109.075 129.855 110.025 129.945 ;
        RECT 100.795 129.035 102.725 129.855 ;
        RECT 102.905 129.035 105.645 129.715 ;
        RECT 106.775 129.035 108.705 129.855 ;
        RECT 109.075 129.035 111.005 129.855 ;
        RECT 111.635 129.035 113.465 129.845 ;
        RECT 113.475 129.035 118.985 129.845 ;
        RECT 118.995 129.035 124.505 129.845 ;
        RECT 124.515 129.035 125.885 129.845 ;
        RECT 78.660 128.845 78.830 129.035 ;
        RECT 74.535 128.825 74.685 128.845 ;
        RECT 37.115 128.115 39.865 128.795 ;
        RECT 37.115 127.915 38.060 128.115 ;
        RECT 39.875 127.915 43.350 128.825 ;
        RECT 43.575 127.915 54.585 128.825 ;
        RECT 54.605 127.915 55.955 128.825 ;
        RECT 56.205 128.145 60.105 128.825 ;
        RECT 59.175 127.915 60.105 128.145 ;
        RECT 61.045 127.955 61.475 128.740 ;
        RECT 62.415 128.045 63.785 128.825 ;
        RECT 63.805 127.915 65.155 128.825 ;
        RECT 65.175 128.015 66.545 128.825 ;
        RECT 66.555 128.015 70.225 128.825 ;
        RECT 70.435 128.005 72.365 128.825 ;
        RECT 72.535 128.015 74.365 128.825 ;
        RECT 74.535 128.005 76.465 128.825 ;
        RECT 70.435 127.915 71.385 128.005 ;
        RECT 75.515 127.915 76.465 128.005 ;
        RECT 76.675 128.795 77.620 128.825 ;
        RECT 79.110 128.795 79.280 129.015 ;
        RECT 81.415 128.845 81.585 129.015 ;
        RECT 81.415 128.825 81.565 128.845 ;
        RECT 82.795 128.825 82.965 129.015 ;
        RECT 86.475 128.825 86.645 129.015 ;
        RECT 87.450 128.875 87.570 128.985 ;
        RECT 88.775 128.825 88.945 129.015 ;
        RECT 89.290 128.875 89.410 128.985 ;
        RECT 91.075 128.825 91.245 129.015 ;
        RECT 92.455 128.845 92.625 129.035 ;
        RECT 92.915 128.845 93.085 129.015 ;
        RECT 93.835 128.845 94.005 129.035 ;
        RECT 95.215 128.845 95.385 129.035 ;
        RECT 96.135 128.845 96.305 129.015 ;
        RECT 96.135 128.825 96.285 128.845 ;
        RECT 96.595 128.825 96.765 129.035 ;
        RECT 99.355 128.845 99.525 129.035 ;
        RECT 102.575 129.015 102.725 129.035 ;
        RECT 100.330 128.875 100.450 128.985 ;
        RECT 102.575 128.845 102.745 129.015 ;
        RECT 105.335 128.845 105.505 129.035 ;
        RECT 108.555 129.015 108.705 129.035 ;
        RECT 110.855 129.015 111.005 129.035 ;
        RECT 106.255 128.880 106.415 128.990 ;
        RECT 107.635 128.845 107.805 129.015 ;
        RECT 108.150 128.875 108.270 128.985 ;
        RECT 108.555 128.845 108.725 129.015 ;
        RECT 110.855 128.845 111.025 129.015 ;
        RECT 111.370 128.875 111.490 128.985 ;
        RECT 107.635 128.825 107.785 128.845 ;
        RECT 111.960 128.825 112.130 129.015 ;
        RECT 113.155 128.845 113.325 129.035 ;
        RECT 113.615 128.870 113.775 128.980 ;
        RECT 118.675 128.845 118.845 129.035 ;
        RECT 123.275 128.825 123.445 129.015 ;
        RECT 124.195 128.845 124.365 129.035 ;
        RECT 125.575 128.825 125.745 129.035 ;
        RECT 76.675 128.115 79.425 128.795 ;
        RECT 76.675 127.915 77.620 128.115 ;
        RECT 79.635 128.005 81.565 128.825 ;
        RECT 81.735 128.015 83.105 128.825 ;
        RECT 83.115 128.015 86.785 128.825 ;
        RECT 79.635 127.915 80.585 128.005 ;
        RECT 86.805 127.955 87.235 128.740 ;
        RECT 87.725 127.915 89.075 128.825 ;
        RECT 89.555 128.015 91.385 128.825 ;
        RECT 91.395 128.145 92.760 128.825 ;
        RECT 94.355 128.005 96.285 128.825 ;
        RECT 96.455 128.145 105.560 128.825 ;
        RECT 105.855 128.005 107.785 128.825 ;
        RECT 108.645 128.145 112.545 128.825 ;
        RECT 94.355 127.915 95.305 128.005 ;
        RECT 105.855 127.915 106.805 128.005 ;
        RECT 111.615 127.915 112.545 128.145 ;
        RECT 112.565 127.955 112.995 128.740 ;
        RECT 114.305 128.145 123.585 128.825 ;
        RECT 114.305 128.025 116.640 128.145 ;
        RECT 114.305 127.915 115.225 128.025 ;
        RECT 121.305 127.925 122.225 128.145 ;
        RECT 124.515 128.015 125.885 128.825 ;
      LAYER nwell ;
        RECT 11.620 124.795 126.080 127.625 ;
      LAYER pwell ;
        RECT 11.815 123.595 13.185 124.405 ;
        RECT 13.195 123.595 16.865 124.405 ;
        RECT 16.885 123.595 18.235 124.505 ;
        RECT 21.455 124.275 22.385 124.505 ;
        RECT 18.485 123.595 22.385 124.275 ;
        RECT 22.405 123.680 22.835 124.465 ;
        RECT 28.135 124.415 29.085 124.505 ;
        RECT 22.855 123.595 24.225 124.375 ;
        RECT 24.235 123.595 26.985 124.405 ;
        RECT 27.155 123.595 29.085 124.415 ;
        RECT 40.760 124.305 41.705 124.505 ;
        RECT 29.380 123.595 38.485 124.275 ;
        RECT 38.955 123.625 41.705 124.305 ;
        RECT 11.955 123.385 12.125 123.595 ;
        RECT 14.255 123.385 14.425 123.575 ;
        RECT 16.555 123.405 16.725 123.595 ;
        RECT 17.015 123.405 17.185 123.595 ;
        RECT 21.800 123.405 21.970 123.595 ;
        RECT 22.995 123.405 23.165 123.595 ;
        RECT 23.915 123.385 24.085 123.575 ;
        RECT 24.835 123.430 24.995 123.540 ;
        RECT 26.675 123.405 26.845 123.595 ;
        RECT 27.155 123.575 27.305 123.595 ;
        RECT 38.175 123.575 38.345 123.595 ;
        RECT 27.135 123.405 27.305 123.575 ;
        RECT 34.495 123.385 34.665 123.575 ;
        RECT 35.010 123.435 35.130 123.545 ;
        RECT 38.170 123.405 38.345 123.575 ;
        RECT 38.635 123.545 38.805 123.575 ;
        RECT 38.635 123.435 38.810 123.545 ;
        RECT 38.170 123.385 38.340 123.405 ;
        RECT 38.635 123.385 38.805 123.435 ;
        RECT 39.100 123.405 39.270 123.625 ;
        RECT 40.760 123.595 41.705 123.625 ;
        RECT 41.715 124.305 42.660 124.505 ;
        RECT 41.715 123.625 44.465 124.305 ;
        RECT 41.715 123.595 42.660 123.625 ;
        RECT 40.070 123.435 40.190 123.545 ;
        RECT 42.315 123.405 42.485 123.575 ;
        RECT 42.775 123.405 42.945 123.575 ;
        RECT 44.150 123.405 44.320 123.625 ;
        RECT 44.475 123.595 47.950 124.505 ;
        RECT 48.165 123.680 48.595 124.465 ;
        RECT 49.535 123.595 53.010 124.505 ;
        RECT 54.135 123.595 57.805 124.405 ;
        RECT 58.185 124.395 59.105 124.505 ;
        RECT 58.185 124.275 60.520 124.395 ;
        RECT 65.185 124.275 66.105 124.495 ;
        RECT 58.185 123.595 67.465 124.275 ;
        RECT 67.935 123.595 70.685 124.405 ;
        RECT 70.695 123.595 73.435 124.275 ;
        RECT 73.925 123.680 74.355 124.465 ;
        RECT 77.795 124.415 78.745 124.505 ;
        RECT 74.835 123.595 77.585 124.405 ;
        RECT 77.795 123.595 79.725 124.415 ;
        RECT 80.355 123.595 84.025 124.405 ;
        RECT 84.120 123.595 93.225 124.275 ;
        RECT 94.155 123.595 99.665 124.405 ;
        RECT 99.685 123.680 100.115 124.465 ;
        RECT 103.335 124.275 104.265 124.505 ;
        RECT 100.365 123.595 104.265 124.275 ;
        RECT 104.735 123.595 106.105 124.375 ;
        RECT 106.115 123.595 107.945 124.405 ;
        RECT 111.155 124.275 112.085 124.505 ;
        RECT 108.185 123.595 112.085 124.275 ;
        RECT 112.465 124.395 113.385 124.505 ;
        RECT 112.465 124.275 114.800 124.395 ;
        RECT 119.465 124.275 120.385 124.495 ;
        RECT 112.465 123.595 121.745 124.275 ;
        RECT 121.755 123.595 123.125 124.375 ;
        RECT 123.135 123.595 124.505 124.375 ;
        RECT 124.515 123.595 125.885 124.405 ;
        RECT 44.620 123.405 44.790 123.595 ;
        RECT 45.130 123.435 45.250 123.545 ;
        RECT 42.315 123.385 42.465 123.405 ;
        RECT 11.815 122.575 13.185 123.385 ;
        RECT 13.195 122.575 14.565 123.385 ;
        RECT 14.945 122.705 24.225 123.385 ;
        RECT 25.525 122.705 34.805 123.385 ;
        RECT 14.945 122.585 17.280 122.705 ;
        RECT 14.945 122.475 15.865 122.585 ;
        RECT 21.945 122.485 22.865 122.705 ;
        RECT 25.525 122.585 27.860 122.705 ;
        RECT 25.525 122.475 26.445 122.585 ;
        RECT 32.525 122.485 33.445 122.705 ;
        RECT 35.285 122.515 35.715 123.300 ;
        RECT 35.875 122.475 38.485 123.385 ;
        RECT 38.495 122.605 39.865 123.385 ;
        RECT 40.535 122.565 42.465 123.385 ;
        RECT 42.795 123.385 42.945 123.405 ;
        RECT 45.535 123.385 45.705 123.575 ;
        RECT 49.215 123.440 49.375 123.550 ;
        RECT 49.680 123.405 49.850 123.595 ;
        RECT 53.815 123.440 53.975 123.550 ;
        RECT 56.115 123.385 56.285 123.575 ;
        RECT 57.495 123.405 57.665 123.595 ;
        RECT 59.980 123.385 60.150 123.575 ;
        RECT 60.770 123.435 60.890 123.545 ;
        RECT 61.635 123.385 61.805 123.575 ;
        RECT 63.070 123.435 63.190 123.545 ;
        RECT 65.775 123.385 65.945 123.575 ;
        RECT 67.155 123.405 67.325 123.595 ;
        RECT 67.670 123.435 67.790 123.545 ;
        RECT 70.375 123.405 70.545 123.595 ;
        RECT 70.835 123.405 71.005 123.595 ;
        RECT 71.295 123.385 71.465 123.575 ;
        RECT 73.650 123.435 73.770 123.545 ;
        RECT 74.570 123.435 74.690 123.545 ;
        RECT 77.275 123.405 77.445 123.595 ;
        RECT 79.575 123.575 79.725 123.595 ;
        RECT 79.575 123.405 79.745 123.575 ;
        RECT 80.090 123.435 80.210 123.545 ;
        RECT 80.955 123.385 81.125 123.575 ;
        RECT 83.715 123.405 83.885 123.595 ;
        RECT 84.820 123.385 84.990 123.575 ;
        RECT 85.555 123.385 85.725 123.575 ;
        RECT 92.915 123.405 93.085 123.595 ;
        RECT 93.835 123.440 93.995 123.550 ;
        RECT 96.595 123.385 96.765 123.575 ;
        RECT 97.515 123.430 97.675 123.540 ;
        RECT 97.975 123.385 98.145 123.575 ;
        RECT 99.355 123.405 99.525 123.595 ;
        RECT 103.680 123.405 103.850 123.595 ;
        RECT 104.470 123.435 104.590 123.545 ;
        RECT 104.875 123.405 105.045 123.595 ;
        RECT 107.635 123.405 107.805 123.595 ;
        RECT 108.555 123.385 108.725 123.575 ;
        RECT 111.500 123.405 111.670 123.595 ;
        RECT 112.235 123.385 112.405 123.575 ;
        RECT 116.560 123.385 116.730 123.575 ;
        RECT 118.215 123.385 118.385 123.575 ;
        RECT 118.675 123.385 118.845 123.575 ;
        RECT 120.515 123.430 120.675 123.540 ;
        RECT 121.435 123.405 121.605 123.595 ;
        RECT 122.815 123.405 122.985 123.595 ;
        RECT 124.195 123.385 124.365 123.595 ;
        RECT 125.575 123.385 125.745 123.595 ;
        RECT 42.795 122.565 44.725 123.385 ;
        RECT 45.395 122.705 54.500 123.385 ;
        RECT 54.595 122.575 56.425 123.385 ;
        RECT 56.665 122.705 60.565 123.385 ;
        RECT 40.535 122.475 41.485 122.565 ;
        RECT 43.775 122.475 44.725 122.565 ;
        RECT 59.635 122.475 60.565 122.705 ;
        RECT 61.045 122.515 61.475 123.300 ;
        RECT 61.495 122.605 62.865 123.385 ;
        RECT 63.335 122.575 66.085 123.385 ;
        RECT 66.095 122.575 71.605 123.385 ;
        RECT 71.985 122.705 81.265 123.385 ;
        RECT 81.505 122.705 85.405 123.385 ;
        RECT 71.985 122.585 74.320 122.705 ;
        RECT 71.985 122.475 72.905 122.585 ;
        RECT 78.985 122.485 79.905 122.705 ;
        RECT 84.475 122.475 85.405 122.705 ;
        RECT 85.425 122.475 86.775 123.385 ;
        RECT 86.805 122.515 87.235 123.300 ;
        RECT 87.625 122.705 96.905 123.385 ;
        RECT 87.625 122.585 89.960 122.705 ;
        RECT 87.625 122.475 88.545 122.585 ;
        RECT 94.625 122.485 95.545 122.705 ;
        RECT 97.845 122.475 99.195 123.385 ;
        RECT 99.585 122.705 108.865 123.385 ;
        RECT 99.585 122.585 101.920 122.705 ;
        RECT 99.585 122.475 100.505 122.585 ;
        RECT 106.585 122.485 107.505 122.705 ;
        RECT 108.875 122.575 112.545 123.385 ;
        RECT 112.565 122.515 112.995 123.300 ;
        RECT 113.245 122.705 117.145 123.385 ;
        RECT 116.215 122.475 117.145 122.705 ;
        RECT 117.165 122.475 118.515 123.385 ;
        RECT 118.545 122.475 119.895 123.385 ;
        RECT 120.835 122.575 124.505 123.385 ;
        RECT 124.515 122.575 125.885 123.385 ;
      LAYER nwell ;
        RECT 11.620 119.355 126.080 122.185 ;
      LAYER pwell ;
        RECT 11.815 118.155 13.185 118.965 ;
        RECT 13.655 118.155 15.485 118.965 ;
        RECT 15.505 118.155 16.855 119.065 ;
        RECT 16.885 118.155 18.235 119.065 ;
        RECT 21.455 118.835 22.385 119.065 ;
        RECT 18.485 118.155 22.385 118.835 ;
        RECT 22.405 118.240 22.835 119.025 ;
        RECT 22.855 118.155 24.225 118.935 ;
        RECT 24.705 118.155 26.055 119.065 ;
        RECT 26.085 118.155 27.435 119.065 ;
        RECT 30.655 118.835 31.585 119.065 ;
        RECT 27.685 118.155 31.585 118.835 ;
        RECT 31.965 118.955 32.885 119.065 ;
        RECT 31.965 118.835 34.300 118.955 ;
        RECT 38.965 118.835 39.885 119.055 ;
        RECT 31.965 118.155 41.245 118.835 ;
        RECT 41.255 118.155 42.625 118.965 ;
        RECT 42.635 118.155 48.145 118.965 ;
        RECT 48.165 118.240 48.595 119.025 ;
        RECT 49.545 118.155 50.895 119.065 ;
        RECT 54.115 118.835 55.045 119.065 ;
        RECT 51.145 118.155 55.045 118.835 ;
        RECT 55.055 118.155 56.425 118.965 ;
        RECT 56.805 118.955 57.725 119.065 ;
        RECT 56.805 118.835 59.140 118.955 ;
        RECT 63.805 118.835 64.725 119.055 ;
        RECT 56.805 118.155 66.085 118.835 ;
        RECT 66.555 118.155 68.385 118.965 ;
        RECT 68.405 118.155 69.755 119.065 ;
        RECT 72.975 118.835 73.905 119.065 ;
        RECT 70.005 118.155 73.905 118.835 ;
        RECT 73.925 118.240 74.355 119.025 ;
        RECT 78.035 118.835 78.965 119.065 ;
        RECT 75.065 118.155 78.965 118.835 ;
        RECT 78.985 118.155 80.335 119.065 ;
        RECT 80.365 118.155 81.715 119.065 ;
        RECT 82.565 118.955 83.485 119.065 ;
        RECT 82.565 118.835 84.900 118.955 ;
        RECT 89.565 118.835 90.485 119.055 ;
        RECT 95.055 118.835 95.985 119.065 ;
        RECT 82.565 118.155 91.845 118.835 ;
        RECT 92.085 118.155 95.985 118.835 ;
        RECT 95.995 118.155 97.365 118.935 ;
        RECT 98.295 118.155 99.665 118.935 ;
        RECT 99.685 118.240 100.115 119.025 ;
        RECT 100.135 118.835 101.065 119.065 ;
        RECT 100.135 118.155 104.035 118.835 ;
        RECT 104.285 118.155 105.635 119.065 ;
        RECT 108.855 118.835 109.785 119.065 ;
        RECT 105.885 118.155 109.785 118.835 ;
        RECT 110.255 118.155 113.005 118.965 ;
        RECT 113.385 118.955 114.305 119.065 ;
        RECT 113.385 118.835 115.720 118.955 ;
        RECT 120.385 118.835 121.305 119.055 ;
        RECT 113.385 118.155 122.665 118.835 ;
        RECT 122.675 118.155 124.505 118.965 ;
        RECT 124.515 118.155 125.885 118.965 ;
        RECT 11.955 117.945 12.125 118.155 ;
        RECT 13.390 117.995 13.510 118.105 ;
        RECT 15.175 117.965 15.345 118.155 ;
        RECT 15.635 117.945 15.805 118.155 ;
        RECT 17.015 117.965 17.185 118.155 ;
        RECT 21.800 117.965 21.970 118.155 ;
        RECT 23.915 117.965 24.085 118.155 ;
        RECT 24.430 117.995 24.550 118.105 ;
        RECT 24.835 117.965 25.005 118.155 ;
        RECT 25.295 117.945 25.465 118.135 ;
        RECT 25.810 117.995 25.930 118.105 ;
        RECT 26.215 117.965 26.385 118.155 ;
        RECT 29.435 117.945 29.605 118.135 ;
        RECT 29.895 117.945 30.065 118.135 ;
        RECT 31.000 117.965 31.170 118.155 ;
        RECT 34.680 117.945 34.850 118.135 ;
        RECT 36.795 117.945 36.965 118.135 ;
        RECT 40.475 117.945 40.645 118.135 ;
        RECT 40.935 117.965 41.105 118.155 ;
        RECT 42.315 117.965 42.485 118.155 ;
        RECT 45.995 117.945 46.165 118.135 ;
        RECT 47.375 117.945 47.545 118.135 ;
        RECT 47.835 117.965 48.005 118.155 ;
        RECT 49.215 118.000 49.375 118.110 ;
        RECT 50.595 117.965 50.765 118.155 ;
        RECT 54.460 117.965 54.630 118.155 ;
        RECT 56.115 117.965 56.285 118.155 ;
        RECT 57.035 117.945 57.205 118.135 ;
        RECT 57.550 117.995 57.670 118.105 ;
        RECT 59.335 117.945 59.505 118.135 ;
        RECT 59.795 117.945 59.965 118.135 ;
        RECT 65.040 117.945 65.210 118.135 ;
        RECT 65.775 117.945 65.945 118.155 ;
        RECT 66.290 117.995 66.410 118.105 ;
        RECT 67.615 117.990 67.775 118.100 ;
        RECT 68.075 117.965 68.245 118.155 ;
        RECT 68.535 117.965 68.705 118.155 ;
        RECT 71.295 117.945 71.465 118.135 ;
        RECT 73.320 117.965 73.490 118.155 ;
        RECT 74.570 117.995 74.690 118.105 ;
        RECT 78.380 117.965 78.550 118.155 ;
        RECT 80.035 117.965 80.205 118.155 ;
        RECT 80.955 117.945 81.125 118.135 ;
        RECT 81.415 117.965 81.585 118.155 ;
        RECT 81.930 117.995 82.050 118.105 ;
        RECT 82.335 117.945 82.505 118.135 ;
        RECT 85.095 117.945 85.265 118.135 ;
        RECT 85.555 117.945 85.725 118.135 ;
        RECT 87.395 117.945 87.565 118.135 ;
        RECT 88.775 117.945 88.945 118.135 ;
        RECT 90.210 117.995 90.330 118.105 ;
        RECT 91.535 117.965 91.705 118.155 ;
        RECT 95.400 117.965 95.570 118.155 ;
        RECT 97.055 117.965 97.225 118.155 ;
        RECT 97.975 118.000 98.135 118.110 ;
        RECT 99.355 117.965 99.525 118.155 ;
        RECT 99.815 117.945 99.985 118.135 ;
        RECT 100.550 117.965 100.720 118.155 ;
        RECT 100.735 117.990 100.895 118.100 ;
        RECT 104.415 117.965 104.585 118.155 ;
        RECT 109.200 117.965 109.370 118.155 ;
        RECT 109.990 117.995 110.110 118.105 ;
        RECT 110.395 117.945 110.565 118.135 ;
        RECT 111.775 117.945 111.945 118.135 ;
        RECT 112.290 117.995 112.410 118.105 ;
        RECT 112.695 117.965 112.865 118.155 ;
        RECT 113.210 117.995 113.330 118.105 ;
        RECT 115.915 117.945 116.085 118.135 ;
        RECT 116.375 117.945 116.545 118.135 ;
        RECT 117.810 117.995 117.930 118.105 ;
        RECT 118.215 117.945 118.385 118.135 ;
        RECT 120.515 117.945 120.685 118.135 ;
        RECT 122.355 117.965 122.525 118.155 ;
        RECT 124.195 117.945 124.365 118.155 ;
        RECT 125.575 117.945 125.745 118.155 ;
        RECT 11.815 117.135 13.185 117.945 ;
        RECT 13.195 117.135 15.945 117.945 ;
        RECT 16.325 117.265 25.605 117.945 ;
        RECT 16.325 117.145 18.660 117.265 ;
        RECT 16.325 117.035 17.245 117.145 ;
        RECT 23.325 117.045 24.245 117.265 ;
        RECT 26.075 117.135 29.745 117.945 ;
        RECT 29.755 117.165 31.125 117.945 ;
        RECT 31.365 117.265 35.265 117.945 ;
        RECT 34.335 117.035 35.265 117.265 ;
        RECT 35.285 117.075 35.715 117.860 ;
        RECT 35.735 117.135 37.105 117.945 ;
        RECT 37.115 117.135 40.785 117.945 ;
        RECT 40.795 117.135 46.305 117.945 ;
        RECT 46.315 117.165 47.685 117.945 ;
        RECT 48.065 117.265 57.345 117.945 ;
        RECT 48.065 117.145 50.400 117.265 ;
        RECT 48.065 117.035 48.985 117.145 ;
        RECT 55.065 117.045 55.985 117.265 ;
        RECT 57.815 117.135 59.645 117.945 ;
        RECT 59.665 117.035 61.015 117.945 ;
        RECT 61.045 117.075 61.475 117.860 ;
        RECT 61.725 117.265 65.625 117.945 ;
        RECT 64.695 117.035 65.625 117.265 ;
        RECT 65.635 117.165 67.005 117.945 ;
        RECT 67.935 117.135 71.605 117.945 ;
        RECT 71.985 117.265 81.265 117.945 ;
        RECT 71.985 117.145 74.320 117.265 ;
        RECT 71.985 117.035 72.905 117.145 ;
        RECT 78.985 117.045 79.905 117.265 ;
        RECT 81.275 117.165 82.645 117.945 ;
        RECT 82.655 117.135 85.405 117.945 ;
        RECT 85.415 117.165 86.785 117.945 ;
        RECT 86.805 117.075 87.235 117.860 ;
        RECT 87.265 117.035 88.615 117.945 ;
        RECT 88.645 117.035 89.995 117.945 ;
        RECT 90.845 117.265 100.125 117.945 ;
        RECT 101.425 117.265 110.705 117.945 ;
        RECT 90.845 117.145 93.180 117.265 ;
        RECT 90.845 117.035 91.765 117.145 ;
        RECT 97.845 117.045 98.765 117.265 ;
        RECT 101.425 117.145 103.760 117.265 ;
        RECT 101.425 117.035 102.345 117.145 ;
        RECT 108.425 117.045 109.345 117.265 ;
        RECT 110.715 117.165 112.085 117.945 ;
        RECT 112.565 117.075 112.995 117.860 ;
        RECT 113.475 117.135 116.225 117.945 ;
        RECT 116.245 117.035 117.595 117.945 ;
        RECT 118.075 117.165 119.445 117.945 ;
        RECT 119.455 117.135 120.825 117.945 ;
        RECT 120.835 117.135 124.505 117.945 ;
        RECT 124.515 117.135 125.885 117.945 ;
      LAYER nwell ;
        RECT 11.620 113.915 126.080 116.745 ;
      LAYER pwell ;
        RECT 11.815 112.715 13.185 113.525 ;
        RECT 13.195 112.715 16.865 113.525 ;
        RECT 16.875 112.715 22.385 113.525 ;
        RECT 22.405 112.800 22.835 113.585 ;
        RECT 22.855 112.715 24.685 113.525 ;
        RECT 24.695 112.715 26.065 113.495 ;
        RECT 26.535 112.715 30.205 113.525 ;
        RECT 30.215 112.715 35.725 113.525 ;
        RECT 35.735 112.715 41.245 113.525 ;
        RECT 41.255 112.715 46.765 113.525 ;
        RECT 46.785 112.715 48.135 113.625 ;
        RECT 48.165 112.800 48.595 113.585 ;
        RECT 49.535 113.395 50.465 113.625 ;
        RECT 49.535 112.715 53.435 113.395 ;
        RECT 54.135 112.715 55.505 113.495 ;
        RECT 55.515 112.715 56.885 113.525 ;
        RECT 56.895 112.715 60.565 113.525 ;
        RECT 60.945 113.515 61.865 113.625 ;
        RECT 60.945 113.395 63.280 113.515 ;
        RECT 67.945 113.395 68.865 113.615 ;
        RECT 60.945 112.715 70.225 113.395 ;
        RECT 70.235 112.715 73.905 113.525 ;
        RECT 73.925 112.800 74.355 113.585 ;
        RECT 74.375 112.715 78.045 113.525 ;
        RECT 78.055 112.715 79.425 113.495 ;
        RECT 79.435 112.715 83.105 113.525 ;
        RECT 83.115 112.715 88.625 113.525 ;
        RECT 88.635 112.715 94.145 113.525 ;
        RECT 94.155 112.715 99.665 113.525 ;
        RECT 99.685 112.800 100.115 113.585 ;
        RECT 100.135 112.715 101.505 113.525 ;
        RECT 101.515 112.715 105.185 113.525 ;
        RECT 105.195 112.715 110.705 113.525 ;
        RECT 110.715 112.715 116.225 113.525 ;
        RECT 116.245 112.715 117.595 113.625 ;
        RECT 117.615 112.715 118.985 113.495 ;
        RECT 118.995 112.715 120.365 113.495 ;
        RECT 120.375 112.715 123.125 113.525 ;
        RECT 123.135 112.715 124.505 113.495 ;
        RECT 124.515 112.715 125.885 113.525 ;
        RECT 11.955 112.505 12.125 112.715 ;
        RECT 16.555 112.505 16.725 112.715 ;
        RECT 22.075 112.525 22.245 112.715 ;
        RECT 24.375 112.525 24.545 112.715 ;
        RECT 24.835 112.525 25.005 112.715 ;
        RECT 26.270 112.555 26.390 112.665 ;
        RECT 27.135 112.505 27.305 112.695 ;
        RECT 28.515 112.505 28.685 112.695 ;
        RECT 29.895 112.505 30.065 112.715 ;
        RECT 31.275 112.505 31.445 112.695 ;
        RECT 32.195 112.550 32.355 112.660 ;
        RECT 33.575 112.505 33.745 112.695 ;
        RECT 34.035 112.505 34.205 112.695 ;
        RECT 35.415 112.525 35.585 112.715 ;
        RECT 35.930 112.555 36.050 112.665 ;
        RECT 38.630 112.505 38.800 112.695 ;
        RECT 39.150 112.555 39.270 112.665 ;
        RECT 39.555 112.505 39.725 112.695 ;
        RECT 40.935 112.525 41.105 112.715 ;
        RECT 41.855 112.505 42.025 112.695 ;
        RECT 42.370 112.555 42.490 112.665 ;
        RECT 42.775 112.505 42.945 112.695 ;
        RECT 44.210 112.555 44.330 112.665 ;
        RECT 44.615 112.505 44.785 112.695 ;
        RECT 46.455 112.525 46.625 112.715 ;
        RECT 46.915 112.525 47.085 112.715 ;
        RECT 49.215 112.560 49.375 112.670 ;
        RECT 49.950 112.525 50.120 112.715 ;
        RECT 53.870 112.555 53.990 112.665 ;
        RECT 54.275 112.525 54.445 112.715 ;
        RECT 55.195 112.505 55.365 112.695 ;
        RECT 56.575 112.525 56.745 112.715 ;
        RECT 60.255 112.525 60.425 112.715 ;
        RECT 60.715 112.505 60.885 112.695 ;
        RECT 61.635 112.505 61.805 112.695 ;
        RECT 63.935 112.505 64.105 112.695 ;
        RECT 65.315 112.505 65.485 112.695 ;
        RECT 65.830 112.555 65.950 112.665 ;
        RECT 68.535 112.505 68.705 112.695 ;
        RECT 69.915 112.525 70.085 112.715 ;
        RECT 73.595 112.525 73.765 112.715 ;
        RECT 74.055 112.505 74.225 112.695 ;
        RECT 74.515 112.505 74.685 112.695 ;
        RECT 75.900 112.505 76.070 112.695 ;
        RECT 77.735 112.525 77.905 112.715 ;
        RECT 78.195 112.525 78.365 112.715 ;
        RECT 80.955 112.505 81.125 112.695 ;
        RECT 82.795 112.525 82.965 112.715 ;
        RECT 86.475 112.505 86.645 112.695 ;
        RECT 87.855 112.550 88.015 112.660 ;
        RECT 88.315 112.525 88.485 112.715 ;
        RECT 91.535 112.505 91.705 112.695 ;
        RECT 93.835 112.525 94.005 112.715 ;
        RECT 97.055 112.505 97.225 112.695 ;
        RECT 97.515 112.505 97.685 112.695 ;
        RECT 99.355 112.525 99.525 112.715 ;
        RECT 101.195 112.505 101.365 112.715 ;
        RECT 101.655 112.505 101.825 112.695 ;
        RECT 103.495 112.550 103.655 112.660 ;
        RECT 103.955 112.505 104.125 112.695 ;
        RECT 104.875 112.525 105.045 112.715 ;
        RECT 106.255 112.505 106.425 112.695 ;
        RECT 106.715 112.505 106.885 112.695 ;
        RECT 108.150 112.555 108.270 112.665 ;
        RECT 110.395 112.525 110.565 112.715 ;
        RECT 110.855 112.505 111.025 112.695 ;
        RECT 111.315 112.505 111.485 112.695 ;
        RECT 113.615 112.550 113.775 112.660 ;
        RECT 114.075 112.505 114.245 112.695 ;
        RECT 115.915 112.525 116.085 112.715 ;
        RECT 116.375 112.525 116.545 112.715 ;
        RECT 118.675 112.525 118.845 112.715 ;
        RECT 119.135 112.525 119.305 112.715 ;
        RECT 122.815 112.525 122.985 112.715 ;
        RECT 124.185 112.525 124.355 112.715 ;
        RECT 125.575 112.505 125.745 112.715 ;
        RECT 11.815 111.695 13.185 112.505 ;
        RECT 13.195 111.695 16.865 112.505 ;
        RECT 17.075 111.825 27.445 112.505 ;
        RECT 17.075 111.595 19.285 111.825 ;
        RECT 22.005 111.605 22.935 111.825 ;
        RECT 27.455 111.695 28.825 112.505 ;
        RECT 28.835 111.725 30.205 112.505 ;
        RECT 30.225 111.595 31.575 112.505 ;
        RECT 32.515 111.725 33.885 112.505 ;
        RECT 33.895 111.725 35.265 112.505 ;
        RECT 35.285 111.635 35.715 112.420 ;
        RECT 36.335 111.595 38.945 112.505 ;
        RECT 39.425 111.595 40.775 112.505 ;
        RECT 40.795 111.725 42.165 112.505 ;
        RECT 42.635 111.725 44.005 112.505 ;
        RECT 44.475 111.825 53.755 112.505 ;
        RECT 45.835 111.605 46.755 111.825 ;
        RECT 51.420 111.705 53.755 111.825 ;
        RECT 52.835 111.595 53.755 111.705 ;
        RECT 54.135 111.695 55.505 112.505 ;
        RECT 55.515 111.695 61.025 112.505 ;
        RECT 61.045 111.635 61.475 112.420 ;
        RECT 61.495 111.725 62.865 112.505 ;
        RECT 62.875 111.695 64.245 112.505 ;
        RECT 64.265 111.595 65.615 112.505 ;
        RECT 66.095 111.695 68.845 112.505 ;
        RECT 68.855 111.695 74.365 112.505 ;
        RECT 74.375 111.725 75.745 112.505 ;
        RECT 75.755 111.595 78.365 112.505 ;
        RECT 78.515 111.695 81.265 112.505 ;
        RECT 81.275 111.695 86.785 112.505 ;
        RECT 86.805 111.635 87.235 112.420 ;
        RECT 88.175 111.695 91.845 112.505 ;
        RECT 91.855 111.695 97.365 112.505 ;
        RECT 97.375 111.725 98.745 112.505 ;
        RECT 98.755 111.695 101.505 112.505 ;
        RECT 101.525 111.595 102.875 112.505 ;
        RECT 103.815 111.725 105.185 112.505 ;
        RECT 105.205 111.595 106.555 112.505 ;
        RECT 106.575 111.725 107.945 112.505 ;
        RECT 108.415 111.695 111.165 112.505 ;
        RECT 111.185 111.595 112.535 112.505 ;
        RECT 112.565 111.635 112.995 112.420 ;
        RECT 113.935 111.825 124.305 112.505 ;
        RECT 118.445 111.605 119.375 111.825 ;
        RECT 122.095 111.595 124.305 111.825 ;
        RECT 124.515 111.695 125.885 112.505 ;
      LAYER nwell ;
        RECT 11.620 108.475 126.080 111.305 ;
      LAYER pwell ;
        RECT 11.815 107.275 13.185 108.085 ;
        RECT 13.195 107.275 18.705 108.085 ;
        RECT 18.725 107.275 20.075 108.185 ;
        RECT 21.025 107.275 22.375 108.185 ;
        RECT 22.405 107.360 22.835 108.145 ;
        RECT 22.855 107.275 24.225 108.085 ;
        RECT 24.245 107.275 25.595 108.185 ;
        RECT 25.815 107.955 28.025 108.185 ;
        RECT 30.745 107.955 31.675 108.175 ;
        RECT 36.395 107.955 38.605 108.185 ;
        RECT 41.325 107.955 42.255 108.175 ;
        RECT 25.815 107.275 36.185 107.955 ;
        RECT 36.395 107.275 46.765 107.955 ;
        RECT 46.775 107.275 48.145 108.055 ;
        RECT 48.165 107.360 48.595 108.145 ;
        RECT 48.615 107.275 50.445 108.085 ;
        RECT 50.455 107.275 51.825 108.055 ;
        RECT 52.295 107.275 55.045 108.085 ;
        RECT 55.065 107.275 56.415 108.185 ;
        RECT 56.635 107.955 58.845 108.185 ;
        RECT 61.565 107.955 62.495 108.175 ;
        RECT 56.635 107.275 67.005 107.955 ;
        RECT 67.015 107.275 68.385 108.055 ;
        RECT 68.855 107.275 72.525 108.085 ;
        RECT 72.535 107.275 73.905 108.055 ;
        RECT 73.925 107.360 74.355 108.145 ;
        RECT 74.575 107.955 76.785 108.185 ;
        RECT 79.505 107.955 80.435 108.175 ;
        RECT 74.575 107.275 84.945 107.955 ;
        RECT 84.955 107.275 86.325 108.055 ;
        RECT 86.335 107.275 87.705 108.085 ;
        RECT 87.715 107.275 89.085 108.055 ;
        RECT 89.295 107.955 91.505 108.185 ;
        RECT 94.225 107.955 95.155 108.175 ;
        RECT 89.295 107.275 99.665 107.955 ;
        RECT 99.685 107.360 100.115 108.145 ;
        RECT 100.795 107.955 103.005 108.185 ;
        RECT 105.725 107.955 106.655 108.175 ;
        RECT 100.795 107.275 111.165 107.955 ;
        RECT 111.175 107.275 112.545 108.055 ;
        RECT 113.675 107.955 115.885 108.185 ;
        RECT 118.605 107.955 119.535 108.175 ;
        RECT 113.675 107.275 124.045 107.955 ;
        RECT 124.515 107.275 125.885 108.085 ;
        RECT 11.955 107.065 12.125 107.275 ;
        RECT 13.795 107.110 13.955 107.220 ;
        RECT 18.395 107.085 18.565 107.275 ;
        RECT 19.775 107.085 19.945 107.275 ;
        RECT 20.695 107.120 20.855 107.230 ;
        RECT 22.075 107.085 22.245 107.275 ;
        RECT 23.915 107.085 24.085 107.275 ;
        RECT 24.375 107.065 24.545 107.255 ;
        RECT 24.835 107.065 25.005 107.255 ;
        RECT 25.295 107.085 25.465 107.275 ;
        RECT 35.875 107.225 36.045 107.275 ;
        RECT 35.875 107.115 36.050 107.225 ;
        RECT 35.875 107.085 36.045 107.115 ;
        RECT 37.255 107.065 37.425 107.255 ;
        RECT 37.770 107.115 37.890 107.225 ;
        RECT 39.555 107.065 39.725 107.255 ;
        RECT 40.015 107.065 40.185 107.255 ;
        RECT 46.455 107.085 46.625 107.275 ;
        RECT 46.915 107.085 47.085 107.275 ;
        RECT 50.135 107.085 50.305 107.275 ;
        RECT 50.595 107.065 50.765 107.275 ;
        RECT 52.030 107.115 52.150 107.225 ;
        RECT 54.735 107.085 54.905 107.275 ;
        RECT 55.195 107.085 55.365 107.275 ;
        RECT 66.695 107.085 66.865 107.275 ;
        RECT 67.155 107.085 67.325 107.275 ;
        RECT 68.590 107.115 68.710 107.225 ;
        RECT 71.755 107.065 71.925 107.255 ;
        RECT 72.215 107.085 72.385 107.275 ;
        RECT 72.675 107.085 72.845 107.275 ;
        RECT 82.335 107.065 82.505 107.255 ;
        RECT 83.715 107.065 83.885 107.255 ;
        RECT 84.635 107.085 84.805 107.275 ;
        RECT 85.095 107.065 85.265 107.255 ;
        RECT 85.555 107.065 85.725 107.255 ;
        RECT 86.015 107.085 86.185 107.275 ;
        RECT 87.395 107.065 87.565 107.275 ;
        RECT 87.855 107.085 88.025 107.275 ;
        RECT 99.355 107.085 99.525 107.275 ;
        RECT 100.330 107.115 100.450 107.225 ;
        RECT 108.095 107.065 108.265 107.255 ;
        RECT 108.610 107.115 108.730 107.225 ;
        RECT 110.855 107.085 111.025 107.275 ;
        RECT 111.315 107.085 111.485 107.275 ;
        RECT 112.235 107.065 112.405 107.255 ;
        RECT 113.155 107.120 113.315 107.230 ;
        RECT 123.275 107.065 123.445 107.255 ;
        RECT 123.735 107.085 123.905 107.275 ;
        RECT 124.250 107.220 124.370 107.225 ;
        RECT 124.195 107.115 124.370 107.220 ;
        RECT 124.195 107.110 124.355 107.115 ;
        RECT 125.575 107.065 125.745 107.275 ;
        RECT 11.815 106.255 13.185 107.065 ;
        RECT 14.315 106.385 24.685 107.065 ;
        RECT 24.695 106.385 35.065 107.065 ;
        RECT 14.315 106.155 16.525 106.385 ;
        RECT 19.245 106.165 20.175 106.385 ;
        RECT 29.205 106.165 30.135 106.385 ;
        RECT 32.855 106.155 35.065 106.385 ;
        RECT 35.285 106.195 35.715 106.980 ;
        RECT 36.205 106.155 37.555 107.065 ;
        RECT 38.035 106.255 39.865 107.065 ;
        RECT 39.875 106.385 50.245 107.065 ;
        RECT 50.455 106.385 60.825 107.065 ;
        RECT 44.385 106.165 45.315 106.385 ;
        RECT 48.035 106.155 50.245 106.385 ;
        RECT 54.965 106.165 55.895 106.385 ;
        RECT 58.615 106.155 60.825 106.385 ;
        RECT 61.045 106.195 61.475 106.980 ;
        RECT 61.695 106.385 72.065 107.065 ;
        RECT 72.275 106.385 82.645 107.065 ;
        RECT 61.695 106.155 63.905 106.385 ;
        RECT 66.625 106.165 67.555 106.385 ;
        RECT 72.275 106.155 74.485 106.385 ;
        RECT 77.205 106.165 78.135 106.385 ;
        RECT 82.655 106.255 84.025 107.065 ;
        RECT 84.045 106.155 85.395 107.065 ;
        RECT 85.425 106.155 86.775 107.065 ;
        RECT 86.805 106.195 87.235 106.980 ;
        RECT 87.255 106.385 97.625 107.065 ;
        RECT 91.765 106.165 92.695 106.385 ;
        RECT 95.415 106.155 97.625 106.385 ;
        RECT 98.035 106.385 108.405 107.065 ;
        RECT 98.035 106.155 100.245 106.385 ;
        RECT 102.965 106.165 103.895 106.385 ;
        RECT 108.875 106.255 112.545 107.065 ;
        RECT 112.565 106.195 112.995 106.980 ;
        RECT 113.215 106.385 123.585 107.065 ;
        RECT 113.215 106.155 115.425 106.385 ;
        RECT 118.145 106.165 119.075 106.385 ;
        RECT 124.515 106.255 125.885 107.065 ;
      LAYER nwell ;
        RECT 11.620 103.035 126.080 105.865 ;
      LAYER pwell ;
        RECT 11.815 101.835 13.185 102.645 ;
        RECT 13.195 101.835 16.865 102.645 ;
        RECT 16.875 101.835 22.385 102.645 ;
        RECT 22.405 101.920 22.835 102.705 ;
        RECT 23.055 102.515 25.265 102.745 ;
        RECT 27.985 102.515 28.915 102.735 ;
        RECT 23.055 101.835 33.425 102.515 ;
        RECT 33.435 101.835 35.265 102.645 ;
        RECT 35.285 101.920 35.715 102.705 ;
        RECT 35.735 101.835 41.245 102.645 ;
        RECT 41.255 101.835 46.765 102.645 ;
        RECT 46.785 101.835 48.135 102.745 ;
        RECT 48.165 101.920 48.595 102.705 ;
        RECT 48.615 101.835 54.125 102.645 ;
        RECT 54.135 101.835 59.645 102.645 ;
        RECT 59.665 101.835 61.015 102.745 ;
        RECT 61.045 101.920 61.475 102.705 ;
        RECT 61.965 101.835 63.315 102.745 ;
        RECT 63.335 101.835 67.005 102.645 ;
        RECT 67.015 101.835 72.525 102.645 ;
        RECT 72.545 101.835 73.895 102.745 ;
        RECT 73.925 101.920 74.355 102.705 ;
        RECT 74.845 101.835 76.195 102.745 ;
        RECT 76.415 102.515 78.625 102.745 ;
        RECT 81.345 102.515 82.275 102.735 ;
        RECT 76.415 101.835 86.785 102.515 ;
        RECT 86.805 101.920 87.235 102.705 ;
        RECT 87.255 101.835 89.085 102.645 ;
        RECT 89.095 101.835 94.605 102.645 ;
        RECT 94.625 101.835 95.975 102.745 ;
        RECT 95.995 101.835 99.665 102.645 ;
        RECT 99.685 101.920 100.115 102.705 ;
        RECT 100.135 101.835 101.505 102.645 ;
        RECT 101.515 101.835 107.025 102.645 ;
        RECT 107.035 101.835 112.545 102.645 ;
        RECT 112.565 101.920 112.995 102.705 ;
        RECT 113.015 101.835 116.685 102.645 ;
        RECT 116.705 101.835 118.055 102.745 ;
        RECT 118.995 101.835 124.505 102.645 ;
        RECT 124.515 101.835 125.885 102.645 ;
        RECT 11.955 101.645 12.125 101.835 ;
        RECT 16.555 101.645 16.725 101.835 ;
        RECT 22.075 101.645 22.245 101.835 ;
        RECT 33.115 101.645 33.285 101.835 ;
        RECT 34.955 101.645 35.125 101.835 ;
        RECT 40.935 101.645 41.105 101.835 ;
        RECT 46.455 101.645 46.625 101.835 ;
        RECT 47.835 101.645 48.005 101.835 ;
        RECT 53.815 101.645 53.985 101.835 ;
        RECT 59.335 101.645 59.505 101.835 ;
        RECT 59.795 101.645 59.965 101.835 ;
        RECT 61.690 101.675 61.810 101.785 ;
        RECT 62.095 101.645 62.265 101.835 ;
        RECT 66.695 101.645 66.865 101.835 ;
        RECT 72.215 101.645 72.385 101.835 ;
        RECT 73.595 101.645 73.765 101.835 ;
        RECT 74.570 101.675 74.690 101.785 ;
        RECT 74.975 101.645 75.145 101.835 ;
        RECT 86.475 101.645 86.645 101.835 ;
        RECT 88.775 101.645 88.945 101.835 ;
        RECT 94.295 101.645 94.465 101.835 ;
        RECT 95.675 101.645 95.845 101.835 ;
        RECT 99.355 101.645 99.525 101.835 ;
        RECT 101.195 101.645 101.365 101.835 ;
        RECT 106.715 101.645 106.885 101.835 ;
        RECT 112.235 101.645 112.405 101.835 ;
        RECT 116.375 101.645 116.545 101.835 ;
        RECT 116.835 101.645 117.005 101.835 ;
        RECT 118.675 101.680 118.835 101.790 ;
        RECT 124.195 101.645 124.365 101.835 ;
        RECT 125.575 101.645 125.745 101.835 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 11.810 215.885 125.890 216.055 ;
        RECT 11.895 215.135 13.105 215.885 ;
        RECT 11.895 214.595 12.415 215.135 ;
        RECT 13.275 215.115 16.785 215.885 ;
        RECT 16.960 215.340 22.305 215.885 ;
        RECT 12.585 214.425 13.105 214.965 ;
        RECT 11.895 213.335 13.105 214.425 ;
        RECT 13.275 214.425 14.965 214.945 ;
        RECT 15.135 214.595 16.785 215.115 ;
        RECT 13.275 213.335 16.785 214.425 ;
        RECT 18.550 213.770 18.900 215.020 ;
        RECT 20.380 214.510 20.720 215.340 ;
        RECT 22.475 215.160 22.765 215.885 ;
        RECT 22.935 215.135 24.145 215.885 ;
        RECT 24.320 215.340 29.665 215.885 ;
        RECT 29.840 215.340 35.185 215.885 ;
        RECT 16.960 213.335 22.305 213.770 ;
        RECT 22.475 213.335 22.765 214.500 ;
        RECT 22.935 214.425 23.455 214.965 ;
        RECT 23.625 214.595 24.145 215.135 ;
        RECT 22.935 213.335 24.145 214.425 ;
        RECT 25.910 213.770 26.260 215.020 ;
        RECT 27.740 214.510 28.080 215.340 ;
        RECT 31.430 213.770 31.780 215.020 ;
        RECT 33.260 214.510 33.600 215.340 ;
        RECT 35.355 215.160 35.645 215.885 ;
        RECT 35.815 215.135 37.025 215.885 ;
        RECT 37.200 215.340 42.545 215.885 ;
        RECT 42.720 215.340 48.065 215.885 ;
        RECT 24.320 213.335 29.665 213.770 ;
        RECT 29.840 213.335 35.185 213.770 ;
        RECT 35.355 213.335 35.645 214.500 ;
        RECT 35.815 214.425 36.335 214.965 ;
        RECT 36.505 214.595 37.025 215.135 ;
        RECT 35.815 213.335 37.025 214.425 ;
        RECT 38.790 213.770 39.140 215.020 ;
        RECT 40.620 214.510 40.960 215.340 ;
        RECT 44.310 213.770 44.660 215.020 ;
        RECT 46.140 214.510 46.480 215.340 ;
        RECT 48.235 215.160 48.525 215.885 ;
        RECT 48.695 215.135 49.905 215.885 ;
        RECT 50.080 215.340 55.425 215.885 ;
        RECT 55.600 215.340 60.945 215.885 ;
        RECT 37.200 213.335 42.545 213.770 ;
        RECT 42.720 213.335 48.065 213.770 ;
        RECT 48.235 213.335 48.525 214.500 ;
        RECT 48.695 214.425 49.215 214.965 ;
        RECT 49.385 214.595 49.905 215.135 ;
        RECT 48.695 213.335 49.905 214.425 ;
        RECT 51.670 213.770 52.020 215.020 ;
        RECT 53.500 214.510 53.840 215.340 ;
        RECT 57.190 213.770 57.540 215.020 ;
        RECT 59.020 214.510 59.360 215.340 ;
        RECT 61.115 215.160 61.405 215.885 ;
        RECT 61.575 215.135 62.785 215.885 ;
        RECT 62.960 215.340 68.305 215.885 ;
        RECT 68.480 215.340 73.825 215.885 ;
        RECT 50.080 213.335 55.425 213.770 ;
        RECT 55.600 213.335 60.945 213.770 ;
        RECT 61.115 213.335 61.405 214.500 ;
        RECT 61.575 214.425 62.095 214.965 ;
        RECT 62.265 214.595 62.785 215.135 ;
        RECT 61.575 213.335 62.785 214.425 ;
        RECT 64.550 213.770 64.900 215.020 ;
        RECT 66.380 214.510 66.720 215.340 ;
        RECT 70.070 213.770 70.420 215.020 ;
        RECT 71.900 214.510 72.240 215.340 ;
        RECT 73.995 215.160 74.285 215.885 ;
        RECT 74.455 215.135 75.665 215.885 ;
        RECT 75.840 215.340 81.185 215.885 ;
        RECT 81.360 215.340 86.705 215.885 ;
        RECT 62.960 213.335 68.305 213.770 ;
        RECT 68.480 213.335 73.825 213.770 ;
        RECT 73.995 213.335 74.285 214.500 ;
        RECT 74.455 214.425 74.975 214.965 ;
        RECT 75.145 214.595 75.665 215.135 ;
        RECT 74.455 213.335 75.665 214.425 ;
        RECT 77.430 213.770 77.780 215.020 ;
        RECT 79.260 214.510 79.600 215.340 ;
        RECT 82.950 213.770 83.300 215.020 ;
        RECT 84.780 214.510 85.120 215.340 ;
        RECT 86.875 215.160 87.165 215.885 ;
        RECT 87.335 215.135 88.545 215.885 ;
        RECT 88.720 215.340 94.065 215.885 ;
        RECT 94.240 215.340 99.585 215.885 ;
        RECT 75.840 213.335 81.185 213.770 ;
        RECT 81.360 213.335 86.705 213.770 ;
        RECT 86.875 213.335 87.165 214.500 ;
        RECT 87.335 214.425 87.855 214.965 ;
        RECT 88.025 214.595 88.545 215.135 ;
        RECT 87.335 213.335 88.545 214.425 ;
        RECT 90.310 213.770 90.660 215.020 ;
        RECT 92.140 214.510 92.480 215.340 ;
        RECT 95.830 213.770 96.180 215.020 ;
        RECT 97.660 214.510 98.000 215.340 ;
        RECT 99.755 215.160 100.045 215.885 ;
        RECT 100.215 215.135 101.425 215.885 ;
        RECT 101.600 215.340 106.945 215.885 ;
        RECT 107.120 215.340 112.465 215.885 ;
        RECT 88.720 213.335 94.065 213.770 ;
        RECT 94.240 213.335 99.585 213.770 ;
        RECT 99.755 213.335 100.045 214.500 ;
        RECT 100.215 214.425 100.735 214.965 ;
        RECT 100.905 214.595 101.425 215.135 ;
        RECT 100.215 213.335 101.425 214.425 ;
        RECT 103.190 213.770 103.540 215.020 ;
        RECT 105.020 214.510 105.360 215.340 ;
        RECT 108.710 213.770 109.060 215.020 ;
        RECT 110.540 214.510 110.880 215.340 ;
        RECT 112.635 215.160 112.925 215.885 ;
        RECT 113.560 215.340 118.905 215.885 ;
        RECT 119.080 215.340 124.425 215.885 ;
        RECT 101.600 213.335 106.945 213.770 ;
        RECT 107.120 213.335 112.465 213.770 ;
        RECT 112.635 213.335 112.925 214.500 ;
        RECT 115.150 213.770 115.500 215.020 ;
        RECT 116.980 214.510 117.320 215.340 ;
        RECT 120.670 213.770 121.020 215.020 ;
        RECT 122.500 214.510 122.840 215.340 ;
        RECT 124.595 215.135 125.805 215.885 ;
        RECT 124.595 214.425 125.115 214.965 ;
        RECT 125.285 214.595 125.805 215.135 ;
        RECT 113.560 213.335 118.905 213.770 ;
        RECT 119.080 213.335 124.425 213.770 ;
        RECT 124.595 213.335 125.805 214.425 ;
        RECT 11.810 213.165 125.890 213.335 ;
        RECT 11.895 212.075 13.105 213.165 ;
        RECT 11.895 211.365 12.415 211.905 ;
        RECT 12.585 211.535 13.105 212.075 ;
        RECT 13.275 212.075 16.785 213.165 ;
        RECT 16.960 212.730 22.305 213.165 ;
        RECT 13.275 211.555 14.965 212.075 ;
        RECT 15.135 211.385 16.785 211.905 ;
        RECT 18.550 211.480 18.900 212.730 ;
        RECT 22.475 212.000 22.765 213.165 ;
        RECT 23.395 212.075 25.985 213.165 ;
        RECT 26.160 212.730 31.505 213.165 ;
        RECT 31.680 212.730 37.025 213.165 ;
        RECT 37.200 212.730 42.545 213.165 ;
        RECT 42.720 212.730 48.065 213.165 ;
        RECT 11.895 210.615 13.105 211.365 ;
        RECT 13.275 210.615 16.785 211.385 ;
        RECT 20.380 211.160 20.720 211.990 ;
        RECT 23.395 211.555 24.605 212.075 ;
        RECT 24.775 211.385 25.985 211.905 ;
        RECT 27.750 211.480 28.100 212.730 ;
        RECT 16.960 210.615 22.305 211.160 ;
        RECT 22.475 210.615 22.765 211.340 ;
        RECT 23.395 210.615 25.985 211.385 ;
        RECT 29.580 211.160 29.920 211.990 ;
        RECT 33.270 211.480 33.620 212.730 ;
        RECT 35.100 211.160 35.440 211.990 ;
        RECT 38.790 211.480 39.140 212.730 ;
        RECT 40.620 211.160 40.960 211.990 ;
        RECT 44.310 211.480 44.660 212.730 ;
        RECT 48.235 212.000 48.525 213.165 ;
        RECT 49.155 212.075 51.745 213.165 ;
        RECT 51.920 212.730 57.265 213.165 ;
        RECT 57.440 212.730 62.785 213.165 ;
        RECT 62.960 212.730 68.305 213.165 ;
        RECT 68.480 212.730 73.825 213.165 ;
        RECT 46.140 211.160 46.480 211.990 ;
        RECT 49.155 211.555 50.365 212.075 ;
        RECT 50.535 211.385 51.745 211.905 ;
        RECT 53.510 211.480 53.860 212.730 ;
        RECT 26.160 210.615 31.505 211.160 ;
        RECT 31.680 210.615 37.025 211.160 ;
        RECT 37.200 210.615 42.545 211.160 ;
        RECT 42.720 210.615 48.065 211.160 ;
        RECT 48.235 210.615 48.525 211.340 ;
        RECT 49.155 210.615 51.745 211.385 ;
        RECT 55.340 211.160 55.680 211.990 ;
        RECT 59.030 211.480 59.380 212.730 ;
        RECT 60.860 211.160 61.200 211.990 ;
        RECT 64.550 211.480 64.900 212.730 ;
        RECT 66.380 211.160 66.720 211.990 ;
        RECT 70.070 211.480 70.420 212.730 ;
        RECT 73.995 212.000 74.285 213.165 ;
        RECT 74.915 212.075 77.505 213.165 ;
        RECT 77.680 212.730 83.025 213.165 ;
        RECT 83.200 212.730 88.545 213.165 ;
        RECT 88.720 212.730 94.065 213.165 ;
        RECT 94.240 212.730 99.585 213.165 ;
        RECT 71.900 211.160 72.240 211.990 ;
        RECT 74.915 211.555 76.125 212.075 ;
        RECT 76.295 211.385 77.505 211.905 ;
        RECT 79.270 211.480 79.620 212.730 ;
        RECT 51.920 210.615 57.265 211.160 ;
        RECT 57.440 210.615 62.785 211.160 ;
        RECT 62.960 210.615 68.305 211.160 ;
        RECT 68.480 210.615 73.825 211.160 ;
        RECT 73.995 210.615 74.285 211.340 ;
        RECT 74.915 210.615 77.505 211.385 ;
        RECT 81.100 211.160 81.440 211.990 ;
        RECT 84.790 211.480 85.140 212.730 ;
        RECT 86.620 211.160 86.960 211.990 ;
        RECT 90.310 211.480 90.660 212.730 ;
        RECT 92.140 211.160 92.480 211.990 ;
        RECT 95.830 211.480 96.180 212.730 ;
        RECT 99.755 212.000 100.045 213.165 ;
        RECT 100.675 212.075 102.345 213.165 ;
        RECT 102.520 212.730 107.865 213.165 ;
        RECT 108.040 212.730 113.385 213.165 ;
        RECT 113.560 212.730 118.905 213.165 ;
        RECT 119.080 212.730 124.425 213.165 ;
        RECT 97.660 211.160 98.000 211.990 ;
        RECT 100.675 211.555 101.425 212.075 ;
        RECT 101.595 211.385 102.345 211.905 ;
        RECT 104.110 211.480 104.460 212.730 ;
        RECT 77.680 210.615 83.025 211.160 ;
        RECT 83.200 210.615 88.545 211.160 ;
        RECT 88.720 210.615 94.065 211.160 ;
        RECT 94.240 210.615 99.585 211.160 ;
        RECT 99.755 210.615 100.045 211.340 ;
        RECT 100.675 210.615 102.345 211.385 ;
        RECT 105.940 211.160 106.280 211.990 ;
        RECT 109.630 211.480 109.980 212.730 ;
        RECT 111.460 211.160 111.800 211.990 ;
        RECT 115.150 211.480 115.500 212.730 ;
        RECT 116.980 211.160 117.320 211.990 ;
        RECT 120.670 211.480 121.020 212.730 ;
        RECT 124.595 212.075 125.805 213.165 ;
        RECT 122.500 211.160 122.840 211.990 ;
        RECT 124.595 211.535 125.115 212.075 ;
        RECT 125.285 211.365 125.805 211.905 ;
        RECT 102.520 210.615 107.865 211.160 ;
        RECT 108.040 210.615 113.385 211.160 ;
        RECT 113.560 210.615 118.905 211.160 ;
        RECT 119.080 210.615 124.425 211.160 ;
        RECT 124.595 210.615 125.805 211.365 ;
        RECT 11.810 210.445 125.890 210.615 ;
        RECT 11.895 209.695 13.105 210.445 ;
        RECT 13.280 209.900 18.625 210.445 ;
        RECT 18.800 209.900 24.145 210.445 ;
        RECT 24.320 209.900 29.665 210.445 ;
        RECT 29.840 209.900 35.185 210.445 ;
        RECT 11.895 209.155 12.415 209.695 ;
        RECT 12.585 208.985 13.105 209.525 ;
        RECT 11.895 207.895 13.105 208.985 ;
        RECT 14.870 208.330 15.220 209.580 ;
        RECT 16.700 209.070 17.040 209.900 ;
        RECT 20.390 208.330 20.740 209.580 ;
        RECT 22.220 209.070 22.560 209.900 ;
        RECT 25.910 208.330 26.260 209.580 ;
        RECT 27.740 209.070 28.080 209.900 ;
        RECT 31.430 208.330 31.780 209.580 ;
        RECT 33.260 209.070 33.600 209.900 ;
        RECT 35.355 209.720 35.645 210.445 ;
        RECT 36.275 209.675 38.865 210.445 ;
        RECT 39.040 209.900 44.385 210.445 ;
        RECT 44.560 209.900 49.905 210.445 ;
        RECT 50.080 209.900 55.425 210.445 ;
        RECT 55.600 209.900 60.945 210.445 ;
        RECT 13.280 207.895 18.625 208.330 ;
        RECT 18.800 207.895 24.145 208.330 ;
        RECT 24.320 207.895 29.665 208.330 ;
        RECT 29.840 207.895 35.185 208.330 ;
        RECT 35.355 207.895 35.645 209.060 ;
        RECT 36.275 208.985 37.485 209.505 ;
        RECT 37.655 209.155 38.865 209.675 ;
        RECT 36.275 207.895 38.865 208.985 ;
        RECT 40.630 208.330 40.980 209.580 ;
        RECT 42.460 209.070 42.800 209.900 ;
        RECT 46.150 208.330 46.500 209.580 ;
        RECT 47.980 209.070 48.320 209.900 ;
        RECT 51.670 208.330 52.020 209.580 ;
        RECT 53.500 209.070 53.840 209.900 ;
        RECT 57.190 208.330 57.540 209.580 ;
        RECT 59.020 209.070 59.360 209.900 ;
        RECT 61.115 209.720 61.405 210.445 ;
        RECT 62.035 209.675 64.625 210.445 ;
        RECT 64.800 209.900 70.145 210.445 ;
        RECT 70.320 209.900 75.665 210.445 ;
        RECT 75.840 209.900 81.185 210.445 ;
        RECT 81.360 209.900 86.705 210.445 ;
        RECT 39.040 207.895 44.385 208.330 ;
        RECT 44.560 207.895 49.905 208.330 ;
        RECT 50.080 207.895 55.425 208.330 ;
        RECT 55.600 207.895 60.945 208.330 ;
        RECT 61.115 207.895 61.405 209.060 ;
        RECT 62.035 208.985 63.245 209.505 ;
        RECT 63.415 209.155 64.625 209.675 ;
        RECT 62.035 207.895 64.625 208.985 ;
        RECT 66.390 208.330 66.740 209.580 ;
        RECT 68.220 209.070 68.560 209.900 ;
        RECT 71.910 208.330 72.260 209.580 ;
        RECT 73.740 209.070 74.080 209.900 ;
        RECT 77.430 208.330 77.780 209.580 ;
        RECT 79.260 209.070 79.600 209.900 ;
        RECT 82.950 208.330 83.300 209.580 ;
        RECT 84.780 209.070 85.120 209.900 ;
        RECT 86.875 209.720 87.165 210.445 ;
        RECT 87.795 209.675 90.385 210.445 ;
        RECT 90.560 209.900 95.905 210.445 ;
        RECT 96.080 209.900 101.425 210.445 ;
        RECT 101.600 209.900 106.945 210.445 ;
        RECT 107.120 209.900 112.465 210.445 ;
        RECT 64.800 207.895 70.145 208.330 ;
        RECT 70.320 207.895 75.665 208.330 ;
        RECT 75.840 207.895 81.185 208.330 ;
        RECT 81.360 207.895 86.705 208.330 ;
        RECT 86.875 207.895 87.165 209.060 ;
        RECT 87.795 208.985 89.005 209.505 ;
        RECT 89.175 209.155 90.385 209.675 ;
        RECT 87.795 207.895 90.385 208.985 ;
        RECT 92.150 208.330 92.500 209.580 ;
        RECT 93.980 209.070 94.320 209.900 ;
        RECT 97.670 208.330 98.020 209.580 ;
        RECT 99.500 209.070 99.840 209.900 ;
        RECT 103.190 208.330 103.540 209.580 ;
        RECT 105.020 209.070 105.360 209.900 ;
        RECT 108.710 208.330 109.060 209.580 ;
        RECT 110.540 209.070 110.880 209.900 ;
        RECT 112.635 209.720 112.925 210.445 ;
        RECT 113.560 209.900 118.905 210.445 ;
        RECT 119.080 209.900 124.425 210.445 ;
        RECT 90.560 207.895 95.905 208.330 ;
        RECT 96.080 207.895 101.425 208.330 ;
        RECT 101.600 207.895 106.945 208.330 ;
        RECT 107.120 207.895 112.465 208.330 ;
        RECT 112.635 207.895 112.925 209.060 ;
        RECT 115.150 208.330 115.500 209.580 ;
        RECT 116.980 209.070 117.320 209.900 ;
        RECT 120.670 208.330 121.020 209.580 ;
        RECT 122.500 209.070 122.840 209.900 ;
        RECT 124.595 209.695 125.805 210.445 ;
        RECT 124.595 208.985 125.115 209.525 ;
        RECT 125.285 209.155 125.805 209.695 ;
        RECT 113.560 207.895 118.905 208.330 ;
        RECT 119.080 207.895 124.425 208.330 ;
        RECT 124.595 207.895 125.805 208.985 ;
        RECT 11.810 207.725 125.890 207.895 ;
        RECT 11.895 206.635 13.105 207.725 ;
        RECT 11.895 205.925 12.415 206.465 ;
        RECT 12.585 206.095 13.105 206.635 ;
        RECT 13.275 206.635 16.785 207.725 ;
        RECT 16.960 207.290 22.305 207.725 ;
        RECT 13.275 206.115 14.965 206.635 ;
        RECT 15.135 205.945 16.785 206.465 ;
        RECT 18.550 206.040 18.900 207.290 ;
        RECT 22.475 206.560 22.765 207.725 ;
        RECT 23.395 206.635 25.985 207.725 ;
        RECT 26.160 207.290 31.505 207.725 ;
        RECT 31.680 207.290 37.025 207.725 ;
        RECT 37.200 207.290 42.545 207.725 ;
        RECT 42.720 207.290 48.065 207.725 ;
        RECT 11.895 205.175 13.105 205.925 ;
        RECT 13.275 205.175 16.785 205.945 ;
        RECT 20.380 205.720 20.720 206.550 ;
        RECT 23.395 206.115 24.605 206.635 ;
        RECT 24.775 205.945 25.985 206.465 ;
        RECT 27.750 206.040 28.100 207.290 ;
        RECT 16.960 205.175 22.305 205.720 ;
        RECT 22.475 205.175 22.765 205.900 ;
        RECT 23.395 205.175 25.985 205.945 ;
        RECT 29.580 205.720 29.920 206.550 ;
        RECT 33.270 206.040 33.620 207.290 ;
        RECT 35.100 205.720 35.440 206.550 ;
        RECT 38.790 206.040 39.140 207.290 ;
        RECT 40.620 205.720 40.960 206.550 ;
        RECT 44.310 206.040 44.660 207.290 ;
        RECT 48.235 206.560 48.525 207.725 ;
        RECT 49.155 206.635 51.745 207.725 ;
        RECT 51.920 207.290 57.265 207.725 ;
        RECT 57.440 207.290 62.785 207.725 ;
        RECT 62.960 207.290 68.305 207.725 ;
        RECT 68.480 207.290 73.825 207.725 ;
        RECT 46.140 205.720 46.480 206.550 ;
        RECT 49.155 206.115 50.365 206.635 ;
        RECT 50.535 205.945 51.745 206.465 ;
        RECT 53.510 206.040 53.860 207.290 ;
        RECT 26.160 205.175 31.505 205.720 ;
        RECT 31.680 205.175 37.025 205.720 ;
        RECT 37.200 205.175 42.545 205.720 ;
        RECT 42.720 205.175 48.065 205.720 ;
        RECT 48.235 205.175 48.525 205.900 ;
        RECT 49.155 205.175 51.745 205.945 ;
        RECT 55.340 205.720 55.680 206.550 ;
        RECT 59.030 206.040 59.380 207.290 ;
        RECT 60.860 205.720 61.200 206.550 ;
        RECT 64.550 206.040 64.900 207.290 ;
        RECT 66.380 205.720 66.720 206.550 ;
        RECT 70.070 206.040 70.420 207.290 ;
        RECT 73.995 206.560 74.285 207.725 ;
        RECT 74.915 206.635 77.505 207.725 ;
        RECT 77.680 207.290 83.025 207.725 ;
        RECT 83.200 207.290 88.545 207.725 ;
        RECT 88.720 207.290 94.065 207.725 ;
        RECT 94.240 207.290 99.585 207.725 ;
        RECT 71.900 205.720 72.240 206.550 ;
        RECT 74.915 206.115 76.125 206.635 ;
        RECT 76.295 205.945 77.505 206.465 ;
        RECT 79.270 206.040 79.620 207.290 ;
        RECT 51.920 205.175 57.265 205.720 ;
        RECT 57.440 205.175 62.785 205.720 ;
        RECT 62.960 205.175 68.305 205.720 ;
        RECT 68.480 205.175 73.825 205.720 ;
        RECT 73.995 205.175 74.285 205.900 ;
        RECT 74.915 205.175 77.505 205.945 ;
        RECT 81.100 205.720 81.440 206.550 ;
        RECT 84.790 206.040 85.140 207.290 ;
        RECT 86.620 205.720 86.960 206.550 ;
        RECT 90.310 206.040 90.660 207.290 ;
        RECT 92.140 205.720 92.480 206.550 ;
        RECT 95.830 206.040 96.180 207.290 ;
        RECT 99.755 206.560 100.045 207.725 ;
        RECT 100.675 206.635 102.345 207.725 ;
        RECT 102.520 207.290 107.865 207.725 ;
        RECT 108.040 207.290 113.385 207.725 ;
        RECT 113.560 207.290 118.905 207.725 ;
        RECT 119.080 207.290 124.425 207.725 ;
        RECT 97.660 205.720 98.000 206.550 ;
        RECT 100.675 206.115 101.425 206.635 ;
        RECT 101.595 205.945 102.345 206.465 ;
        RECT 104.110 206.040 104.460 207.290 ;
        RECT 77.680 205.175 83.025 205.720 ;
        RECT 83.200 205.175 88.545 205.720 ;
        RECT 88.720 205.175 94.065 205.720 ;
        RECT 94.240 205.175 99.585 205.720 ;
        RECT 99.755 205.175 100.045 205.900 ;
        RECT 100.675 205.175 102.345 205.945 ;
        RECT 105.940 205.720 106.280 206.550 ;
        RECT 109.630 206.040 109.980 207.290 ;
        RECT 111.460 205.720 111.800 206.550 ;
        RECT 115.150 206.040 115.500 207.290 ;
        RECT 116.980 205.720 117.320 206.550 ;
        RECT 120.670 206.040 121.020 207.290 ;
        RECT 124.595 206.635 125.805 207.725 ;
        RECT 122.500 205.720 122.840 206.550 ;
        RECT 124.595 206.095 125.115 206.635 ;
        RECT 125.285 205.925 125.805 206.465 ;
        RECT 102.520 205.175 107.865 205.720 ;
        RECT 108.040 205.175 113.385 205.720 ;
        RECT 113.560 205.175 118.905 205.720 ;
        RECT 119.080 205.175 124.425 205.720 ;
        RECT 124.595 205.175 125.805 205.925 ;
        RECT 11.810 205.005 125.890 205.175 ;
        RECT 11.895 204.255 13.105 205.005 ;
        RECT 13.280 204.460 18.625 205.005 ;
        RECT 18.800 204.460 24.145 205.005 ;
        RECT 24.320 204.460 29.665 205.005 ;
        RECT 29.840 204.460 35.185 205.005 ;
        RECT 11.895 203.715 12.415 204.255 ;
        RECT 12.585 203.545 13.105 204.085 ;
        RECT 11.895 202.455 13.105 203.545 ;
        RECT 14.870 202.890 15.220 204.140 ;
        RECT 16.700 203.630 17.040 204.460 ;
        RECT 20.390 202.890 20.740 204.140 ;
        RECT 22.220 203.630 22.560 204.460 ;
        RECT 25.910 202.890 26.260 204.140 ;
        RECT 27.740 203.630 28.080 204.460 ;
        RECT 31.430 202.890 31.780 204.140 ;
        RECT 33.260 203.630 33.600 204.460 ;
        RECT 35.355 204.280 35.645 205.005 ;
        RECT 36.275 204.235 38.865 205.005 ;
        RECT 39.040 204.460 44.385 205.005 ;
        RECT 44.560 204.460 49.905 205.005 ;
        RECT 50.080 204.460 55.425 205.005 ;
        RECT 55.600 204.460 60.945 205.005 ;
        RECT 13.280 202.455 18.625 202.890 ;
        RECT 18.800 202.455 24.145 202.890 ;
        RECT 24.320 202.455 29.665 202.890 ;
        RECT 29.840 202.455 35.185 202.890 ;
        RECT 35.355 202.455 35.645 203.620 ;
        RECT 36.275 203.545 37.485 204.065 ;
        RECT 37.655 203.715 38.865 204.235 ;
        RECT 36.275 202.455 38.865 203.545 ;
        RECT 40.630 202.890 40.980 204.140 ;
        RECT 42.460 203.630 42.800 204.460 ;
        RECT 46.150 202.890 46.500 204.140 ;
        RECT 47.980 203.630 48.320 204.460 ;
        RECT 51.670 202.890 52.020 204.140 ;
        RECT 53.500 203.630 53.840 204.460 ;
        RECT 57.190 202.890 57.540 204.140 ;
        RECT 59.020 203.630 59.360 204.460 ;
        RECT 61.115 204.280 61.405 205.005 ;
        RECT 62.035 204.235 64.625 205.005 ;
        RECT 64.800 204.460 70.145 205.005 ;
        RECT 70.320 204.460 75.665 205.005 ;
        RECT 75.840 204.460 81.185 205.005 ;
        RECT 81.360 204.460 86.705 205.005 ;
        RECT 39.040 202.455 44.385 202.890 ;
        RECT 44.560 202.455 49.905 202.890 ;
        RECT 50.080 202.455 55.425 202.890 ;
        RECT 55.600 202.455 60.945 202.890 ;
        RECT 61.115 202.455 61.405 203.620 ;
        RECT 62.035 203.545 63.245 204.065 ;
        RECT 63.415 203.715 64.625 204.235 ;
        RECT 62.035 202.455 64.625 203.545 ;
        RECT 66.390 202.890 66.740 204.140 ;
        RECT 68.220 203.630 68.560 204.460 ;
        RECT 71.910 202.890 72.260 204.140 ;
        RECT 73.740 203.630 74.080 204.460 ;
        RECT 77.430 202.890 77.780 204.140 ;
        RECT 79.260 203.630 79.600 204.460 ;
        RECT 82.950 202.890 83.300 204.140 ;
        RECT 84.780 203.630 85.120 204.460 ;
        RECT 86.875 204.280 87.165 205.005 ;
        RECT 87.795 204.235 90.385 205.005 ;
        RECT 90.560 204.460 95.905 205.005 ;
        RECT 96.080 204.460 101.425 205.005 ;
        RECT 101.600 204.460 106.945 205.005 ;
        RECT 107.120 204.460 112.465 205.005 ;
        RECT 64.800 202.455 70.145 202.890 ;
        RECT 70.320 202.455 75.665 202.890 ;
        RECT 75.840 202.455 81.185 202.890 ;
        RECT 81.360 202.455 86.705 202.890 ;
        RECT 86.875 202.455 87.165 203.620 ;
        RECT 87.795 203.545 89.005 204.065 ;
        RECT 89.175 203.715 90.385 204.235 ;
        RECT 87.795 202.455 90.385 203.545 ;
        RECT 92.150 202.890 92.500 204.140 ;
        RECT 93.980 203.630 94.320 204.460 ;
        RECT 97.670 202.890 98.020 204.140 ;
        RECT 99.500 203.630 99.840 204.460 ;
        RECT 103.190 202.890 103.540 204.140 ;
        RECT 105.020 203.630 105.360 204.460 ;
        RECT 108.710 202.890 109.060 204.140 ;
        RECT 110.540 203.630 110.880 204.460 ;
        RECT 112.635 204.280 112.925 205.005 ;
        RECT 113.560 204.460 118.905 205.005 ;
        RECT 119.080 204.460 124.425 205.005 ;
        RECT 90.560 202.455 95.905 202.890 ;
        RECT 96.080 202.455 101.425 202.890 ;
        RECT 101.600 202.455 106.945 202.890 ;
        RECT 107.120 202.455 112.465 202.890 ;
        RECT 112.635 202.455 112.925 203.620 ;
        RECT 115.150 202.890 115.500 204.140 ;
        RECT 116.980 203.630 117.320 204.460 ;
        RECT 120.670 202.890 121.020 204.140 ;
        RECT 122.500 203.630 122.840 204.460 ;
        RECT 124.595 204.255 125.805 205.005 ;
        RECT 124.595 203.545 125.115 204.085 ;
        RECT 125.285 203.715 125.805 204.255 ;
        RECT 113.560 202.455 118.905 202.890 ;
        RECT 119.080 202.455 124.425 202.890 ;
        RECT 124.595 202.455 125.805 203.545 ;
        RECT 11.810 202.285 125.890 202.455 ;
        RECT 11.895 201.195 13.105 202.285 ;
        RECT 11.895 200.485 12.415 201.025 ;
        RECT 12.585 200.655 13.105 201.195 ;
        RECT 13.275 201.195 16.785 202.285 ;
        RECT 16.960 201.850 22.305 202.285 ;
        RECT 13.275 200.675 14.965 201.195 ;
        RECT 15.135 200.505 16.785 201.025 ;
        RECT 18.550 200.600 18.900 201.850 ;
        RECT 22.475 201.120 22.765 202.285 ;
        RECT 23.395 201.195 25.985 202.285 ;
        RECT 26.160 201.850 31.505 202.285 ;
        RECT 31.680 201.850 37.025 202.285 ;
        RECT 37.200 201.850 42.545 202.285 ;
        RECT 42.720 201.850 48.065 202.285 ;
        RECT 11.895 199.735 13.105 200.485 ;
        RECT 13.275 199.735 16.785 200.505 ;
        RECT 20.380 200.280 20.720 201.110 ;
        RECT 23.395 200.675 24.605 201.195 ;
        RECT 24.775 200.505 25.985 201.025 ;
        RECT 27.750 200.600 28.100 201.850 ;
        RECT 16.960 199.735 22.305 200.280 ;
        RECT 22.475 199.735 22.765 200.460 ;
        RECT 23.395 199.735 25.985 200.505 ;
        RECT 29.580 200.280 29.920 201.110 ;
        RECT 33.270 200.600 33.620 201.850 ;
        RECT 35.100 200.280 35.440 201.110 ;
        RECT 38.790 200.600 39.140 201.850 ;
        RECT 40.620 200.280 40.960 201.110 ;
        RECT 44.310 200.600 44.660 201.850 ;
        RECT 48.235 201.120 48.525 202.285 ;
        RECT 49.155 201.195 51.745 202.285 ;
        RECT 51.920 201.850 57.265 202.285 ;
        RECT 57.440 201.850 62.785 202.285 ;
        RECT 62.960 201.850 68.305 202.285 ;
        RECT 68.480 201.850 73.825 202.285 ;
        RECT 46.140 200.280 46.480 201.110 ;
        RECT 49.155 200.675 50.365 201.195 ;
        RECT 50.535 200.505 51.745 201.025 ;
        RECT 53.510 200.600 53.860 201.850 ;
        RECT 26.160 199.735 31.505 200.280 ;
        RECT 31.680 199.735 37.025 200.280 ;
        RECT 37.200 199.735 42.545 200.280 ;
        RECT 42.720 199.735 48.065 200.280 ;
        RECT 48.235 199.735 48.525 200.460 ;
        RECT 49.155 199.735 51.745 200.505 ;
        RECT 55.340 200.280 55.680 201.110 ;
        RECT 59.030 200.600 59.380 201.850 ;
        RECT 60.860 200.280 61.200 201.110 ;
        RECT 64.550 200.600 64.900 201.850 ;
        RECT 66.380 200.280 66.720 201.110 ;
        RECT 70.070 200.600 70.420 201.850 ;
        RECT 73.995 201.120 74.285 202.285 ;
        RECT 74.915 201.195 77.505 202.285 ;
        RECT 77.680 201.850 83.025 202.285 ;
        RECT 83.200 201.850 88.545 202.285 ;
        RECT 88.720 201.850 94.065 202.285 ;
        RECT 94.240 201.850 99.585 202.285 ;
        RECT 71.900 200.280 72.240 201.110 ;
        RECT 74.915 200.675 76.125 201.195 ;
        RECT 76.295 200.505 77.505 201.025 ;
        RECT 79.270 200.600 79.620 201.850 ;
        RECT 51.920 199.735 57.265 200.280 ;
        RECT 57.440 199.735 62.785 200.280 ;
        RECT 62.960 199.735 68.305 200.280 ;
        RECT 68.480 199.735 73.825 200.280 ;
        RECT 73.995 199.735 74.285 200.460 ;
        RECT 74.915 199.735 77.505 200.505 ;
        RECT 81.100 200.280 81.440 201.110 ;
        RECT 84.790 200.600 85.140 201.850 ;
        RECT 86.620 200.280 86.960 201.110 ;
        RECT 90.310 200.600 90.660 201.850 ;
        RECT 92.140 200.280 92.480 201.110 ;
        RECT 95.830 200.600 96.180 201.850 ;
        RECT 99.755 201.120 100.045 202.285 ;
        RECT 100.675 201.195 102.345 202.285 ;
        RECT 102.520 201.850 107.865 202.285 ;
        RECT 108.040 201.850 113.385 202.285 ;
        RECT 113.560 201.850 118.905 202.285 ;
        RECT 119.080 201.850 124.425 202.285 ;
        RECT 97.660 200.280 98.000 201.110 ;
        RECT 100.675 200.675 101.425 201.195 ;
        RECT 101.595 200.505 102.345 201.025 ;
        RECT 104.110 200.600 104.460 201.850 ;
        RECT 77.680 199.735 83.025 200.280 ;
        RECT 83.200 199.735 88.545 200.280 ;
        RECT 88.720 199.735 94.065 200.280 ;
        RECT 94.240 199.735 99.585 200.280 ;
        RECT 99.755 199.735 100.045 200.460 ;
        RECT 100.675 199.735 102.345 200.505 ;
        RECT 105.940 200.280 106.280 201.110 ;
        RECT 109.630 200.600 109.980 201.850 ;
        RECT 111.460 200.280 111.800 201.110 ;
        RECT 115.150 200.600 115.500 201.850 ;
        RECT 116.980 200.280 117.320 201.110 ;
        RECT 120.670 200.600 121.020 201.850 ;
        RECT 124.595 201.195 125.805 202.285 ;
        RECT 122.500 200.280 122.840 201.110 ;
        RECT 124.595 200.655 125.115 201.195 ;
        RECT 125.285 200.485 125.805 201.025 ;
        RECT 102.520 199.735 107.865 200.280 ;
        RECT 108.040 199.735 113.385 200.280 ;
        RECT 113.560 199.735 118.905 200.280 ;
        RECT 119.080 199.735 124.425 200.280 ;
        RECT 124.595 199.735 125.805 200.485 ;
        RECT 11.810 199.565 125.890 199.735 ;
        RECT 11.895 198.815 13.105 199.565 ;
        RECT 13.280 199.020 18.625 199.565 ;
        RECT 18.800 199.020 24.145 199.565 ;
        RECT 24.320 199.020 29.665 199.565 ;
        RECT 29.840 199.020 35.185 199.565 ;
        RECT 11.895 198.275 12.415 198.815 ;
        RECT 12.585 198.105 13.105 198.645 ;
        RECT 11.895 197.015 13.105 198.105 ;
        RECT 14.870 197.450 15.220 198.700 ;
        RECT 16.700 198.190 17.040 199.020 ;
        RECT 20.390 197.450 20.740 198.700 ;
        RECT 22.220 198.190 22.560 199.020 ;
        RECT 25.910 197.450 26.260 198.700 ;
        RECT 27.740 198.190 28.080 199.020 ;
        RECT 31.430 197.450 31.780 198.700 ;
        RECT 33.260 198.190 33.600 199.020 ;
        RECT 35.355 198.840 35.645 199.565 ;
        RECT 36.275 198.795 38.865 199.565 ;
        RECT 39.040 199.020 44.385 199.565 ;
        RECT 44.560 199.020 49.905 199.565 ;
        RECT 50.080 199.020 55.425 199.565 ;
        RECT 55.600 199.020 60.945 199.565 ;
        RECT 13.280 197.015 18.625 197.450 ;
        RECT 18.800 197.015 24.145 197.450 ;
        RECT 24.320 197.015 29.665 197.450 ;
        RECT 29.840 197.015 35.185 197.450 ;
        RECT 35.355 197.015 35.645 198.180 ;
        RECT 36.275 198.105 37.485 198.625 ;
        RECT 37.655 198.275 38.865 198.795 ;
        RECT 36.275 197.015 38.865 198.105 ;
        RECT 40.630 197.450 40.980 198.700 ;
        RECT 42.460 198.190 42.800 199.020 ;
        RECT 46.150 197.450 46.500 198.700 ;
        RECT 47.980 198.190 48.320 199.020 ;
        RECT 51.670 197.450 52.020 198.700 ;
        RECT 53.500 198.190 53.840 199.020 ;
        RECT 57.190 197.450 57.540 198.700 ;
        RECT 59.020 198.190 59.360 199.020 ;
        RECT 61.115 198.840 61.405 199.565 ;
        RECT 61.575 198.815 62.785 199.565 ;
        RECT 39.040 197.015 44.385 197.450 ;
        RECT 44.560 197.015 49.905 197.450 ;
        RECT 50.080 197.015 55.425 197.450 ;
        RECT 55.600 197.015 60.945 197.450 ;
        RECT 61.115 197.015 61.405 198.180 ;
        RECT 61.575 198.105 62.095 198.645 ;
        RECT 62.265 198.275 62.785 198.815 ;
        RECT 62.960 198.855 63.215 199.385 ;
        RECT 63.385 199.105 63.690 199.565 ;
        RECT 63.935 199.185 65.005 199.355 ;
        RECT 62.960 198.205 63.170 198.855 ;
        RECT 63.935 198.830 64.255 199.185 ;
        RECT 63.930 198.655 64.255 198.830 ;
        RECT 63.340 198.355 64.255 198.655 ;
        RECT 64.425 198.615 64.665 199.015 ;
        RECT 64.835 198.955 65.005 199.185 ;
        RECT 65.175 199.125 65.365 199.565 ;
        RECT 65.535 199.115 66.485 199.395 ;
        RECT 66.705 199.205 67.055 199.375 ;
        RECT 64.835 198.785 65.365 198.955 ;
        RECT 63.340 198.325 64.080 198.355 ;
        RECT 61.575 197.015 62.785 198.105 ;
        RECT 62.960 197.325 63.215 198.205 ;
        RECT 63.385 197.015 63.690 198.155 ;
        RECT 63.910 197.735 64.080 198.325 ;
        RECT 64.425 198.245 64.965 198.615 ;
        RECT 65.145 198.505 65.365 198.785 ;
        RECT 65.535 198.335 65.705 199.115 ;
        RECT 65.300 198.165 65.705 198.335 ;
        RECT 65.875 198.325 66.225 198.945 ;
        RECT 65.300 198.075 65.470 198.165 ;
        RECT 66.395 198.155 66.605 198.945 ;
        RECT 64.250 197.905 65.470 198.075 ;
        RECT 65.930 197.995 66.605 198.155 ;
        RECT 63.910 197.565 64.710 197.735 ;
        RECT 64.030 197.015 64.360 197.395 ;
        RECT 64.540 197.275 64.710 197.565 ;
        RECT 65.300 197.525 65.470 197.905 ;
        RECT 65.640 197.985 66.605 197.995 ;
        RECT 66.795 198.815 67.055 199.205 ;
        RECT 67.265 199.105 67.595 199.565 ;
        RECT 68.470 199.175 69.325 199.345 ;
        RECT 69.530 199.175 70.025 199.345 ;
        RECT 70.195 199.205 70.525 199.565 ;
        RECT 66.795 198.125 66.965 198.815 ;
        RECT 67.135 198.465 67.305 198.645 ;
        RECT 67.475 198.635 68.265 198.885 ;
        RECT 68.470 198.465 68.640 199.175 ;
        RECT 68.810 198.665 69.165 198.885 ;
        RECT 67.135 198.295 68.825 198.465 ;
        RECT 65.640 197.695 66.100 197.985 ;
        RECT 66.795 197.955 68.295 198.125 ;
        RECT 66.795 197.815 66.965 197.955 ;
        RECT 66.405 197.645 66.965 197.815 ;
        RECT 64.880 197.015 65.130 197.475 ;
        RECT 65.300 197.185 66.170 197.525 ;
        RECT 66.405 197.185 66.575 197.645 ;
        RECT 67.410 197.615 68.485 197.785 ;
        RECT 66.745 197.015 67.115 197.475 ;
        RECT 67.410 197.275 67.580 197.615 ;
        RECT 67.750 197.015 68.080 197.445 ;
        RECT 68.315 197.275 68.485 197.615 ;
        RECT 68.655 197.515 68.825 198.295 ;
        RECT 68.995 198.075 69.165 198.665 ;
        RECT 69.335 198.265 69.685 198.885 ;
        RECT 68.995 197.685 69.460 198.075 ;
        RECT 69.855 197.815 70.025 199.175 ;
        RECT 70.195 197.985 70.655 199.035 ;
        RECT 69.630 197.645 70.025 197.815 ;
        RECT 69.630 197.515 69.800 197.645 ;
        RECT 68.655 197.185 69.335 197.515 ;
        RECT 69.550 197.185 69.800 197.515 ;
        RECT 69.970 197.015 70.220 197.475 ;
        RECT 70.390 197.200 70.715 197.985 ;
        RECT 70.885 197.185 71.055 199.305 ;
        RECT 71.225 199.185 71.555 199.565 ;
        RECT 71.725 199.015 71.980 199.305 ;
        RECT 71.230 198.845 71.980 199.015 ;
        RECT 71.230 197.855 71.460 198.845 ;
        RECT 72.155 198.795 75.665 199.565 ;
        RECT 75.840 199.020 81.185 199.565 ;
        RECT 81.360 199.020 86.705 199.565 ;
        RECT 71.630 198.025 71.980 198.675 ;
        RECT 72.155 198.105 73.845 198.625 ;
        RECT 74.015 198.275 75.665 198.795 ;
        RECT 71.230 197.685 71.980 197.855 ;
        RECT 71.225 197.015 71.555 197.515 ;
        RECT 71.725 197.185 71.980 197.685 ;
        RECT 72.155 197.015 75.665 198.105 ;
        RECT 77.430 197.450 77.780 198.700 ;
        RECT 79.260 198.190 79.600 199.020 ;
        RECT 82.950 197.450 83.300 198.700 ;
        RECT 84.780 198.190 85.120 199.020 ;
        RECT 86.875 198.840 87.165 199.565 ;
        RECT 87.795 198.795 90.385 199.565 ;
        RECT 90.560 199.020 95.905 199.565 ;
        RECT 96.080 199.020 101.425 199.565 ;
        RECT 101.600 199.020 106.945 199.565 ;
        RECT 107.120 199.020 112.465 199.565 ;
        RECT 75.840 197.015 81.185 197.450 ;
        RECT 81.360 197.015 86.705 197.450 ;
        RECT 86.875 197.015 87.165 198.180 ;
        RECT 87.795 198.105 89.005 198.625 ;
        RECT 89.175 198.275 90.385 198.795 ;
        RECT 87.795 197.015 90.385 198.105 ;
        RECT 92.150 197.450 92.500 198.700 ;
        RECT 93.980 198.190 94.320 199.020 ;
        RECT 97.670 197.450 98.020 198.700 ;
        RECT 99.500 198.190 99.840 199.020 ;
        RECT 103.190 197.450 103.540 198.700 ;
        RECT 105.020 198.190 105.360 199.020 ;
        RECT 108.710 197.450 109.060 198.700 ;
        RECT 110.540 198.190 110.880 199.020 ;
        RECT 112.635 198.840 112.925 199.565 ;
        RECT 113.560 199.020 118.905 199.565 ;
        RECT 119.080 199.020 124.425 199.565 ;
        RECT 90.560 197.015 95.905 197.450 ;
        RECT 96.080 197.015 101.425 197.450 ;
        RECT 101.600 197.015 106.945 197.450 ;
        RECT 107.120 197.015 112.465 197.450 ;
        RECT 112.635 197.015 112.925 198.180 ;
        RECT 115.150 197.450 115.500 198.700 ;
        RECT 116.980 198.190 117.320 199.020 ;
        RECT 120.670 197.450 121.020 198.700 ;
        RECT 122.500 198.190 122.840 199.020 ;
        RECT 124.595 198.815 125.805 199.565 ;
        RECT 124.595 198.105 125.115 198.645 ;
        RECT 125.285 198.275 125.805 198.815 ;
        RECT 113.560 197.015 118.905 197.450 ;
        RECT 119.080 197.015 124.425 197.450 ;
        RECT 124.595 197.015 125.805 198.105 ;
        RECT 11.810 196.845 125.890 197.015 ;
        RECT 11.895 195.755 13.105 196.845 ;
        RECT 11.895 195.045 12.415 195.585 ;
        RECT 12.585 195.215 13.105 195.755 ;
        RECT 13.275 195.755 16.785 196.845 ;
        RECT 16.960 196.410 22.305 196.845 ;
        RECT 13.275 195.235 14.965 195.755 ;
        RECT 15.135 195.065 16.785 195.585 ;
        RECT 18.550 195.160 18.900 196.410 ;
        RECT 22.475 195.680 22.765 196.845 ;
        RECT 23.395 195.755 25.985 196.845 ;
        RECT 26.160 196.410 31.505 196.845 ;
        RECT 31.680 196.410 37.025 196.845 ;
        RECT 37.200 196.410 42.545 196.845 ;
        RECT 42.720 196.410 48.065 196.845 ;
        RECT 11.895 194.295 13.105 195.045 ;
        RECT 13.275 194.295 16.785 195.065 ;
        RECT 20.380 194.840 20.720 195.670 ;
        RECT 23.395 195.235 24.605 195.755 ;
        RECT 24.775 195.065 25.985 195.585 ;
        RECT 27.750 195.160 28.100 196.410 ;
        RECT 16.960 194.295 22.305 194.840 ;
        RECT 22.475 194.295 22.765 195.020 ;
        RECT 23.395 194.295 25.985 195.065 ;
        RECT 29.580 194.840 29.920 195.670 ;
        RECT 33.270 195.160 33.620 196.410 ;
        RECT 35.100 194.840 35.440 195.670 ;
        RECT 38.790 195.160 39.140 196.410 ;
        RECT 40.620 194.840 40.960 195.670 ;
        RECT 44.310 195.160 44.660 196.410 ;
        RECT 48.235 195.680 48.525 196.845 ;
        RECT 49.155 195.755 52.665 196.845 ;
        RECT 52.840 196.410 58.185 196.845 ;
        RECT 46.140 194.840 46.480 195.670 ;
        RECT 49.155 195.235 50.845 195.755 ;
        RECT 51.015 195.065 52.665 195.585 ;
        RECT 54.430 195.160 54.780 196.410 ;
        RECT 58.360 196.175 58.615 196.675 ;
        RECT 58.785 196.345 59.115 196.845 ;
        RECT 58.360 196.005 59.110 196.175 ;
        RECT 26.160 194.295 31.505 194.840 ;
        RECT 31.680 194.295 37.025 194.840 ;
        RECT 37.200 194.295 42.545 194.840 ;
        RECT 42.720 194.295 48.065 194.840 ;
        RECT 48.235 194.295 48.525 195.020 ;
        RECT 49.155 194.295 52.665 195.065 ;
        RECT 56.260 194.840 56.600 195.670 ;
        RECT 58.360 195.185 58.710 195.835 ;
        RECT 58.880 195.015 59.110 196.005 ;
        RECT 58.360 194.845 59.110 195.015 ;
        RECT 52.840 194.295 58.185 194.840 ;
        RECT 58.360 194.555 58.615 194.845 ;
        RECT 58.785 194.295 59.115 194.675 ;
        RECT 59.285 194.555 59.455 196.675 ;
        RECT 59.625 195.875 59.950 196.660 ;
        RECT 60.120 196.385 60.370 196.845 ;
        RECT 60.540 196.345 60.790 196.675 ;
        RECT 61.005 196.345 61.685 196.675 ;
        RECT 60.540 196.215 60.710 196.345 ;
        RECT 60.315 196.045 60.710 196.215 ;
        RECT 59.685 194.825 60.145 195.875 ;
        RECT 60.315 194.685 60.485 196.045 ;
        RECT 60.880 195.785 61.345 196.175 ;
        RECT 60.655 194.975 61.005 195.595 ;
        RECT 61.175 195.195 61.345 195.785 ;
        RECT 61.515 195.565 61.685 196.345 ;
        RECT 61.855 196.245 62.025 196.585 ;
        RECT 62.260 196.415 62.590 196.845 ;
        RECT 62.760 196.245 62.930 196.585 ;
        RECT 63.225 196.385 63.595 196.845 ;
        RECT 61.855 196.075 62.930 196.245 ;
        RECT 63.765 196.215 63.935 196.675 ;
        RECT 64.170 196.335 65.040 196.675 ;
        RECT 65.210 196.385 65.460 196.845 ;
        RECT 63.375 196.045 63.935 196.215 ;
        RECT 63.375 195.905 63.545 196.045 ;
        RECT 62.045 195.735 63.545 195.905 ;
        RECT 64.240 195.875 64.700 196.165 ;
        RECT 61.515 195.395 63.205 195.565 ;
        RECT 61.175 194.975 61.530 195.195 ;
        RECT 61.700 194.685 61.870 195.395 ;
        RECT 62.075 194.975 62.865 195.225 ;
        RECT 63.035 195.215 63.205 195.395 ;
        RECT 63.375 195.045 63.545 195.735 ;
        RECT 59.815 194.295 60.145 194.655 ;
        RECT 60.315 194.515 60.810 194.685 ;
        RECT 61.015 194.515 61.870 194.685 ;
        RECT 62.745 194.295 63.075 194.755 ;
        RECT 63.285 194.655 63.545 195.045 ;
        RECT 63.735 195.865 64.700 195.875 ;
        RECT 64.870 195.955 65.040 196.335 ;
        RECT 65.630 196.295 65.800 196.585 ;
        RECT 65.980 196.465 66.310 196.845 ;
        RECT 65.630 196.125 66.430 196.295 ;
        RECT 63.735 195.705 64.410 195.865 ;
        RECT 64.870 195.785 66.090 195.955 ;
        RECT 63.735 194.915 63.945 195.705 ;
        RECT 64.870 195.695 65.040 195.785 ;
        RECT 64.115 194.915 64.465 195.535 ;
        RECT 64.635 195.525 65.040 195.695 ;
        RECT 64.635 194.745 64.805 195.525 ;
        RECT 64.975 195.075 65.195 195.355 ;
        RECT 65.375 195.245 65.915 195.615 ;
        RECT 66.260 195.505 66.430 196.125 ;
        RECT 66.605 195.785 66.775 196.845 ;
        RECT 66.985 195.835 67.275 196.675 ;
        RECT 67.445 196.005 67.615 196.845 ;
        RECT 67.825 195.835 68.075 196.675 ;
        RECT 68.285 196.005 68.455 196.845 ;
        RECT 66.985 195.665 68.710 195.835 ;
        RECT 68.995 195.705 69.205 196.845 ;
        RECT 64.975 194.905 65.505 195.075 ;
        RECT 63.285 194.485 63.635 194.655 ;
        RECT 63.855 194.465 64.805 194.745 ;
        RECT 64.975 194.295 65.165 194.735 ;
        RECT 65.335 194.675 65.505 194.905 ;
        RECT 65.675 194.845 65.915 195.245 ;
        RECT 66.085 195.495 66.430 195.505 ;
        RECT 66.085 195.285 68.115 195.495 ;
        RECT 66.085 195.030 66.410 195.285 ;
        RECT 68.300 195.115 68.710 195.665 ;
        RECT 69.375 195.695 69.705 196.675 ;
        RECT 69.875 195.705 70.105 196.845 ;
        RECT 70.315 195.755 73.825 196.845 ;
        RECT 66.085 194.675 66.405 195.030 ;
        RECT 65.335 194.505 66.405 194.675 ;
        RECT 66.605 194.295 66.775 195.105 ;
        RECT 66.945 194.945 68.710 195.115 ;
        RECT 66.945 194.465 67.275 194.945 ;
        RECT 67.445 194.295 67.615 194.765 ;
        RECT 67.785 194.465 68.115 194.945 ;
        RECT 68.285 194.295 68.455 194.765 ;
        RECT 68.995 194.295 69.205 195.115 ;
        RECT 69.375 195.095 69.625 195.695 ;
        RECT 69.795 195.285 70.125 195.535 ;
        RECT 70.315 195.235 72.005 195.755 ;
        RECT 73.995 195.680 74.285 196.845 ;
        RECT 74.495 195.705 74.725 196.845 ;
        RECT 74.895 195.695 75.225 196.675 ;
        RECT 75.395 195.705 75.605 196.845 ;
        RECT 69.375 194.465 69.705 195.095 ;
        RECT 69.875 194.295 70.105 195.115 ;
        RECT 72.175 195.065 73.825 195.585 ;
        RECT 74.475 195.285 74.805 195.535 ;
        RECT 70.315 194.295 73.825 195.065 ;
        RECT 73.995 194.295 74.285 195.020 ;
        RECT 74.495 194.295 74.725 195.115 ;
        RECT 74.975 195.095 75.225 195.695 ;
        RECT 75.840 195.655 76.095 196.535 ;
        RECT 76.265 195.705 76.570 196.845 ;
        RECT 76.910 196.465 77.240 196.845 ;
        RECT 77.420 196.295 77.590 196.585 ;
        RECT 77.760 196.385 78.010 196.845 ;
        RECT 76.790 196.125 77.590 196.295 ;
        RECT 78.180 196.335 79.050 196.675 ;
        RECT 74.895 194.465 75.225 195.095 ;
        RECT 75.395 194.295 75.605 195.115 ;
        RECT 75.840 195.005 76.050 195.655 ;
        RECT 76.790 195.535 76.960 196.125 ;
        RECT 78.180 195.955 78.350 196.335 ;
        RECT 79.285 196.215 79.455 196.675 ;
        RECT 79.625 196.385 79.995 196.845 ;
        RECT 80.290 196.245 80.460 196.585 ;
        RECT 80.630 196.415 80.960 196.845 ;
        RECT 81.195 196.245 81.365 196.585 ;
        RECT 77.130 195.785 78.350 195.955 ;
        RECT 78.520 195.875 78.980 196.165 ;
        RECT 79.285 196.045 79.845 196.215 ;
        RECT 80.290 196.075 81.365 196.245 ;
        RECT 81.535 196.345 82.215 196.675 ;
        RECT 82.430 196.345 82.680 196.675 ;
        RECT 82.850 196.385 83.100 196.845 ;
        RECT 79.675 195.905 79.845 196.045 ;
        RECT 78.520 195.865 79.485 195.875 ;
        RECT 78.180 195.695 78.350 195.785 ;
        RECT 78.810 195.705 79.485 195.865 ;
        RECT 76.220 195.505 76.960 195.535 ;
        RECT 76.220 195.205 77.135 195.505 ;
        RECT 76.810 195.030 77.135 195.205 ;
        RECT 75.840 194.475 76.095 195.005 ;
        RECT 76.265 194.295 76.570 194.755 ;
        RECT 76.815 194.675 77.135 195.030 ;
        RECT 77.305 195.245 77.845 195.615 ;
        RECT 78.180 195.525 78.585 195.695 ;
        RECT 77.305 194.845 77.545 195.245 ;
        RECT 78.025 195.075 78.245 195.355 ;
        RECT 77.715 194.905 78.245 195.075 ;
        RECT 77.715 194.675 77.885 194.905 ;
        RECT 78.415 194.745 78.585 195.525 ;
        RECT 78.755 194.915 79.105 195.535 ;
        RECT 79.275 194.915 79.485 195.705 ;
        RECT 79.675 195.735 81.175 195.905 ;
        RECT 79.675 195.045 79.845 195.735 ;
        RECT 81.535 195.565 81.705 196.345 ;
        RECT 82.510 196.215 82.680 196.345 ;
        RECT 80.015 195.395 81.705 195.565 ;
        RECT 81.875 195.785 82.340 196.175 ;
        RECT 82.510 196.045 82.905 196.215 ;
        RECT 80.015 195.215 80.185 195.395 ;
        RECT 76.815 194.505 77.885 194.675 ;
        RECT 78.055 194.295 78.245 194.735 ;
        RECT 78.415 194.465 79.365 194.745 ;
        RECT 79.675 194.655 79.935 195.045 ;
        RECT 80.355 194.975 81.145 195.225 ;
        RECT 79.585 194.485 79.935 194.655 ;
        RECT 80.145 194.295 80.475 194.755 ;
        RECT 81.350 194.685 81.520 195.395 ;
        RECT 81.875 195.195 82.045 195.785 ;
        RECT 81.690 194.975 82.045 195.195 ;
        RECT 82.215 194.975 82.565 195.595 ;
        RECT 82.735 194.685 82.905 196.045 ;
        RECT 83.270 195.875 83.595 196.660 ;
        RECT 83.075 194.825 83.535 195.875 ;
        RECT 81.350 194.515 82.205 194.685 ;
        RECT 82.410 194.515 82.905 194.685 ;
        RECT 83.075 194.295 83.405 194.655 ;
        RECT 83.765 194.555 83.935 196.675 ;
        RECT 84.105 196.345 84.435 196.845 ;
        RECT 84.605 196.175 84.860 196.675 ;
        RECT 84.110 196.005 84.860 196.175 ;
        RECT 84.110 195.015 84.340 196.005 ;
        RECT 84.510 195.185 84.860 195.835 ;
        RECT 85.035 195.755 88.545 196.845 ;
        RECT 88.720 196.410 94.065 196.845 ;
        RECT 94.240 196.410 99.585 196.845 ;
        RECT 85.035 195.235 86.725 195.755 ;
        RECT 86.895 195.065 88.545 195.585 ;
        RECT 90.310 195.160 90.660 196.410 ;
        RECT 84.110 194.845 84.860 195.015 ;
        RECT 84.105 194.295 84.435 194.675 ;
        RECT 84.605 194.555 84.860 194.845 ;
        RECT 85.035 194.295 88.545 195.065 ;
        RECT 92.140 194.840 92.480 195.670 ;
        RECT 95.830 195.160 96.180 196.410 ;
        RECT 99.755 195.680 100.045 196.845 ;
        RECT 100.675 195.755 102.345 196.845 ;
        RECT 102.520 196.410 107.865 196.845 ;
        RECT 108.040 196.410 113.385 196.845 ;
        RECT 113.560 196.410 118.905 196.845 ;
        RECT 119.080 196.410 124.425 196.845 ;
        RECT 97.660 194.840 98.000 195.670 ;
        RECT 100.675 195.235 101.425 195.755 ;
        RECT 101.595 195.065 102.345 195.585 ;
        RECT 104.110 195.160 104.460 196.410 ;
        RECT 88.720 194.295 94.065 194.840 ;
        RECT 94.240 194.295 99.585 194.840 ;
        RECT 99.755 194.295 100.045 195.020 ;
        RECT 100.675 194.295 102.345 195.065 ;
        RECT 105.940 194.840 106.280 195.670 ;
        RECT 109.630 195.160 109.980 196.410 ;
        RECT 111.460 194.840 111.800 195.670 ;
        RECT 115.150 195.160 115.500 196.410 ;
        RECT 116.980 194.840 117.320 195.670 ;
        RECT 120.670 195.160 121.020 196.410 ;
        RECT 124.595 195.755 125.805 196.845 ;
        RECT 122.500 194.840 122.840 195.670 ;
        RECT 124.595 195.215 125.115 195.755 ;
        RECT 125.285 195.045 125.805 195.585 ;
        RECT 102.520 194.295 107.865 194.840 ;
        RECT 108.040 194.295 113.385 194.840 ;
        RECT 113.560 194.295 118.905 194.840 ;
        RECT 119.080 194.295 124.425 194.840 ;
        RECT 124.595 194.295 125.805 195.045 ;
        RECT 11.810 194.125 125.890 194.295 ;
        RECT 11.895 193.375 13.105 194.125 ;
        RECT 13.280 193.580 18.625 194.125 ;
        RECT 18.800 193.580 24.145 194.125 ;
        RECT 24.320 193.580 29.665 194.125 ;
        RECT 29.840 193.580 35.185 194.125 ;
        RECT 11.895 192.835 12.415 193.375 ;
        RECT 12.585 192.665 13.105 193.205 ;
        RECT 11.895 191.575 13.105 192.665 ;
        RECT 14.870 192.010 15.220 193.260 ;
        RECT 16.700 192.750 17.040 193.580 ;
        RECT 20.390 192.010 20.740 193.260 ;
        RECT 22.220 192.750 22.560 193.580 ;
        RECT 25.910 192.010 26.260 193.260 ;
        RECT 27.740 192.750 28.080 193.580 ;
        RECT 31.430 192.010 31.780 193.260 ;
        RECT 33.260 192.750 33.600 193.580 ;
        RECT 35.355 193.400 35.645 194.125 ;
        RECT 36.275 193.355 38.865 194.125 ;
        RECT 39.040 193.580 44.385 194.125 ;
        RECT 44.560 193.580 49.905 194.125 ;
        RECT 50.080 193.580 55.425 194.125 ;
        RECT 55.600 193.580 60.945 194.125 ;
        RECT 13.280 191.575 18.625 192.010 ;
        RECT 18.800 191.575 24.145 192.010 ;
        RECT 24.320 191.575 29.665 192.010 ;
        RECT 29.840 191.575 35.185 192.010 ;
        RECT 35.355 191.575 35.645 192.740 ;
        RECT 36.275 192.665 37.485 193.185 ;
        RECT 37.655 192.835 38.865 193.355 ;
        RECT 36.275 191.575 38.865 192.665 ;
        RECT 40.630 192.010 40.980 193.260 ;
        RECT 42.460 192.750 42.800 193.580 ;
        RECT 46.150 192.010 46.500 193.260 ;
        RECT 47.980 192.750 48.320 193.580 ;
        RECT 51.670 192.010 52.020 193.260 ;
        RECT 53.500 192.750 53.840 193.580 ;
        RECT 57.190 192.010 57.540 193.260 ;
        RECT 59.020 192.750 59.360 193.580 ;
        RECT 61.115 193.400 61.405 194.125 ;
        RECT 61.575 193.355 63.245 194.125 ;
        RECT 39.040 191.575 44.385 192.010 ;
        RECT 44.560 191.575 49.905 192.010 ;
        RECT 50.080 191.575 55.425 192.010 ;
        RECT 55.600 191.575 60.945 192.010 ;
        RECT 61.115 191.575 61.405 192.740 ;
        RECT 61.575 192.665 62.325 193.185 ;
        RECT 62.495 192.835 63.245 193.355 ;
        RECT 63.455 193.305 63.685 194.125 ;
        RECT 63.855 193.325 64.185 193.955 ;
        RECT 63.435 192.885 63.765 193.135 ;
        RECT 63.935 192.725 64.185 193.325 ;
        RECT 64.355 193.305 64.565 194.125 ;
        RECT 65.805 193.575 65.975 193.955 ;
        RECT 66.190 193.745 66.520 194.125 ;
        RECT 65.805 193.405 66.520 193.575 ;
        RECT 65.715 192.855 66.070 193.225 ;
        RECT 66.350 193.215 66.520 193.405 ;
        RECT 66.690 193.380 66.945 193.955 ;
        RECT 66.350 192.885 66.605 193.215 ;
        RECT 61.575 191.575 63.245 192.665 ;
        RECT 63.455 191.575 63.685 192.715 ;
        RECT 63.855 191.745 64.185 192.725 ;
        RECT 64.355 191.575 64.565 192.715 ;
        RECT 66.350 192.675 66.520 192.885 ;
        RECT 65.805 192.505 66.520 192.675 ;
        RECT 66.775 192.650 66.945 193.380 ;
        RECT 67.120 193.285 67.380 194.125 ;
        RECT 67.565 193.400 67.895 193.910 ;
        RECT 68.065 193.725 68.395 194.125 ;
        RECT 69.445 193.555 69.775 193.895 ;
        RECT 69.945 193.725 70.275 194.125 ;
        RECT 65.805 191.745 65.975 192.505 ;
        RECT 66.190 191.575 66.520 192.335 ;
        RECT 66.690 191.745 66.945 192.650 ;
        RECT 67.120 191.575 67.380 192.725 ;
        RECT 67.565 192.635 67.755 193.400 ;
        RECT 68.065 193.385 70.430 193.555 ;
        RECT 68.065 193.215 68.235 193.385 ;
        RECT 67.925 192.885 68.235 193.215 ;
        RECT 68.405 192.885 68.710 193.215 ;
        RECT 67.565 191.785 67.895 192.635 ;
        RECT 68.065 191.575 68.315 192.715 ;
        RECT 68.495 192.555 68.710 192.885 ;
        RECT 68.885 192.555 69.170 193.215 ;
        RECT 69.365 192.555 69.630 193.215 ;
        RECT 69.845 192.555 70.090 193.215 ;
        RECT 70.260 192.385 70.430 193.385 ;
        RECT 68.505 192.215 69.795 192.385 ;
        RECT 68.505 191.795 68.755 192.215 ;
        RECT 68.985 191.575 69.315 192.045 ;
        RECT 69.545 191.795 69.795 192.215 ;
        RECT 69.975 192.215 70.430 192.385 ;
        RECT 71.695 193.385 72.015 193.865 ;
        RECT 72.185 193.555 72.415 193.955 ;
        RECT 72.585 193.735 72.935 194.125 ;
        RECT 72.185 193.475 72.695 193.555 ;
        RECT 73.105 193.475 73.435 193.955 ;
        RECT 72.185 193.385 73.435 193.475 ;
        RECT 71.695 192.455 71.865 193.385 ;
        RECT 72.525 193.305 73.435 193.385 ;
        RECT 73.605 193.305 73.775 194.125 ;
        RECT 74.280 193.385 74.745 193.930 ;
        RECT 72.035 192.795 72.205 193.215 ;
        RECT 72.435 192.965 73.035 193.135 ;
        RECT 72.035 192.625 72.695 192.795 ;
        RECT 71.695 192.255 72.355 192.455 ;
        RECT 72.525 192.425 72.695 192.625 ;
        RECT 72.865 192.765 73.035 192.965 ;
        RECT 73.205 192.935 73.900 193.135 ;
        RECT 74.160 192.765 74.405 193.215 ;
        RECT 72.865 192.595 74.405 192.765 ;
        RECT 74.575 192.425 74.745 193.385 ;
        RECT 72.525 192.255 74.745 192.425 ;
        RECT 74.920 193.415 75.175 193.945 ;
        RECT 75.345 193.665 75.650 194.125 ;
        RECT 75.895 193.745 76.965 193.915 ;
        RECT 74.920 192.765 75.130 193.415 ;
        RECT 75.895 193.390 76.215 193.745 ;
        RECT 75.890 193.215 76.215 193.390 ;
        RECT 75.300 192.915 76.215 193.215 ;
        RECT 76.385 193.175 76.625 193.575 ;
        RECT 76.795 193.515 76.965 193.745 ;
        RECT 77.135 193.685 77.325 194.125 ;
        RECT 77.495 193.675 78.445 193.955 ;
        RECT 78.665 193.765 79.015 193.935 ;
        RECT 76.795 193.345 77.325 193.515 ;
        RECT 75.300 192.885 76.040 192.915 ;
        RECT 69.975 191.785 70.305 192.215 ;
        RECT 72.185 192.085 72.355 192.255 ;
        RECT 71.715 191.575 72.015 192.085 ;
        RECT 72.185 191.915 72.565 192.085 ;
        RECT 73.145 191.575 73.775 192.085 ;
        RECT 73.945 191.745 74.275 192.255 ;
        RECT 74.445 191.575 74.745 192.085 ;
        RECT 74.920 191.885 75.175 192.765 ;
        RECT 75.345 191.575 75.650 192.715 ;
        RECT 75.870 192.295 76.040 192.885 ;
        RECT 76.385 192.805 76.925 193.175 ;
        RECT 77.105 193.065 77.325 193.345 ;
        RECT 77.495 192.895 77.665 193.675 ;
        RECT 77.260 192.725 77.665 192.895 ;
        RECT 77.835 192.885 78.185 193.505 ;
        RECT 77.260 192.635 77.430 192.725 ;
        RECT 78.355 192.715 78.565 193.505 ;
        RECT 76.210 192.465 77.430 192.635 ;
        RECT 77.890 192.555 78.565 192.715 ;
        RECT 75.870 192.125 76.670 192.295 ;
        RECT 75.990 191.575 76.320 191.955 ;
        RECT 76.500 191.835 76.670 192.125 ;
        RECT 77.260 192.085 77.430 192.465 ;
        RECT 77.600 192.545 78.565 192.555 ;
        RECT 78.755 193.375 79.015 193.765 ;
        RECT 79.225 193.665 79.555 194.125 ;
        RECT 80.430 193.735 81.285 193.905 ;
        RECT 81.490 193.735 81.985 193.905 ;
        RECT 82.155 193.765 82.485 194.125 ;
        RECT 78.755 192.685 78.925 193.375 ;
        RECT 79.095 193.025 79.265 193.205 ;
        RECT 79.435 193.195 80.225 193.445 ;
        RECT 80.430 193.025 80.600 193.735 ;
        RECT 80.770 193.225 81.125 193.445 ;
        RECT 79.095 192.855 80.785 193.025 ;
        RECT 77.600 192.255 78.060 192.545 ;
        RECT 78.755 192.515 80.255 192.685 ;
        RECT 78.755 192.375 78.925 192.515 ;
        RECT 78.365 192.205 78.925 192.375 ;
        RECT 76.840 191.575 77.090 192.035 ;
        RECT 77.260 191.745 78.130 192.085 ;
        RECT 78.365 191.745 78.535 192.205 ;
        RECT 79.370 192.175 80.445 192.345 ;
        RECT 78.705 191.575 79.075 192.035 ;
        RECT 79.370 191.835 79.540 192.175 ;
        RECT 79.710 191.575 80.040 192.005 ;
        RECT 80.275 191.835 80.445 192.175 ;
        RECT 80.615 192.075 80.785 192.855 ;
        RECT 80.955 192.635 81.125 193.225 ;
        RECT 81.295 192.825 81.645 193.445 ;
        RECT 80.955 192.245 81.420 192.635 ;
        RECT 81.815 192.375 81.985 193.735 ;
        RECT 82.155 192.545 82.615 193.595 ;
        RECT 81.590 192.205 81.985 192.375 ;
        RECT 81.590 192.075 81.760 192.205 ;
        RECT 80.615 191.745 81.295 192.075 ;
        RECT 81.510 191.745 81.760 192.075 ;
        RECT 81.930 191.575 82.180 192.035 ;
        RECT 82.350 191.760 82.675 192.545 ;
        RECT 82.845 191.745 83.015 193.865 ;
        RECT 83.185 193.745 83.515 194.125 ;
        RECT 83.685 193.575 83.940 193.865 ;
        RECT 83.190 193.405 83.940 193.575 ;
        RECT 83.190 192.415 83.420 193.405 ;
        RECT 84.175 193.305 84.385 194.125 ;
        RECT 84.555 193.325 84.885 193.955 ;
        RECT 83.590 192.585 83.940 193.235 ;
        RECT 84.555 192.725 84.805 193.325 ;
        RECT 85.055 193.305 85.285 194.125 ;
        RECT 85.495 193.375 86.705 194.125 ;
        RECT 86.875 193.400 87.165 194.125 ;
        RECT 84.975 192.885 85.305 193.135 ;
        RECT 83.190 192.245 83.940 192.415 ;
        RECT 83.185 191.575 83.515 192.075 ;
        RECT 83.685 191.745 83.940 192.245 ;
        RECT 84.175 191.575 84.385 192.715 ;
        RECT 84.555 191.745 84.885 192.725 ;
        RECT 85.055 191.575 85.285 192.715 ;
        RECT 85.495 192.665 86.015 193.205 ;
        RECT 86.185 192.835 86.705 193.375 ;
        RECT 87.335 193.355 90.845 194.125 ;
        RECT 91.020 193.580 96.365 194.125 ;
        RECT 85.495 191.575 86.705 192.665 ;
        RECT 86.875 191.575 87.165 192.740 ;
        RECT 87.335 192.665 89.025 193.185 ;
        RECT 89.195 192.835 90.845 193.355 ;
        RECT 87.335 191.575 90.845 192.665 ;
        RECT 92.610 192.010 92.960 193.260 ;
        RECT 94.440 192.750 94.780 193.580 ;
        RECT 96.540 193.415 96.795 193.945 ;
        RECT 96.965 193.665 97.270 194.125 ;
        RECT 97.515 193.745 98.585 193.915 ;
        RECT 96.540 192.765 96.750 193.415 ;
        RECT 97.515 193.390 97.835 193.745 ;
        RECT 97.510 193.215 97.835 193.390 ;
        RECT 96.920 192.915 97.835 193.215 ;
        RECT 98.005 193.175 98.245 193.575 ;
        RECT 98.415 193.515 98.585 193.745 ;
        RECT 98.755 193.685 98.945 194.125 ;
        RECT 99.115 193.675 100.065 193.955 ;
        RECT 100.285 193.765 100.635 193.935 ;
        RECT 98.415 193.345 98.945 193.515 ;
        RECT 96.920 192.885 97.660 192.915 ;
        RECT 91.020 191.575 96.365 192.010 ;
        RECT 96.540 191.885 96.795 192.765 ;
        RECT 96.965 191.575 97.270 192.715 ;
        RECT 97.490 192.295 97.660 192.885 ;
        RECT 98.005 192.805 98.545 193.175 ;
        RECT 98.725 193.065 98.945 193.345 ;
        RECT 99.115 192.895 99.285 193.675 ;
        RECT 98.880 192.725 99.285 192.895 ;
        RECT 99.455 192.885 99.805 193.505 ;
        RECT 98.880 192.635 99.050 192.725 ;
        RECT 99.975 192.715 100.185 193.505 ;
        RECT 97.830 192.465 99.050 192.635 ;
        RECT 99.510 192.555 100.185 192.715 ;
        RECT 97.490 192.125 98.290 192.295 ;
        RECT 97.610 191.575 97.940 191.955 ;
        RECT 98.120 191.835 98.290 192.125 ;
        RECT 98.880 192.085 99.050 192.465 ;
        RECT 99.220 192.545 100.185 192.555 ;
        RECT 100.375 193.375 100.635 193.765 ;
        RECT 100.845 193.665 101.175 194.125 ;
        RECT 102.050 193.735 102.905 193.905 ;
        RECT 103.110 193.735 103.605 193.905 ;
        RECT 103.775 193.765 104.105 194.125 ;
        RECT 100.375 192.685 100.545 193.375 ;
        RECT 100.715 193.025 100.885 193.205 ;
        RECT 101.055 193.195 101.845 193.445 ;
        RECT 102.050 193.025 102.220 193.735 ;
        RECT 102.390 193.225 102.745 193.445 ;
        RECT 100.715 192.855 102.405 193.025 ;
        RECT 99.220 192.255 99.680 192.545 ;
        RECT 100.375 192.515 101.875 192.685 ;
        RECT 100.375 192.375 100.545 192.515 ;
        RECT 99.985 192.205 100.545 192.375 ;
        RECT 98.460 191.575 98.710 192.035 ;
        RECT 98.880 191.745 99.750 192.085 ;
        RECT 99.985 191.745 100.155 192.205 ;
        RECT 100.990 192.175 102.065 192.345 ;
        RECT 100.325 191.575 100.695 192.035 ;
        RECT 100.990 191.835 101.160 192.175 ;
        RECT 101.330 191.575 101.660 192.005 ;
        RECT 101.895 191.835 102.065 192.175 ;
        RECT 102.235 192.075 102.405 192.855 ;
        RECT 102.575 192.635 102.745 193.225 ;
        RECT 102.915 192.825 103.265 193.445 ;
        RECT 102.575 192.245 103.040 192.635 ;
        RECT 103.435 192.375 103.605 193.735 ;
        RECT 103.775 192.545 104.235 193.595 ;
        RECT 103.210 192.205 103.605 192.375 ;
        RECT 103.210 192.075 103.380 192.205 ;
        RECT 102.235 191.745 102.915 192.075 ;
        RECT 103.130 191.745 103.380 192.075 ;
        RECT 103.550 191.575 103.800 192.035 ;
        RECT 103.970 191.760 104.295 192.545 ;
        RECT 104.465 191.745 104.635 193.865 ;
        RECT 104.805 193.745 105.135 194.125 ;
        RECT 105.305 193.575 105.560 193.865 ;
        RECT 104.810 193.405 105.560 193.575 ;
        RECT 104.810 192.415 105.040 193.405 ;
        RECT 105.775 193.305 106.005 194.125 ;
        RECT 106.175 193.325 106.505 193.955 ;
        RECT 105.210 192.585 105.560 193.235 ;
        RECT 105.755 192.885 106.085 193.135 ;
        RECT 106.255 192.725 106.505 193.325 ;
        RECT 106.675 193.305 106.885 194.125 ;
        RECT 107.665 193.575 107.835 193.955 ;
        RECT 108.015 193.745 108.345 194.125 ;
        RECT 107.665 193.405 108.330 193.575 ;
        RECT 108.525 193.450 108.785 193.955 ;
        RECT 107.595 192.855 107.925 193.225 ;
        RECT 108.160 193.150 108.330 193.405 ;
        RECT 104.810 192.245 105.560 192.415 ;
        RECT 104.805 191.575 105.135 192.075 ;
        RECT 105.305 191.745 105.560 192.245 ;
        RECT 105.775 191.575 106.005 192.715 ;
        RECT 106.175 191.745 106.505 192.725 ;
        RECT 108.160 192.820 108.445 193.150 ;
        RECT 106.675 191.575 106.885 192.715 ;
        RECT 108.160 192.675 108.330 192.820 ;
        RECT 107.665 192.505 108.330 192.675 ;
        RECT 108.615 192.650 108.785 193.450 ;
        RECT 108.955 193.355 112.465 194.125 ;
        RECT 112.635 193.400 112.925 194.125 ;
        RECT 113.560 193.580 118.905 194.125 ;
        RECT 119.080 193.580 124.425 194.125 ;
        RECT 107.665 191.745 107.835 192.505 ;
        RECT 108.015 191.575 108.345 192.335 ;
        RECT 108.515 191.745 108.785 192.650 ;
        RECT 108.955 192.665 110.645 193.185 ;
        RECT 110.815 192.835 112.465 193.355 ;
        RECT 108.955 191.575 112.465 192.665 ;
        RECT 112.635 191.575 112.925 192.740 ;
        RECT 115.150 192.010 115.500 193.260 ;
        RECT 116.980 192.750 117.320 193.580 ;
        RECT 120.670 192.010 121.020 193.260 ;
        RECT 122.500 192.750 122.840 193.580 ;
        RECT 124.595 193.375 125.805 194.125 ;
        RECT 124.595 192.665 125.115 193.205 ;
        RECT 125.285 192.835 125.805 193.375 ;
        RECT 113.560 191.575 118.905 192.010 ;
        RECT 119.080 191.575 124.425 192.010 ;
        RECT 124.595 191.575 125.805 192.665 ;
        RECT 11.810 191.405 125.890 191.575 ;
        RECT 11.895 190.315 13.105 191.405 ;
        RECT 11.895 189.605 12.415 190.145 ;
        RECT 12.585 189.775 13.105 190.315 ;
        RECT 13.275 190.315 16.785 191.405 ;
        RECT 16.960 190.970 22.305 191.405 ;
        RECT 13.275 189.795 14.965 190.315 ;
        RECT 15.135 189.625 16.785 190.145 ;
        RECT 18.550 189.720 18.900 190.970 ;
        RECT 22.475 190.240 22.765 191.405 ;
        RECT 23.395 190.315 25.985 191.405 ;
        RECT 26.160 190.970 31.505 191.405 ;
        RECT 31.680 190.970 37.025 191.405 ;
        RECT 37.200 190.970 42.545 191.405 ;
        RECT 42.720 190.970 48.065 191.405 ;
        RECT 11.895 188.855 13.105 189.605 ;
        RECT 13.275 188.855 16.785 189.625 ;
        RECT 20.380 189.400 20.720 190.230 ;
        RECT 23.395 189.795 24.605 190.315 ;
        RECT 24.775 189.625 25.985 190.145 ;
        RECT 27.750 189.720 28.100 190.970 ;
        RECT 16.960 188.855 22.305 189.400 ;
        RECT 22.475 188.855 22.765 189.580 ;
        RECT 23.395 188.855 25.985 189.625 ;
        RECT 29.580 189.400 29.920 190.230 ;
        RECT 33.270 189.720 33.620 190.970 ;
        RECT 35.100 189.400 35.440 190.230 ;
        RECT 38.790 189.720 39.140 190.970 ;
        RECT 40.620 189.400 40.960 190.230 ;
        RECT 44.310 189.720 44.660 190.970 ;
        RECT 48.235 190.240 48.525 191.405 ;
        RECT 49.155 190.315 52.665 191.405 ;
        RECT 52.840 190.970 58.185 191.405 ;
        RECT 58.360 190.970 63.705 191.405 ;
        RECT 46.140 189.400 46.480 190.230 ;
        RECT 49.155 189.795 50.845 190.315 ;
        RECT 51.015 189.625 52.665 190.145 ;
        RECT 54.430 189.720 54.780 190.970 ;
        RECT 26.160 188.855 31.505 189.400 ;
        RECT 31.680 188.855 37.025 189.400 ;
        RECT 37.200 188.855 42.545 189.400 ;
        RECT 42.720 188.855 48.065 189.400 ;
        RECT 48.235 188.855 48.525 189.580 ;
        RECT 49.155 188.855 52.665 189.625 ;
        RECT 56.260 189.400 56.600 190.230 ;
        RECT 59.950 189.720 60.300 190.970 ;
        RECT 63.875 190.435 64.145 191.205 ;
        RECT 64.315 190.625 64.645 191.405 ;
        RECT 64.850 190.800 65.035 191.205 ;
        RECT 65.205 190.980 65.540 191.405 ;
        RECT 64.850 190.625 65.515 190.800 ;
        RECT 63.875 190.265 65.005 190.435 ;
        RECT 61.780 189.400 62.120 190.230 ;
        RECT 52.840 188.855 58.185 189.400 ;
        RECT 58.360 188.855 63.705 189.400 ;
        RECT 63.875 189.355 64.045 190.265 ;
        RECT 64.215 189.515 64.575 190.095 ;
        RECT 64.755 189.765 65.005 190.265 ;
        RECT 65.175 189.595 65.515 190.625 ;
        RECT 65.800 190.785 65.975 191.235 ;
        RECT 66.145 190.965 66.475 191.405 ;
        RECT 66.780 190.815 66.950 191.235 ;
        RECT 67.185 190.995 67.855 191.405 ;
        RECT 68.070 190.815 68.240 191.235 ;
        RECT 68.440 190.995 68.770 191.405 ;
        RECT 65.800 190.615 66.430 190.785 ;
        RECT 65.715 189.765 66.080 190.445 ;
        RECT 66.260 190.095 66.430 190.615 ;
        RECT 66.780 190.645 68.795 190.815 ;
        RECT 66.260 189.765 66.610 190.095 ;
        RECT 66.260 189.595 66.430 189.765 ;
        RECT 64.830 189.425 65.515 189.595 ;
        RECT 65.800 189.425 66.430 189.595 ;
        RECT 63.875 189.025 64.135 189.355 ;
        RECT 64.345 188.855 64.620 189.335 ;
        RECT 64.830 189.025 65.035 189.425 ;
        RECT 65.205 188.855 65.540 189.255 ;
        RECT 65.800 189.025 65.975 189.425 ;
        RECT 66.780 189.355 66.950 190.645 ;
        RECT 66.145 188.855 66.475 189.235 ;
        RECT 66.720 189.025 66.950 189.355 ;
        RECT 67.150 189.190 67.430 190.465 ;
        RECT 67.655 189.365 67.925 190.465 ;
        RECT 68.115 189.435 68.455 190.465 ;
        RECT 68.625 190.095 68.795 190.645 ;
        RECT 68.965 190.265 69.225 191.235 ;
        RECT 68.625 189.765 68.885 190.095 ;
        RECT 69.055 189.575 69.225 190.265 ;
        RECT 67.615 189.195 67.925 189.365 ;
        RECT 67.655 189.190 67.925 189.195 ;
        RECT 68.385 188.855 68.715 189.235 ;
        RECT 68.885 189.110 69.225 189.575 ;
        RECT 69.395 190.905 69.655 191.235 ;
        RECT 69.965 191.025 70.295 191.405 ;
        RECT 69.395 190.225 69.565 190.905 ;
        RECT 70.535 190.855 70.725 191.235 ;
        RECT 70.975 191.025 71.305 191.405 ;
        RECT 71.515 190.855 71.685 191.235 ;
        RECT 71.880 191.025 72.210 191.405 ;
        RECT 72.470 190.855 72.640 191.235 ;
        RECT 73.065 191.025 73.395 191.405 ;
        RECT 69.735 190.395 70.085 190.725 ;
        RECT 70.535 190.685 71.275 190.855 ;
        RECT 70.355 190.345 70.935 190.515 ;
        RECT 70.355 190.225 70.525 190.345 ;
        RECT 69.395 190.055 70.525 190.225 ;
        RECT 71.105 190.175 71.275 190.685 ;
        RECT 69.395 189.355 69.565 190.055 ;
        RECT 70.705 190.005 71.275 190.175 ;
        RECT 71.445 190.685 73.395 190.855 ;
        RECT 69.915 189.715 70.535 189.885 ;
        RECT 69.915 189.535 70.125 189.715 ;
        RECT 70.705 189.525 70.875 190.005 ;
        RECT 71.445 189.695 71.615 190.685 ;
        RECT 72.205 190.095 72.390 190.405 ;
        RECT 72.660 190.095 72.855 190.405 ;
        RECT 68.885 189.065 69.220 189.110 ;
        RECT 69.395 189.025 69.655 189.355 ;
        RECT 69.965 188.855 70.295 189.235 ;
        RECT 70.475 189.195 70.875 189.525 ;
        RECT 71.065 189.365 71.615 189.695 ;
        RECT 71.785 189.195 71.955 190.095 ;
        RECT 70.475 189.025 71.955 189.195 ;
        RECT 72.205 189.765 72.435 190.095 ;
        RECT 72.660 189.765 72.915 190.095 ;
        RECT 73.225 189.765 73.395 190.685 ;
        RECT 72.205 189.185 72.390 189.765 ;
        RECT 72.660 189.190 72.855 189.765 ;
        RECT 73.065 188.855 73.395 189.235 ;
        RECT 73.565 189.025 73.825 191.235 ;
        RECT 73.995 190.240 74.285 191.405 ;
        RECT 74.490 190.615 75.025 191.235 ;
        RECT 74.490 189.595 74.805 190.615 ;
        RECT 75.195 190.605 75.525 191.405 ;
        RECT 76.010 190.435 76.400 190.610 ;
        RECT 74.975 190.265 76.400 190.435 ;
        RECT 76.755 190.435 77.025 191.205 ;
        RECT 77.195 190.625 77.525 191.405 ;
        RECT 77.730 190.800 77.915 191.205 ;
        RECT 78.085 190.980 78.420 191.405 ;
        RECT 77.730 190.625 78.395 190.800 ;
        RECT 76.755 190.265 77.885 190.435 ;
        RECT 74.975 189.765 75.145 190.265 ;
        RECT 73.995 188.855 74.285 189.580 ;
        RECT 74.490 189.025 75.105 189.595 ;
        RECT 75.395 189.535 75.660 190.095 ;
        RECT 75.830 189.365 76.000 190.265 ;
        RECT 76.170 189.535 76.525 190.095 ;
        RECT 75.275 188.855 75.490 189.365 ;
        RECT 75.720 189.035 76.000 189.365 ;
        RECT 76.180 188.855 76.420 189.365 ;
        RECT 76.755 189.355 76.925 190.265 ;
        RECT 77.095 189.515 77.455 190.095 ;
        RECT 77.635 189.765 77.885 190.265 ;
        RECT 78.055 189.595 78.395 190.625 ;
        RECT 79.095 190.265 79.325 191.405 ;
        RECT 79.495 190.255 79.825 191.235 ;
        RECT 79.995 190.265 80.205 191.405 ;
        RECT 80.525 190.475 80.695 191.235 ;
        RECT 80.875 190.645 81.205 191.405 ;
        RECT 80.525 190.305 81.190 190.475 ;
        RECT 81.375 190.330 81.645 191.235 ;
        RECT 79.075 189.845 79.405 190.095 ;
        RECT 77.710 189.425 78.395 189.595 ;
        RECT 76.755 189.025 77.015 189.355 ;
        RECT 77.225 188.855 77.500 189.335 ;
        RECT 77.710 189.025 77.915 189.425 ;
        RECT 78.085 188.855 78.420 189.255 ;
        RECT 79.095 188.855 79.325 189.675 ;
        RECT 79.575 189.655 79.825 190.255 ;
        RECT 81.020 190.160 81.190 190.305 ;
        RECT 80.455 189.755 80.785 190.125 ;
        RECT 81.020 189.830 81.305 190.160 ;
        RECT 79.495 189.025 79.825 189.655 ;
        RECT 79.995 188.855 80.205 189.675 ;
        RECT 81.020 189.575 81.190 189.830 ;
        RECT 80.525 189.405 81.190 189.575 ;
        RECT 81.475 189.530 81.645 190.330 ;
        RECT 81.815 190.315 84.405 191.405 ;
        RECT 84.580 190.970 89.925 191.405 ;
        RECT 81.815 189.795 83.025 190.315 ;
        RECT 83.195 189.625 84.405 190.145 ;
        RECT 86.170 189.720 86.520 190.970 ;
        RECT 90.155 190.265 90.365 191.405 ;
        RECT 90.535 190.255 90.865 191.235 ;
        RECT 91.035 190.265 91.265 191.405 ;
        RECT 92.485 190.475 92.655 191.235 ;
        RECT 92.835 190.645 93.165 191.405 ;
        RECT 92.485 190.305 93.150 190.475 ;
        RECT 93.335 190.330 93.605 191.235 ;
        RECT 80.525 189.025 80.695 189.405 ;
        RECT 80.875 188.855 81.205 189.235 ;
        RECT 81.385 189.025 81.645 189.530 ;
        RECT 81.815 188.855 84.405 189.625 ;
        RECT 88.000 189.400 88.340 190.230 ;
        RECT 84.580 188.855 89.925 189.400 ;
        RECT 90.155 188.855 90.365 189.675 ;
        RECT 90.535 189.655 90.785 190.255 ;
        RECT 92.980 190.160 93.150 190.305 ;
        RECT 90.955 189.845 91.285 190.095 ;
        RECT 92.415 189.755 92.745 190.125 ;
        RECT 92.980 189.830 93.265 190.160 ;
        RECT 90.535 189.025 90.865 189.655 ;
        RECT 91.035 188.855 91.265 189.675 ;
        RECT 92.980 189.575 93.150 189.830 ;
        RECT 92.485 189.405 93.150 189.575 ;
        RECT 93.435 189.530 93.605 190.330 ;
        RECT 94.695 190.315 98.205 191.405 ;
        RECT 94.695 189.795 96.385 190.315 ;
        RECT 98.415 190.265 98.645 191.405 ;
        RECT 98.815 190.255 99.145 191.235 ;
        RECT 99.315 190.265 99.525 191.405 ;
        RECT 96.555 189.625 98.205 190.145 ;
        RECT 98.395 189.845 98.725 190.095 ;
        RECT 92.485 189.025 92.655 189.405 ;
        RECT 92.835 188.855 93.165 189.235 ;
        RECT 93.345 189.025 93.605 189.530 ;
        RECT 94.695 188.855 98.205 189.625 ;
        RECT 98.415 188.855 98.645 189.675 ;
        RECT 98.895 189.655 99.145 190.255 ;
        RECT 99.755 190.240 100.045 191.405 ;
        RECT 100.675 190.315 102.345 191.405 ;
        RECT 100.675 189.795 101.425 190.315 ;
        RECT 102.520 190.215 102.775 191.095 ;
        RECT 102.945 190.265 103.250 191.405 ;
        RECT 103.590 191.025 103.920 191.405 ;
        RECT 104.100 190.855 104.270 191.145 ;
        RECT 104.440 190.945 104.690 191.405 ;
        RECT 103.470 190.685 104.270 190.855 ;
        RECT 104.860 190.895 105.730 191.235 ;
        RECT 98.815 189.025 99.145 189.655 ;
        RECT 99.315 188.855 99.525 189.675 ;
        RECT 101.595 189.625 102.345 190.145 ;
        RECT 99.755 188.855 100.045 189.580 ;
        RECT 100.675 188.855 102.345 189.625 ;
        RECT 102.520 189.565 102.730 190.215 ;
        RECT 103.470 190.095 103.640 190.685 ;
        RECT 104.860 190.515 105.030 190.895 ;
        RECT 105.965 190.775 106.135 191.235 ;
        RECT 106.305 190.945 106.675 191.405 ;
        RECT 106.970 190.805 107.140 191.145 ;
        RECT 107.310 190.975 107.640 191.405 ;
        RECT 107.875 190.805 108.045 191.145 ;
        RECT 103.810 190.345 105.030 190.515 ;
        RECT 105.200 190.435 105.660 190.725 ;
        RECT 105.965 190.605 106.525 190.775 ;
        RECT 106.970 190.635 108.045 190.805 ;
        RECT 108.215 190.905 108.895 191.235 ;
        RECT 109.110 190.905 109.360 191.235 ;
        RECT 109.530 190.945 109.780 191.405 ;
        RECT 106.355 190.465 106.525 190.605 ;
        RECT 105.200 190.425 106.165 190.435 ;
        RECT 104.860 190.255 105.030 190.345 ;
        RECT 105.490 190.265 106.165 190.425 ;
        RECT 102.900 190.065 103.640 190.095 ;
        RECT 102.900 189.765 103.815 190.065 ;
        RECT 103.490 189.590 103.815 189.765 ;
        RECT 102.520 189.035 102.775 189.565 ;
        RECT 102.945 188.855 103.250 189.315 ;
        RECT 103.495 189.235 103.815 189.590 ;
        RECT 103.985 189.805 104.525 190.175 ;
        RECT 104.860 190.085 105.265 190.255 ;
        RECT 103.985 189.405 104.225 189.805 ;
        RECT 104.705 189.635 104.925 189.915 ;
        RECT 104.395 189.465 104.925 189.635 ;
        RECT 104.395 189.235 104.565 189.465 ;
        RECT 105.095 189.305 105.265 190.085 ;
        RECT 105.435 189.475 105.785 190.095 ;
        RECT 105.955 189.475 106.165 190.265 ;
        RECT 106.355 190.295 107.855 190.465 ;
        RECT 106.355 189.605 106.525 190.295 ;
        RECT 108.215 190.125 108.385 190.905 ;
        RECT 109.190 190.775 109.360 190.905 ;
        RECT 106.695 189.955 108.385 190.125 ;
        RECT 108.555 190.345 109.020 190.735 ;
        RECT 109.190 190.605 109.585 190.775 ;
        RECT 106.695 189.775 106.865 189.955 ;
        RECT 103.495 189.065 104.565 189.235 ;
        RECT 104.735 188.855 104.925 189.295 ;
        RECT 105.095 189.025 106.045 189.305 ;
        RECT 106.355 189.215 106.615 189.605 ;
        RECT 107.035 189.535 107.825 189.785 ;
        RECT 106.265 189.045 106.615 189.215 ;
        RECT 106.825 188.855 107.155 189.315 ;
        RECT 108.030 189.245 108.200 189.955 ;
        RECT 108.555 189.755 108.725 190.345 ;
        RECT 108.370 189.535 108.725 189.755 ;
        RECT 108.895 189.535 109.245 190.155 ;
        RECT 109.415 189.245 109.585 190.605 ;
        RECT 109.950 190.435 110.275 191.220 ;
        RECT 109.755 189.385 110.215 190.435 ;
        RECT 108.030 189.075 108.885 189.245 ;
        RECT 109.090 189.075 109.585 189.245 ;
        RECT 109.755 188.855 110.085 189.215 ;
        RECT 110.445 189.115 110.615 191.235 ;
        RECT 110.785 190.905 111.115 191.405 ;
        RECT 111.285 190.735 111.540 191.235 ;
        RECT 110.790 190.565 111.540 190.735 ;
        RECT 110.790 189.575 111.020 190.565 ;
        RECT 111.190 189.745 111.540 190.395 ;
        RECT 111.715 190.315 113.385 191.405 ;
        RECT 113.560 190.970 118.905 191.405 ;
        RECT 119.080 190.970 124.425 191.405 ;
        RECT 111.715 189.795 112.465 190.315 ;
        RECT 112.635 189.625 113.385 190.145 ;
        RECT 115.150 189.720 115.500 190.970 ;
        RECT 110.790 189.405 111.540 189.575 ;
        RECT 110.785 188.855 111.115 189.235 ;
        RECT 111.285 189.115 111.540 189.405 ;
        RECT 111.715 188.855 113.385 189.625 ;
        RECT 116.980 189.400 117.320 190.230 ;
        RECT 120.670 189.720 121.020 190.970 ;
        RECT 124.595 190.315 125.805 191.405 ;
        RECT 122.500 189.400 122.840 190.230 ;
        RECT 124.595 189.775 125.115 190.315 ;
        RECT 125.285 189.605 125.805 190.145 ;
        RECT 113.560 188.855 118.905 189.400 ;
        RECT 119.080 188.855 124.425 189.400 ;
        RECT 124.595 188.855 125.805 189.605 ;
        RECT 11.810 188.685 125.890 188.855 ;
        RECT 11.895 187.935 13.105 188.685 ;
        RECT 13.280 188.140 18.625 188.685 ;
        RECT 18.800 188.140 24.145 188.685 ;
        RECT 24.320 188.140 29.665 188.685 ;
        RECT 29.840 188.140 35.185 188.685 ;
        RECT 11.895 187.395 12.415 187.935 ;
        RECT 12.585 187.225 13.105 187.765 ;
        RECT 11.895 186.135 13.105 187.225 ;
        RECT 14.870 186.570 15.220 187.820 ;
        RECT 16.700 187.310 17.040 188.140 ;
        RECT 20.390 186.570 20.740 187.820 ;
        RECT 22.220 187.310 22.560 188.140 ;
        RECT 25.910 186.570 26.260 187.820 ;
        RECT 27.740 187.310 28.080 188.140 ;
        RECT 31.430 186.570 31.780 187.820 ;
        RECT 33.260 187.310 33.600 188.140 ;
        RECT 35.355 187.960 35.645 188.685 ;
        RECT 35.815 187.915 38.405 188.685 ;
        RECT 13.280 186.135 18.625 186.570 ;
        RECT 18.800 186.135 24.145 186.570 ;
        RECT 24.320 186.135 29.665 186.570 ;
        RECT 29.840 186.135 35.185 186.570 ;
        RECT 35.355 186.135 35.645 187.300 ;
        RECT 35.815 187.225 37.025 187.745 ;
        RECT 37.195 187.395 38.405 187.915 ;
        RECT 38.615 187.865 38.845 188.685 ;
        RECT 39.015 187.885 39.345 188.515 ;
        RECT 38.595 187.445 38.925 187.695 ;
        RECT 39.095 187.285 39.345 187.885 ;
        RECT 39.515 187.865 39.725 188.685 ;
        RECT 39.960 187.975 40.215 188.505 ;
        RECT 40.385 188.225 40.690 188.685 ;
        RECT 40.935 188.305 42.005 188.475 ;
        RECT 35.815 186.135 38.405 187.225 ;
        RECT 38.615 186.135 38.845 187.275 ;
        RECT 39.015 186.305 39.345 187.285 ;
        RECT 39.960 187.325 40.170 187.975 ;
        RECT 40.935 187.950 41.255 188.305 ;
        RECT 40.930 187.775 41.255 187.950 ;
        RECT 40.340 187.475 41.255 187.775 ;
        RECT 41.425 187.735 41.665 188.135 ;
        RECT 41.835 188.075 42.005 188.305 ;
        RECT 42.175 188.245 42.365 188.685 ;
        RECT 42.535 188.235 43.485 188.515 ;
        RECT 43.705 188.325 44.055 188.495 ;
        RECT 41.835 187.905 42.365 188.075 ;
        RECT 40.340 187.445 41.080 187.475 ;
        RECT 39.515 186.135 39.725 187.275 ;
        RECT 39.960 186.445 40.215 187.325 ;
        RECT 40.385 186.135 40.690 187.275 ;
        RECT 40.910 186.855 41.080 187.445 ;
        RECT 41.425 187.365 41.965 187.735 ;
        RECT 42.145 187.625 42.365 187.905 ;
        RECT 42.535 187.455 42.705 188.235 ;
        RECT 42.300 187.285 42.705 187.455 ;
        RECT 42.875 187.445 43.225 188.065 ;
        RECT 42.300 187.195 42.470 187.285 ;
        RECT 43.395 187.275 43.605 188.065 ;
        RECT 41.250 187.025 42.470 187.195 ;
        RECT 42.930 187.115 43.605 187.275 ;
        RECT 40.910 186.685 41.710 186.855 ;
        RECT 41.030 186.135 41.360 186.515 ;
        RECT 41.540 186.395 41.710 186.685 ;
        RECT 42.300 186.645 42.470 187.025 ;
        RECT 42.640 187.105 43.605 187.115 ;
        RECT 43.795 187.935 44.055 188.325 ;
        RECT 44.265 188.225 44.595 188.685 ;
        RECT 45.470 188.295 46.325 188.465 ;
        RECT 46.530 188.295 47.025 188.465 ;
        RECT 47.195 188.325 47.525 188.685 ;
        RECT 43.795 187.245 43.965 187.935 ;
        RECT 44.135 187.585 44.305 187.765 ;
        RECT 44.475 187.755 45.265 188.005 ;
        RECT 45.470 187.585 45.640 188.295 ;
        RECT 45.810 187.785 46.165 188.005 ;
        RECT 44.135 187.415 45.825 187.585 ;
        RECT 42.640 186.815 43.100 187.105 ;
        RECT 43.795 187.075 45.295 187.245 ;
        RECT 43.795 186.935 43.965 187.075 ;
        RECT 43.405 186.765 43.965 186.935 ;
        RECT 41.880 186.135 42.130 186.595 ;
        RECT 42.300 186.305 43.170 186.645 ;
        RECT 43.405 186.305 43.575 186.765 ;
        RECT 44.410 186.735 45.485 186.905 ;
        RECT 43.745 186.135 44.115 186.595 ;
        RECT 44.410 186.395 44.580 186.735 ;
        RECT 44.750 186.135 45.080 186.565 ;
        RECT 45.315 186.395 45.485 186.735 ;
        RECT 45.655 186.635 45.825 187.415 ;
        RECT 45.995 187.195 46.165 187.785 ;
        RECT 46.335 187.385 46.685 188.005 ;
        RECT 45.995 186.805 46.460 187.195 ;
        RECT 46.855 186.935 47.025 188.295 ;
        RECT 47.195 187.105 47.655 188.155 ;
        RECT 46.630 186.765 47.025 186.935 ;
        RECT 46.630 186.635 46.800 186.765 ;
        RECT 45.655 186.305 46.335 186.635 ;
        RECT 46.550 186.305 46.800 186.635 ;
        RECT 46.970 186.135 47.220 186.595 ;
        RECT 47.390 186.320 47.715 187.105 ;
        RECT 47.885 186.305 48.055 188.425 ;
        RECT 48.225 188.305 48.555 188.685 ;
        RECT 48.725 188.135 48.980 188.425 ;
        RECT 48.230 187.965 48.980 188.135 ;
        RECT 48.230 186.975 48.460 187.965 ;
        RECT 49.155 187.935 50.365 188.685 ;
        RECT 48.630 187.145 48.980 187.795 ;
        RECT 49.155 187.225 49.675 187.765 ;
        RECT 49.845 187.395 50.365 187.935 ;
        RECT 50.575 187.865 50.805 188.685 ;
        RECT 50.975 187.885 51.305 188.515 ;
        RECT 50.555 187.445 50.885 187.695 ;
        RECT 51.055 187.285 51.305 187.885 ;
        RECT 51.475 187.865 51.685 188.685 ;
        RECT 52.465 188.135 52.635 188.515 ;
        RECT 52.815 188.305 53.145 188.685 ;
        RECT 52.465 187.965 53.130 188.135 ;
        RECT 53.325 188.010 53.585 188.515 ;
        RECT 52.395 187.415 52.725 187.785 ;
        RECT 52.960 187.710 53.130 187.965 ;
        RECT 48.230 186.805 48.980 186.975 ;
        RECT 48.225 186.135 48.555 186.635 ;
        RECT 48.725 186.305 48.980 186.805 ;
        RECT 49.155 186.135 50.365 187.225 ;
        RECT 50.575 186.135 50.805 187.275 ;
        RECT 50.975 186.305 51.305 187.285 ;
        RECT 52.960 187.380 53.245 187.710 ;
        RECT 51.475 186.135 51.685 187.275 ;
        RECT 52.960 187.235 53.130 187.380 ;
        RECT 52.465 187.065 53.130 187.235 ;
        RECT 53.415 187.210 53.585 188.010 ;
        RECT 53.815 187.865 54.025 188.685 ;
        RECT 54.195 187.885 54.525 188.515 ;
        RECT 54.195 187.285 54.445 187.885 ;
        RECT 54.695 187.865 54.925 188.685 ;
        RECT 55.600 188.140 60.945 188.685 ;
        RECT 54.615 187.445 54.945 187.695 ;
        RECT 52.465 186.305 52.635 187.065 ;
        RECT 52.815 186.135 53.145 186.895 ;
        RECT 53.315 186.305 53.585 187.210 ;
        RECT 53.815 186.135 54.025 187.275 ;
        RECT 54.195 186.305 54.525 187.285 ;
        RECT 54.695 186.135 54.925 187.275 ;
        RECT 57.190 186.570 57.540 187.820 ;
        RECT 59.020 187.310 59.360 188.140 ;
        RECT 61.115 187.960 61.405 188.685 ;
        RECT 61.575 187.915 65.085 188.685 ;
        RECT 55.600 186.135 60.945 186.570 ;
        RECT 61.115 186.135 61.405 187.300 ;
        RECT 61.575 187.225 63.265 187.745 ;
        RECT 63.435 187.395 65.085 187.915 ;
        RECT 65.255 188.010 65.515 188.515 ;
        RECT 65.695 188.305 66.025 188.685 ;
        RECT 66.205 188.135 66.375 188.515 ;
        RECT 61.575 186.135 65.085 187.225 ;
        RECT 65.255 187.210 65.425 188.010 ;
        RECT 65.710 187.965 66.375 188.135 ;
        RECT 66.635 188.035 66.895 188.515 ;
        RECT 67.065 188.145 67.315 188.685 ;
        RECT 65.710 187.710 65.880 187.965 ;
        RECT 65.595 187.380 65.880 187.710 ;
        RECT 66.115 187.415 66.445 187.785 ;
        RECT 65.710 187.235 65.880 187.380 ;
        RECT 65.255 186.305 65.525 187.210 ;
        RECT 65.710 187.065 66.375 187.235 ;
        RECT 65.695 186.135 66.025 186.895 ;
        RECT 66.205 186.305 66.375 187.065 ;
        RECT 66.635 187.005 66.805 188.035 ;
        RECT 67.485 187.980 67.705 188.465 ;
        RECT 66.975 187.385 67.205 187.780 ;
        RECT 67.375 187.555 67.705 187.980 ;
        RECT 67.875 188.305 68.765 188.475 ;
        RECT 67.875 187.580 68.045 188.305 ;
        RECT 68.215 187.750 68.765 188.135 ;
        RECT 68.935 187.865 69.195 188.685 ;
        RECT 69.365 187.865 69.695 188.285 ;
        RECT 69.875 188.115 70.135 188.515 ;
        RECT 70.305 188.285 70.635 188.685 ;
        RECT 70.805 188.115 70.975 188.465 ;
        RECT 71.145 188.285 71.520 188.685 ;
        RECT 69.875 187.945 71.540 188.115 ;
        RECT 71.710 188.010 71.985 188.355 ;
        RECT 73.075 188.305 73.965 188.475 ;
        RECT 69.445 187.775 69.695 187.865 ;
        RECT 71.370 187.775 71.540 187.945 ;
        RECT 67.875 187.510 68.765 187.580 ;
        RECT 67.870 187.485 68.765 187.510 ;
        RECT 67.860 187.470 68.765 187.485 ;
        RECT 67.855 187.455 68.765 187.470 ;
        RECT 67.845 187.450 68.765 187.455 ;
        RECT 67.840 187.440 68.765 187.450 ;
        RECT 68.940 187.445 69.275 187.695 ;
        RECT 69.445 187.445 70.160 187.775 ;
        RECT 70.375 187.445 71.200 187.775 ;
        RECT 71.370 187.445 71.645 187.775 ;
        RECT 67.835 187.430 68.765 187.440 ;
        RECT 67.825 187.425 68.765 187.430 ;
        RECT 67.815 187.415 68.765 187.425 ;
        RECT 67.805 187.410 68.765 187.415 ;
        RECT 67.805 187.405 68.140 187.410 ;
        RECT 67.790 187.400 68.140 187.405 ;
        RECT 67.775 187.390 68.140 187.400 ;
        RECT 67.750 187.385 68.140 187.390 ;
        RECT 66.975 187.380 68.140 187.385 ;
        RECT 66.975 187.345 68.110 187.380 ;
        RECT 66.975 187.320 68.075 187.345 ;
        RECT 66.975 187.290 68.045 187.320 ;
        RECT 66.975 187.260 68.025 187.290 ;
        RECT 66.975 187.230 68.005 187.260 ;
        RECT 66.975 187.220 67.935 187.230 ;
        RECT 66.975 187.210 67.910 187.220 ;
        RECT 66.975 187.195 67.890 187.210 ;
        RECT 66.975 187.180 67.870 187.195 ;
        RECT 67.080 187.170 67.865 187.180 ;
        RECT 67.080 187.135 67.850 187.170 ;
        RECT 66.635 186.305 66.910 187.005 ;
        RECT 67.080 186.885 67.835 187.135 ;
        RECT 68.005 186.815 68.335 187.060 ;
        RECT 68.505 186.960 68.765 187.410 ;
        RECT 68.150 186.790 68.335 186.815 ;
        RECT 68.150 186.690 68.765 186.790 ;
        RECT 67.080 186.135 67.335 186.680 ;
        RECT 67.505 186.305 67.985 186.645 ;
        RECT 68.160 186.135 68.765 186.690 ;
        RECT 68.935 186.135 69.195 187.275 ;
        RECT 69.445 186.885 69.615 187.445 ;
        RECT 69.875 186.985 70.205 187.275 ;
        RECT 70.375 187.155 70.620 187.445 ;
        RECT 71.370 187.275 71.540 187.445 ;
        RECT 71.815 187.275 71.985 188.010 ;
        RECT 73.075 187.750 73.625 188.135 ;
        RECT 73.795 187.580 73.965 188.305 ;
        RECT 70.880 187.105 71.540 187.275 ;
        RECT 70.880 186.985 71.050 187.105 ;
        RECT 69.875 186.815 71.050 186.985 ;
        RECT 69.435 186.315 71.050 186.645 ;
        RECT 71.220 186.135 71.500 186.935 ;
        RECT 71.710 186.305 71.985 187.275 ;
        RECT 73.075 187.510 73.965 187.580 ;
        RECT 74.135 187.980 74.355 188.465 ;
        RECT 74.525 188.145 74.775 188.685 ;
        RECT 74.945 188.035 75.205 188.515 ;
        RECT 74.135 187.555 74.465 187.980 ;
        RECT 73.075 187.485 73.970 187.510 ;
        RECT 73.075 187.470 73.980 187.485 ;
        RECT 73.075 187.455 73.985 187.470 ;
        RECT 73.075 187.450 73.995 187.455 ;
        RECT 73.075 187.440 74.000 187.450 ;
        RECT 73.075 187.430 74.005 187.440 ;
        RECT 73.075 187.425 74.015 187.430 ;
        RECT 73.075 187.415 74.025 187.425 ;
        RECT 73.075 187.410 74.035 187.415 ;
        RECT 73.075 186.960 73.335 187.410 ;
        RECT 73.700 187.405 74.035 187.410 ;
        RECT 73.700 187.400 74.050 187.405 ;
        RECT 73.700 187.390 74.065 187.400 ;
        RECT 73.700 187.385 74.090 187.390 ;
        RECT 74.635 187.385 74.865 187.780 ;
        RECT 73.700 187.380 74.865 187.385 ;
        RECT 73.730 187.345 74.865 187.380 ;
        RECT 73.765 187.320 74.865 187.345 ;
        RECT 73.795 187.290 74.865 187.320 ;
        RECT 73.815 187.260 74.865 187.290 ;
        RECT 73.835 187.230 74.865 187.260 ;
        RECT 73.905 187.220 74.865 187.230 ;
        RECT 73.930 187.210 74.865 187.220 ;
        RECT 73.950 187.195 74.865 187.210 ;
        RECT 73.970 187.180 74.865 187.195 ;
        RECT 73.975 187.170 74.760 187.180 ;
        RECT 73.990 187.135 74.760 187.170 ;
        RECT 73.505 186.815 73.835 187.060 ;
        RECT 74.005 186.885 74.760 187.135 ;
        RECT 75.035 187.005 75.205 188.035 ;
        RECT 75.375 187.885 76.070 188.515 ;
        RECT 76.275 187.885 76.585 188.685 ;
        RECT 77.675 187.915 81.185 188.685 ;
        RECT 81.360 188.140 86.705 188.685 ;
        RECT 75.895 187.835 76.070 187.885 ;
        RECT 75.395 187.445 75.730 187.695 ;
        RECT 75.900 187.285 76.070 187.835 ;
        RECT 76.240 187.445 76.575 187.715 ;
        RECT 73.505 186.790 73.690 186.815 ;
        RECT 73.075 186.690 73.690 186.790 ;
        RECT 73.075 186.135 73.680 186.690 ;
        RECT 73.855 186.305 74.335 186.645 ;
        RECT 74.505 186.135 74.760 186.680 ;
        RECT 74.930 186.305 75.205 187.005 ;
        RECT 75.375 186.135 75.635 187.275 ;
        RECT 75.805 186.305 76.135 187.285 ;
        RECT 76.305 186.135 76.585 187.275 ;
        RECT 77.675 187.225 79.365 187.745 ;
        RECT 79.535 187.395 81.185 187.915 ;
        RECT 77.675 186.135 81.185 187.225 ;
        RECT 82.950 186.570 83.300 187.820 ;
        RECT 84.780 187.310 85.120 188.140 ;
        RECT 86.875 187.960 87.165 188.685 ;
        RECT 87.340 187.975 87.595 188.505 ;
        RECT 87.765 188.225 88.070 188.685 ;
        RECT 88.315 188.305 89.385 188.475 ;
        RECT 87.340 187.325 87.550 187.975 ;
        RECT 88.315 187.950 88.635 188.305 ;
        RECT 88.310 187.775 88.635 187.950 ;
        RECT 87.720 187.475 88.635 187.775 ;
        RECT 88.805 187.735 89.045 188.135 ;
        RECT 89.215 188.075 89.385 188.305 ;
        RECT 89.555 188.245 89.745 188.685 ;
        RECT 89.915 188.235 90.865 188.515 ;
        RECT 91.085 188.325 91.435 188.495 ;
        RECT 89.215 187.905 89.745 188.075 ;
        RECT 87.720 187.445 88.460 187.475 ;
        RECT 81.360 186.135 86.705 186.570 ;
        RECT 86.875 186.135 87.165 187.300 ;
        RECT 87.340 186.445 87.595 187.325 ;
        RECT 87.765 186.135 88.070 187.275 ;
        RECT 88.290 186.855 88.460 187.445 ;
        RECT 88.805 187.365 89.345 187.735 ;
        RECT 89.525 187.625 89.745 187.905 ;
        RECT 89.915 187.455 90.085 188.235 ;
        RECT 89.680 187.285 90.085 187.455 ;
        RECT 90.255 187.445 90.605 188.065 ;
        RECT 89.680 187.195 89.850 187.285 ;
        RECT 90.775 187.275 90.985 188.065 ;
        RECT 88.630 187.025 89.850 187.195 ;
        RECT 90.310 187.115 90.985 187.275 ;
        RECT 88.290 186.685 89.090 186.855 ;
        RECT 88.410 186.135 88.740 186.515 ;
        RECT 88.920 186.395 89.090 186.685 ;
        RECT 89.680 186.645 89.850 187.025 ;
        RECT 90.020 187.105 90.985 187.115 ;
        RECT 91.175 187.935 91.435 188.325 ;
        RECT 91.645 188.225 91.975 188.685 ;
        RECT 92.850 188.295 93.705 188.465 ;
        RECT 93.910 188.295 94.405 188.465 ;
        RECT 94.575 188.325 94.905 188.685 ;
        RECT 91.175 187.245 91.345 187.935 ;
        RECT 91.515 187.585 91.685 187.765 ;
        RECT 91.855 187.755 92.645 188.005 ;
        RECT 92.850 187.585 93.020 188.295 ;
        RECT 93.190 187.785 93.545 188.005 ;
        RECT 91.515 187.415 93.205 187.585 ;
        RECT 90.020 186.815 90.480 187.105 ;
        RECT 91.175 187.075 92.675 187.245 ;
        RECT 91.175 186.935 91.345 187.075 ;
        RECT 90.785 186.765 91.345 186.935 ;
        RECT 89.260 186.135 89.510 186.595 ;
        RECT 89.680 186.305 90.550 186.645 ;
        RECT 90.785 186.305 90.955 186.765 ;
        RECT 91.790 186.735 92.865 186.905 ;
        RECT 91.125 186.135 91.495 186.595 ;
        RECT 91.790 186.395 91.960 186.735 ;
        RECT 92.130 186.135 92.460 186.565 ;
        RECT 92.695 186.395 92.865 186.735 ;
        RECT 93.035 186.635 93.205 187.415 ;
        RECT 93.375 187.195 93.545 187.785 ;
        RECT 93.715 187.385 94.065 188.005 ;
        RECT 93.375 186.805 93.840 187.195 ;
        RECT 94.235 186.935 94.405 188.295 ;
        RECT 94.575 187.105 95.035 188.155 ;
        RECT 94.010 186.765 94.405 186.935 ;
        RECT 94.010 186.635 94.180 186.765 ;
        RECT 93.035 186.305 93.715 186.635 ;
        RECT 93.930 186.305 94.180 186.635 ;
        RECT 94.350 186.135 94.600 186.595 ;
        RECT 94.770 186.320 95.095 187.105 ;
        RECT 95.265 186.305 95.435 188.425 ;
        RECT 95.605 188.305 95.935 188.685 ;
        RECT 96.105 188.135 96.360 188.425 ;
        RECT 95.610 187.965 96.360 188.135 ;
        RECT 95.610 186.975 95.840 187.965 ;
        RECT 96.535 187.915 98.205 188.685 ;
        RECT 96.010 187.145 96.360 187.795 ;
        RECT 96.535 187.225 97.285 187.745 ;
        RECT 97.455 187.395 98.205 187.915 ;
        RECT 98.650 187.875 98.895 188.480 ;
        RECT 99.115 188.150 99.625 188.685 ;
        RECT 98.375 187.705 99.605 187.875 ;
        RECT 95.610 186.805 96.360 186.975 ;
        RECT 95.605 186.135 95.935 186.635 ;
        RECT 96.105 186.305 96.360 186.805 ;
        RECT 96.535 186.135 98.205 187.225 ;
        RECT 98.375 186.895 98.715 187.705 ;
        RECT 98.885 187.140 99.635 187.330 ;
        RECT 98.375 186.485 98.890 186.895 ;
        RECT 99.125 186.135 99.295 186.895 ;
        RECT 99.465 186.475 99.635 187.140 ;
        RECT 99.805 187.155 99.995 188.515 ;
        RECT 100.165 188.005 100.440 188.515 ;
        RECT 100.630 188.150 101.160 188.515 ;
        RECT 101.585 188.285 101.915 188.685 ;
        RECT 100.985 188.115 101.160 188.150 ;
        RECT 100.165 187.835 100.445 188.005 ;
        RECT 100.165 187.355 100.440 187.835 ;
        RECT 100.645 187.155 100.815 187.955 ;
        RECT 99.805 186.985 100.815 187.155 ;
        RECT 100.985 187.945 101.915 188.115 ;
        RECT 102.085 187.945 102.340 188.515 ;
        RECT 100.985 186.815 101.155 187.945 ;
        RECT 101.745 187.775 101.915 187.945 ;
        RECT 100.030 186.645 101.155 186.815 ;
        RECT 101.325 187.445 101.520 187.775 ;
        RECT 101.745 187.445 102.000 187.775 ;
        RECT 101.325 186.475 101.495 187.445 ;
        RECT 102.170 187.275 102.340 187.945 ;
        RECT 102.790 187.875 103.035 188.480 ;
        RECT 103.255 188.150 103.765 188.685 ;
        RECT 99.465 186.305 101.495 186.475 ;
        RECT 101.665 186.135 101.835 187.275 ;
        RECT 102.005 186.305 102.340 187.275 ;
        RECT 102.515 187.705 103.745 187.875 ;
        RECT 102.515 186.895 102.855 187.705 ;
        RECT 103.025 187.140 103.775 187.330 ;
        RECT 102.515 186.485 103.030 186.895 ;
        RECT 103.265 186.135 103.435 186.895 ;
        RECT 103.605 186.475 103.775 187.140 ;
        RECT 103.945 187.155 104.135 188.515 ;
        RECT 104.305 188.005 104.580 188.515 ;
        RECT 104.770 188.150 105.300 188.515 ;
        RECT 105.725 188.285 106.055 188.685 ;
        RECT 105.125 188.115 105.300 188.150 ;
        RECT 104.305 187.835 104.585 188.005 ;
        RECT 104.305 187.355 104.580 187.835 ;
        RECT 104.785 187.155 104.955 187.955 ;
        RECT 103.945 186.985 104.955 187.155 ;
        RECT 105.125 187.945 106.055 188.115 ;
        RECT 106.225 187.945 106.480 188.515 ;
        RECT 105.125 186.815 105.295 187.945 ;
        RECT 105.885 187.775 106.055 187.945 ;
        RECT 104.170 186.645 105.295 186.815 ;
        RECT 105.465 187.445 105.660 187.775 ;
        RECT 105.885 187.445 106.140 187.775 ;
        RECT 105.465 186.475 105.635 187.445 ;
        RECT 106.310 187.275 106.480 187.945 ;
        RECT 107.115 187.915 109.705 188.685 ;
        RECT 109.965 188.135 110.135 188.515 ;
        RECT 110.315 188.305 110.645 188.685 ;
        RECT 109.965 187.965 110.630 188.135 ;
        RECT 110.825 188.010 111.085 188.515 ;
        RECT 103.605 186.305 105.635 186.475 ;
        RECT 105.805 186.135 105.975 187.275 ;
        RECT 106.145 186.305 106.480 187.275 ;
        RECT 107.115 187.225 108.325 187.745 ;
        RECT 108.495 187.395 109.705 187.915 ;
        RECT 109.895 187.415 110.225 187.785 ;
        RECT 110.460 187.710 110.630 187.965 ;
        RECT 110.460 187.380 110.745 187.710 ;
        RECT 110.460 187.235 110.630 187.380 ;
        RECT 107.115 186.135 109.705 187.225 ;
        RECT 109.965 187.065 110.630 187.235 ;
        RECT 110.915 187.210 111.085 188.010 ;
        RECT 111.255 187.935 112.465 188.685 ;
        RECT 112.635 187.960 112.925 188.685 ;
        RECT 113.560 188.140 118.905 188.685 ;
        RECT 119.080 188.140 124.425 188.685 ;
        RECT 109.965 186.305 110.135 187.065 ;
        RECT 110.315 186.135 110.645 186.895 ;
        RECT 110.815 186.305 111.085 187.210 ;
        RECT 111.255 187.225 111.775 187.765 ;
        RECT 111.945 187.395 112.465 187.935 ;
        RECT 111.255 186.135 112.465 187.225 ;
        RECT 112.635 186.135 112.925 187.300 ;
        RECT 115.150 186.570 115.500 187.820 ;
        RECT 116.980 187.310 117.320 188.140 ;
        RECT 120.670 186.570 121.020 187.820 ;
        RECT 122.500 187.310 122.840 188.140 ;
        RECT 124.595 187.935 125.805 188.685 ;
        RECT 124.595 187.225 125.115 187.765 ;
        RECT 125.285 187.395 125.805 187.935 ;
        RECT 113.560 186.135 118.905 186.570 ;
        RECT 119.080 186.135 124.425 186.570 ;
        RECT 124.595 186.135 125.805 187.225 ;
        RECT 11.810 185.965 125.890 186.135 ;
        RECT 11.895 184.875 13.105 185.965 ;
        RECT 11.895 184.165 12.415 184.705 ;
        RECT 12.585 184.335 13.105 184.875 ;
        RECT 13.275 184.875 16.785 185.965 ;
        RECT 16.960 185.530 22.305 185.965 ;
        RECT 13.275 184.355 14.965 184.875 ;
        RECT 15.135 184.185 16.785 184.705 ;
        RECT 18.550 184.280 18.900 185.530 ;
        RECT 22.475 184.800 22.765 185.965 ;
        RECT 23.395 184.875 26.905 185.965 ;
        RECT 27.080 185.530 32.425 185.965 ;
        RECT 11.895 183.415 13.105 184.165 ;
        RECT 13.275 183.415 16.785 184.185 ;
        RECT 20.380 183.960 20.720 184.790 ;
        RECT 23.395 184.355 25.085 184.875 ;
        RECT 25.255 184.185 26.905 184.705 ;
        RECT 28.670 184.280 29.020 185.530 ;
        RECT 32.635 184.825 32.865 185.965 ;
        RECT 33.035 184.815 33.365 185.795 ;
        RECT 33.535 184.825 33.745 185.965 ;
        RECT 33.980 185.295 34.235 185.795 ;
        RECT 34.405 185.465 34.735 185.965 ;
        RECT 33.980 185.125 34.730 185.295 ;
        RECT 16.960 183.415 22.305 183.960 ;
        RECT 22.475 183.415 22.765 184.140 ;
        RECT 23.395 183.415 26.905 184.185 ;
        RECT 30.500 183.960 30.840 184.790 ;
        RECT 32.615 184.405 32.945 184.655 ;
        RECT 27.080 183.415 32.425 183.960 ;
        RECT 32.635 183.415 32.865 184.235 ;
        RECT 33.115 184.215 33.365 184.815 ;
        RECT 33.980 184.305 34.330 184.955 ;
        RECT 33.035 183.585 33.365 184.215 ;
        RECT 33.535 183.415 33.745 184.235 ;
        RECT 34.500 184.135 34.730 185.125 ;
        RECT 33.980 183.965 34.730 184.135 ;
        RECT 33.980 183.675 34.235 183.965 ;
        RECT 34.405 183.415 34.735 183.795 ;
        RECT 34.905 183.675 35.075 185.795 ;
        RECT 35.245 184.995 35.570 185.780 ;
        RECT 35.740 185.505 35.990 185.965 ;
        RECT 36.160 185.465 36.410 185.795 ;
        RECT 36.625 185.465 37.305 185.795 ;
        RECT 36.160 185.335 36.330 185.465 ;
        RECT 35.935 185.165 36.330 185.335 ;
        RECT 35.305 183.945 35.765 184.995 ;
        RECT 35.935 183.805 36.105 185.165 ;
        RECT 36.500 184.905 36.965 185.295 ;
        RECT 36.275 184.095 36.625 184.715 ;
        RECT 36.795 184.315 36.965 184.905 ;
        RECT 37.135 184.685 37.305 185.465 ;
        RECT 37.475 185.365 37.645 185.705 ;
        RECT 37.880 185.535 38.210 185.965 ;
        RECT 38.380 185.365 38.550 185.705 ;
        RECT 38.845 185.505 39.215 185.965 ;
        RECT 37.475 185.195 38.550 185.365 ;
        RECT 39.385 185.335 39.555 185.795 ;
        RECT 39.790 185.455 40.660 185.795 ;
        RECT 40.830 185.505 41.080 185.965 ;
        RECT 38.995 185.165 39.555 185.335 ;
        RECT 38.995 185.025 39.165 185.165 ;
        RECT 37.665 184.855 39.165 185.025 ;
        RECT 39.860 184.995 40.320 185.285 ;
        RECT 37.135 184.515 38.825 184.685 ;
        RECT 36.795 184.095 37.150 184.315 ;
        RECT 37.320 183.805 37.490 184.515 ;
        RECT 37.695 184.095 38.485 184.345 ;
        RECT 38.655 184.335 38.825 184.515 ;
        RECT 38.995 184.165 39.165 184.855 ;
        RECT 35.435 183.415 35.765 183.775 ;
        RECT 35.935 183.635 36.430 183.805 ;
        RECT 36.635 183.635 37.490 183.805 ;
        RECT 38.365 183.415 38.695 183.875 ;
        RECT 38.905 183.775 39.165 184.165 ;
        RECT 39.355 184.985 40.320 184.995 ;
        RECT 40.490 185.075 40.660 185.455 ;
        RECT 41.250 185.415 41.420 185.705 ;
        RECT 41.600 185.585 41.930 185.965 ;
        RECT 41.250 185.245 42.050 185.415 ;
        RECT 39.355 184.825 40.030 184.985 ;
        RECT 40.490 184.905 41.710 185.075 ;
        RECT 39.355 184.035 39.565 184.825 ;
        RECT 40.490 184.815 40.660 184.905 ;
        RECT 39.735 184.035 40.085 184.655 ;
        RECT 40.255 184.645 40.660 184.815 ;
        RECT 40.255 183.865 40.425 184.645 ;
        RECT 40.595 184.195 40.815 184.475 ;
        RECT 40.995 184.365 41.535 184.735 ;
        RECT 41.880 184.655 42.050 185.245 ;
        RECT 42.270 184.825 42.575 185.965 ;
        RECT 42.745 184.775 43.000 185.655 ;
        RECT 41.880 184.625 42.620 184.655 ;
        RECT 40.595 184.025 41.125 184.195 ;
        RECT 38.905 183.605 39.255 183.775 ;
        RECT 39.475 183.585 40.425 183.865 ;
        RECT 40.595 183.415 40.785 183.855 ;
        RECT 40.955 183.795 41.125 184.025 ;
        RECT 41.295 183.965 41.535 184.365 ;
        RECT 41.705 184.325 42.620 184.625 ;
        RECT 41.705 184.150 42.030 184.325 ;
        RECT 41.705 183.795 42.025 184.150 ;
        RECT 42.790 184.125 43.000 184.775 ;
        RECT 40.955 183.625 42.025 183.795 ;
        RECT 42.270 183.415 42.575 183.875 ;
        RECT 42.745 183.595 43.000 184.125 ;
        RECT 44.100 184.825 44.435 185.795 ;
        RECT 44.605 184.825 44.775 185.965 ;
        RECT 44.945 185.625 46.975 185.795 ;
        RECT 44.100 184.155 44.270 184.825 ;
        RECT 44.945 184.655 45.115 185.625 ;
        RECT 44.440 184.325 44.695 184.655 ;
        RECT 44.920 184.325 45.115 184.655 ;
        RECT 45.285 185.285 46.410 185.455 ;
        RECT 44.525 184.155 44.695 184.325 ;
        RECT 45.285 184.155 45.455 185.285 ;
        RECT 44.100 183.585 44.355 184.155 ;
        RECT 44.525 183.985 45.455 184.155 ;
        RECT 45.625 184.945 46.635 185.115 ;
        RECT 45.625 184.145 45.795 184.945 ;
        RECT 46.000 184.265 46.275 184.745 ;
        RECT 45.995 184.095 46.275 184.265 ;
        RECT 45.280 183.950 45.455 183.985 ;
        RECT 44.525 183.415 44.855 183.815 ;
        RECT 45.280 183.585 45.810 183.950 ;
        RECT 46.000 183.585 46.275 184.095 ;
        RECT 46.445 183.585 46.635 184.945 ;
        RECT 46.805 184.960 46.975 185.625 ;
        RECT 47.145 185.205 47.315 185.965 ;
        RECT 47.550 185.205 48.065 185.615 ;
        RECT 46.805 184.770 47.555 184.960 ;
        RECT 47.725 184.395 48.065 185.205 ;
        RECT 48.235 184.800 48.525 185.965 ;
        RECT 46.835 184.225 48.065 184.395 ;
        RECT 48.700 184.775 48.955 185.655 ;
        RECT 49.125 184.825 49.430 185.965 ;
        RECT 49.770 185.585 50.100 185.965 ;
        RECT 50.280 185.415 50.450 185.705 ;
        RECT 50.620 185.505 50.870 185.965 ;
        RECT 49.650 185.245 50.450 185.415 ;
        RECT 51.040 185.455 51.910 185.795 ;
        RECT 46.815 183.415 47.325 183.950 ;
        RECT 47.545 183.620 47.790 184.225 ;
        RECT 48.235 183.415 48.525 184.140 ;
        RECT 48.700 184.125 48.910 184.775 ;
        RECT 49.650 184.655 49.820 185.245 ;
        RECT 51.040 185.075 51.210 185.455 ;
        RECT 52.145 185.335 52.315 185.795 ;
        RECT 52.485 185.505 52.855 185.965 ;
        RECT 53.150 185.365 53.320 185.705 ;
        RECT 53.490 185.535 53.820 185.965 ;
        RECT 54.055 185.365 54.225 185.705 ;
        RECT 49.990 184.905 51.210 185.075 ;
        RECT 51.380 184.995 51.840 185.285 ;
        RECT 52.145 185.165 52.705 185.335 ;
        RECT 53.150 185.195 54.225 185.365 ;
        RECT 54.395 185.465 55.075 185.795 ;
        RECT 55.290 185.465 55.540 185.795 ;
        RECT 55.710 185.505 55.960 185.965 ;
        RECT 52.535 185.025 52.705 185.165 ;
        RECT 51.380 184.985 52.345 184.995 ;
        RECT 51.040 184.815 51.210 184.905 ;
        RECT 51.670 184.825 52.345 184.985 ;
        RECT 49.080 184.625 49.820 184.655 ;
        RECT 49.080 184.325 49.995 184.625 ;
        RECT 49.670 184.150 49.995 184.325 ;
        RECT 48.700 183.595 48.955 184.125 ;
        RECT 49.125 183.415 49.430 183.875 ;
        RECT 49.675 183.795 49.995 184.150 ;
        RECT 50.165 184.365 50.705 184.735 ;
        RECT 51.040 184.645 51.445 184.815 ;
        RECT 50.165 183.965 50.405 184.365 ;
        RECT 50.885 184.195 51.105 184.475 ;
        RECT 50.575 184.025 51.105 184.195 ;
        RECT 50.575 183.795 50.745 184.025 ;
        RECT 51.275 183.865 51.445 184.645 ;
        RECT 51.615 184.035 51.965 184.655 ;
        RECT 52.135 184.035 52.345 184.825 ;
        RECT 52.535 184.855 54.035 185.025 ;
        RECT 52.535 184.165 52.705 184.855 ;
        RECT 54.395 184.685 54.565 185.465 ;
        RECT 55.370 185.335 55.540 185.465 ;
        RECT 52.875 184.515 54.565 184.685 ;
        RECT 54.735 184.905 55.200 185.295 ;
        RECT 55.370 185.165 55.765 185.335 ;
        RECT 52.875 184.335 53.045 184.515 ;
        RECT 49.675 183.625 50.745 183.795 ;
        RECT 50.915 183.415 51.105 183.855 ;
        RECT 51.275 183.585 52.225 183.865 ;
        RECT 52.535 183.775 52.795 184.165 ;
        RECT 53.215 184.095 54.005 184.345 ;
        RECT 52.445 183.605 52.795 183.775 ;
        RECT 53.005 183.415 53.335 183.875 ;
        RECT 54.210 183.805 54.380 184.515 ;
        RECT 54.735 184.315 54.905 184.905 ;
        RECT 54.550 184.095 54.905 184.315 ;
        RECT 55.075 184.095 55.425 184.715 ;
        RECT 55.595 183.805 55.765 185.165 ;
        RECT 56.130 184.995 56.455 185.780 ;
        RECT 55.935 183.945 56.395 184.995 ;
        RECT 54.210 183.635 55.065 183.805 ;
        RECT 55.270 183.635 55.765 183.805 ;
        RECT 55.935 183.415 56.265 183.775 ;
        RECT 56.625 183.675 56.795 185.795 ;
        RECT 56.965 185.465 57.295 185.965 ;
        RECT 57.465 185.295 57.720 185.795 ;
        RECT 56.970 185.125 57.720 185.295 ;
        RECT 56.970 184.135 57.200 185.125 ;
        RECT 57.370 184.305 57.720 184.955 ;
        RECT 58.355 184.875 61.865 185.965 ;
        RECT 58.355 184.355 60.045 184.875 ;
        RECT 62.095 184.825 62.305 185.965 ;
        RECT 62.475 184.815 62.805 185.795 ;
        RECT 62.975 184.825 63.205 185.965 ;
        RECT 63.530 185.335 63.815 185.795 ;
        RECT 63.985 185.505 64.255 185.965 ;
        RECT 63.530 185.115 64.485 185.335 ;
        RECT 60.215 184.185 61.865 184.705 ;
        RECT 56.970 183.965 57.720 184.135 ;
        RECT 56.965 183.415 57.295 183.795 ;
        RECT 57.465 183.675 57.720 183.965 ;
        RECT 58.355 183.415 61.865 184.185 ;
        RECT 62.095 183.415 62.305 184.235 ;
        RECT 62.475 184.215 62.725 184.815 ;
        RECT 62.895 184.405 63.225 184.655 ;
        RECT 63.415 184.385 64.105 184.945 ;
        RECT 62.475 183.585 62.805 184.215 ;
        RECT 62.975 183.415 63.205 184.235 ;
        RECT 64.275 184.215 64.485 185.115 ;
        RECT 63.530 184.045 64.485 184.215 ;
        RECT 64.655 184.945 65.055 185.795 ;
        RECT 65.245 185.335 65.525 185.795 ;
        RECT 66.045 185.505 66.370 185.965 ;
        RECT 65.245 185.115 66.370 185.335 ;
        RECT 64.655 184.385 65.750 184.945 ;
        RECT 65.920 184.655 66.370 185.115 ;
        RECT 66.540 184.825 66.925 185.795 ;
        RECT 68.015 184.825 68.275 185.965 ;
        RECT 68.515 185.455 70.130 185.785 ;
        RECT 63.530 183.585 63.815 184.045 ;
        RECT 63.985 183.415 64.255 183.875 ;
        RECT 64.655 183.585 65.055 184.385 ;
        RECT 65.920 184.325 66.475 184.655 ;
        RECT 65.920 184.215 66.370 184.325 ;
        RECT 65.245 184.045 66.370 184.215 ;
        RECT 66.645 184.155 66.925 184.825 ;
        RECT 68.525 184.655 68.695 185.215 ;
        RECT 68.955 185.115 70.130 185.285 ;
        RECT 70.300 185.165 70.580 185.965 ;
        RECT 68.955 184.825 69.285 185.115 ;
        RECT 69.960 184.995 70.130 185.115 ;
        RECT 69.455 184.655 69.700 184.945 ;
        RECT 69.960 184.825 70.620 184.995 ;
        RECT 70.790 184.825 71.065 185.795 ;
        RECT 71.255 185.165 71.535 185.965 ;
        RECT 71.735 184.995 72.065 185.795 ;
        RECT 72.265 185.165 72.435 185.965 ;
        RECT 72.605 184.995 72.935 185.795 ;
        RECT 70.450 184.655 70.620 184.825 ;
        RECT 68.020 184.405 68.355 184.655 ;
        RECT 68.525 184.325 69.240 184.655 ;
        RECT 69.455 184.325 70.280 184.655 ;
        RECT 70.450 184.325 70.725 184.655 ;
        RECT 68.525 184.235 68.775 184.325 ;
        RECT 65.245 183.585 65.525 184.045 ;
        RECT 66.045 183.415 66.370 183.875 ;
        RECT 66.540 183.585 66.925 184.155 ;
        RECT 68.015 183.415 68.275 184.235 ;
        RECT 68.445 183.815 68.775 184.235 ;
        RECT 70.450 184.155 70.620 184.325 ;
        RECT 68.955 183.985 70.620 184.155 ;
        RECT 70.895 184.090 71.065 184.825 ;
        RECT 71.235 184.325 71.475 184.995 ;
        RECT 71.655 184.825 72.935 184.995 ;
        RECT 73.105 184.825 73.365 185.965 ;
        RECT 71.655 184.155 71.825 184.825 ;
        RECT 73.995 184.800 74.285 185.965 ;
        RECT 74.915 184.875 76.585 185.965 ;
        RECT 76.760 185.530 82.105 185.965 ;
        RECT 71.995 184.325 72.305 184.655 ;
        RECT 72.475 184.325 72.855 184.655 ;
        RECT 73.055 184.325 73.340 184.655 ;
        RECT 74.915 184.355 75.665 184.875 ;
        RECT 72.100 184.155 72.305 184.325 ;
        RECT 68.955 183.585 69.215 183.985 ;
        RECT 69.385 183.415 69.715 183.815 ;
        RECT 69.885 183.635 70.055 183.985 ;
        RECT 70.225 183.415 70.600 183.815 ;
        RECT 70.790 183.745 71.065 184.090 ;
        RECT 71.235 183.585 71.930 184.155 ;
        RECT 72.100 183.630 72.450 184.155 ;
        RECT 72.640 183.630 72.855 184.325 ;
        RECT 75.835 184.185 76.585 184.705 ;
        RECT 78.350 184.280 78.700 185.530 ;
        RECT 82.335 184.825 82.545 185.965 ;
        RECT 82.715 184.815 83.045 185.795 ;
        RECT 83.215 184.825 83.445 185.965 ;
        RECT 84.175 184.825 84.385 185.965 ;
        RECT 84.555 184.815 84.885 185.795 ;
        RECT 85.055 184.825 85.285 185.965 ;
        RECT 85.495 184.875 88.085 185.965 ;
        RECT 88.255 185.205 88.770 185.615 ;
        RECT 89.005 185.205 89.175 185.965 ;
        RECT 89.345 185.625 91.375 185.795 ;
        RECT 73.025 183.415 73.360 184.155 ;
        RECT 73.995 183.415 74.285 184.140 ;
        RECT 74.915 183.415 76.585 184.185 ;
        RECT 80.180 183.960 80.520 184.790 ;
        RECT 76.760 183.415 82.105 183.960 ;
        RECT 82.335 183.415 82.545 184.235 ;
        RECT 82.715 184.215 82.965 184.815 ;
        RECT 83.135 184.405 83.465 184.655 ;
        RECT 82.715 183.585 83.045 184.215 ;
        RECT 83.215 183.415 83.445 184.235 ;
        RECT 84.175 183.415 84.385 184.235 ;
        RECT 84.555 184.215 84.805 184.815 ;
        RECT 84.975 184.405 85.305 184.655 ;
        RECT 85.495 184.355 86.705 184.875 ;
        RECT 84.555 183.585 84.885 184.215 ;
        RECT 85.055 183.415 85.285 184.235 ;
        RECT 86.875 184.185 88.085 184.705 ;
        RECT 88.255 184.395 88.595 185.205 ;
        RECT 89.345 184.960 89.515 185.625 ;
        RECT 89.910 185.285 91.035 185.455 ;
        RECT 88.765 184.770 89.515 184.960 ;
        RECT 89.685 184.945 90.695 185.115 ;
        RECT 88.255 184.225 89.485 184.395 ;
        RECT 85.495 183.415 88.085 184.185 ;
        RECT 88.530 183.620 88.775 184.225 ;
        RECT 88.995 183.415 89.505 183.950 ;
        RECT 89.685 183.585 89.875 184.945 ;
        RECT 90.045 184.265 90.320 184.745 ;
        RECT 90.045 184.095 90.325 184.265 ;
        RECT 90.525 184.145 90.695 184.945 ;
        RECT 90.865 184.155 91.035 185.285 ;
        RECT 91.205 184.655 91.375 185.625 ;
        RECT 91.545 184.825 91.715 185.965 ;
        RECT 91.885 184.825 92.220 185.795 ;
        RECT 91.205 184.325 91.400 184.655 ;
        RECT 91.625 184.325 91.880 184.655 ;
        RECT 91.625 184.155 91.795 184.325 ;
        RECT 92.050 184.155 92.220 184.825 ;
        RECT 92.395 184.875 94.065 185.965 ;
        RECT 94.240 185.530 99.585 185.965 ;
        RECT 92.395 184.355 93.145 184.875 ;
        RECT 93.315 184.185 94.065 184.705 ;
        RECT 95.830 184.280 96.180 185.530 ;
        RECT 99.755 184.800 100.045 185.965 ;
        RECT 100.675 184.875 102.345 185.965 ;
        RECT 102.605 185.035 102.775 185.795 ;
        RECT 102.955 185.205 103.285 185.965 ;
        RECT 90.045 183.585 90.320 184.095 ;
        RECT 90.865 183.985 91.795 184.155 ;
        RECT 90.865 183.950 91.040 183.985 ;
        RECT 90.510 183.585 91.040 183.950 ;
        RECT 91.465 183.415 91.795 183.815 ;
        RECT 91.965 183.585 92.220 184.155 ;
        RECT 92.395 183.415 94.065 184.185 ;
        RECT 97.660 183.960 98.000 184.790 ;
        RECT 100.675 184.355 101.425 184.875 ;
        RECT 102.605 184.865 103.270 185.035 ;
        RECT 103.455 184.890 103.725 185.795 ;
        RECT 103.100 184.720 103.270 184.865 ;
        RECT 101.595 184.185 102.345 184.705 ;
        RECT 102.535 184.315 102.865 184.685 ;
        RECT 103.100 184.390 103.385 184.720 ;
        RECT 94.240 183.415 99.585 183.960 ;
        RECT 99.755 183.415 100.045 184.140 ;
        RECT 100.675 183.415 102.345 184.185 ;
        RECT 103.100 184.135 103.270 184.390 ;
        RECT 102.605 183.965 103.270 184.135 ;
        RECT 103.555 184.090 103.725 184.890 ;
        RECT 103.935 184.825 104.165 185.965 ;
        RECT 104.335 184.815 104.665 185.795 ;
        RECT 104.835 184.825 105.045 185.965 ;
        RECT 103.915 184.405 104.245 184.655 ;
        RECT 102.605 183.585 102.775 183.965 ;
        RECT 102.955 183.415 103.285 183.795 ;
        RECT 103.465 183.585 103.725 184.090 ;
        RECT 103.935 183.415 104.165 184.235 ;
        RECT 104.415 184.215 104.665 184.815 ;
        RECT 105.280 184.775 105.535 185.655 ;
        RECT 105.705 184.825 106.010 185.965 ;
        RECT 106.350 185.585 106.680 185.965 ;
        RECT 106.860 185.415 107.030 185.705 ;
        RECT 107.200 185.505 107.450 185.965 ;
        RECT 106.230 185.245 107.030 185.415 ;
        RECT 107.620 185.455 108.490 185.795 ;
        RECT 104.335 183.585 104.665 184.215 ;
        RECT 104.835 183.415 105.045 184.235 ;
        RECT 105.280 184.125 105.490 184.775 ;
        RECT 106.230 184.655 106.400 185.245 ;
        RECT 107.620 185.075 107.790 185.455 ;
        RECT 108.725 185.335 108.895 185.795 ;
        RECT 109.065 185.505 109.435 185.965 ;
        RECT 109.730 185.365 109.900 185.705 ;
        RECT 110.070 185.535 110.400 185.965 ;
        RECT 110.635 185.365 110.805 185.705 ;
        RECT 106.570 184.905 107.790 185.075 ;
        RECT 107.960 184.995 108.420 185.285 ;
        RECT 108.725 185.165 109.285 185.335 ;
        RECT 109.730 185.195 110.805 185.365 ;
        RECT 110.975 185.465 111.655 185.795 ;
        RECT 111.870 185.465 112.120 185.795 ;
        RECT 112.290 185.505 112.540 185.965 ;
        RECT 109.115 185.025 109.285 185.165 ;
        RECT 107.960 184.985 108.925 184.995 ;
        RECT 107.620 184.815 107.790 184.905 ;
        RECT 108.250 184.825 108.925 184.985 ;
        RECT 105.660 184.625 106.400 184.655 ;
        RECT 105.660 184.325 106.575 184.625 ;
        RECT 106.250 184.150 106.575 184.325 ;
        RECT 105.280 183.595 105.535 184.125 ;
        RECT 105.705 183.415 106.010 183.875 ;
        RECT 106.255 183.795 106.575 184.150 ;
        RECT 106.745 184.365 107.285 184.735 ;
        RECT 107.620 184.645 108.025 184.815 ;
        RECT 106.745 183.965 106.985 184.365 ;
        RECT 107.465 184.195 107.685 184.475 ;
        RECT 107.155 184.025 107.685 184.195 ;
        RECT 107.155 183.795 107.325 184.025 ;
        RECT 107.855 183.865 108.025 184.645 ;
        RECT 108.195 184.035 108.545 184.655 ;
        RECT 108.715 184.035 108.925 184.825 ;
        RECT 109.115 184.855 110.615 185.025 ;
        RECT 109.115 184.165 109.285 184.855 ;
        RECT 110.975 184.685 111.145 185.465 ;
        RECT 111.950 185.335 112.120 185.465 ;
        RECT 109.455 184.515 111.145 184.685 ;
        RECT 111.315 184.905 111.780 185.295 ;
        RECT 111.950 185.165 112.345 185.335 ;
        RECT 109.455 184.335 109.625 184.515 ;
        RECT 106.255 183.625 107.325 183.795 ;
        RECT 107.495 183.415 107.685 183.855 ;
        RECT 107.855 183.585 108.805 183.865 ;
        RECT 109.115 183.775 109.375 184.165 ;
        RECT 109.795 184.095 110.585 184.345 ;
        RECT 109.025 183.605 109.375 183.775 ;
        RECT 109.585 183.415 109.915 183.875 ;
        RECT 110.790 183.805 110.960 184.515 ;
        RECT 111.315 184.315 111.485 184.905 ;
        RECT 111.130 184.095 111.485 184.315 ;
        RECT 111.655 184.095 112.005 184.715 ;
        RECT 112.175 183.805 112.345 185.165 ;
        RECT 112.710 184.995 113.035 185.780 ;
        RECT 112.515 183.945 112.975 184.995 ;
        RECT 110.790 183.635 111.645 183.805 ;
        RECT 111.850 183.635 112.345 183.805 ;
        RECT 112.515 183.415 112.845 183.775 ;
        RECT 113.205 183.675 113.375 185.795 ;
        RECT 113.545 185.465 113.875 185.965 ;
        RECT 114.045 185.295 114.300 185.795 ;
        RECT 113.550 185.125 114.300 185.295 ;
        RECT 113.550 184.135 113.780 185.125 ;
        RECT 113.950 184.305 114.300 184.955 ;
        RECT 115.395 184.875 118.905 185.965 ;
        RECT 119.080 185.530 124.425 185.965 ;
        RECT 115.395 184.355 117.085 184.875 ;
        RECT 117.255 184.185 118.905 184.705 ;
        RECT 120.670 184.280 121.020 185.530 ;
        RECT 124.595 184.875 125.805 185.965 ;
        RECT 113.550 183.965 114.300 184.135 ;
        RECT 113.545 183.415 113.875 183.795 ;
        RECT 114.045 183.675 114.300 183.965 ;
        RECT 115.395 183.415 118.905 184.185 ;
        RECT 122.500 183.960 122.840 184.790 ;
        RECT 124.595 184.335 125.115 184.875 ;
        RECT 125.285 184.165 125.805 184.705 ;
        RECT 119.080 183.415 124.425 183.960 ;
        RECT 124.595 183.415 125.805 184.165 ;
        RECT 11.810 183.245 125.890 183.415 ;
        RECT 11.895 182.495 13.105 183.245 ;
        RECT 13.280 182.700 18.625 183.245 ;
        RECT 18.800 182.700 24.145 183.245 ;
        RECT 24.320 182.700 29.665 183.245 ;
        RECT 29.840 182.700 35.185 183.245 ;
        RECT 11.895 181.955 12.415 182.495 ;
        RECT 12.585 181.785 13.105 182.325 ;
        RECT 11.895 180.695 13.105 181.785 ;
        RECT 14.870 181.130 15.220 182.380 ;
        RECT 16.700 181.870 17.040 182.700 ;
        RECT 20.390 181.130 20.740 182.380 ;
        RECT 22.220 181.870 22.560 182.700 ;
        RECT 25.910 181.130 26.260 182.380 ;
        RECT 27.740 181.870 28.080 182.700 ;
        RECT 31.430 181.130 31.780 182.380 ;
        RECT 33.260 181.870 33.600 182.700 ;
        RECT 35.355 182.520 35.645 183.245 ;
        RECT 35.815 182.475 39.325 183.245 ;
        RECT 13.280 180.695 18.625 181.130 ;
        RECT 18.800 180.695 24.145 181.130 ;
        RECT 24.320 180.695 29.665 181.130 ;
        RECT 29.840 180.695 35.185 181.130 ;
        RECT 35.355 180.695 35.645 181.860 ;
        RECT 35.815 181.785 37.505 182.305 ;
        RECT 37.675 181.955 39.325 182.475 ;
        RECT 39.495 182.570 39.755 183.075 ;
        RECT 39.935 182.865 40.265 183.245 ;
        RECT 40.445 182.695 40.615 183.075 ;
        RECT 35.815 180.695 39.325 181.785 ;
        RECT 39.495 181.770 39.665 182.570 ;
        RECT 39.950 182.525 40.615 182.695 ;
        RECT 39.950 182.270 40.120 182.525 ;
        RECT 40.880 182.505 41.135 183.075 ;
        RECT 41.305 182.845 41.635 183.245 ;
        RECT 42.060 182.710 42.590 183.075 ;
        RECT 42.060 182.675 42.235 182.710 ;
        RECT 41.305 182.505 42.235 182.675 ;
        RECT 42.780 182.565 43.055 183.075 ;
        RECT 39.835 181.940 40.120 182.270 ;
        RECT 40.355 181.975 40.685 182.345 ;
        RECT 39.950 181.795 40.120 181.940 ;
        RECT 40.880 181.835 41.050 182.505 ;
        RECT 41.305 182.335 41.475 182.505 ;
        RECT 41.220 182.005 41.475 182.335 ;
        RECT 41.700 182.005 41.895 182.335 ;
        RECT 39.495 180.865 39.765 181.770 ;
        RECT 39.950 181.625 40.615 181.795 ;
        RECT 39.935 180.695 40.265 181.455 ;
        RECT 40.445 180.865 40.615 181.625 ;
        RECT 40.880 180.865 41.215 181.835 ;
        RECT 41.385 180.695 41.555 181.835 ;
        RECT 41.725 181.035 41.895 182.005 ;
        RECT 42.065 181.375 42.235 182.505 ;
        RECT 42.405 181.715 42.575 182.515 ;
        RECT 42.775 182.395 43.055 182.565 ;
        RECT 42.780 181.915 43.055 182.395 ;
        RECT 43.225 181.715 43.415 183.075 ;
        RECT 43.595 182.710 44.105 183.245 ;
        RECT 44.325 182.435 44.570 183.040 ;
        RECT 45.565 182.695 45.735 183.075 ;
        RECT 45.915 182.865 46.245 183.245 ;
        RECT 45.565 182.525 46.230 182.695 ;
        RECT 46.425 182.570 46.685 183.075 ;
        RECT 43.615 182.265 44.845 182.435 ;
        RECT 42.405 181.545 43.415 181.715 ;
        RECT 43.585 181.700 44.335 181.890 ;
        RECT 42.065 181.205 43.190 181.375 ;
        RECT 43.585 181.035 43.755 181.700 ;
        RECT 44.505 181.455 44.845 182.265 ;
        RECT 45.495 181.975 45.825 182.345 ;
        RECT 46.060 182.270 46.230 182.525 ;
        RECT 46.060 181.940 46.345 182.270 ;
        RECT 46.060 181.795 46.230 181.940 ;
        RECT 41.725 180.865 43.755 181.035 ;
        RECT 43.925 180.695 44.095 181.455 ;
        RECT 44.330 181.045 44.845 181.455 ;
        RECT 45.565 181.625 46.230 181.795 ;
        RECT 46.515 181.770 46.685 182.570 ;
        RECT 47.130 182.435 47.375 183.040 ;
        RECT 47.595 182.710 48.105 183.245 ;
        RECT 45.565 180.865 45.735 181.625 ;
        RECT 45.915 180.695 46.245 181.455 ;
        RECT 46.415 180.865 46.685 181.770 ;
        RECT 46.855 182.265 48.085 182.435 ;
        RECT 46.855 181.455 47.195 182.265 ;
        RECT 47.365 181.700 48.115 181.890 ;
        RECT 46.855 181.045 47.370 181.455 ;
        RECT 47.605 180.695 47.775 181.455 ;
        RECT 47.945 181.035 48.115 181.700 ;
        RECT 48.285 181.715 48.475 183.075 ;
        RECT 48.645 182.225 48.920 183.075 ;
        RECT 49.110 182.710 49.640 183.075 ;
        RECT 50.065 182.845 50.395 183.245 ;
        RECT 49.465 182.675 49.640 182.710 ;
        RECT 48.645 182.055 48.925 182.225 ;
        RECT 48.645 181.915 48.920 182.055 ;
        RECT 49.125 181.715 49.295 182.515 ;
        RECT 48.285 181.545 49.295 181.715 ;
        RECT 49.465 182.505 50.395 182.675 ;
        RECT 50.565 182.505 50.820 183.075 ;
        RECT 49.465 181.375 49.635 182.505 ;
        RECT 50.225 182.335 50.395 182.505 ;
        RECT 48.510 181.205 49.635 181.375 ;
        RECT 49.805 182.005 50.000 182.335 ;
        RECT 50.225 182.005 50.480 182.335 ;
        RECT 49.805 181.035 49.975 182.005 ;
        RECT 50.650 181.835 50.820 182.505 ;
        RECT 47.945 180.865 49.975 181.035 ;
        RECT 50.145 180.695 50.315 181.835 ;
        RECT 50.485 180.865 50.820 181.835 ;
        RECT 51.000 182.535 51.255 183.065 ;
        RECT 51.425 182.785 51.730 183.245 ;
        RECT 51.975 182.865 53.045 183.035 ;
        RECT 51.000 181.885 51.210 182.535 ;
        RECT 51.975 182.510 52.295 182.865 ;
        RECT 51.970 182.335 52.295 182.510 ;
        RECT 51.380 182.035 52.295 182.335 ;
        RECT 52.465 182.295 52.705 182.695 ;
        RECT 52.875 182.635 53.045 182.865 ;
        RECT 53.215 182.805 53.405 183.245 ;
        RECT 53.575 182.795 54.525 183.075 ;
        RECT 54.745 182.885 55.095 183.055 ;
        RECT 52.875 182.465 53.405 182.635 ;
        RECT 51.380 182.005 52.120 182.035 ;
        RECT 51.000 181.005 51.255 181.885 ;
        RECT 51.425 180.695 51.730 181.835 ;
        RECT 51.950 181.415 52.120 182.005 ;
        RECT 52.465 181.925 53.005 182.295 ;
        RECT 53.185 182.185 53.405 182.465 ;
        RECT 53.575 182.015 53.745 182.795 ;
        RECT 53.340 181.845 53.745 182.015 ;
        RECT 53.915 182.005 54.265 182.625 ;
        RECT 53.340 181.755 53.510 181.845 ;
        RECT 54.435 181.835 54.645 182.625 ;
        RECT 52.290 181.585 53.510 181.755 ;
        RECT 53.970 181.675 54.645 181.835 ;
        RECT 51.950 181.245 52.750 181.415 ;
        RECT 52.070 180.695 52.400 181.075 ;
        RECT 52.580 180.955 52.750 181.245 ;
        RECT 53.340 181.205 53.510 181.585 ;
        RECT 53.680 181.665 54.645 181.675 ;
        RECT 54.835 182.495 55.095 182.885 ;
        RECT 55.305 182.785 55.635 183.245 ;
        RECT 56.510 182.855 57.365 183.025 ;
        RECT 57.570 182.855 58.065 183.025 ;
        RECT 58.235 182.885 58.565 183.245 ;
        RECT 54.835 181.805 55.005 182.495 ;
        RECT 55.175 182.145 55.345 182.325 ;
        RECT 55.515 182.315 56.305 182.565 ;
        RECT 56.510 182.145 56.680 182.855 ;
        RECT 56.850 182.345 57.205 182.565 ;
        RECT 55.175 181.975 56.865 182.145 ;
        RECT 53.680 181.375 54.140 181.665 ;
        RECT 54.835 181.635 56.335 181.805 ;
        RECT 54.835 181.495 55.005 181.635 ;
        RECT 54.445 181.325 55.005 181.495 ;
        RECT 52.920 180.695 53.170 181.155 ;
        RECT 53.340 180.865 54.210 181.205 ;
        RECT 54.445 180.865 54.615 181.325 ;
        RECT 55.450 181.295 56.525 181.465 ;
        RECT 54.785 180.695 55.155 181.155 ;
        RECT 55.450 180.955 55.620 181.295 ;
        RECT 55.790 180.695 56.120 181.125 ;
        RECT 56.355 180.955 56.525 181.295 ;
        RECT 56.695 181.195 56.865 181.975 ;
        RECT 57.035 181.755 57.205 182.345 ;
        RECT 57.375 181.945 57.725 182.565 ;
        RECT 57.035 181.365 57.500 181.755 ;
        RECT 57.895 181.495 58.065 182.855 ;
        RECT 58.235 181.665 58.695 182.715 ;
        RECT 57.670 181.325 58.065 181.495 ;
        RECT 57.670 181.195 57.840 181.325 ;
        RECT 56.695 180.865 57.375 181.195 ;
        RECT 57.590 180.865 57.840 181.195 ;
        RECT 58.010 180.695 58.260 181.155 ;
        RECT 58.430 180.880 58.755 181.665 ;
        RECT 58.925 180.865 59.095 182.985 ;
        RECT 59.265 182.865 59.595 183.245 ;
        RECT 59.765 182.695 60.020 182.985 ;
        RECT 59.270 182.525 60.020 182.695 ;
        RECT 59.270 181.535 59.500 182.525 ;
        RECT 61.115 182.520 61.405 183.245 ;
        RECT 61.580 182.535 61.835 183.065 ;
        RECT 62.005 182.785 62.310 183.245 ;
        RECT 62.555 182.865 63.625 183.035 ;
        RECT 59.670 181.705 60.020 182.355 ;
        RECT 61.580 181.885 61.790 182.535 ;
        RECT 62.555 182.510 62.875 182.865 ;
        RECT 62.550 182.335 62.875 182.510 ;
        RECT 61.960 182.035 62.875 182.335 ;
        RECT 63.045 182.295 63.285 182.695 ;
        RECT 63.455 182.635 63.625 182.865 ;
        RECT 63.795 182.805 63.985 183.245 ;
        RECT 64.155 182.795 65.105 183.075 ;
        RECT 65.325 182.885 65.675 183.055 ;
        RECT 63.455 182.465 63.985 182.635 ;
        RECT 61.960 182.005 62.700 182.035 ;
        RECT 59.270 181.365 60.020 181.535 ;
        RECT 59.265 180.695 59.595 181.195 ;
        RECT 59.765 180.865 60.020 181.365 ;
        RECT 61.115 180.695 61.405 181.860 ;
        RECT 61.580 181.005 61.835 181.885 ;
        RECT 62.005 180.695 62.310 181.835 ;
        RECT 62.530 181.415 62.700 182.005 ;
        RECT 63.045 181.925 63.585 182.295 ;
        RECT 63.765 182.185 63.985 182.465 ;
        RECT 64.155 182.015 64.325 182.795 ;
        RECT 63.920 181.845 64.325 182.015 ;
        RECT 64.495 182.005 64.845 182.625 ;
        RECT 63.920 181.755 64.090 181.845 ;
        RECT 65.015 181.835 65.225 182.625 ;
        RECT 62.870 181.585 64.090 181.755 ;
        RECT 64.550 181.675 65.225 181.835 ;
        RECT 62.530 181.245 63.330 181.415 ;
        RECT 62.650 180.695 62.980 181.075 ;
        RECT 63.160 180.955 63.330 181.245 ;
        RECT 63.920 181.205 64.090 181.585 ;
        RECT 64.260 181.665 65.225 181.675 ;
        RECT 65.415 182.495 65.675 182.885 ;
        RECT 65.885 182.785 66.215 183.245 ;
        RECT 67.090 182.855 67.945 183.025 ;
        RECT 68.150 182.855 68.645 183.025 ;
        RECT 68.815 182.885 69.145 183.245 ;
        RECT 65.415 181.805 65.585 182.495 ;
        RECT 65.755 182.145 65.925 182.325 ;
        RECT 66.095 182.315 66.885 182.565 ;
        RECT 67.090 182.145 67.260 182.855 ;
        RECT 67.430 182.345 67.785 182.565 ;
        RECT 65.755 181.975 67.445 182.145 ;
        RECT 64.260 181.375 64.720 181.665 ;
        RECT 65.415 181.635 66.915 181.805 ;
        RECT 65.415 181.495 65.585 181.635 ;
        RECT 65.025 181.325 65.585 181.495 ;
        RECT 63.500 180.695 63.750 181.155 ;
        RECT 63.920 180.865 64.790 181.205 ;
        RECT 65.025 180.865 65.195 181.325 ;
        RECT 66.030 181.295 67.105 181.465 ;
        RECT 65.365 180.695 65.735 181.155 ;
        RECT 66.030 180.955 66.200 181.295 ;
        RECT 66.370 180.695 66.700 181.125 ;
        RECT 66.935 180.955 67.105 181.295 ;
        RECT 67.275 181.195 67.445 181.975 ;
        RECT 67.615 181.755 67.785 182.345 ;
        RECT 67.955 181.945 68.305 182.565 ;
        RECT 67.615 181.365 68.080 181.755 ;
        RECT 68.475 181.495 68.645 182.855 ;
        RECT 68.815 181.665 69.275 182.715 ;
        RECT 68.250 181.325 68.645 181.495 ;
        RECT 68.250 181.195 68.420 181.325 ;
        RECT 67.275 180.865 67.955 181.195 ;
        RECT 68.170 180.865 68.420 181.195 ;
        RECT 68.590 180.695 68.840 181.155 ;
        RECT 69.010 180.880 69.335 181.665 ;
        RECT 69.505 180.865 69.675 182.985 ;
        RECT 69.845 182.865 70.175 183.245 ;
        RECT 70.345 182.695 70.600 182.985 ;
        RECT 69.850 182.525 70.600 182.695 ;
        RECT 69.850 181.535 70.080 182.525 ;
        RECT 70.775 182.505 71.095 182.985 ;
        RECT 71.265 182.675 71.495 183.075 ;
        RECT 71.665 182.855 72.015 183.245 ;
        RECT 71.265 182.595 71.775 182.675 ;
        RECT 72.185 182.595 72.515 183.075 ;
        RECT 71.265 182.505 72.515 182.595 ;
        RECT 70.250 181.705 70.600 182.355 ;
        RECT 70.775 181.575 70.945 182.505 ;
        RECT 71.605 182.425 72.515 182.505 ;
        RECT 72.685 182.425 72.855 183.245 ;
        RECT 73.360 182.505 73.825 183.050 ;
        RECT 71.115 181.915 71.285 182.335 ;
        RECT 71.515 182.085 72.115 182.255 ;
        RECT 71.115 181.745 71.775 181.915 ;
        RECT 69.850 181.365 70.600 181.535 ;
        RECT 70.775 181.375 71.435 181.575 ;
        RECT 71.605 181.545 71.775 181.745 ;
        RECT 71.945 181.885 72.115 182.085 ;
        RECT 72.285 182.055 72.980 182.255 ;
        RECT 73.240 181.885 73.485 182.335 ;
        RECT 71.945 181.715 73.485 181.885 ;
        RECT 73.655 181.545 73.825 182.505 ;
        RECT 74.455 182.475 77.045 183.245 ;
        RECT 71.605 181.375 73.825 181.545 ;
        RECT 74.455 181.785 75.665 182.305 ;
        RECT 75.835 181.955 77.045 182.475 ;
        RECT 77.590 182.535 77.845 183.065 ;
        RECT 78.025 182.785 78.310 183.245 ;
        RECT 69.845 180.695 70.175 181.195 ;
        RECT 70.345 180.865 70.600 181.365 ;
        RECT 71.265 181.205 71.435 181.375 ;
        RECT 70.795 180.695 71.095 181.205 ;
        RECT 71.265 181.035 71.645 181.205 ;
        RECT 72.225 180.695 72.855 181.205 ;
        RECT 73.025 180.865 73.355 181.375 ;
        RECT 73.525 180.695 73.825 181.205 ;
        RECT 74.455 180.695 77.045 181.785 ;
        RECT 77.590 181.675 77.770 182.535 ;
        RECT 78.490 182.335 78.740 182.985 ;
        RECT 77.940 182.005 78.740 182.335 ;
        RECT 77.590 181.205 77.845 181.675 ;
        RECT 77.505 181.035 77.845 181.205 ;
        RECT 77.590 181.005 77.845 181.035 ;
        RECT 78.025 180.695 78.310 181.495 ;
        RECT 78.490 181.415 78.740 182.005 ;
        RECT 78.940 182.650 79.260 182.980 ;
        RECT 79.440 182.765 80.100 183.245 ;
        RECT 80.300 182.855 81.150 183.025 ;
        RECT 78.940 181.755 79.130 182.650 ;
        RECT 79.450 182.325 80.110 182.595 ;
        RECT 79.780 182.265 80.110 182.325 ;
        RECT 79.300 182.095 79.630 182.155 ;
        RECT 80.300 182.095 80.470 182.855 ;
        RECT 81.710 182.785 82.030 183.245 ;
        RECT 82.230 182.605 82.480 183.035 ;
        RECT 82.770 182.805 83.180 183.245 ;
        RECT 83.350 182.865 84.365 183.065 ;
        RECT 80.640 182.435 81.890 182.605 ;
        RECT 80.640 182.315 80.970 182.435 ;
        RECT 79.300 181.925 81.200 182.095 ;
        RECT 78.940 181.585 80.860 181.755 ;
        RECT 78.940 181.565 79.260 181.585 ;
        RECT 78.490 180.905 78.820 181.415 ;
        RECT 79.090 180.955 79.260 181.565 ;
        RECT 81.030 181.415 81.200 181.925 ;
        RECT 81.370 181.855 81.550 182.265 ;
        RECT 81.720 181.675 81.890 182.435 ;
        RECT 79.430 180.695 79.760 181.385 ;
        RECT 79.990 181.245 81.200 181.415 ;
        RECT 81.370 181.365 81.890 181.675 ;
        RECT 82.060 182.265 82.480 182.605 ;
        RECT 82.770 182.265 83.180 182.595 ;
        RECT 82.060 181.495 82.250 182.265 ;
        RECT 83.350 182.135 83.520 182.865 ;
        RECT 84.665 182.695 84.835 183.025 ;
        RECT 85.005 182.865 85.335 183.245 ;
        RECT 83.690 182.315 84.040 182.685 ;
        RECT 83.350 182.095 83.770 182.135 ;
        RECT 82.420 181.925 83.770 182.095 ;
        RECT 82.420 181.765 82.670 181.925 ;
        RECT 83.180 181.495 83.430 181.755 ;
        RECT 82.060 181.245 83.430 181.495 ;
        RECT 79.990 180.955 80.230 181.245 ;
        RECT 81.030 181.165 81.200 181.245 ;
        RECT 80.430 180.695 80.850 181.075 ;
        RECT 81.030 180.915 81.660 181.165 ;
        RECT 82.130 180.695 82.460 181.075 ;
        RECT 82.630 180.955 82.800 181.245 ;
        RECT 83.600 181.080 83.770 181.925 ;
        RECT 84.220 181.755 84.440 182.625 ;
        RECT 84.665 182.505 85.360 182.695 ;
        RECT 83.940 181.375 84.440 181.755 ;
        RECT 84.610 181.705 85.020 182.325 ;
        RECT 85.190 181.535 85.360 182.505 ;
        RECT 84.665 181.365 85.360 181.535 ;
        RECT 82.980 180.695 83.360 181.075 ;
        RECT 83.600 180.910 84.430 181.080 ;
        RECT 84.665 180.865 84.835 181.365 ;
        RECT 85.005 180.695 85.335 181.195 ;
        RECT 85.550 180.865 85.775 182.985 ;
        RECT 85.945 182.865 86.275 183.245 ;
        RECT 86.445 182.695 86.615 182.985 ;
        RECT 85.950 182.525 86.615 182.695 ;
        RECT 85.950 181.535 86.180 182.525 ;
        RECT 86.875 182.520 87.165 183.245 ;
        RECT 87.335 182.570 87.595 183.075 ;
        RECT 87.775 182.865 88.105 183.245 ;
        RECT 88.285 182.695 88.455 183.075 ;
        RECT 86.350 181.705 86.700 182.355 ;
        RECT 85.950 181.365 86.615 181.535 ;
        RECT 85.945 180.695 86.275 181.195 ;
        RECT 86.445 180.865 86.615 181.365 ;
        RECT 86.875 180.695 87.165 181.860 ;
        RECT 87.335 181.770 87.505 182.570 ;
        RECT 87.790 182.525 88.455 182.695 ;
        RECT 87.790 182.270 87.960 182.525 ;
        RECT 89.175 182.475 91.765 183.245 ;
        RECT 91.940 182.700 97.285 183.245 ;
        RECT 87.675 181.940 87.960 182.270 ;
        RECT 88.195 181.975 88.525 182.345 ;
        RECT 87.790 181.795 87.960 181.940 ;
        RECT 87.335 180.865 87.605 181.770 ;
        RECT 87.790 181.625 88.455 181.795 ;
        RECT 87.775 180.695 88.105 181.455 ;
        RECT 88.285 180.865 88.455 181.625 ;
        RECT 89.175 181.785 90.385 182.305 ;
        RECT 90.555 181.955 91.765 182.475 ;
        RECT 89.175 180.695 91.765 181.785 ;
        RECT 93.530 181.130 93.880 182.380 ;
        RECT 95.360 181.870 95.700 182.700 ;
        RECT 97.515 182.425 97.725 183.245 ;
        RECT 97.895 182.445 98.225 183.075 ;
        RECT 97.895 181.845 98.145 182.445 ;
        RECT 98.395 182.425 98.625 183.245 ;
        RECT 99.295 182.475 101.885 183.245 ;
        RECT 98.315 182.005 98.645 182.255 ;
        RECT 91.940 180.695 97.285 181.130 ;
        RECT 97.515 180.695 97.725 181.835 ;
        RECT 97.895 180.865 98.225 181.845 ;
        RECT 98.395 180.695 98.625 181.835 ;
        RECT 99.295 181.785 100.505 182.305 ;
        RECT 100.675 181.955 101.885 182.475 ;
        RECT 102.095 182.425 102.325 183.245 ;
        RECT 102.495 182.445 102.825 183.075 ;
        RECT 102.075 182.005 102.405 182.255 ;
        RECT 102.575 181.845 102.825 182.445 ;
        RECT 102.995 182.425 103.205 183.245 ;
        RECT 103.710 182.435 103.955 183.040 ;
        RECT 104.175 182.710 104.685 183.245 ;
        RECT 99.295 180.695 101.885 181.785 ;
        RECT 102.095 180.695 102.325 181.835 ;
        RECT 102.495 180.865 102.825 181.845 ;
        RECT 103.435 182.265 104.665 182.435 ;
        RECT 102.995 180.695 103.205 181.835 ;
        RECT 103.435 181.455 103.775 182.265 ;
        RECT 103.945 181.700 104.695 181.890 ;
        RECT 103.435 181.045 103.950 181.455 ;
        RECT 104.185 180.695 104.355 181.455 ;
        RECT 104.525 181.035 104.695 181.700 ;
        RECT 104.865 181.715 105.055 183.075 ;
        RECT 105.225 182.225 105.500 183.075 ;
        RECT 105.690 182.710 106.220 183.075 ;
        RECT 106.645 182.845 106.975 183.245 ;
        RECT 106.045 182.675 106.220 182.710 ;
        RECT 105.225 182.055 105.505 182.225 ;
        RECT 105.225 181.915 105.500 182.055 ;
        RECT 105.705 181.715 105.875 182.515 ;
        RECT 104.865 181.545 105.875 181.715 ;
        RECT 106.045 182.505 106.975 182.675 ;
        RECT 107.145 182.505 107.400 183.075 ;
        RECT 106.045 181.375 106.215 182.505 ;
        RECT 106.805 182.335 106.975 182.505 ;
        RECT 105.090 181.205 106.215 181.375 ;
        RECT 106.385 182.005 106.580 182.335 ;
        RECT 106.805 182.005 107.060 182.335 ;
        RECT 106.385 181.035 106.555 182.005 ;
        RECT 107.230 181.835 107.400 182.505 ;
        RECT 107.850 182.435 108.095 183.040 ;
        RECT 108.315 182.710 108.825 183.245 ;
        RECT 104.525 180.865 106.555 181.035 ;
        RECT 106.725 180.695 106.895 181.835 ;
        RECT 107.065 180.865 107.400 181.835 ;
        RECT 107.575 182.265 108.805 182.435 ;
        RECT 107.575 181.455 107.915 182.265 ;
        RECT 108.085 181.700 108.835 181.890 ;
        RECT 107.575 181.045 108.090 181.455 ;
        RECT 108.325 180.695 108.495 181.455 ;
        RECT 108.665 181.035 108.835 181.700 ;
        RECT 109.005 181.715 109.195 183.075 ;
        RECT 109.365 182.565 109.640 183.075 ;
        RECT 109.830 182.710 110.360 183.075 ;
        RECT 110.785 182.845 111.115 183.245 ;
        RECT 110.185 182.675 110.360 182.710 ;
        RECT 109.365 182.395 109.645 182.565 ;
        RECT 109.365 181.915 109.640 182.395 ;
        RECT 109.845 181.715 110.015 182.515 ;
        RECT 109.005 181.545 110.015 181.715 ;
        RECT 110.185 182.505 111.115 182.675 ;
        RECT 111.285 182.505 111.540 183.075 ;
        RECT 112.635 182.520 112.925 183.245 ;
        RECT 113.560 182.700 118.905 183.245 ;
        RECT 119.080 182.700 124.425 183.245 ;
        RECT 110.185 181.375 110.355 182.505 ;
        RECT 110.945 182.335 111.115 182.505 ;
        RECT 109.230 181.205 110.355 181.375 ;
        RECT 110.525 182.005 110.720 182.335 ;
        RECT 110.945 182.005 111.200 182.335 ;
        RECT 110.525 181.035 110.695 182.005 ;
        RECT 111.370 181.835 111.540 182.505 ;
        RECT 108.665 180.865 110.695 181.035 ;
        RECT 110.865 180.695 111.035 181.835 ;
        RECT 111.205 180.865 111.540 181.835 ;
        RECT 112.635 180.695 112.925 181.860 ;
        RECT 115.150 181.130 115.500 182.380 ;
        RECT 116.980 181.870 117.320 182.700 ;
        RECT 120.670 181.130 121.020 182.380 ;
        RECT 122.500 181.870 122.840 182.700 ;
        RECT 124.595 182.495 125.805 183.245 ;
        RECT 124.595 181.785 125.115 182.325 ;
        RECT 125.285 181.955 125.805 182.495 ;
        RECT 113.560 180.695 118.905 181.130 ;
        RECT 119.080 180.695 124.425 181.130 ;
        RECT 124.595 180.695 125.805 181.785 ;
        RECT 11.810 180.525 125.890 180.695 ;
        RECT 11.895 179.435 13.105 180.525 ;
        RECT 11.895 178.725 12.415 179.265 ;
        RECT 12.585 178.895 13.105 179.435 ;
        RECT 13.275 179.435 16.785 180.525 ;
        RECT 16.960 180.090 22.305 180.525 ;
        RECT 13.275 178.915 14.965 179.435 ;
        RECT 15.135 178.745 16.785 179.265 ;
        RECT 18.550 178.840 18.900 180.090 ;
        RECT 22.475 179.360 22.765 180.525 ;
        RECT 22.935 179.435 24.145 180.525 ;
        RECT 24.315 179.435 27.825 180.525 ;
        RECT 28.000 180.090 33.345 180.525 ;
        RECT 33.520 180.090 38.865 180.525 ;
        RECT 11.895 177.975 13.105 178.725 ;
        RECT 13.275 177.975 16.785 178.745 ;
        RECT 20.380 178.520 20.720 179.350 ;
        RECT 22.935 178.895 23.455 179.435 ;
        RECT 23.625 178.725 24.145 179.265 ;
        RECT 24.315 178.915 26.005 179.435 ;
        RECT 26.175 178.745 27.825 179.265 ;
        RECT 29.590 178.840 29.940 180.090 ;
        RECT 16.960 177.975 22.305 178.520 ;
        RECT 22.475 177.975 22.765 178.700 ;
        RECT 22.935 177.975 24.145 178.725 ;
        RECT 24.315 177.975 27.825 178.745 ;
        RECT 31.420 178.520 31.760 179.350 ;
        RECT 35.110 178.840 35.460 180.090 ;
        RECT 39.150 179.895 39.435 180.355 ;
        RECT 39.605 180.065 39.875 180.525 ;
        RECT 39.150 179.675 40.105 179.895 ;
        RECT 36.940 178.520 37.280 179.350 ;
        RECT 39.035 178.945 39.725 179.505 ;
        RECT 39.895 178.775 40.105 179.675 ;
        RECT 39.150 178.605 40.105 178.775 ;
        RECT 40.275 179.505 40.675 180.355 ;
        RECT 40.865 179.895 41.145 180.355 ;
        RECT 41.665 180.065 41.990 180.525 ;
        RECT 40.865 179.675 41.990 179.895 ;
        RECT 40.275 178.945 41.370 179.505 ;
        RECT 41.540 179.215 41.990 179.675 ;
        RECT 42.160 179.385 42.545 180.355 ;
        RECT 28.000 177.975 33.345 178.520 ;
        RECT 33.520 177.975 38.865 178.520 ;
        RECT 39.150 178.145 39.435 178.605 ;
        RECT 39.605 177.975 39.875 178.435 ;
        RECT 40.275 178.145 40.675 178.945 ;
        RECT 41.540 178.885 42.095 179.215 ;
        RECT 41.540 178.775 41.990 178.885 ;
        RECT 40.865 178.605 41.990 178.775 ;
        RECT 42.265 178.715 42.545 179.385 ;
        RECT 42.715 179.765 43.230 180.175 ;
        RECT 43.465 179.765 43.635 180.525 ;
        RECT 43.805 180.185 45.835 180.355 ;
        RECT 42.715 178.955 43.055 179.765 ;
        RECT 43.805 179.520 43.975 180.185 ;
        RECT 44.370 179.845 45.495 180.015 ;
        RECT 43.225 179.330 43.975 179.520 ;
        RECT 44.145 179.505 45.155 179.675 ;
        RECT 42.715 178.785 43.945 178.955 ;
        RECT 40.865 178.145 41.145 178.605 ;
        RECT 41.665 177.975 41.990 178.435 ;
        RECT 42.160 178.145 42.545 178.715 ;
        RECT 42.990 178.180 43.235 178.785 ;
        RECT 43.455 177.975 43.965 178.510 ;
        RECT 44.145 178.145 44.335 179.505 ;
        RECT 44.505 179.165 44.780 179.305 ;
        RECT 44.505 178.995 44.785 179.165 ;
        RECT 44.505 178.145 44.780 178.995 ;
        RECT 44.985 178.705 45.155 179.505 ;
        RECT 45.325 178.715 45.495 179.845 ;
        RECT 45.665 179.215 45.835 180.185 ;
        RECT 46.005 179.385 46.175 180.525 ;
        RECT 46.345 179.385 46.680 180.355 ;
        RECT 45.665 178.885 45.860 179.215 ;
        RECT 46.085 178.885 46.340 179.215 ;
        RECT 46.085 178.715 46.255 178.885 ;
        RECT 46.510 178.715 46.680 179.385 ;
        RECT 46.855 179.435 48.065 180.525 ;
        RECT 46.855 178.895 47.375 179.435 ;
        RECT 48.235 179.360 48.525 180.525 ;
        RECT 49.155 179.435 51.745 180.525 ;
        RECT 51.915 179.765 52.430 180.175 ;
        RECT 52.665 179.765 52.835 180.525 ;
        RECT 53.005 180.185 55.035 180.355 ;
        RECT 47.545 178.725 48.065 179.265 ;
        RECT 49.155 178.915 50.365 179.435 ;
        RECT 50.535 178.745 51.745 179.265 ;
        RECT 51.915 178.955 52.255 179.765 ;
        RECT 53.005 179.520 53.175 180.185 ;
        RECT 53.570 179.845 54.695 180.015 ;
        RECT 52.425 179.330 53.175 179.520 ;
        RECT 53.345 179.505 54.355 179.675 ;
        RECT 51.915 178.785 53.145 178.955 ;
        RECT 45.325 178.545 46.255 178.715 ;
        RECT 45.325 178.510 45.500 178.545 ;
        RECT 44.970 178.145 45.500 178.510 ;
        RECT 45.925 177.975 46.255 178.375 ;
        RECT 46.425 178.145 46.680 178.715 ;
        RECT 46.855 177.975 48.065 178.725 ;
        RECT 48.235 177.975 48.525 178.700 ;
        RECT 49.155 177.975 51.745 178.745 ;
        RECT 52.190 178.180 52.435 178.785 ;
        RECT 52.655 177.975 53.165 178.510 ;
        RECT 53.345 178.145 53.535 179.505 ;
        RECT 53.705 178.485 53.980 179.305 ;
        RECT 54.185 178.705 54.355 179.505 ;
        RECT 54.525 178.715 54.695 179.845 ;
        RECT 54.865 179.215 55.035 180.185 ;
        RECT 55.205 179.385 55.375 180.525 ;
        RECT 55.545 179.385 55.880 180.355 ;
        RECT 56.605 179.595 56.775 180.355 ;
        RECT 56.955 179.765 57.285 180.525 ;
        RECT 56.605 179.425 57.270 179.595 ;
        RECT 57.455 179.450 57.725 180.355 ;
        RECT 54.865 178.885 55.060 179.215 ;
        RECT 55.285 178.885 55.540 179.215 ;
        RECT 55.285 178.715 55.455 178.885 ;
        RECT 55.710 178.715 55.880 179.385 ;
        RECT 57.100 179.280 57.270 179.425 ;
        RECT 56.535 178.875 56.865 179.245 ;
        RECT 57.100 178.950 57.385 179.280 ;
        RECT 54.525 178.545 55.455 178.715 ;
        RECT 54.525 178.510 54.700 178.545 ;
        RECT 53.705 178.315 53.985 178.485 ;
        RECT 53.705 178.145 53.980 178.315 ;
        RECT 54.170 178.145 54.700 178.510 ;
        RECT 55.125 177.975 55.455 178.375 ;
        RECT 55.625 178.145 55.880 178.715 ;
        RECT 57.100 178.695 57.270 178.950 ;
        RECT 56.605 178.525 57.270 178.695 ;
        RECT 57.555 178.650 57.725 179.450 ;
        RECT 57.895 179.435 60.485 180.525 ;
        RECT 60.660 180.090 66.005 180.525 ;
        RECT 57.895 178.915 59.105 179.435 ;
        RECT 59.275 178.745 60.485 179.265 ;
        RECT 62.250 178.840 62.600 180.090 ;
        RECT 66.185 179.545 66.515 180.355 ;
        RECT 66.685 179.725 66.925 180.525 ;
        RECT 66.185 179.375 66.900 179.545 ;
        RECT 56.605 178.145 56.775 178.525 ;
        RECT 56.955 177.975 57.285 178.355 ;
        RECT 57.465 178.145 57.725 178.650 ;
        RECT 57.895 177.975 60.485 178.745 ;
        RECT 64.080 178.520 64.420 179.350 ;
        RECT 66.180 178.965 66.560 179.205 ;
        RECT 66.730 179.135 66.900 179.375 ;
        RECT 67.105 179.505 67.275 180.355 ;
        RECT 67.445 179.725 67.775 180.525 ;
        RECT 67.945 179.505 68.115 180.355 ;
        RECT 67.105 179.335 68.115 179.505 ;
        RECT 68.285 179.375 68.615 180.525 ;
        RECT 68.935 179.435 70.145 180.525 ;
        RECT 70.315 179.435 73.825 180.525 ;
        RECT 66.730 178.965 67.230 179.135 ;
        RECT 66.730 178.795 66.900 178.965 ;
        RECT 67.620 178.795 68.115 179.335 ;
        RECT 68.935 178.895 69.455 179.435 ;
        RECT 66.265 178.625 66.900 178.795 ;
        RECT 67.105 178.625 68.115 178.795 ;
        RECT 60.660 177.975 66.005 178.520 ;
        RECT 66.265 178.145 66.435 178.625 ;
        RECT 66.615 177.975 66.855 178.455 ;
        RECT 67.105 178.145 67.275 178.625 ;
        RECT 67.445 177.975 67.775 178.455 ;
        RECT 67.945 178.145 68.115 178.625 ;
        RECT 68.285 177.975 68.615 178.775 ;
        RECT 69.625 178.725 70.145 179.265 ;
        RECT 70.315 178.915 72.005 179.435 ;
        RECT 73.995 179.360 74.285 180.525 ;
        RECT 74.455 179.765 74.970 180.175 ;
        RECT 75.205 179.765 75.375 180.525 ;
        RECT 75.545 180.185 77.575 180.355 ;
        RECT 72.175 178.745 73.825 179.265 ;
        RECT 74.455 178.955 74.795 179.765 ;
        RECT 75.545 179.520 75.715 180.185 ;
        RECT 76.110 179.845 77.235 180.015 ;
        RECT 74.965 179.330 75.715 179.520 ;
        RECT 75.885 179.505 76.895 179.675 ;
        RECT 74.455 178.785 75.685 178.955 ;
        RECT 68.935 177.975 70.145 178.725 ;
        RECT 70.315 177.975 73.825 178.745 ;
        RECT 73.995 177.975 74.285 178.700 ;
        RECT 74.730 178.180 74.975 178.785 ;
        RECT 75.195 177.975 75.705 178.510 ;
        RECT 75.885 178.145 76.075 179.505 ;
        RECT 76.245 178.485 76.520 179.305 ;
        RECT 76.725 178.705 76.895 179.505 ;
        RECT 77.065 178.715 77.235 179.845 ;
        RECT 77.405 179.215 77.575 180.185 ;
        RECT 77.745 179.385 77.915 180.525 ;
        RECT 78.085 179.385 78.420 180.355 ;
        RECT 77.405 178.885 77.600 179.215 ;
        RECT 77.825 178.885 78.080 179.215 ;
        RECT 77.825 178.715 77.995 178.885 ;
        RECT 78.250 178.715 78.420 179.385 ;
        RECT 77.065 178.545 77.995 178.715 ;
        RECT 77.065 178.510 77.240 178.545 ;
        RECT 76.245 178.315 76.525 178.485 ;
        RECT 76.245 178.145 76.520 178.315 ;
        RECT 76.710 178.145 77.240 178.510 ;
        RECT 77.665 177.975 77.995 178.375 ;
        RECT 78.165 178.145 78.420 178.715 ;
        RECT 78.970 179.545 79.225 180.215 ;
        RECT 79.405 179.725 79.690 180.525 ;
        RECT 79.870 179.805 80.200 180.315 ;
        RECT 78.970 178.685 79.150 179.545 ;
        RECT 79.870 179.215 80.120 179.805 ;
        RECT 80.470 179.655 80.640 180.265 ;
        RECT 80.810 179.835 81.140 180.525 ;
        RECT 81.370 179.975 81.610 180.265 ;
        RECT 81.810 180.145 82.230 180.525 ;
        RECT 82.410 180.055 83.040 180.305 ;
        RECT 83.510 180.145 83.840 180.525 ;
        RECT 82.410 179.975 82.580 180.055 ;
        RECT 84.010 179.975 84.180 180.265 ;
        RECT 84.360 180.145 84.740 180.525 ;
        RECT 84.980 180.140 85.810 180.310 ;
        RECT 81.370 179.805 82.580 179.975 ;
        RECT 79.320 178.885 80.120 179.215 ;
        RECT 78.970 178.485 79.225 178.685 ;
        RECT 78.885 178.315 79.225 178.485 ;
        RECT 78.970 178.155 79.225 178.315 ;
        RECT 79.405 177.975 79.690 178.435 ;
        RECT 79.870 178.235 80.120 178.885 ;
        RECT 80.320 179.635 80.640 179.655 ;
        RECT 80.320 179.465 82.240 179.635 ;
        RECT 80.320 178.570 80.510 179.465 ;
        RECT 82.410 179.295 82.580 179.805 ;
        RECT 82.750 179.545 83.270 179.855 ;
        RECT 80.680 179.125 82.580 179.295 ;
        RECT 80.680 179.065 81.010 179.125 ;
        RECT 81.160 178.895 81.490 178.955 ;
        RECT 80.830 178.625 81.490 178.895 ;
        RECT 80.320 178.240 80.640 178.570 ;
        RECT 80.820 177.975 81.480 178.455 ;
        RECT 81.680 178.365 81.850 179.125 ;
        RECT 82.750 178.955 82.930 179.365 ;
        RECT 82.020 178.785 82.350 178.905 ;
        RECT 83.100 178.785 83.270 179.545 ;
        RECT 82.020 178.615 83.270 178.785 ;
        RECT 83.440 179.725 84.810 179.975 ;
        RECT 83.440 178.955 83.630 179.725 ;
        RECT 84.560 179.465 84.810 179.725 ;
        RECT 83.800 179.295 84.050 179.455 ;
        RECT 84.980 179.295 85.150 180.140 ;
        RECT 86.045 179.855 86.215 180.355 ;
        RECT 86.385 180.025 86.715 180.525 ;
        RECT 85.320 179.465 85.820 179.845 ;
        RECT 86.045 179.685 86.740 179.855 ;
        RECT 83.800 179.125 85.150 179.295 ;
        RECT 84.730 179.085 85.150 179.125 ;
        RECT 83.440 178.615 83.860 178.955 ;
        RECT 84.150 178.625 84.560 178.955 ;
        RECT 81.680 178.195 82.530 178.365 ;
        RECT 83.090 177.975 83.410 178.435 ;
        RECT 83.610 178.185 83.860 178.615 ;
        RECT 84.150 177.975 84.560 178.415 ;
        RECT 84.730 178.355 84.900 179.085 ;
        RECT 85.070 178.535 85.420 178.905 ;
        RECT 85.600 178.595 85.820 179.465 ;
        RECT 85.990 178.895 86.400 179.515 ;
        RECT 86.570 178.715 86.740 179.685 ;
        RECT 86.045 178.525 86.740 178.715 ;
        RECT 84.730 178.155 85.745 178.355 ;
        RECT 86.045 178.195 86.215 178.525 ;
        RECT 86.385 177.975 86.715 178.355 ;
        RECT 86.930 178.235 87.155 180.355 ;
        RECT 87.325 180.025 87.655 180.525 ;
        RECT 87.825 179.855 87.995 180.355 ;
        RECT 87.330 179.685 87.995 179.855 ;
        RECT 87.330 178.695 87.560 179.685 ;
        RECT 87.730 178.865 88.080 179.515 ;
        RECT 88.715 179.435 90.385 180.525 ;
        RECT 90.560 179.855 90.815 180.355 ;
        RECT 90.985 180.025 91.315 180.525 ;
        RECT 90.560 179.685 91.310 179.855 ;
        RECT 88.715 178.915 89.465 179.435 ;
        RECT 89.635 178.745 90.385 179.265 ;
        RECT 90.560 178.865 90.910 179.515 ;
        RECT 87.330 178.525 87.995 178.695 ;
        RECT 87.325 177.975 87.655 178.355 ;
        RECT 87.825 178.235 87.995 178.525 ;
        RECT 88.715 177.975 90.385 178.745 ;
        RECT 91.080 178.695 91.310 179.685 ;
        RECT 90.560 178.525 91.310 178.695 ;
        RECT 90.560 178.235 90.815 178.525 ;
        RECT 90.985 177.975 91.315 178.355 ;
        RECT 91.485 178.235 91.655 180.355 ;
        RECT 91.825 179.555 92.150 180.340 ;
        RECT 92.320 180.065 92.570 180.525 ;
        RECT 92.740 180.025 92.990 180.355 ;
        RECT 93.205 180.025 93.885 180.355 ;
        RECT 92.740 179.895 92.910 180.025 ;
        RECT 92.515 179.725 92.910 179.895 ;
        RECT 91.885 178.505 92.345 179.555 ;
        RECT 92.515 178.365 92.685 179.725 ;
        RECT 93.080 179.465 93.545 179.855 ;
        RECT 92.855 178.655 93.205 179.275 ;
        RECT 93.375 178.875 93.545 179.465 ;
        RECT 93.715 179.245 93.885 180.025 ;
        RECT 94.055 179.925 94.225 180.265 ;
        RECT 94.460 180.095 94.790 180.525 ;
        RECT 94.960 179.925 95.130 180.265 ;
        RECT 95.425 180.065 95.795 180.525 ;
        RECT 94.055 179.755 95.130 179.925 ;
        RECT 95.965 179.895 96.135 180.355 ;
        RECT 96.370 180.015 97.240 180.355 ;
        RECT 97.410 180.065 97.660 180.525 ;
        RECT 95.575 179.725 96.135 179.895 ;
        RECT 95.575 179.585 95.745 179.725 ;
        RECT 94.245 179.415 95.745 179.585 ;
        RECT 96.440 179.555 96.900 179.845 ;
        RECT 93.715 179.075 95.405 179.245 ;
        RECT 93.375 178.655 93.730 178.875 ;
        RECT 93.900 178.365 94.070 179.075 ;
        RECT 94.275 178.655 95.065 178.905 ;
        RECT 95.235 178.895 95.405 179.075 ;
        RECT 95.575 178.725 95.745 179.415 ;
        RECT 92.015 177.975 92.345 178.335 ;
        RECT 92.515 178.195 93.010 178.365 ;
        RECT 93.215 178.195 94.070 178.365 ;
        RECT 94.945 177.975 95.275 178.435 ;
        RECT 95.485 178.335 95.745 178.725 ;
        RECT 95.935 179.545 96.900 179.555 ;
        RECT 97.070 179.635 97.240 180.015 ;
        RECT 97.830 179.975 98.000 180.265 ;
        RECT 98.180 180.145 98.510 180.525 ;
        RECT 97.830 179.805 98.630 179.975 ;
        RECT 95.935 179.385 96.610 179.545 ;
        RECT 97.070 179.465 98.290 179.635 ;
        RECT 95.935 178.595 96.145 179.385 ;
        RECT 97.070 179.375 97.240 179.465 ;
        RECT 96.315 178.595 96.665 179.215 ;
        RECT 96.835 179.205 97.240 179.375 ;
        RECT 96.835 178.425 97.005 179.205 ;
        RECT 97.175 178.755 97.395 179.035 ;
        RECT 97.575 178.925 98.115 179.295 ;
        RECT 98.460 179.215 98.630 179.805 ;
        RECT 98.850 179.385 99.155 180.525 ;
        RECT 99.325 179.335 99.580 180.215 ;
        RECT 99.755 179.360 100.045 180.525 ;
        RECT 100.675 179.435 103.265 180.525 ;
        RECT 98.460 179.185 99.200 179.215 ;
        RECT 97.175 178.585 97.705 178.755 ;
        RECT 95.485 178.165 95.835 178.335 ;
        RECT 96.055 178.145 97.005 178.425 ;
        RECT 97.175 177.975 97.365 178.415 ;
        RECT 97.535 178.355 97.705 178.585 ;
        RECT 97.875 178.525 98.115 178.925 ;
        RECT 98.285 178.885 99.200 179.185 ;
        RECT 98.285 178.710 98.610 178.885 ;
        RECT 98.285 178.355 98.605 178.710 ;
        RECT 99.370 178.685 99.580 179.335 ;
        RECT 100.675 178.915 101.885 179.435 ;
        RECT 103.440 179.335 103.695 180.215 ;
        RECT 103.865 179.385 104.170 180.525 ;
        RECT 104.510 180.145 104.840 180.525 ;
        RECT 105.020 179.975 105.190 180.265 ;
        RECT 105.360 180.065 105.610 180.525 ;
        RECT 104.390 179.805 105.190 179.975 ;
        RECT 105.780 180.015 106.650 180.355 ;
        RECT 102.055 178.745 103.265 179.265 ;
        RECT 97.535 178.185 98.605 178.355 ;
        RECT 98.850 177.975 99.155 178.435 ;
        RECT 99.325 178.155 99.580 178.685 ;
        RECT 99.755 177.975 100.045 178.700 ;
        RECT 100.675 177.975 103.265 178.745 ;
        RECT 103.440 178.685 103.650 179.335 ;
        RECT 104.390 179.215 104.560 179.805 ;
        RECT 105.780 179.635 105.950 180.015 ;
        RECT 106.885 179.895 107.055 180.355 ;
        RECT 107.225 180.065 107.595 180.525 ;
        RECT 107.890 179.925 108.060 180.265 ;
        RECT 108.230 180.095 108.560 180.525 ;
        RECT 108.795 179.925 108.965 180.265 ;
        RECT 104.730 179.465 105.950 179.635 ;
        RECT 106.120 179.555 106.580 179.845 ;
        RECT 106.885 179.725 107.445 179.895 ;
        RECT 107.890 179.755 108.965 179.925 ;
        RECT 109.135 180.025 109.815 180.355 ;
        RECT 110.030 180.025 110.280 180.355 ;
        RECT 110.450 180.065 110.700 180.525 ;
        RECT 107.275 179.585 107.445 179.725 ;
        RECT 106.120 179.545 107.085 179.555 ;
        RECT 105.780 179.375 105.950 179.465 ;
        RECT 106.410 179.385 107.085 179.545 ;
        RECT 103.820 179.185 104.560 179.215 ;
        RECT 103.820 178.885 104.735 179.185 ;
        RECT 104.410 178.710 104.735 178.885 ;
        RECT 103.440 178.155 103.695 178.685 ;
        RECT 103.865 177.975 104.170 178.435 ;
        RECT 104.415 178.355 104.735 178.710 ;
        RECT 104.905 178.925 105.445 179.295 ;
        RECT 105.780 179.205 106.185 179.375 ;
        RECT 104.905 178.525 105.145 178.925 ;
        RECT 105.625 178.755 105.845 179.035 ;
        RECT 105.315 178.585 105.845 178.755 ;
        RECT 105.315 178.355 105.485 178.585 ;
        RECT 106.015 178.425 106.185 179.205 ;
        RECT 106.355 178.595 106.705 179.215 ;
        RECT 106.875 178.595 107.085 179.385 ;
        RECT 107.275 179.415 108.775 179.585 ;
        RECT 107.275 178.725 107.445 179.415 ;
        RECT 109.135 179.245 109.305 180.025 ;
        RECT 110.110 179.895 110.280 180.025 ;
        RECT 107.615 179.075 109.305 179.245 ;
        RECT 109.475 179.465 109.940 179.855 ;
        RECT 110.110 179.725 110.505 179.895 ;
        RECT 107.615 178.895 107.785 179.075 ;
        RECT 104.415 178.185 105.485 178.355 ;
        RECT 105.655 177.975 105.845 178.415 ;
        RECT 106.015 178.145 106.965 178.425 ;
        RECT 107.275 178.335 107.535 178.725 ;
        RECT 107.955 178.655 108.745 178.905 ;
        RECT 107.185 178.165 107.535 178.335 ;
        RECT 107.745 177.975 108.075 178.435 ;
        RECT 108.950 178.365 109.120 179.075 ;
        RECT 109.475 178.875 109.645 179.465 ;
        RECT 109.290 178.655 109.645 178.875 ;
        RECT 109.815 178.655 110.165 179.275 ;
        RECT 110.335 178.365 110.505 179.725 ;
        RECT 110.870 179.555 111.195 180.340 ;
        RECT 110.675 178.505 111.135 179.555 ;
        RECT 108.950 178.195 109.805 178.365 ;
        RECT 110.010 178.195 110.505 178.365 ;
        RECT 110.675 177.975 111.005 178.335 ;
        RECT 111.365 178.235 111.535 180.355 ;
        RECT 111.705 180.025 112.035 180.525 ;
        RECT 112.205 179.855 112.460 180.355 ;
        RECT 113.560 180.090 118.905 180.525 ;
        RECT 119.080 180.090 124.425 180.525 ;
        RECT 111.710 179.685 112.460 179.855 ;
        RECT 111.710 178.695 111.940 179.685 ;
        RECT 112.110 178.865 112.460 179.515 ;
        RECT 115.150 178.840 115.500 180.090 ;
        RECT 111.710 178.525 112.460 178.695 ;
        RECT 111.705 177.975 112.035 178.355 ;
        RECT 112.205 178.235 112.460 178.525 ;
        RECT 116.980 178.520 117.320 179.350 ;
        RECT 120.670 178.840 121.020 180.090 ;
        RECT 124.595 179.435 125.805 180.525 ;
        RECT 122.500 178.520 122.840 179.350 ;
        RECT 124.595 178.895 125.115 179.435 ;
        RECT 125.285 178.725 125.805 179.265 ;
        RECT 113.560 177.975 118.905 178.520 ;
        RECT 119.080 177.975 124.425 178.520 ;
        RECT 124.595 177.975 125.805 178.725 ;
        RECT 11.810 177.805 125.890 177.975 ;
        RECT 11.895 177.055 13.105 177.805 ;
        RECT 13.740 177.260 19.085 177.805 ;
        RECT 19.260 177.260 24.605 177.805 ;
        RECT 24.780 177.260 30.125 177.805 ;
        RECT 11.895 176.515 12.415 177.055 ;
        RECT 12.585 176.345 13.105 176.885 ;
        RECT 11.895 175.255 13.105 176.345 ;
        RECT 15.330 175.690 15.680 176.940 ;
        RECT 17.160 176.430 17.500 177.260 ;
        RECT 20.850 175.690 21.200 176.940 ;
        RECT 22.680 176.430 23.020 177.260 ;
        RECT 26.370 175.690 26.720 176.940 ;
        RECT 28.200 176.430 28.540 177.260 ;
        RECT 30.335 176.985 30.565 177.805 ;
        RECT 30.735 177.005 31.065 177.635 ;
        RECT 30.315 176.565 30.645 176.815 ;
        RECT 30.815 176.405 31.065 177.005 ;
        RECT 31.235 176.985 31.445 177.805 ;
        RECT 31.675 177.035 35.185 177.805 ;
        RECT 35.355 177.080 35.645 177.805 ;
        RECT 36.275 177.035 37.945 177.805 ;
        RECT 13.740 175.255 19.085 175.690 ;
        RECT 19.260 175.255 24.605 175.690 ;
        RECT 24.780 175.255 30.125 175.690 ;
        RECT 30.335 175.255 30.565 176.395 ;
        RECT 30.735 175.425 31.065 176.405 ;
        RECT 31.235 175.255 31.445 176.395 ;
        RECT 31.675 176.345 33.365 176.865 ;
        RECT 33.535 176.515 35.185 177.035 ;
        RECT 31.675 175.255 35.185 176.345 ;
        RECT 35.355 175.255 35.645 176.420 ;
        RECT 36.275 176.345 37.025 176.865 ;
        RECT 37.195 176.515 37.945 177.035 ;
        RECT 38.155 176.985 38.385 177.805 ;
        RECT 38.555 177.005 38.885 177.635 ;
        RECT 38.135 176.565 38.465 176.815 ;
        RECT 38.635 176.405 38.885 177.005 ;
        RECT 39.055 176.985 39.265 177.805 ;
        RECT 39.500 177.095 39.755 177.625 ;
        RECT 39.925 177.345 40.230 177.805 ;
        RECT 40.475 177.425 41.545 177.595 ;
        RECT 36.275 175.255 37.945 176.345 ;
        RECT 38.155 175.255 38.385 176.395 ;
        RECT 38.555 175.425 38.885 176.405 ;
        RECT 39.500 176.445 39.710 177.095 ;
        RECT 40.475 177.070 40.795 177.425 ;
        RECT 40.470 176.895 40.795 177.070 ;
        RECT 39.880 176.595 40.795 176.895 ;
        RECT 40.965 176.855 41.205 177.255 ;
        RECT 41.375 177.195 41.545 177.425 ;
        RECT 41.715 177.365 41.905 177.805 ;
        RECT 42.075 177.355 43.025 177.635 ;
        RECT 43.245 177.445 43.595 177.615 ;
        RECT 41.375 177.025 41.905 177.195 ;
        RECT 39.880 176.565 40.620 176.595 ;
        RECT 39.055 175.255 39.265 176.395 ;
        RECT 39.500 175.565 39.755 176.445 ;
        RECT 39.925 175.255 40.230 176.395 ;
        RECT 40.450 175.975 40.620 176.565 ;
        RECT 40.965 176.485 41.505 176.855 ;
        RECT 41.685 176.745 41.905 177.025 ;
        RECT 42.075 176.575 42.245 177.355 ;
        RECT 41.840 176.405 42.245 176.575 ;
        RECT 42.415 176.565 42.765 177.185 ;
        RECT 41.840 176.315 42.010 176.405 ;
        RECT 42.935 176.395 43.145 177.185 ;
        RECT 40.790 176.145 42.010 176.315 ;
        RECT 42.470 176.235 43.145 176.395 ;
        RECT 40.450 175.805 41.250 175.975 ;
        RECT 40.570 175.255 40.900 175.635 ;
        RECT 41.080 175.515 41.250 175.805 ;
        RECT 41.840 175.765 42.010 176.145 ;
        RECT 42.180 176.225 43.145 176.235 ;
        RECT 43.335 177.055 43.595 177.445 ;
        RECT 43.805 177.345 44.135 177.805 ;
        RECT 45.010 177.415 45.865 177.585 ;
        RECT 46.070 177.415 46.565 177.585 ;
        RECT 46.735 177.445 47.065 177.805 ;
        RECT 43.335 176.365 43.505 177.055 ;
        RECT 43.675 176.705 43.845 176.885 ;
        RECT 44.015 176.875 44.805 177.125 ;
        RECT 45.010 176.705 45.180 177.415 ;
        RECT 45.350 176.905 45.705 177.125 ;
        RECT 43.675 176.535 45.365 176.705 ;
        RECT 42.180 175.935 42.640 176.225 ;
        RECT 43.335 176.195 44.835 176.365 ;
        RECT 43.335 176.055 43.505 176.195 ;
        RECT 42.945 175.885 43.505 176.055 ;
        RECT 41.420 175.255 41.670 175.715 ;
        RECT 41.840 175.425 42.710 175.765 ;
        RECT 42.945 175.425 43.115 175.885 ;
        RECT 43.950 175.855 45.025 176.025 ;
        RECT 43.285 175.255 43.655 175.715 ;
        RECT 43.950 175.515 44.120 175.855 ;
        RECT 44.290 175.255 44.620 175.685 ;
        RECT 44.855 175.515 45.025 175.855 ;
        RECT 45.195 175.755 45.365 176.535 ;
        RECT 45.535 176.315 45.705 176.905 ;
        RECT 45.875 176.505 46.225 177.125 ;
        RECT 45.535 175.925 46.000 176.315 ;
        RECT 46.395 176.055 46.565 177.415 ;
        RECT 46.735 176.225 47.195 177.275 ;
        RECT 46.170 175.885 46.565 176.055 ;
        RECT 46.170 175.755 46.340 175.885 ;
        RECT 45.195 175.425 45.875 175.755 ;
        RECT 46.090 175.425 46.340 175.755 ;
        RECT 46.510 175.255 46.760 175.715 ;
        RECT 46.930 175.440 47.255 176.225 ;
        RECT 47.425 175.425 47.595 177.545 ;
        RECT 47.765 177.425 48.095 177.805 ;
        RECT 48.265 177.255 48.520 177.545 ;
        RECT 47.770 177.085 48.520 177.255 ;
        RECT 47.770 176.095 48.000 177.085 ;
        RECT 48.695 177.055 49.905 177.805 ;
        RECT 50.080 177.260 55.425 177.805 ;
        RECT 48.170 176.265 48.520 176.915 ;
        RECT 48.695 176.345 49.215 176.885 ;
        RECT 49.385 176.515 49.905 177.055 ;
        RECT 47.770 175.925 48.520 176.095 ;
        RECT 47.765 175.255 48.095 175.755 ;
        RECT 48.265 175.425 48.520 175.925 ;
        RECT 48.695 175.255 49.905 176.345 ;
        RECT 51.670 175.690 52.020 176.940 ;
        RECT 53.500 176.430 53.840 177.260 ;
        RECT 55.655 176.985 55.865 177.805 ;
        RECT 56.035 177.005 56.365 177.635 ;
        RECT 56.035 176.405 56.285 177.005 ;
        RECT 56.535 176.985 56.765 177.805 ;
        RECT 57.435 177.035 60.945 177.805 ;
        RECT 61.115 177.080 61.405 177.805 ;
        RECT 61.575 177.035 64.165 177.805 ;
        RECT 64.340 177.260 69.685 177.805 ;
        RECT 70.125 177.410 70.455 177.805 ;
        RECT 56.455 176.565 56.785 176.815 ;
        RECT 50.080 175.255 55.425 175.690 ;
        RECT 55.655 175.255 55.865 176.395 ;
        RECT 56.035 175.425 56.365 176.405 ;
        RECT 56.535 175.255 56.765 176.395 ;
        RECT 57.435 176.345 59.125 176.865 ;
        RECT 59.295 176.515 60.945 177.035 ;
        RECT 57.435 175.255 60.945 176.345 ;
        RECT 61.115 175.255 61.405 176.420 ;
        RECT 61.575 176.345 62.785 176.865 ;
        RECT 62.955 176.515 64.165 177.035 ;
        RECT 61.575 175.255 64.165 176.345 ;
        RECT 65.930 175.690 66.280 176.940 ;
        RECT 67.760 176.430 68.100 177.260 ;
        RECT 70.625 177.235 70.825 177.590 ;
        RECT 70.995 177.405 71.325 177.805 ;
        RECT 71.495 177.235 71.695 177.580 ;
        RECT 69.855 177.065 71.695 177.235 ;
        RECT 71.865 177.065 72.195 177.805 ;
        RECT 72.430 177.235 72.600 177.485 ;
        RECT 72.430 177.065 72.905 177.235 ;
        RECT 64.340 175.255 69.685 175.690 ;
        RECT 69.855 175.440 70.115 177.065 ;
        RECT 70.295 176.095 70.515 176.895 ;
        RECT 70.755 176.275 71.055 176.895 ;
        RECT 71.225 176.275 71.555 176.895 ;
        RECT 71.725 176.275 72.045 176.895 ;
        RECT 72.215 176.275 72.565 176.895 ;
        RECT 72.735 176.095 72.905 177.065 ;
        RECT 73.075 177.055 74.285 177.805 ;
        RECT 70.295 175.885 72.905 176.095 ;
        RECT 73.075 176.345 73.595 176.885 ;
        RECT 73.765 176.515 74.285 177.055 ;
        RECT 74.545 177.155 74.715 177.635 ;
        RECT 74.895 177.325 75.135 177.805 ;
        RECT 75.385 177.155 75.555 177.635 ;
        RECT 75.725 177.325 76.055 177.805 ;
        RECT 76.225 177.155 76.395 177.635 ;
        RECT 74.545 176.985 75.180 177.155 ;
        RECT 75.385 176.985 76.395 177.155 ;
        RECT 76.565 177.005 76.895 177.805 ;
        RECT 77.490 176.995 77.735 177.600 ;
        RECT 77.955 177.270 78.465 177.805 ;
        RECT 75.010 176.815 75.180 176.985 ;
        RECT 74.460 176.575 74.840 176.815 ;
        RECT 75.010 176.645 75.510 176.815 ;
        RECT 75.010 176.405 75.180 176.645 ;
        RECT 75.900 176.445 76.395 176.985 ;
        RECT 71.865 175.255 72.195 175.705 ;
        RECT 73.075 175.255 74.285 176.345 ;
        RECT 74.465 176.235 75.180 176.405 ;
        RECT 75.385 176.275 76.395 176.445 ;
        RECT 77.215 176.825 78.445 176.995 ;
        RECT 74.465 175.425 74.795 176.235 ;
        RECT 74.965 175.255 75.205 176.055 ;
        RECT 75.385 175.425 75.555 176.275 ;
        RECT 75.725 175.255 76.055 176.055 ;
        RECT 76.225 175.425 76.395 176.275 ;
        RECT 76.565 175.255 76.895 176.405 ;
        RECT 77.215 176.015 77.555 176.825 ;
        RECT 77.725 176.260 78.475 176.450 ;
        RECT 77.215 175.605 77.730 176.015 ;
        RECT 77.965 175.255 78.135 176.015 ;
        RECT 78.305 175.595 78.475 176.260 ;
        RECT 78.645 176.275 78.835 177.635 ;
        RECT 79.005 176.785 79.280 177.635 ;
        RECT 79.470 177.270 80.000 177.635 ;
        RECT 80.425 177.405 80.755 177.805 ;
        RECT 79.825 177.235 80.000 177.270 ;
        RECT 79.005 176.615 79.285 176.785 ;
        RECT 79.005 176.475 79.280 176.615 ;
        RECT 79.485 176.275 79.655 177.075 ;
        RECT 78.645 176.105 79.655 176.275 ;
        RECT 79.825 177.065 80.755 177.235 ;
        RECT 80.925 177.065 81.180 177.635 ;
        RECT 79.825 175.935 79.995 177.065 ;
        RECT 80.585 176.895 80.755 177.065 ;
        RECT 78.870 175.765 79.995 175.935 ;
        RECT 80.165 176.565 80.360 176.895 ;
        RECT 80.585 176.565 80.840 176.895 ;
        RECT 80.165 175.595 80.335 176.565 ;
        RECT 81.010 176.395 81.180 177.065 ;
        RECT 81.630 176.995 81.875 177.600 ;
        RECT 82.095 177.270 82.605 177.805 ;
        RECT 78.305 175.425 80.335 175.595 ;
        RECT 80.505 175.255 80.675 176.395 ;
        RECT 80.845 175.425 81.180 176.395 ;
        RECT 81.355 176.825 82.585 176.995 ;
        RECT 81.355 176.015 81.695 176.825 ;
        RECT 81.865 176.260 82.615 176.450 ;
        RECT 81.355 175.605 81.870 176.015 ;
        RECT 82.105 175.255 82.275 176.015 ;
        RECT 82.445 175.595 82.615 176.260 ;
        RECT 82.785 176.275 82.975 177.635 ;
        RECT 83.145 177.125 83.420 177.635 ;
        RECT 83.610 177.270 84.140 177.635 ;
        RECT 84.565 177.405 84.895 177.805 ;
        RECT 83.965 177.235 84.140 177.270 ;
        RECT 83.145 176.955 83.425 177.125 ;
        RECT 83.145 176.475 83.420 176.955 ;
        RECT 83.625 176.275 83.795 177.075 ;
        RECT 82.785 176.105 83.795 176.275 ;
        RECT 83.965 177.065 84.895 177.235 ;
        RECT 85.065 177.065 85.320 177.635 ;
        RECT 85.585 177.255 85.755 177.635 ;
        RECT 85.935 177.425 86.265 177.805 ;
        RECT 85.585 177.085 86.250 177.255 ;
        RECT 86.445 177.130 86.705 177.635 ;
        RECT 83.965 175.935 84.135 177.065 ;
        RECT 84.725 176.895 84.895 177.065 ;
        RECT 83.010 175.765 84.135 175.935 ;
        RECT 84.305 176.565 84.500 176.895 ;
        RECT 84.725 176.565 84.980 176.895 ;
        RECT 84.305 175.595 84.475 176.565 ;
        RECT 85.150 176.395 85.320 177.065 ;
        RECT 85.515 176.535 85.845 176.905 ;
        RECT 86.080 176.830 86.250 177.085 ;
        RECT 82.445 175.425 84.475 175.595 ;
        RECT 84.645 175.255 84.815 176.395 ;
        RECT 84.985 175.425 85.320 176.395 ;
        RECT 86.080 176.500 86.365 176.830 ;
        RECT 86.080 176.355 86.250 176.500 ;
        RECT 85.585 176.185 86.250 176.355 ;
        RECT 86.535 176.330 86.705 177.130 ;
        RECT 86.875 177.080 87.165 177.805 ;
        RECT 87.335 177.055 88.545 177.805 ;
        RECT 85.585 175.425 85.755 176.185 ;
        RECT 85.935 175.255 86.265 176.015 ;
        RECT 86.435 175.425 86.705 176.330 ;
        RECT 86.875 175.255 87.165 176.420 ;
        RECT 87.335 176.345 87.855 176.885 ;
        RECT 88.025 176.515 88.545 177.055 ;
        RECT 88.755 176.985 88.985 177.805 ;
        RECT 89.155 177.005 89.485 177.635 ;
        RECT 88.735 176.565 89.065 176.815 ;
        RECT 89.235 176.405 89.485 177.005 ;
        RECT 89.655 176.985 89.865 177.805 ;
        RECT 90.100 177.095 90.355 177.625 ;
        RECT 90.525 177.345 90.830 177.805 ;
        RECT 91.075 177.425 92.145 177.595 ;
        RECT 87.335 175.255 88.545 176.345 ;
        RECT 88.755 175.255 88.985 176.395 ;
        RECT 89.155 175.425 89.485 176.405 ;
        RECT 90.100 176.445 90.310 177.095 ;
        RECT 91.075 177.070 91.395 177.425 ;
        RECT 91.070 176.895 91.395 177.070 ;
        RECT 90.480 176.595 91.395 176.895 ;
        RECT 91.565 176.855 91.805 177.255 ;
        RECT 91.975 177.195 92.145 177.425 ;
        RECT 92.315 177.365 92.505 177.805 ;
        RECT 92.675 177.355 93.625 177.635 ;
        RECT 93.845 177.445 94.195 177.615 ;
        RECT 91.975 177.025 92.505 177.195 ;
        RECT 90.480 176.565 91.220 176.595 ;
        RECT 89.655 175.255 89.865 176.395 ;
        RECT 90.100 175.565 90.355 176.445 ;
        RECT 90.525 175.255 90.830 176.395 ;
        RECT 91.050 175.975 91.220 176.565 ;
        RECT 91.565 176.485 92.105 176.855 ;
        RECT 92.285 176.745 92.505 177.025 ;
        RECT 92.675 176.575 92.845 177.355 ;
        RECT 92.440 176.405 92.845 176.575 ;
        RECT 93.015 176.565 93.365 177.185 ;
        RECT 92.440 176.315 92.610 176.405 ;
        RECT 93.535 176.395 93.745 177.185 ;
        RECT 91.390 176.145 92.610 176.315 ;
        RECT 93.070 176.235 93.745 176.395 ;
        RECT 91.050 175.805 91.850 175.975 ;
        RECT 91.170 175.255 91.500 175.635 ;
        RECT 91.680 175.515 91.850 175.805 ;
        RECT 92.440 175.765 92.610 176.145 ;
        RECT 92.780 176.225 93.745 176.235 ;
        RECT 93.935 177.055 94.195 177.445 ;
        RECT 94.405 177.345 94.735 177.805 ;
        RECT 95.610 177.415 96.465 177.585 ;
        RECT 96.670 177.415 97.165 177.585 ;
        RECT 97.335 177.445 97.665 177.805 ;
        RECT 93.935 176.365 94.105 177.055 ;
        RECT 94.275 176.705 94.445 176.885 ;
        RECT 94.615 176.875 95.405 177.125 ;
        RECT 95.610 176.705 95.780 177.415 ;
        RECT 95.950 176.905 96.305 177.125 ;
        RECT 94.275 176.535 95.965 176.705 ;
        RECT 92.780 175.935 93.240 176.225 ;
        RECT 93.935 176.195 95.435 176.365 ;
        RECT 93.935 176.055 94.105 176.195 ;
        RECT 93.545 175.885 94.105 176.055 ;
        RECT 92.020 175.255 92.270 175.715 ;
        RECT 92.440 175.425 93.310 175.765 ;
        RECT 93.545 175.425 93.715 175.885 ;
        RECT 94.550 175.855 95.625 176.025 ;
        RECT 93.885 175.255 94.255 175.715 ;
        RECT 94.550 175.515 94.720 175.855 ;
        RECT 94.890 175.255 95.220 175.685 ;
        RECT 95.455 175.515 95.625 175.855 ;
        RECT 95.795 175.755 95.965 176.535 ;
        RECT 96.135 176.315 96.305 176.905 ;
        RECT 96.475 176.505 96.825 177.125 ;
        RECT 96.135 175.925 96.600 176.315 ;
        RECT 96.995 176.055 97.165 177.415 ;
        RECT 97.335 176.225 97.795 177.275 ;
        RECT 96.770 175.885 97.165 176.055 ;
        RECT 96.770 175.755 96.940 175.885 ;
        RECT 95.795 175.425 96.475 175.755 ;
        RECT 96.690 175.425 96.940 175.755 ;
        RECT 97.110 175.255 97.360 175.715 ;
        RECT 97.530 175.440 97.855 176.225 ;
        RECT 98.025 175.425 98.195 177.545 ;
        RECT 98.365 177.425 98.695 177.805 ;
        RECT 98.865 177.255 99.120 177.545 ;
        RECT 98.370 177.085 99.120 177.255 ;
        RECT 98.370 176.095 98.600 177.085 ;
        RECT 99.570 176.995 99.815 177.600 ;
        RECT 100.035 177.270 100.545 177.805 ;
        RECT 98.770 176.265 99.120 176.915 ;
        RECT 99.295 176.825 100.525 176.995 ;
        RECT 98.370 175.925 99.120 176.095 ;
        RECT 98.365 175.255 98.695 175.755 ;
        RECT 98.865 175.425 99.120 175.925 ;
        RECT 99.295 176.015 99.635 176.825 ;
        RECT 99.805 176.260 100.555 176.450 ;
        RECT 99.295 175.605 99.810 176.015 ;
        RECT 100.045 175.255 100.215 176.015 ;
        RECT 100.385 175.595 100.555 176.260 ;
        RECT 100.725 176.275 100.915 177.635 ;
        RECT 101.085 177.125 101.360 177.635 ;
        RECT 101.550 177.270 102.080 177.635 ;
        RECT 102.505 177.405 102.835 177.805 ;
        RECT 101.905 177.235 102.080 177.270 ;
        RECT 101.085 176.955 101.365 177.125 ;
        RECT 101.085 176.475 101.360 176.955 ;
        RECT 101.565 176.275 101.735 177.075 ;
        RECT 100.725 176.105 101.735 176.275 ;
        RECT 101.905 177.065 102.835 177.235 ;
        RECT 103.005 177.065 103.260 177.635 ;
        RECT 101.905 175.935 102.075 177.065 ;
        RECT 102.665 176.895 102.835 177.065 ;
        RECT 100.950 175.765 102.075 175.935 ;
        RECT 102.245 176.565 102.440 176.895 ;
        RECT 102.665 176.565 102.920 176.895 ;
        RECT 102.245 175.595 102.415 176.565 ;
        RECT 103.090 176.395 103.260 177.065 ;
        RECT 100.385 175.425 102.415 175.595 ;
        RECT 102.585 175.255 102.755 176.395 ;
        RECT 102.925 175.425 103.260 176.395 ;
        RECT 103.435 177.065 103.820 177.635 ;
        RECT 103.990 177.345 104.315 177.805 ;
        RECT 104.835 177.175 105.115 177.635 ;
        RECT 103.435 176.395 103.715 177.065 ;
        RECT 103.990 177.005 105.115 177.175 ;
        RECT 103.990 176.895 104.440 177.005 ;
        RECT 103.885 176.565 104.440 176.895 ;
        RECT 105.305 176.835 105.705 177.635 ;
        RECT 106.105 177.345 106.375 177.805 ;
        RECT 106.545 177.175 106.830 177.635 ;
        RECT 103.435 175.425 103.820 176.395 ;
        RECT 103.990 176.105 104.440 176.565 ;
        RECT 104.610 176.275 105.705 176.835 ;
        RECT 103.990 175.885 105.115 176.105 ;
        RECT 103.990 175.255 104.315 175.715 ;
        RECT 104.835 175.425 105.115 175.885 ;
        RECT 105.305 175.425 105.705 176.275 ;
        RECT 105.875 177.005 106.830 177.175 ;
        RECT 107.115 177.055 108.325 177.805 ;
        RECT 108.585 177.255 108.755 177.635 ;
        RECT 108.935 177.425 109.265 177.805 ;
        RECT 108.585 177.085 109.250 177.255 ;
        RECT 109.445 177.130 109.705 177.635 ;
        RECT 105.875 176.105 106.085 177.005 ;
        RECT 106.255 176.275 106.945 176.835 ;
        RECT 107.115 176.345 107.635 176.885 ;
        RECT 107.805 176.515 108.325 177.055 ;
        RECT 108.515 176.535 108.845 176.905 ;
        RECT 109.080 176.830 109.250 177.085 ;
        RECT 109.080 176.500 109.365 176.830 ;
        RECT 109.080 176.355 109.250 176.500 ;
        RECT 105.875 175.885 106.830 176.105 ;
        RECT 106.105 175.255 106.375 175.715 ;
        RECT 106.545 175.425 106.830 175.885 ;
        RECT 107.115 175.255 108.325 176.345 ;
        RECT 108.585 176.185 109.250 176.355 ;
        RECT 109.535 176.330 109.705 177.130 ;
        RECT 109.875 177.055 111.085 177.805 ;
        RECT 108.585 175.425 108.755 176.185 ;
        RECT 108.935 175.255 109.265 176.015 ;
        RECT 109.435 175.425 109.705 176.330 ;
        RECT 109.875 176.345 110.395 176.885 ;
        RECT 110.565 176.515 111.085 177.055 ;
        RECT 111.295 176.985 111.525 177.805 ;
        RECT 111.695 177.005 112.025 177.635 ;
        RECT 111.275 176.565 111.605 176.815 ;
        RECT 111.775 176.405 112.025 177.005 ;
        RECT 112.195 176.985 112.405 177.805 ;
        RECT 112.635 177.080 112.925 177.805 ;
        RECT 114.020 177.095 114.275 177.625 ;
        RECT 114.445 177.345 114.750 177.805 ;
        RECT 114.995 177.425 116.065 177.595 ;
        RECT 114.020 176.445 114.230 177.095 ;
        RECT 114.995 177.070 115.315 177.425 ;
        RECT 114.990 176.895 115.315 177.070 ;
        RECT 114.400 176.595 115.315 176.895 ;
        RECT 115.485 176.855 115.725 177.255 ;
        RECT 115.895 177.195 116.065 177.425 ;
        RECT 116.235 177.365 116.425 177.805 ;
        RECT 116.595 177.355 117.545 177.635 ;
        RECT 117.765 177.445 118.115 177.615 ;
        RECT 115.895 177.025 116.425 177.195 ;
        RECT 114.400 176.565 115.140 176.595 ;
        RECT 109.875 175.255 111.085 176.345 ;
        RECT 111.295 175.255 111.525 176.395 ;
        RECT 111.695 175.425 112.025 176.405 ;
        RECT 112.195 175.255 112.405 176.395 ;
        RECT 112.635 175.255 112.925 176.420 ;
        RECT 114.020 175.565 114.275 176.445 ;
        RECT 114.445 175.255 114.750 176.395 ;
        RECT 114.970 175.975 115.140 176.565 ;
        RECT 115.485 176.485 116.025 176.855 ;
        RECT 116.205 176.745 116.425 177.025 ;
        RECT 116.595 176.575 116.765 177.355 ;
        RECT 116.360 176.405 116.765 176.575 ;
        RECT 116.935 176.565 117.285 177.185 ;
        RECT 116.360 176.315 116.530 176.405 ;
        RECT 117.455 176.395 117.665 177.185 ;
        RECT 115.310 176.145 116.530 176.315 ;
        RECT 116.990 176.235 117.665 176.395 ;
        RECT 114.970 175.805 115.770 175.975 ;
        RECT 115.090 175.255 115.420 175.635 ;
        RECT 115.600 175.515 115.770 175.805 ;
        RECT 116.360 175.765 116.530 176.145 ;
        RECT 116.700 176.225 117.665 176.235 ;
        RECT 117.855 177.055 118.115 177.445 ;
        RECT 118.325 177.345 118.655 177.805 ;
        RECT 119.530 177.415 120.385 177.585 ;
        RECT 120.590 177.415 121.085 177.585 ;
        RECT 121.255 177.445 121.585 177.805 ;
        RECT 117.855 176.365 118.025 177.055 ;
        RECT 118.195 176.705 118.365 176.885 ;
        RECT 118.535 176.875 119.325 177.125 ;
        RECT 119.530 176.705 119.700 177.415 ;
        RECT 119.870 176.905 120.225 177.125 ;
        RECT 118.195 176.535 119.885 176.705 ;
        RECT 116.700 175.935 117.160 176.225 ;
        RECT 117.855 176.195 119.355 176.365 ;
        RECT 117.855 176.055 118.025 176.195 ;
        RECT 117.465 175.885 118.025 176.055 ;
        RECT 115.940 175.255 116.190 175.715 ;
        RECT 116.360 175.425 117.230 175.765 ;
        RECT 117.465 175.425 117.635 175.885 ;
        RECT 118.470 175.855 119.545 176.025 ;
        RECT 117.805 175.255 118.175 175.715 ;
        RECT 118.470 175.515 118.640 175.855 ;
        RECT 118.810 175.255 119.140 175.685 ;
        RECT 119.375 175.515 119.545 175.855 ;
        RECT 119.715 175.755 119.885 176.535 ;
        RECT 120.055 176.315 120.225 176.905 ;
        RECT 120.395 176.505 120.745 177.125 ;
        RECT 120.055 175.925 120.520 176.315 ;
        RECT 120.915 176.055 121.085 177.415 ;
        RECT 121.255 176.225 121.715 177.275 ;
        RECT 120.690 175.885 121.085 176.055 ;
        RECT 120.690 175.755 120.860 175.885 ;
        RECT 119.715 175.425 120.395 175.755 ;
        RECT 120.610 175.425 120.860 175.755 ;
        RECT 121.030 175.255 121.280 175.715 ;
        RECT 121.450 175.440 121.775 176.225 ;
        RECT 121.945 175.425 122.115 177.545 ;
        RECT 122.285 177.425 122.615 177.805 ;
        RECT 122.785 177.255 123.040 177.545 ;
        RECT 122.290 177.085 123.040 177.255 ;
        RECT 122.290 176.095 122.520 177.085 ;
        RECT 123.215 177.055 124.425 177.805 ;
        RECT 124.595 177.055 125.805 177.805 ;
        RECT 122.690 176.265 123.040 176.915 ;
        RECT 123.215 176.345 123.735 176.885 ;
        RECT 123.905 176.515 124.425 177.055 ;
        RECT 124.595 176.345 125.115 176.885 ;
        RECT 125.285 176.515 125.805 177.055 ;
        RECT 122.290 175.925 123.040 176.095 ;
        RECT 122.285 175.255 122.615 175.755 ;
        RECT 122.785 175.425 123.040 175.925 ;
        RECT 123.215 175.255 124.425 176.345 ;
        RECT 124.595 175.255 125.805 176.345 ;
        RECT 11.810 175.085 125.890 175.255 ;
        RECT 11.895 173.995 13.105 175.085 ;
        RECT 11.895 173.285 12.415 173.825 ;
        RECT 12.585 173.455 13.105 173.995 ;
        RECT 13.275 173.995 16.785 175.085 ;
        RECT 16.960 174.650 22.305 175.085 ;
        RECT 13.275 173.475 14.965 173.995 ;
        RECT 15.135 173.305 16.785 173.825 ;
        RECT 18.550 173.400 18.900 174.650 ;
        RECT 22.475 173.920 22.765 175.085 ;
        RECT 23.895 173.945 24.125 175.085 ;
        RECT 24.295 173.935 24.625 174.915 ;
        RECT 24.795 173.945 25.005 175.085 ;
        RECT 25.275 173.945 25.505 175.085 ;
        RECT 25.675 173.935 26.005 174.915 ;
        RECT 26.175 173.945 26.385 175.085 ;
        RECT 26.705 174.155 26.875 174.915 ;
        RECT 27.055 174.325 27.385 175.085 ;
        RECT 26.705 173.985 27.370 174.155 ;
        RECT 27.555 174.010 27.825 174.915 ;
        RECT 11.895 172.535 13.105 173.285 ;
        RECT 13.275 172.535 16.785 173.305 ;
        RECT 20.380 173.080 20.720 173.910 ;
        RECT 23.875 173.525 24.205 173.775 ;
        RECT 16.960 172.535 22.305 173.080 ;
        RECT 22.475 172.535 22.765 173.260 ;
        RECT 23.895 172.535 24.125 173.355 ;
        RECT 24.375 173.335 24.625 173.935 ;
        RECT 25.255 173.525 25.585 173.775 ;
        RECT 24.295 172.705 24.625 173.335 ;
        RECT 24.795 172.535 25.005 173.355 ;
        RECT 25.275 172.535 25.505 173.355 ;
        RECT 25.755 173.335 26.005 173.935 ;
        RECT 27.200 173.840 27.370 173.985 ;
        RECT 26.635 173.435 26.965 173.805 ;
        RECT 27.200 173.510 27.485 173.840 ;
        RECT 25.675 172.705 26.005 173.335 ;
        RECT 26.175 172.535 26.385 173.355 ;
        RECT 27.200 173.255 27.370 173.510 ;
        RECT 26.705 173.085 27.370 173.255 ;
        RECT 27.655 173.210 27.825 174.010 ;
        RECT 26.705 172.705 26.875 173.085 ;
        RECT 27.055 172.535 27.385 172.915 ;
        RECT 27.565 172.705 27.825 173.210 ;
        RECT 28.000 173.895 28.255 174.775 ;
        RECT 28.425 173.945 28.730 175.085 ;
        RECT 29.070 174.705 29.400 175.085 ;
        RECT 29.580 174.535 29.750 174.825 ;
        RECT 29.920 174.625 30.170 175.085 ;
        RECT 28.950 174.365 29.750 174.535 ;
        RECT 30.340 174.575 31.210 174.915 ;
        RECT 28.000 173.245 28.210 173.895 ;
        RECT 28.950 173.775 29.120 174.365 ;
        RECT 30.340 174.195 30.510 174.575 ;
        RECT 31.445 174.455 31.615 174.915 ;
        RECT 31.785 174.625 32.155 175.085 ;
        RECT 32.450 174.485 32.620 174.825 ;
        RECT 32.790 174.655 33.120 175.085 ;
        RECT 33.355 174.485 33.525 174.825 ;
        RECT 29.290 174.025 30.510 174.195 ;
        RECT 30.680 174.115 31.140 174.405 ;
        RECT 31.445 174.285 32.005 174.455 ;
        RECT 32.450 174.315 33.525 174.485 ;
        RECT 33.695 174.585 34.375 174.915 ;
        RECT 34.590 174.585 34.840 174.915 ;
        RECT 35.010 174.625 35.260 175.085 ;
        RECT 31.835 174.145 32.005 174.285 ;
        RECT 30.680 174.105 31.645 174.115 ;
        RECT 30.340 173.935 30.510 174.025 ;
        RECT 30.970 173.945 31.645 174.105 ;
        RECT 28.380 173.745 29.120 173.775 ;
        RECT 28.380 173.445 29.295 173.745 ;
        RECT 28.970 173.270 29.295 173.445 ;
        RECT 28.000 172.715 28.255 173.245 ;
        RECT 28.425 172.535 28.730 172.995 ;
        RECT 28.975 172.915 29.295 173.270 ;
        RECT 29.465 173.485 30.005 173.855 ;
        RECT 30.340 173.765 30.745 173.935 ;
        RECT 29.465 173.085 29.705 173.485 ;
        RECT 30.185 173.315 30.405 173.595 ;
        RECT 29.875 173.145 30.405 173.315 ;
        RECT 29.875 172.915 30.045 173.145 ;
        RECT 30.575 172.985 30.745 173.765 ;
        RECT 30.915 173.155 31.265 173.775 ;
        RECT 31.435 173.155 31.645 173.945 ;
        RECT 31.835 173.975 33.335 174.145 ;
        RECT 31.835 173.285 32.005 173.975 ;
        RECT 33.695 173.805 33.865 174.585 ;
        RECT 34.670 174.455 34.840 174.585 ;
        RECT 32.175 173.635 33.865 173.805 ;
        RECT 34.035 174.025 34.500 174.415 ;
        RECT 34.670 174.285 35.065 174.455 ;
        RECT 32.175 173.455 32.345 173.635 ;
        RECT 28.975 172.745 30.045 172.915 ;
        RECT 30.215 172.535 30.405 172.975 ;
        RECT 30.575 172.705 31.525 172.985 ;
        RECT 31.835 172.895 32.095 173.285 ;
        RECT 32.515 173.215 33.305 173.465 ;
        RECT 31.745 172.725 32.095 172.895 ;
        RECT 32.305 172.535 32.635 172.995 ;
        RECT 33.510 172.925 33.680 173.635 ;
        RECT 34.035 173.435 34.205 174.025 ;
        RECT 33.850 173.215 34.205 173.435 ;
        RECT 34.375 173.215 34.725 173.835 ;
        RECT 34.895 172.925 35.065 174.285 ;
        RECT 35.430 174.115 35.755 174.900 ;
        RECT 35.235 173.065 35.695 174.115 ;
        RECT 33.510 172.755 34.365 172.925 ;
        RECT 34.570 172.755 35.065 172.925 ;
        RECT 35.235 172.535 35.565 172.895 ;
        RECT 35.925 172.795 36.095 174.915 ;
        RECT 36.265 174.585 36.595 175.085 ;
        RECT 36.765 174.415 37.020 174.915 ;
        RECT 36.270 174.245 37.020 174.415 ;
        RECT 36.270 173.255 36.500 174.245 ;
        RECT 36.670 173.425 37.020 174.075 ;
        RECT 37.195 174.010 37.465 174.915 ;
        RECT 37.635 174.325 37.965 175.085 ;
        RECT 38.145 174.155 38.315 174.915 ;
        RECT 36.270 173.085 37.020 173.255 ;
        RECT 36.265 172.535 36.595 172.915 ;
        RECT 36.765 172.795 37.020 173.085 ;
        RECT 37.195 173.210 37.365 174.010 ;
        RECT 37.650 173.985 38.315 174.155 ;
        RECT 38.575 173.995 40.245 175.085 ;
        RECT 40.420 174.650 45.765 175.085 ;
        RECT 37.650 173.840 37.820 173.985 ;
        RECT 37.535 173.510 37.820 173.840 ;
        RECT 37.650 173.255 37.820 173.510 ;
        RECT 38.055 173.435 38.385 173.805 ;
        RECT 38.575 173.475 39.325 173.995 ;
        RECT 39.495 173.305 40.245 173.825 ;
        RECT 42.010 173.400 42.360 174.650 ;
        RECT 46.025 174.155 46.195 174.915 ;
        RECT 46.375 174.325 46.705 175.085 ;
        RECT 46.025 173.985 46.690 174.155 ;
        RECT 46.875 174.010 47.145 174.915 ;
        RECT 37.195 172.705 37.455 173.210 ;
        RECT 37.650 173.085 38.315 173.255 ;
        RECT 37.635 172.535 37.965 172.915 ;
        RECT 38.145 172.705 38.315 173.085 ;
        RECT 38.575 172.535 40.245 173.305 ;
        RECT 43.840 173.080 44.180 173.910 ;
        RECT 46.520 173.840 46.690 173.985 ;
        RECT 45.955 173.435 46.285 173.805 ;
        RECT 46.520 173.510 46.805 173.840 ;
        RECT 46.520 173.255 46.690 173.510 ;
        RECT 46.025 173.085 46.690 173.255 ;
        RECT 46.975 173.210 47.145 174.010 ;
        RECT 48.235 173.920 48.525 175.085 ;
        RECT 48.695 173.995 50.365 175.085 ;
        RECT 48.695 173.475 49.445 173.995 ;
        RECT 50.595 173.945 50.805 175.085 ;
        RECT 50.975 173.935 51.305 174.915 ;
        RECT 51.475 173.945 51.705 175.085 ;
        RECT 52.290 174.105 52.545 174.775 ;
        RECT 52.725 174.285 53.010 175.085 ;
        RECT 53.190 174.365 53.520 174.875 ;
        RECT 49.615 173.305 50.365 173.825 ;
        RECT 40.420 172.535 45.765 173.080 ;
        RECT 46.025 172.705 46.195 173.085 ;
        RECT 46.375 172.535 46.705 172.915 ;
        RECT 46.885 172.705 47.145 173.210 ;
        RECT 48.235 172.535 48.525 173.260 ;
        RECT 48.695 172.535 50.365 173.305 ;
        RECT 50.595 172.535 50.805 173.355 ;
        RECT 50.975 173.335 51.225 173.935 ;
        RECT 51.395 173.525 51.725 173.775 ;
        RECT 50.975 172.705 51.305 173.335 ;
        RECT 51.475 172.535 51.705 173.355 ;
        RECT 52.290 173.245 52.470 174.105 ;
        RECT 53.190 173.775 53.440 174.365 ;
        RECT 53.790 174.215 53.960 174.825 ;
        RECT 54.130 174.395 54.460 175.085 ;
        RECT 54.690 174.535 54.930 174.825 ;
        RECT 55.130 174.705 55.550 175.085 ;
        RECT 55.730 174.615 56.360 174.865 ;
        RECT 56.830 174.705 57.160 175.085 ;
        RECT 55.730 174.535 55.900 174.615 ;
        RECT 57.330 174.535 57.500 174.825 ;
        RECT 57.680 174.705 58.060 175.085 ;
        RECT 58.300 174.700 59.130 174.870 ;
        RECT 54.690 174.365 55.900 174.535 ;
        RECT 52.640 173.445 53.440 173.775 ;
        RECT 52.290 173.045 52.545 173.245 ;
        RECT 52.205 172.875 52.545 173.045 ;
        RECT 52.290 172.715 52.545 172.875 ;
        RECT 52.725 172.535 53.010 172.995 ;
        RECT 53.190 172.795 53.440 173.445 ;
        RECT 53.640 174.195 53.960 174.215 ;
        RECT 53.640 174.025 55.560 174.195 ;
        RECT 53.640 173.130 53.830 174.025 ;
        RECT 55.730 173.855 55.900 174.365 ;
        RECT 56.070 174.105 56.590 174.415 ;
        RECT 54.000 173.685 55.900 173.855 ;
        RECT 54.000 173.625 54.330 173.685 ;
        RECT 54.480 173.455 54.810 173.515 ;
        RECT 54.150 173.185 54.810 173.455 ;
        RECT 53.640 172.800 53.960 173.130 ;
        RECT 54.140 172.535 54.800 173.015 ;
        RECT 55.000 172.925 55.170 173.685 ;
        RECT 56.070 173.515 56.250 173.925 ;
        RECT 55.340 173.345 55.670 173.465 ;
        RECT 56.420 173.345 56.590 174.105 ;
        RECT 55.340 173.175 56.590 173.345 ;
        RECT 56.760 174.285 58.130 174.535 ;
        RECT 56.760 173.515 56.950 174.285 ;
        RECT 57.880 174.025 58.130 174.285 ;
        RECT 57.120 173.855 57.370 174.015 ;
        RECT 58.300 173.855 58.470 174.700 ;
        RECT 59.365 174.415 59.535 174.915 ;
        RECT 59.705 174.585 60.035 175.085 ;
        RECT 58.640 174.025 59.140 174.405 ;
        RECT 59.365 174.245 60.060 174.415 ;
        RECT 57.120 173.685 58.470 173.855 ;
        RECT 58.050 173.645 58.470 173.685 ;
        RECT 56.760 173.175 57.180 173.515 ;
        RECT 57.470 173.185 57.880 173.515 ;
        RECT 55.000 172.755 55.850 172.925 ;
        RECT 56.410 172.535 56.730 172.995 ;
        RECT 56.930 172.745 57.180 173.175 ;
        RECT 57.470 172.535 57.880 172.975 ;
        RECT 58.050 172.915 58.220 173.645 ;
        RECT 58.390 173.095 58.740 173.465 ;
        RECT 58.920 173.155 59.140 174.025 ;
        RECT 59.310 173.455 59.720 174.075 ;
        RECT 59.890 173.275 60.060 174.245 ;
        RECT 59.365 173.085 60.060 173.275 ;
        RECT 58.050 172.715 59.065 172.915 ;
        RECT 59.365 172.755 59.535 173.085 ;
        RECT 59.705 172.535 60.035 172.915 ;
        RECT 60.250 172.795 60.475 174.915 ;
        RECT 60.645 174.585 60.975 175.085 ;
        RECT 61.145 174.415 61.315 174.915 ;
        RECT 60.650 174.245 61.315 174.415 ;
        RECT 60.650 173.255 60.880 174.245 ;
        RECT 61.050 173.425 61.400 174.075 ;
        RECT 62.495 173.995 66.005 175.085 ;
        RECT 62.495 173.475 64.185 173.995 ;
        RECT 64.355 173.305 66.005 173.825 ;
        RECT 60.650 173.085 61.315 173.255 ;
        RECT 60.645 172.535 60.975 172.915 ;
        RECT 61.145 172.795 61.315 173.085 ;
        RECT 62.495 172.535 66.005 173.305 ;
        RECT 66.175 173.275 66.435 174.900 ;
        RECT 68.185 174.635 68.515 175.085 ;
        RECT 69.395 174.585 69.655 174.915 ;
        RECT 69.965 174.705 70.295 175.085 ;
        RECT 66.615 174.245 69.225 174.455 ;
        RECT 66.615 173.445 66.835 174.245 ;
        RECT 67.075 173.445 67.375 174.065 ;
        RECT 67.545 173.445 67.875 174.065 ;
        RECT 68.045 173.445 68.365 174.065 ;
        RECT 68.535 173.445 68.885 174.065 ;
        RECT 69.055 173.275 69.225 174.245 ;
        RECT 66.175 173.105 68.015 173.275 ;
        RECT 66.445 172.535 66.775 172.930 ;
        RECT 66.945 172.750 67.145 173.105 ;
        RECT 67.315 172.535 67.645 172.935 ;
        RECT 67.815 172.760 68.015 173.105 ;
        RECT 68.185 172.535 68.515 173.275 ;
        RECT 68.750 173.105 69.225 173.275 ;
        RECT 69.395 173.905 69.565 174.585 ;
        RECT 70.535 174.535 70.725 174.915 ;
        RECT 70.975 174.705 71.305 175.085 ;
        RECT 71.515 174.535 71.685 174.915 ;
        RECT 71.880 174.705 72.210 175.085 ;
        RECT 72.470 174.535 72.640 174.915 ;
        RECT 73.065 174.705 73.395 175.085 ;
        RECT 69.735 174.075 70.085 174.405 ;
        RECT 70.535 174.365 71.275 174.535 ;
        RECT 70.355 174.025 70.935 174.195 ;
        RECT 70.355 173.905 70.525 174.025 ;
        RECT 69.395 173.735 70.525 173.905 ;
        RECT 71.105 173.855 71.275 174.365 ;
        RECT 68.750 172.855 68.920 173.105 ;
        RECT 69.395 173.035 69.565 173.735 ;
        RECT 70.705 173.685 71.275 173.855 ;
        RECT 71.445 174.365 73.395 174.535 ;
        RECT 69.915 173.395 70.535 173.565 ;
        RECT 69.915 173.215 70.125 173.395 ;
        RECT 70.705 173.205 70.875 173.685 ;
        RECT 71.445 173.375 71.615 174.365 ;
        RECT 72.205 173.775 72.390 174.085 ;
        RECT 72.660 173.775 72.855 174.085 ;
        RECT 69.395 172.705 69.655 173.035 ;
        RECT 69.965 172.535 70.295 172.915 ;
        RECT 70.475 172.875 70.875 173.205 ;
        RECT 71.065 173.045 71.615 173.375 ;
        RECT 71.785 172.875 71.955 173.775 ;
        RECT 70.475 172.705 71.955 172.875 ;
        RECT 72.205 173.445 72.435 173.775 ;
        RECT 72.660 173.445 72.915 173.775 ;
        RECT 73.225 173.445 73.395 174.365 ;
        RECT 72.205 172.865 72.390 173.445 ;
        RECT 72.660 172.870 72.855 173.445 ;
        RECT 73.065 172.535 73.395 172.915 ;
        RECT 73.565 172.705 73.825 174.915 ;
        RECT 73.995 173.920 74.285 175.085 ;
        RECT 74.455 173.275 74.715 174.900 ;
        RECT 76.465 174.635 76.795 175.085 ;
        RECT 74.895 174.245 77.505 174.455 ;
        RECT 74.895 173.445 75.115 174.245 ;
        RECT 75.355 173.445 75.655 174.065 ;
        RECT 75.825 173.445 76.155 174.065 ;
        RECT 76.325 173.445 76.645 174.065 ;
        RECT 76.815 173.445 77.165 174.065 ;
        RECT 77.335 173.275 77.505 174.245 ;
        RECT 78.175 173.945 78.405 175.085 ;
        RECT 78.575 173.935 78.905 174.915 ;
        RECT 79.075 173.945 79.285 175.085 ;
        RECT 78.155 173.525 78.485 173.775 ;
        RECT 73.995 172.535 74.285 173.260 ;
        RECT 74.455 173.105 76.295 173.275 ;
        RECT 74.725 172.535 75.055 172.930 ;
        RECT 75.225 172.750 75.425 173.105 ;
        RECT 75.595 172.535 75.925 172.935 ;
        RECT 76.095 172.760 76.295 173.105 ;
        RECT 76.465 172.535 76.795 173.275 ;
        RECT 77.030 173.105 77.505 173.275 ;
        RECT 77.030 172.855 77.200 173.105 ;
        RECT 78.175 172.535 78.405 173.355 ;
        RECT 78.655 173.335 78.905 173.935 ;
        RECT 79.520 173.895 79.775 174.775 ;
        RECT 79.945 173.945 80.250 175.085 ;
        RECT 80.590 174.705 80.920 175.085 ;
        RECT 81.100 174.535 81.270 174.825 ;
        RECT 81.440 174.625 81.690 175.085 ;
        RECT 80.470 174.365 81.270 174.535 ;
        RECT 81.860 174.575 82.730 174.915 ;
        RECT 78.575 172.705 78.905 173.335 ;
        RECT 79.075 172.535 79.285 173.355 ;
        RECT 79.520 173.245 79.730 173.895 ;
        RECT 80.470 173.775 80.640 174.365 ;
        RECT 81.860 174.195 82.030 174.575 ;
        RECT 82.965 174.455 83.135 174.915 ;
        RECT 83.305 174.625 83.675 175.085 ;
        RECT 83.970 174.485 84.140 174.825 ;
        RECT 84.310 174.655 84.640 175.085 ;
        RECT 84.875 174.485 85.045 174.825 ;
        RECT 80.810 174.025 82.030 174.195 ;
        RECT 82.200 174.115 82.660 174.405 ;
        RECT 82.965 174.285 83.525 174.455 ;
        RECT 83.970 174.315 85.045 174.485 ;
        RECT 85.215 174.585 85.895 174.915 ;
        RECT 86.110 174.585 86.360 174.915 ;
        RECT 86.530 174.625 86.780 175.085 ;
        RECT 83.355 174.145 83.525 174.285 ;
        RECT 82.200 174.105 83.165 174.115 ;
        RECT 81.860 173.935 82.030 174.025 ;
        RECT 82.490 173.945 83.165 174.105 ;
        RECT 79.900 173.745 80.640 173.775 ;
        RECT 79.900 173.445 80.815 173.745 ;
        RECT 80.490 173.270 80.815 173.445 ;
        RECT 79.520 172.715 79.775 173.245 ;
        RECT 79.945 172.535 80.250 172.995 ;
        RECT 80.495 172.915 80.815 173.270 ;
        RECT 80.985 173.485 81.525 173.855 ;
        RECT 81.860 173.765 82.265 173.935 ;
        RECT 80.985 173.085 81.225 173.485 ;
        RECT 81.705 173.315 81.925 173.595 ;
        RECT 81.395 173.145 81.925 173.315 ;
        RECT 81.395 172.915 81.565 173.145 ;
        RECT 82.095 172.985 82.265 173.765 ;
        RECT 82.435 173.155 82.785 173.775 ;
        RECT 82.955 173.155 83.165 173.945 ;
        RECT 83.355 173.975 84.855 174.145 ;
        RECT 83.355 173.285 83.525 173.975 ;
        RECT 85.215 173.805 85.385 174.585 ;
        RECT 86.190 174.455 86.360 174.585 ;
        RECT 83.695 173.635 85.385 173.805 ;
        RECT 85.555 174.025 86.020 174.415 ;
        RECT 86.190 174.285 86.585 174.455 ;
        RECT 83.695 173.455 83.865 173.635 ;
        RECT 80.495 172.745 81.565 172.915 ;
        RECT 81.735 172.535 81.925 172.975 ;
        RECT 82.095 172.705 83.045 172.985 ;
        RECT 83.355 172.895 83.615 173.285 ;
        RECT 84.035 173.215 84.825 173.465 ;
        RECT 83.265 172.725 83.615 172.895 ;
        RECT 83.825 172.535 84.155 172.995 ;
        RECT 85.030 172.925 85.200 173.635 ;
        RECT 85.555 173.435 85.725 174.025 ;
        RECT 85.370 173.215 85.725 173.435 ;
        RECT 85.895 173.215 86.245 173.835 ;
        RECT 86.415 172.925 86.585 174.285 ;
        RECT 86.950 174.115 87.275 174.900 ;
        RECT 86.755 173.065 87.215 174.115 ;
        RECT 85.030 172.755 85.885 172.925 ;
        RECT 86.090 172.755 86.585 172.925 ;
        RECT 86.755 172.535 87.085 172.895 ;
        RECT 87.445 172.795 87.615 174.915 ;
        RECT 87.785 174.585 88.115 175.085 ;
        RECT 88.285 174.415 88.540 174.915 ;
        RECT 87.790 174.245 88.540 174.415 ;
        RECT 87.790 173.255 88.020 174.245 ;
        RECT 88.190 173.425 88.540 174.075 ;
        RECT 89.175 173.995 92.685 175.085 ;
        RECT 92.855 174.325 93.370 174.735 ;
        RECT 93.605 174.325 93.775 175.085 ;
        RECT 93.945 174.745 95.975 174.915 ;
        RECT 89.175 173.475 90.865 173.995 ;
        RECT 91.035 173.305 92.685 173.825 ;
        RECT 92.855 173.515 93.195 174.325 ;
        RECT 93.945 174.080 94.115 174.745 ;
        RECT 94.510 174.405 95.635 174.575 ;
        RECT 93.365 173.890 94.115 174.080 ;
        RECT 94.285 174.065 95.295 174.235 ;
        RECT 92.855 173.345 94.085 173.515 ;
        RECT 87.790 173.085 88.540 173.255 ;
        RECT 87.785 172.535 88.115 172.915 ;
        RECT 88.285 172.795 88.540 173.085 ;
        RECT 89.175 172.535 92.685 173.305 ;
        RECT 93.130 172.740 93.375 173.345 ;
        RECT 93.595 172.535 94.105 173.070 ;
        RECT 94.285 172.705 94.475 174.065 ;
        RECT 94.645 173.725 94.920 173.865 ;
        RECT 94.645 173.555 94.925 173.725 ;
        RECT 94.645 172.705 94.920 173.555 ;
        RECT 95.125 173.265 95.295 174.065 ;
        RECT 95.465 173.275 95.635 174.405 ;
        RECT 95.805 173.775 95.975 174.745 ;
        RECT 96.145 173.945 96.315 175.085 ;
        RECT 96.485 173.945 96.820 174.915 ;
        RECT 97.085 174.155 97.255 174.915 ;
        RECT 97.435 174.325 97.765 175.085 ;
        RECT 97.085 173.985 97.750 174.155 ;
        RECT 97.935 174.010 98.205 174.915 ;
        RECT 95.805 173.445 96.000 173.775 ;
        RECT 96.225 173.445 96.480 173.775 ;
        RECT 96.225 173.275 96.395 173.445 ;
        RECT 96.650 173.275 96.820 173.945 ;
        RECT 97.580 173.840 97.750 173.985 ;
        RECT 97.015 173.435 97.345 173.805 ;
        RECT 97.580 173.510 97.865 173.840 ;
        RECT 95.465 173.105 96.395 173.275 ;
        RECT 95.465 173.070 95.640 173.105 ;
        RECT 95.110 172.705 95.640 173.070 ;
        RECT 96.065 172.535 96.395 172.935 ;
        RECT 96.565 172.705 96.820 173.275 ;
        RECT 97.580 173.255 97.750 173.510 ;
        RECT 97.085 173.085 97.750 173.255 ;
        RECT 98.035 173.210 98.205 174.010 ;
        RECT 98.375 173.995 99.585 175.085 ;
        RECT 98.375 173.455 98.895 173.995 ;
        RECT 99.755 173.920 100.045 175.085 ;
        RECT 100.675 173.995 103.265 175.085 ;
        RECT 103.435 174.010 103.705 174.915 ;
        RECT 103.875 174.325 104.205 175.085 ;
        RECT 104.385 174.155 104.555 174.915 ;
        RECT 105.740 174.650 111.085 175.085 ;
        RECT 99.065 173.285 99.585 173.825 ;
        RECT 100.675 173.475 101.885 173.995 ;
        RECT 102.055 173.305 103.265 173.825 ;
        RECT 97.085 172.705 97.255 173.085 ;
        RECT 97.435 172.535 97.765 172.915 ;
        RECT 97.945 172.705 98.205 173.210 ;
        RECT 98.375 172.535 99.585 173.285 ;
        RECT 99.755 172.535 100.045 173.260 ;
        RECT 100.675 172.535 103.265 173.305 ;
        RECT 103.435 173.210 103.605 174.010 ;
        RECT 103.890 173.985 104.555 174.155 ;
        RECT 103.890 173.840 104.060 173.985 ;
        RECT 103.775 173.510 104.060 173.840 ;
        RECT 103.890 173.255 104.060 173.510 ;
        RECT 104.295 173.435 104.625 173.805 ;
        RECT 107.330 173.400 107.680 174.650 ;
        RECT 111.295 173.945 111.525 175.085 ;
        RECT 111.695 173.935 112.025 174.915 ;
        RECT 112.195 173.945 112.405 175.085 ;
        RECT 103.435 172.705 103.695 173.210 ;
        RECT 103.890 173.085 104.555 173.255 ;
        RECT 103.875 172.535 104.205 172.915 ;
        RECT 104.385 172.705 104.555 173.085 ;
        RECT 109.160 173.080 109.500 173.910 ;
        RECT 111.275 173.525 111.605 173.775 ;
        RECT 105.740 172.535 111.085 173.080 ;
        RECT 111.295 172.535 111.525 173.355 ;
        RECT 111.775 173.335 112.025 173.935 ;
        RECT 112.640 173.895 112.895 174.775 ;
        RECT 113.065 173.945 113.370 175.085 ;
        RECT 113.710 174.705 114.040 175.085 ;
        RECT 114.220 174.535 114.390 174.825 ;
        RECT 114.560 174.625 114.810 175.085 ;
        RECT 113.590 174.365 114.390 174.535 ;
        RECT 114.980 174.575 115.850 174.915 ;
        RECT 111.695 172.705 112.025 173.335 ;
        RECT 112.195 172.535 112.405 173.355 ;
        RECT 112.640 173.245 112.850 173.895 ;
        RECT 113.590 173.775 113.760 174.365 ;
        RECT 114.980 174.195 115.150 174.575 ;
        RECT 116.085 174.455 116.255 174.915 ;
        RECT 116.425 174.625 116.795 175.085 ;
        RECT 117.090 174.485 117.260 174.825 ;
        RECT 117.430 174.655 117.760 175.085 ;
        RECT 117.995 174.485 118.165 174.825 ;
        RECT 113.930 174.025 115.150 174.195 ;
        RECT 115.320 174.115 115.780 174.405 ;
        RECT 116.085 174.285 116.645 174.455 ;
        RECT 117.090 174.315 118.165 174.485 ;
        RECT 118.335 174.585 119.015 174.915 ;
        RECT 119.230 174.585 119.480 174.915 ;
        RECT 119.650 174.625 119.900 175.085 ;
        RECT 116.475 174.145 116.645 174.285 ;
        RECT 115.320 174.105 116.285 174.115 ;
        RECT 114.980 173.935 115.150 174.025 ;
        RECT 115.610 173.945 116.285 174.105 ;
        RECT 113.020 173.745 113.760 173.775 ;
        RECT 113.020 173.445 113.935 173.745 ;
        RECT 113.610 173.270 113.935 173.445 ;
        RECT 112.640 172.715 112.895 173.245 ;
        RECT 113.065 172.535 113.370 172.995 ;
        RECT 113.615 172.915 113.935 173.270 ;
        RECT 114.105 173.485 114.645 173.855 ;
        RECT 114.980 173.765 115.385 173.935 ;
        RECT 114.105 173.085 114.345 173.485 ;
        RECT 114.825 173.315 115.045 173.595 ;
        RECT 114.515 173.145 115.045 173.315 ;
        RECT 114.515 172.915 114.685 173.145 ;
        RECT 115.215 172.985 115.385 173.765 ;
        RECT 115.555 173.155 115.905 173.775 ;
        RECT 116.075 173.155 116.285 173.945 ;
        RECT 116.475 173.975 117.975 174.145 ;
        RECT 116.475 173.285 116.645 173.975 ;
        RECT 118.335 173.805 118.505 174.585 ;
        RECT 119.310 174.455 119.480 174.585 ;
        RECT 116.815 173.635 118.505 173.805 ;
        RECT 118.675 174.025 119.140 174.415 ;
        RECT 119.310 174.285 119.705 174.455 ;
        RECT 116.815 173.455 116.985 173.635 ;
        RECT 113.615 172.745 114.685 172.915 ;
        RECT 114.855 172.535 115.045 172.975 ;
        RECT 115.215 172.705 116.165 172.985 ;
        RECT 116.475 172.895 116.735 173.285 ;
        RECT 117.155 173.215 117.945 173.465 ;
        RECT 116.385 172.725 116.735 172.895 ;
        RECT 116.945 172.535 117.275 172.995 ;
        RECT 118.150 172.925 118.320 173.635 ;
        RECT 118.675 173.435 118.845 174.025 ;
        RECT 118.490 173.215 118.845 173.435 ;
        RECT 119.015 173.215 119.365 173.835 ;
        RECT 119.535 172.925 119.705 174.285 ;
        RECT 120.070 174.115 120.395 174.900 ;
        RECT 119.875 173.065 120.335 174.115 ;
        RECT 118.150 172.755 119.005 172.925 ;
        RECT 119.210 172.755 119.705 172.925 ;
        RECT 119.875 172.535 120.205 172.895 ;
        RECT 120.565 172.795 120.735 174.915 ;
        RECT 120.905 174.585 121.235 175.085 ;
        RECT 121.405 174.415 121.660 174.915 ;
        RECT 121.840 174.660 122.175 175.085 ;
        RECT 122.345 174.480 122.530 174.885 ;
        RECT 120.910 174.245 121.660 174.415 ;
        RECT 121.865 174.305 122.530 174.480 ;
        RECT 122.735 174.305 123.065 175.085 ;
        RECT 120.910 173.255 121.140 174.245 ;
        RECT 121.310 173.425 121.660 174.075 ;
        RECT 121.865 173.275 122.205 174.305 ;
        RECT 123.235 174.115 123.505 174.885 ;
        RECT 122.375 173.945 123.505 174.115 ;
        RECT 122.375 173.445 122.625 173.945 ;
        RECT 120.910 173.085 121.660 173.255 ;
        RECT 121.865 173.105 122.550 173.275 ;
        RECT 122.805 173.195 123.165 173.775 ;
        RECT 120.905 172.535 121.235 172.915 ;
        RECT 121.405 172.795 121.660 173.085 ;
        RECT 121.840 172.535 122.175 172.935 ;
        RECT 122.345 172.705 122.550 173.105 ;
        RECT 123.335 173.035 123.505 173.945 ;
        RECT 124.595 173.995 125.805 175.085 ;
        RECT 124.595 173.455 125.115 173.995 ;
        RECT 125.285 173.285 125.805 173.825 ;
        RECT 122.760 172.535 123.035 173.015 ;
        RECT 123.245 172.705 123.505 173.035 ;
        RECT 124.595 172.535 125.805 173.285 ;
        RECT 11.810 172.365 125.890 172.535 ;
        RECT 11.895 171.615 13.105 172.365 ;
        RECT 11.895 171.075 12.415 171.615 ;
        RECT 13.735 171.595 17.245 172.365 ;
        RECT 12.585 170.905 13.105 171.445 ;
        RECT 11.895 169.815 13.105 170.905 ;
        RECT 13.735 170.905 15.425 171.425 ;
        RECT 15.595 171.075 17.245 171.595 ;
        RECT 17.790 171.655 18.045 172.185 ;
        RECT 18.225 171.905 18.510 172.365 ;
        RECT 13.735 169.815 17.245 170.905 ;
        RECT 17.790 170.795 17.970 171.655 ;
        RECT 18.690 171.455 18.940 172.105 ;
        RECT 18.140 171.125 18.940 171.455 ;
        RECT 17.790 170.325 18.045 170.795 ;
        RECT 17.705 170.155 18.045 170.325 ;
        RECT 17.790 170.125 18.045 170.155 ;
        RECT 18.225 169.815 18.510 170.615 ;
        RECT 18.690 170.535 18.940 171.125 ;
        RECT 19.140 171.770 19.460 172.100 ;
        RECT 19.640 171.885 20.300 172.365 ;
        RECT 20.500 171.975 21.350 172.145 ;
        RECT 19.140 170.875 19.330 171.770 ;
        RECT 19.650 171.445 20.310 171.715 ;
        RECT 19.980 171.385 20.310 171.445 ;
        RECT 19.500 171.215 19.830 171.275 ;
        RECT 20.500 171.215 20.670 171.975 ;
        RECT 21.910 171.905 22.230 172.365 ;
        RECT 22.430 171.725 22.680 172.155 ;
        RECT 22.970 171.925 23.380 172.365 ;
        RECT 23.550 171.985 24.565 172.185 ;
        RECT 20.840 171.555 22.090 171.725 ;
        RECT 20.840 171.435 21.170 171.555 ;
        RECT 19.500 171.045 21.400 171.215 ;
        RECT 19.140 170.705 21.060 170.875 ;
        RECT 19.140 170.685 19.460 170.705 ;
        RECT 18.690 170.025 19.020 170.535 ;
        RECT 19.290 170.075 19.460 170.685 ;
        RECT 21.230 170.535 21.400 171.045 ;
        RECT 21.570 170.975 21.750 171.385 ;
        RECT 21.920 170.795 22.090 171.555 ;
        RECT 19.630 169.815 19.960 170.505 ;
        RECT 20.190 170.365 21.400 170.535 ;
        RECT 21.570 170.485 22.090 170.795 ;
        RECT 22.260 171.385 22.680 171.725 ;
        RECT 22.970 171.385 23.380 171.715 ;
        RECT 22.260 170.615 22.450 171.385 ;
        RECT 23.550 171.255 23.720 171.985 ;
        RECT 24.865 171.815 25.035 172.145 ;
        RECT 25.205 171.985 25.535 172.365 ;
        RECT 23.890 171.435 24.240 171.805 ;
        RECT 23.550 171.215 23.970 171.255 ;
        RECT 22.620 171.045 23.970 171.215 ;
        RECT 22.620 170.885 22.870 171.045 ;
        RECT 23.380 170.615 23.630 170.875 ;
        RECT 22.260 170.365 23.630 170.615 ;
        RECT 20.190 170.075 20.430 170.365 ;
        RECT 21.230 170.285 21.400 170.365 ;
        RECT 20.630 169.815 21.050 170.195 ;
        RECT 21.230 170.035 21.860 170.285 ;
        RECT 22.330 169.815 22.660 170.195 ;
        RECT 22.830 170.075 23.000 170.365 ;
        RECT 23.800 170.200 23.970 171.045 ;
        RECT 24.420 170.875 24.640 171.745 ;
        RECT 24.865 171.625 25.560 171.815 ;
        RECT 24.140 170.495 24.640 170.875 ;
        RECT 24.810 170.825 25.220 171.445 ;
        RECT 25.390 170.655 25.560 171.625 ;
        RECT 24.865 170.485 25.560 170.655 ;
        RECT 23.180 169.815 23.560 170.195 ;
        RECT 23.800 170.030 24.630 170.200 ;
        RECT 24.865 169.985 25.035 170.485 ;
        RECT 25.205 169.815 25.535 170.315 ;
        RECT 25.750 169.985 25.975 172.105 ;
        RECT 26.145 171.985 26.475 172.365 ;
        RECT 26.645 171.815 26.815 172.105 ;
        RECT 26.150 171.645 26.815 171.815 ;
        RECT 27.650 171.735 27.935 172.195 ;
        RECT 28.105 171.905 28.375 172.365 ;
        RECT 26.150 170.655 26.380 171.645 ;
        RECT 27.650 171.565 28.605 171.735 ;
        RECT 26.550 170.825 26.900 171.475 ;
        RECT 27.535 170.835 28.225 171.395 ;
        RECT 28.395 170.665 28.605 171.565 ;
        RECT 26.150 170.485 26.815 170.655 ;
        RECT 26.145 169.815 26.475 170.315 ;
        RECT 26.645 169.985 26.815 170.485 ;
        RECT 27.650 170.445 28.605 170.665 ;
        RECT 28.775 171.395 29.175 172.195 ;
        RECT 29.365 171.735 29.645 172.195 ;
        RECT 30.165 171.905 30.490 172.365 ;
        RECT 29.365 171.565 30.490 171.735 ;
        RECT 30.660 171.625 31.045 172.195 ;
        RECT 30.040 171.455 30.490 171.565 ;
        RECT 28.775 170.835 29.870 171.395 ;
        RECT 30.040 171.125 30.595 171.455 ;
        RECT 27.650 169.985 27.935 170.445 ;
        RECT 28.105 169.815 28.375 170.275 ;
        RECT 28.775 169.985 29.175 170.835 ;
        RECT 30.040 170.665 30.490 171.125 ;
        RECT 30.765 170.955 31.045 171.625 ;
        RECT 31.490 171.555 31.735 172.160 ;
        RECT 31.955 171.830 32.465 172.365 ;
        RECT 29.365 170.445 30.490 170.665 ;
        RECT 29.365 169.985 29.645 170.445 ;
        RECT 30.165 169.815 30.490 170.275 ;
        RECT 30.660 169.985 31.045 170.955 ;
        RECT 31.215 171.385 32.445 171.555 ;
        RECT 31.215 170.575 31.555 171.385 ;
        RECT 31.725 170.820 32.475 171.010 ;
        RECT 31.215 170.165 31.730 170.575 ;
        RECT 31.965 169.815 32.135 170.575 ;
        RECT 32.305 170.155 32.475 170.820 ;
        RECT 32.645 170.835 32.835 172.195 ;
        RECT 33.005 171.685 33.280 172.195 ;
        RECT 33.470 171.830 34.000 172.195 ;
        RECT 34.425 171.965 34.755 172.365 ;
        RECT 33.825 171.795 34.000 171.830 ;
        RECT 33.005 171.515 33.285 171.685 ;
        RECT 33.005 171.035 33.280 171.515 ;
        RECT 33.485 170.835 33.655 171.635 ;
        RECT 32.645 170.665 33.655 170.835 ;
        RECT 33.825 171.625 34.755 171.795 ;
        RECT 34.925 171.625 35.180 172.195 ;
        RECT 35.355 171.640 35.645 172.365 ;
        RECT 35.820 171.655 36.075 172.185 ;
        RECT 36.245 171.905 36.550 172.365 ;
        RECT 36.795 171.985 37.865 172.155 ;
        RECT 33.825 170.495 33.995 171.625 ;
        RECT 34.585 171.455 34.755 171.625 ;
        RECT 32.870 170.325 33.995 170.495 ;
        RECT 34.165 171.125 34.360 171.455 ;
        RECT 34.585 171.125 34.840 171.455 ;
        RECT 34.165 170.155 34.335 171.125 ;
        RECT 35.010 170.955 35.180 171.625 ;
        RECT 35.820 171.005 36.030 171.655 ;
        RECT 36.795 171.630 37.115 171.985 ;
        RECT 36.790 171.455 37.115 171.630 ;
        RECT 36.200 171.155 37.115 171.455 ;
        RECT 37.285 171.415 37.525 171.815 ;
        RECT 37.695 171.755 37.865 171.985 ;
        RECT 38.035 171.925 38.225 172.365 ;
        RECT 38.395 171.915 39.345 172.195 ;
        RECT 39.565 172.005 39.915 172.175 ;
        RECT 37.695 171.585 38.225 171.755 ;
        RECT 36.200 171.125 36.940 171.155 ;
        RECT 32.305 169.985 34.335 170.155 ;
        RECT 34.505 169.815 34.675 170.955 ;
        RECT 34.845 169.985 35.180 170.955 ;
        RECT 35.355 169.815 35.645 170.980 ;
        RECT 35.820 170.125 36.075 171.005 ;
        RECT 36.245 169.815 36.550 170.955 ;
        RECT 36.770 170.535 36.940 171.125 ;
        RECT 37.285 171.045 37.825 171.415 ;
        RECT 38.005 171.305 38.225 171.585 ;
        RECT 38.395 171.135 38.565 171.915 ;
        RECT 38.160 170.965 38.565 171.135 ;
        RECT 38.735 171.125 39.085 171.745 ;
        RECT 38.160 170.875 38.330 170.965 ;
        RECT 39.255 170.955 39.465 171.745 ;
        RECT 37.110 170.705 38.330 170.875 ;
        RECT 38.790 170.795 39.465 170.955 ;
        RECT 36.770 170.365 37.570 170.535 ;
        RECT 36.890 169.815 37.220 170.195 ;
        RECT 37.400 170.075 37.570 170.365 ;
        RECT 38.160 170.325 38.330 170.705 ;
        RECT 38.500 170.785 39.465 170.795 ;
        RECT 39.655 171.615 39.915 172.005 ;
        RECT 40.125 171.905 40.455 172.365 ;
        RECT 41.330 171.975 42.185 172.145 ;
        RECT 42.390 171.975 42.885 172.145 ;
        RECT 43.055 172.005 43.385 172.365 ;
        RECT 39.655 170.925 39.825 171.615 ;
        RECT 39.995 171.265 40.165 171.445 ;
        RECT 40.335 171.435 41.125 171.685 ;
        RECT 41.330 171.265 41.500 171.975 ;
        RECT 41.670 171.465 42.025 171.685 ;
        RECT 39.995 171.095 41.685 171.265 ;
        RECT 38.500 170.495 38.960 170.785 ;
        RECT 39.655 170.755 41.155 170.925 ;
        RECT 39.655 170.615 39.825 170.755 ;
        RECT 39.265 170.445 39.825 170.615 ;
        RECT 37.740 169.815 37.990 170.275 ;
        RECT 38.160 169.985 39.030 170.325 ;
        RECT 39.265 169.985 39.435 170.445 ;
        RECT 40.270 170.415 41.345 170.585 ;
        RECT 39.605 169.815 39.975 170.275 ;
        RECT 40.270 170.075 40.440 170.415 ;
        RECT 40.610 169.815 40.940 170.245 ;
        RECT 41.175 170.075 41.345 170.415 ;
        RECT 41.515 170.315 41.685 171.095 ;
        RECT 41.855 170.875 42.025 171.465 ;
        RECT 42.195 171.065 42.545 171.685 ;
        RECT 41.855 170.485 42.320 170.875 ;
        RECT 42.715 170.615 42.885 171.975 ;
        RECT 43.055 170.785 43.515 171.835 ;
        RECT 42.490 170.445 42.885 170.615 ;
        RECT 42.490 170.315 42.660 170.445 ;
        RECT 41.515 169.985 42.195 170.315 ;
        RECT 42.410 169.985 42.660 170.315 ;
        RECT 42.830 169.815 43.080 170.275 ;
        RECT 43.250 170.000 43.575 170.785 ;
        RECT 43.745 169.985 43.915 172.105 ;
        RECT 44.085 171.985 44.415 172.365 ;
        RECT 44.585 171.815 44.840 172.105 ;
        RECT 44.090 171.645 44.840 171.815 ;
        RECT 46.310 171.655 46.565 172.185 ;
        RECT 46.745 171.905 47.030 172.365 ;
        RECT 44.090 170.655 44.320 171.645 ;
        RECT 44.490 170.825 44.840 171.475 ;
        RECT 46.310 171.345 46.490 171.655 ;
        RECT 47.210 171.455 47.460 172.105 ;
        RECT 46.225 171.175 46.490 171.345 ;
        RECT 46.310 170.795 46.490 171.175 ;
        RECT 46.660 171.125 47.460 171.455 ;
        RECT 44.090 170.485 44.840 170.655 ;
        RECT 44.085 169.815 44.415 170.315 ;
        RECT 44.585 169.985 44.840 170.485 ;
        RECT 46.310 170.125 46.565 170.795 ;
        RECT 46.745 169.815 47.030 170.615 ;
        RECT 47.210 170.535 47.460 171.125 ;
        RECT 47.660 171.770 47.980 172.100 ;
        RECT 48.160 171.885 48.820 172.365 ;
        RECT 49.020 171.975 49.870 172.145 ;
        RECT 47.660 170.875 47.850 171.770 ;
        RECT 48.170 171.445 48.830 171.715 ;
        RECT 48.500 171.385 48.830 171.445 ;
        RECT 48.020 171.215 48.350 171.275 ;
        RECT 49.020 171.215 49.190 171.975 ;
        RECT 50.430 171.905 50.750 172.365 ;
        RECT 50.950 171.725 51.200 172.155 ;
        RECT 51.490 171.925 51.900 172.365 ;
        RECT 52.070 171.985 53.085 172.185 ;
        RECT 49.360 171.555 50.610 171.725 ;
        RECT 49.360 171.435 49.690 171.555 ;
        RECT 48.020 171.045 49.920 171.215 ;
        RECT 47.660 170.705 49.580 170.875 ;
        RECT 47.660 170.685 47.980 170.705 ;
        RECT 47.210 170.025 47.540 170.535 ;
        RECT 47.810 170.075 47.980 170.685 ;
        RECT 49.750 170.535 49.920 171.045 ;
        RECT 50.090 170.975 50.270 171.385 ;
        RECT 50.440 170.795 50.610 171.555 ;
        RECT 48.150 169.815 48.480 170.505 ;
        RECT 48.710 170.365 49.920 170.535 ;
        RECT 50.090 170.485 50.610 170.795 ;
        RECT 50.780 171.385 51.200 171.725 ;
        RECT 51.490 171.385 51.900 171.715 ;
        RECT 50.780 170.615 50.970 171.385 ;
        RECT 52.070 171.255 52.240 171.985 ;
        RECT 53.385 171.815 53.555 172.145 ;
        RECT 53.725 171.985 54.055 172.365 ;
        RECT 52.410 171.435 52.760 171.805 ;
        RECT 52.070 171.215 52.490 171.255 ;
        RECT 51.140 171.045 52.490 171.215 ;
        RECT 51.140 170.885 51.390 171.045 ;
        RECT 51.900 170.615 52.150 170.875 ;
        RECT 50.780 170.365 52.150 170.615 ;
        RECT 48.710 170.075 48.950 170.365 ;
        RECT 49.750 170.285 49.920 170.365 ;
        RECT 49.150 169.815 49.570 170.195 ;
        RECT 49.750 170.035 50.380 170.285 ;
        RECT 50.850 169.815 51.180 170.195 ;
        RECT 51.350 170.075 51.520 170.365 ;
        RECT 52.320 170.200 52.490 171.045 ;
        RECT 52.940 170.875 53.160 171.745 ;
        RECT 53.385 171.625 54.080 171.815 ;
        RECT 52.660 170.495 53.160 170.875 ;
        RECT 53.330 170.825 53.740 171.445 ;
        RECT 53.910 170.655 54.080 171.625 ;
        RECT 53.385 170.485 54.080 170.655 ;
        RECT 51.700 169.815 52.080 170.195 ;
        RECT 52.320 170.030 53.150 170.200 ;
        RECT 53.385 169.985 53.555 170.485 ;
        RECT 53.725 169.815 54.055 170.315 ;
        RECT 54.270 169.985 54.495 172.105 ;
        RECT 54.665 171.985 54.995 172.365 ;
        RECT 55.165 171.815 55.335 172.105 ;
        RECT 54.670 171.645 55.335 171.815 ;
        RECT 54.670 170.655 54.900 171.645 ;
        RECT 55.870 171.555 56.115 172.160 ;
        RECT 56.335 171.830 56.845 172.365 ;
        RECT 55.070 170.825 55.420 171.475 ;
        RECT 55.595 171.385 56.825 171.555 ;
        RECT 54.670 170.485 55.335 170.655 ;
        RECT 54.665 169.815 54.995 170.315 ;
        RECT 55.165 169.985 55.335 170.485 ;
        RECT 55.595 170.575 55.935 171.385 ;
        RECT 56.105 170.820 56.855 171.010 ;
        RECT 55.595 170.165 56.110 170.575 ;
        RECT 56.345 169.815 56.515 170.575 ;
        RECT 56.685 170.155 56.855 170.820 ;
        RECT 57.025 170.835 57.215 172.195 ;
        RECT 57.385 171.345 57.660 172.195 ;
        RECT 57.850 171.830 58.380 172.195 ;
        RECT 58.805 171.965 59.135 172.365 ;
        RECT 58.205 171.795 58.380 171.830 ;
        RECT 57.385 171.175 57.665 171.345 ;
        RECT 57.385 171.035 57.660 171.175 ;
        RECT 57.865 170.835 58.035 171.635 ;
        RECT 57.025 170.665 58.035 170.835 ;
        RECT 58.205 171.625 59.135 171.795 ;
        RECT 59.305 171.625 59.560 172.195 ;
        RECT 58.205 170.495 58.375 171.625 ;
        RECT 58.965 171.455 59.135 171.625 ;
        RECT 57.250 170.325 58.375 170.495 ;
        RECT 58.545 171.125 58.740 171.455 ;
        RECT 58.965 171.125 59.220 171.455 ;
        RECT 58.545 170.155 58.715 171.125 ;
        RECT 59.390 170.955 59.560 171.625 ;
        RECT 56.685 169.985 58.715 170.155 ;
        RECT 58.885 169.815 59.055 170.955 ;
        RECT 59.225 169.985 59.560 170.955 ;
        RECT 59.735 171.690 59.995 172.195 ;
        RECT 60.175 171.985 60.505 172.365 ;
        RECT 60.685 171.815 60.855 172.195 ;
        RECT 59.735 170.890 59.905 171.690 ;
        RECT 60.190 171.645 60.855 171.815 ;
        RECT 60.190 171.390 60.360 171.645 ;
        RECT 61.115 171.640 61.405 172.365 ;
        RECT 61.635 171.885 61.915 172.365 ;
        RECT 62.085 171.715 62.345 172.105 ;
        RECT 62.520 171.885 62.775 172.365 ;
        RECT 62.945 171.715 63.240 172.105 ;
        RECT 63.420 171.885 63.695 172.365 ;
        RECT 63.865 171.865 64.165 172.195 ;
        RECT 61.590 171.545 63.240 171.715 ;
        RECT 60.075 171.060 60.360 171.390 ;
        RECT 60.595 171.095 60.925 171.465 ;
        RECT 60.190 170.915 60.360 171.060 ;
        RECT 61.590 171.035 61.995 171.545 ;
        RECT 62.165 171.205 63.305 171.375 ;
        RECT 59.735 169.985 60.005 170.890 ;
        RECT 60.190 170.745 60.855 170.915 ;
        RECT 60.175 169.815 60.505 170.575 ;
        RECT 60.685 169.985 60.855 170.745 ;
        RECT 61.115 169.815 61.405 170.980 ;
        RECT 61.590 170.865 62.345 171.035 ;
        RECT 61.630 169.815 61.915 170.685 ;
        RECT 62.085 170.615 62.345 170.865 ;
        RECT 63.135 170.955 63.305 171.205 ;
        RECT 63.475 171.125 63.825 171.695 ;
        RECT 63.995 170.955 64.165 171.865 ;
        RECT 65.255 171.595 68.765 172.365 ;
        RECT 63.135 170.785 64.165 170.955 ;
        RECT 62.555 170.615 62.725 170.665 ;
        RECT 62.085 170.445 63.205 170.615 ;
        RECT 62.085 169.985 62.345 170.445 ;
        RECT 62.520 169.815 62.775 170.275 ;
        RECT 62.945 169.985 63.205 170.445 ;
        RECT 63.375 169.815 63.685 170.615 ;
        RECT 63.855 169.985 64.165 170.785 ;
        RECT 65.255 170.905 66.945 171.425 ;
        RECT 67.115 171.075 68.765 171.595 ;
        RECT 68.975 171.545 69.205 172.365 ;
        RECT 69.375 171.565 69.705 172.195 ;
        RECT 68.955 171.125 69.285 171.375 ;
        RECT 69.455 170.965 69.705 171.565 ;
        RECT 69.875 171.545 70.085 172.365 ;
        RECT 70.620 171.795 70.790 172.045 ;
        RECT 70.315 171.625 70.790 171.795 ;
        RECT 71.025 171.625 71.355 172.365 ;
        RECT 71.525 171.795 71.725 172.140 ;
        RECT 71.895 171.965 72.225 172.365 ;
        RECT 72.395 171.795 72.595 172.150 ;
        RECT 72.765 171.970 73.095 172.365 ;
        RECT 73.535 171.865 73.835 172.195 ;
        RECT 74.005 171.885 74.280 172.365 ;
        RECT 71.525 171.625 73.365 171.795 ;
        RECT 65.255 169.815 68.765 170.905 ;
        RECT 68.975 169.815 69.205 170.955 ;
        RECT 69.375 169.985 69.705 170.965 ;
        RECT 69.875 169.815 70.085 170.955 ;
        RECT 70.315 170.655 70.485 171.625 ;
        RECT 70.655 170.835 71.005 171.455 ;
        RECT 71.175 170.835 71.495 171.455 ;
        RECT 71.665 170.835 71.995 171.455 ;
        RECT 72.165 170.835 72.465 171.455 ;
        RECT 72.705 170.655 72.925 171.455 ;
        RECT 70.315 170.445 72.925 170.655 ;
        RECT 71.025 169.815 71.355 170.265 ;
        RECT 73.105 170.000 73.365 171.625 ;
        RECT 73.535 170.955 73.705 171.865 ;
        RECT 74.460 171.715 74.755 172.105 ;
        RECT 74.925 171.885 75.180 172.365 ;
        RECT 75.355 171.715 75.615 172.105 ;
        RECT 75.785 171.885 76.065 172.365 ;
        RECT 73.875 171.125 74.225 171.695 ;
        RECT 74.460 171.545 76.110 171.715 ;
        RECT 76.755 171.595 79.345 172.365 ;
        RECT 79.520 171.820 84.865 172.365 ;
        RECT 74.395 171.205 75.535 171.375 ;
        RECT 74.395 170.955 74.565 171.205 ;
        RECT 75.705 171.035 76.110 171.545 ;
        RECT 73.535 170.785 74.565 170.955 ;
        RECT 75.355 170.865 76.110 171.035 ;
        RECT 76.755 170.905 77.965 171.425 ;
        RECT 78.135 171.075 79.345 171.595 ;
        RECT 73.535 169.985 73.845 170.785 ;
        RECT 75.355 170.615 75.615 170.865 ;
        RECT 74.015 169.815 74.325 170.615 ;
        RECT 74.495 170.445 75.615 170.615 ;
        RECT 74.495 169.985 74.755 170.445 ;
        RECT 74.925 169.815 75.180 170.275 ;
        RECT 75.355 169.985 75.615 170.445 ;
        RECT 75.785 169.815 76.070 170.685 ;
        RECT 76.755 169.815 79.345 170.905 ;
        RECT 81.110 170.250 81.460 171.500 ;
        RECT 82.940 170.990 83.280 171.820 ;
        RECT 85.125 171.815 85.295 172.195 ;
        RECT 85.475 171.985 85.805 172.365 ;
        RECT 85.125 171.645 85.790 171.815 ;
        RECT 85.985 171.690 86.245 172.195 ;
        RECT 85.055 171.095 85.385 171.465 ;
        RECT 85.620 171.390 85.790 171.645 ;
        RECT 85.620 171.060 85.905 171.390 ;
        RECT 85.620 170.915 85.790 171.060 ;
        RECT 85.125 170.745 85.790 170.915 ;
        RECT 86.075 170.890 86.245 171.690 ;
        RECT 86.875 171.640 87.165 172.365 ;
        RECT 87.395 171.545 87.605 172.365 ;
        RECT 87.775 171.565 88.105 172.195 ;
        RECT 79.520 169.815 84.865 170.250 ;
        RECT 85.125 169.985 85.295 170.745 ;
        RECT 85.475 169.815 85.805 170.575 ;
        RECT 85.975 169.985 86.245 170.890 ;
        RECT 86.875 169.815 87.165 170.980 ;
        RECT 87.775 170.965 88.025 171.565 ;
        RECT 88.275 171.545 88.505 172.365 ;
        RECT 89.175 171.595 90.845 172.365 ;
        RECT 88.195 171.125 88.525 171.375 ;
        RECT 87.395 169.815 87.605 170.955 ;
        RECT 87.775 169.985 88.105 170.965 ;
        RECT 88.275 169.815 88.505 170.955 ;
        RECT 89.175 170.905 89.925 171.425 ;
        RECT 90.095 171.075 90.845 171.595 ;
        RECT 91.220 171.585 91.720 172.195 ;
        RECT 91.015 171.125 91.365 171.375 ;
        RECT 91.550 170.955 91.720 171.585 ;
        RECT 92.350 171.715 92.680 172.195 ;
        RECT 92.850 171.905 93.075 172.365 ;
        RECT 93.245 171.715 93.575 172.195 ;
        RECT 92.350 171.545 93.575 171.715 ;
        RECT 93.765 171.565 94.015 172.365 ;
        RECT 94.185 171.565 94.525 172.195 ;
        RECT 94.695 171.615 95.905 172.365 ;
        RECT 91.890 171.175 92.220 171.375 ;
        RECT 92.390 171.175 92.720 171.375 ;
        RECT 92.890 171.175 93.310 171.375 ;
        RECT 93.485 171.205 94.180 171.375 ;
        RECT 93.485 170.955 93.655 171.205 ;
        RECT 94.350 170.955 94.525 171.565 ;
        RECT 89.175 169.815 90.845 170.905 ;
        RECT 91.220 170.785 93.655 170.955 ;
        RECT 91.220 169.985 91.550 170.785 ;
        RECT 91.720 169.815 92.050 170.615 ;
        RECT 92.350 169.985 92.680 170.785 ;
        RECT 93.325 169.815 93.575 170.615 ;
        RECT 93.845 169.815 94.015 170.955 ;
        RECT 94.185 169.985 94.525 170.955 ;
        RECT 94.695 170.905 95.215 171.445 ;
        RECT 95.385 171.075 95.905 171.615 ;
        RECT 96.075 171.595 99.585 172.365 ;
        RECT 96.075 170.905 97.765 171.425 ;
        RECT 97.935 171.075 99.585 171.595 ;
        RECT 99.755 171.690 100.015 172.195 ;
        RECT 100.195 171.985 100.525 172.365 ;
        RECT 100.705 171.815 100.875 172.195 ;
        RECT 94.695 169.815 95.905 170.905 ;
        RECT 96.075 169.815 99.585 170.905 ;
        RECT 99.755 170.890 99.925 171.690 ;
        RECT 100.210 171.645 100.875 171.815 ;
        RECT 100.210 171.390 100.380 171.645 ;
        RECT 101.135 171.595 103.725 172.365 ;
        RECT 100.095 171.060 100.380 171.390 ;
        RECT 100.615 171.095 100.945 171.465 ;
        RECT 100.210 170.915 100.380 171.060 ;
        RECT 99.755 169.985 100.025 170.890 ;
        RECT 100.210 170.745 100.875 170.915 ;
        RECT 100.195 169.815 100.525 170.575 ;
        RECT 100.705 169.985 100.875 170.745 ;
        RECT 101.135 170.905 102.345 171.425 ;
        RECT 102.515 171.075 103.725 171.595 ;
        RECT 103.895 171.565 104.235 172.195 ;
        RECT 104.405 171.565 104.655 172.365 ;
        RECT 104.845 171.715 105.175 172.195 ;
        RECT 105.345 171.905 105.570 172.365 ;
        RECT 105.740 171.715 106.070 172.195 ;
        RECT 103.895 170.955 104.070 171.565 ;
        RECT 104.845 171.545 106.070 171.715 ;
        RECT 106.700 171.585 107.200 172.195 ;
        RECT 104.240 171.205 104.935 171.375 ;
        RECT 104.765 170.955 104.935 171.205 ;
        RECT 105.110 171.175 105.530 171.375 ;
        RECT 105.700 171.175 106.030 171.375 ;
        RECT 106.200 171.175 106.530 171.375 ;
        RECT 106.700 170.955 106.870 171.585 ;
        RECT 108.770 171.555 109.015 172.160 ;
        RECT 109.235 171.830 109.745 172.365 ;
        RECT 108.495 171.385 109.725 171.555 ;
        RECT 107.055 171.125 107.405 171.375 ;
        RECT 101.135 169.815 103.725 170.905 ;
        RECT 103.895 169.985 104.235 170.955 ;
        RECT 104.405 169.815 104.575 170.955 ;
        RECT 104.765 170.785 107.200 170.955 ;
        RECT 104.845 169.815 105.095 170.615 ;
        RECT 105.740 169.985 106.070 170.785 ;
        RECT 106.370 169.815 106.700 170.615 ;
        RECT 106.870 169.985 107.200 170.785 ;
        RECT 108.495 170.575 108.835 171.385 ;
        RECT 109.005 170.820 109.755 171.010 ;
        RECT 108.495 170.165 109.010 170.575 ;
        RECT 109.245 169.815 109.415 170.575 ;
        RECT 109.585 170.155 109.755 170.820 ;
        RECT 109.925 170.835 110.115 172.195 ;
        RECT 110.285 171.345 110.560 172.195 ;
        RECT 110.750 171.830 111.280 172.195 ;
        RECT 111.705 171.965 112.035 172.365 ;
        RECT 111.105 171.795 111.280 171.830 ;
        RECT 110.285 171.175 110.565 171.345 ;
        RECT 110.285 171.035 110.560 171.175 ;
        RECT 110.765 170.835 110.935 171.635 ;
        RECT 109.925 170.665 110.935 170.835 ;
        RECT 111.105 171.625 112.035 171.795 ;
        RECT 112.205 171.625 112.460 172.195 ;
        RECT 112.635 171.640 112.925 172.365 ;
        RECT 111.105 170.495 111.275 171.625 ;
        RECT 111.865 171.455 112.035 171.625 ;
        RECT 110.150 170.325 111.275 170.495 ;
        RECT 111.445 171.125 111.640 171.455 ;
        RECT 111.865 171.125 112.120 171.455 ;
        RECT 111.445 170.155 111.615 171.125 ;
        RECT 112.290 170.955 112.460 171.625 ;
        RECT 113.370 171.555 113.615 172.160 ;
        RECT 113.835 171.830 114.345 172.365 ;
        RECT 113.095 171.385 114.325 171.555 ;
        RECT 109.585 169.985 111.615 170.155 ;
        RECT 111.785 169.815 111.955 170.955 ;
        RECT 112.125 169.985 112.460 170.955 ;
        RECT 112.635 169.815 112.925 170.980 ;
        RECT 113.095 170.575 113.435 171.385 ;
        RECT 113.605 170.820 114.355 171.010 ;
        RECT 113.095 170.165 113.610 170.575 ;
        RECT 113.845 169.815 114.015 170.575 ;
        RECT 114.185 170.155 114.355 170.820 ;
        RECT 114.525 170.835 114.715 172.195 ;
        RECT 114.885 171.685 115.160 172.195 ;
        RECT 115.350 171.830 115.880 172.195 ;
        RECT 116.305 171.965 116.635 172.365 ;
        RECT 115.705 171.795 115.880 171.830 ;
        RECT 114.885 171.515 115.165 171.685 ;
        RECT 114.885 171.035 115.160 171.515 ;
        RECT 115.365 170.835 115.535 171.635 ;
        RECT 114.525 170.665 115.535 170.835 ;
        RECT 115.705 171.625 116.635 171.795 ;
        RECT 116.805 171.625 117.060 172.195 ;
        RECT 117.325 171.815 117.495 172.195 ;
        RECT 117.675 171.985 118.005 172.365 ;
        RECT 117.325 171.645 117.990 171.815 ;
        RECT 118.185 171.690 118.445 172.195 ;
        RECT 115.705 170.495 115.875 171.625 ;
        RECT 116.465 171.455 116.635 171.625 ;
        RECT 114.750 170.325 115.875 170.495 ;
        RECT 116.045 171.125 116.240 171.455 ;
        RECT 116.465 171.125 116.720 171.455 ;
        RECT 116.045 170.155 116.215 171.125 ;
        RECT 116.890 170.955 117.060 171.625 ;
        RECT 117.255 171.095 117.585 171.465 ;
        RECT 117.820 171.390 117.990 171.645 ;
        RECT 114.185 169.985 116.215 170.155 ;
        RECT 116.385 169.815 116.555 170.955 ;
        RECT 116.725 169.985 117.060 170.955 ;
        RECT 117.820 171.060 118.105 171.390 ;
        RECT 117.820 170.915 117.990 171.060 ;
        RECT 117.325 170.745 117.990 170.915 ;
        RECT 118.275 170.890 118.445 171.690 ;
        RECT 119.165 171.815 119.335 172.195 ;
        RECT 119.515 171.985 119.845 172.365 ;
        RECT 119.165 171.645 119.830 171.815 ;
        RECT 120.025 171.690 120.285 172.195 ;
        RECT 119.095 171.095 119.425 171.465 ;
        RECT 119.660 171.390 119.830 171.645 ;
        RECT 119.660 171.060 119.945 171.390 ;
        RECT 119.660 170.915 119.830 171.060 ;
        RECT 117.325 169.985 117.495 170.745 ;
        RECT 117.675 169.815 118.005 170.575 ;
        RECT 118.175 169.985 118.445 170.890 ;
        RECT 119.165 170.745 119.830 170.915 ;
        RECT 120.115 170.890 120.285 171.690 ;
        RECT 120.915 171.595 124.425 172.365 ;
        RECT 124.595 171.615 125.805 172.365 ;
        RECT 119.165 169.985 119.335 170.745 ;
        RECT 119.515 169.815 119.845 170.575 ;
        RECT 120.015 169.985 120.285 170.890 ;
        RECT 120.915 170.905 122.605 171.425 ;
        RECT 122.775 171.075 124.425 171.595 ;
        RECT 124.595 170.905 125.115 171.445 ;
        RECT 125.285 171.075 125.805 171.615 ;
        RECT 120.915 169.815 124.425 170.905 ;
        RECT 124.595 169.815 125.805 170.905 ;
        RECT 11.810 169.645 125.890 169.815 ;
        RECT 11.895 168.555 13.105 169.645 ;
        RECT 11.895 167.845 12.415 168.385 ;
        RECT 12.585 168.015 13.105 168.555 ;
        RECT 13.275 168.555 16.785 169.645 ;
        RECT 13.275 168.035 14.965 168.555 ;
        RECT 17.015 168.505 17.225 169.645 ;
        RECT 17.395 168.495 17.725 169.475 ;
        RECT 17.895 168.505 18.125 169.645 ;
        RECT 18.335 168.885 18.850 169.295 ;
        RECT 19.085 168.885 19.255 169.645 ;
        RECT 19.425 169.305 21.455 169.475 ;
        RECT 15.135 167.865 16.785 168.385 ;
        RECT 11.895 167.095 13.105 167.845 ;
        RECT 13.275 167.095 16.785 167.865 ;
        RECT 17.015 167.095 17.225 167.915 ;
        RECT 17.395 167.895 17.645 168.495 ;
        RECT 17.815 168.085 18.145 168.335 ;
        RECT 18.335 168.075 18.675 168.885 ;
        RECT 19.425 168.640 19.595 169.305 ;
        RECT 19.990 168.965 21.115 169.135 ;
        RECT 18.845 168.450 19.595 168.640 ;
        RECT 19.765 168.625 20.775 168.795 ;
        RECT 17.395 167.265 17.725 167.895 ;
        RECT 17.895 167.095 18.125 167.915 ;
        RECT 18.335 167.905 19.565 168.075 ;
        RECT 18.610 167.300 18.855 167.905 ;
        RECT 19.075 167.095 19.585 167.630 ;
        RECT 19.765 167.265 19.955 168.625 ;
        RECT 20.125 167.945 20.400 168.425 ;
        RECT 20.125 167.775 20.405 167.945 ;
        RECT 20.605 167.825 20.775 168.625 ;
        RECT 20.945 167.835 21.115 168.965 ;
        RECT 21.285 168.335 21.455 169.305 ;
        RECT 21.625 168.505 21.795 169.645 ;
        RECT 21.965 168.505 22.300 169.475 ;
        RECT 21.285 168.005 21.480 168.335 ;
        RECT 21.705 168.005 21.960 168.335 ;
        RECT 21.705 167.835 21.875 168.005 ;
        RECT 22.130 167.835 22.300 168.505 ;
        RECT 22.475 168.480 22.765 169.645 ;
        RECT 20.125 167.265 20.400 167.775 ;
        RECT 20.945 167.665 21.875 167.835 ;
        RECT 20.945 167.630 21.120 167.665 ;
        RECT 20.590 167.265 21.120 167.630 ;
        RECT 21.545 167.095 21.875 167.495 ;
        RECT 22.045 167.265 22.300 167.835 ;
        RECT 22.940 168.455 23.195 169.335 ;
        RECT 23.365 168.505 23.670 169.645 ;
        RECT 24.010 169.265 24.340 169.645 ;
        RECT 24.520 169.095 24.690 169.385 ;
        RECT 24.860 169.185 25.110 169.645 ;
        RECT 23.890 168.925 24.690 169.095 ;
        RECT 25.280 169.135 26.150 169.475 ;
        RECT 22.475 167.095 22.765 167.820 ;
        RECT 22.940 167.805 23.150 168.455 ;
        RECT 23.890 168.335 24.060 168.925 ;
        RECT 25.280 168.755 25.450 169.135 ;
        RECT 26.385 169.015 26.555 169.475 ;
        RECT 26.725 169.185 27.095 169.645 ;
        RECT 27.390 169.045 27.560 169.385 ;
        RECT 27.730 169.215 28.060 169.645 ;
        RECT 28.295 169.045 28.465 169.385 ;
        RECT 24.230 168.585 25.450 168.755 ;
        RECT 25.620 168.675 26.080 168.965 ;
        RECT 26.385 168.845 26.945 169.015 ;
        RECT 27.390 168.875 28.465 169.045 ;
        RECT 28.635 169.145 29.315 169.475 ;
        RECT 29.530 169.145 29.780 169.475 ;
        RECT 29.950 169.185 30.200 169.645 ;
        RECT 26.775 168.705 26.945 168.845 ;
        RECT 25.620 168.665 26.585 168.675 ;
        RECT 25.280 168.495 25.450 168.585 ;
        RECT 25.910 168.505 26.585 168.665 ;
        RECT 23.320 168.305 24.060 168.335 ;
        RECT 23.320 168.005 24.235 168.305 ;
        RECT 23.910 167.830 24.235 168.005 ;
        RECT 22.940 167.275 23.195 167.805 ;
        RECT 23.365 167.095 23.670 167.555 ;
        RECT 23.915 167.475 24.235 167.830 ;
        RECT 24.405 168.045 24.945 168.415 ;
        RECT 25.280 168.325 25.685 168.495 ;
        RECT 24.405 167.645 24.645 168.045 ;
        RECT 25.125 167.875 25.345 168.155 ;
        RECT 24.815 167.705 25.345 167.875 ;
        RECT 24.815 167.475 24.985 167.705 ;
        RECT 25.515 167.545 25.685 168.325 ;
        RECT 25.855 167.715 26.205 168.335 ;
        RECT 26.375 167.715 26.585 168.505 ;
        RECT 26.775 168.535 28.275 168.705 ;
        RECT 26.775 167.845 26.945 168.535 ;
        RECT 28.635 168.365 28.805 169.145 ;
        RECT 29.610 169.015 29.780 169.145 ;
        RECT 27.115 168.195 28.805 168.365 ;
        RECT 28.975 168.585 29.440 168.975 ;
        RECT 29.610 168.845 30.005 169.015 ;
        RECT 27.115 168.015 27.285 168.195 ;
        RECT 23.915 167.305 24.985 167.475 ;
        RECT 25.155 167.095 25.345 167.535 ;
        RECT 25.515 167.265 26.465 167.545 ;
        RECT 26.775 167.455 27.035 167.845 ;
        RECT 27.455 167.775 28.245 168.025 ;
        RECT 26.685 167.285 27.035 167.455 ;
        RECT 27.245 167.095 27.575 167.555 ;
        RECT 28.450 167.485 28.620 168.195 ;
        RECT 28.975 167.995 29.145 168.585 ;
        RECT 28.790 167.775 29.145 167.995 ;
        RECT 29.315 167.775 29.665 168.395 ;
        RECT 29.835 167.485 30.005 168.845 ;
        RECT 30.370 168.675 30.695 169.460 ;
        RECT 30.175 167.625 30.635 168.675 ;
        RECT 28.450 167.315 29.305 167.485 ;
        RECT 29.510 167.315 30.005 167.485 ;
        RECT 30.175 167.095 30.505 167.455 ;
        RECT 30.865 167.355 31.035 169.475 ;
        RECT 31.205 169.145 31.535 169.645 ;
        RECT 31.705 168.975 31.960 169.475 ;
        RECT 31.210 168.805 31.960 168.975 ;
        RECT 31.210 167.815 31.440 168.805 ;
        RECT 31.610 167.985 31.960 168.635 ;
        RECT 32.135 168.555 35.645 169.645 ;
        RECT 32.135 168.035 33.825 168.555 ;
        RECT 35.855 168.505 36.085 169.645 ;
        RECT 36.255 168.495 36.585 169.475 ;
        RECT 36.755 168.505 36.965 169.645 ;
        RECT 37.195 168.885 37.710 169.295 ;
        RECT 37.945 168.885 38.115 169.645 ;
        RECT 38.285 169.305 40.315 169.475 ;
        RECT 33.995 167.865 35.645 168.385 ;
        RECT 35.835 168.085 36.165 168.335 ;
        RECT 31.210 167.645 31.960 167.815 ;
        RECT 31.205 167.095 31.535 167.475 ;
        RECT 31.705 167.355 31.960 167.645 ;
        RECT 32.135 167.095 35.645 167.865 ;
        RECT 35.855 167.095 36.085 167.915 ;
        RECT 36.335 167.895 36.585 168.495 ;
        RECT 37.195 168.075 37.535 168.885 ;
        RECT 38.285 168.640 38.455 169.305 ;
        RECT 38.850 168.965 39.975 169.135 ;
        RECT 37.705 168.450 38.455 168.640 ;
        RECT 38.625 168.625 39.635 168.795 ;
        RECT 36.255 167.265 36.585 167.895 ;
        RECT 36.755 167.095 36.965 167.915 ;
        RECT 37.195 167.905 38.425 168.075 ;
        RECT 37.470 167.300 37.715 167.905 ;
        RECT 37.935 167.095 38.445 167.630 ;
        RECT 38.625 167.265 38.815 168.625 ;
        RECT 38.985 167.605 39.260 168.425 ;
        RECT 39.465 167.825 39.635 168.625 ;
        RECT 39.805 167.835 39.975 168.965 ;
        RECT 40.145 168.335 40.315 169.305 ;
        RECT 40.485 168.505 40.655 169.645 ;
        RECT 40.825 168.505 41.160 169.475 ;
        RECT 41.425 168.715 41.595 169.475 ;
        RECT 41.775 168.885 42.105 169.645 ;
        RECT 41.425 168.545 42.090 168.715 ;
        RECT 42.275 168.570 42.545 169.475 ;
        RECT 40.145 168.005 40.340 168.335 ;
        RECT 40.565 168.005 40.820 168.335 ;
        RECT 40.565 167.835 40.735 168.005 ;
        RECT 40.990 167.835 41.160 168.505 ;
        RECT 41.920 168.400 42.090 168.545 ;
        RECT 41.355 167.995 41.685 168.365 ;
        RECT 41.920 168.070 42.205 168.400 ;
        RECT 39.805 167.665 40.735 167.835 ;
        RECT 39.805 167.630 39.980 167.665 ;
        RECT 38.985 167.435 39.265 167.605 ;
        RECT 38.985 167.265 39.260 167.435 ;
        RECT 39.450 167.265 39.980 167.630 ;
        RECT 40.405 167.095 40.735 167.495 ;
        RECT 40.905 167.265 41.160 167.835 ;
        RECT 41.920 167.815 42.090 168.070 ;
        RECT 41.425 167.645 42.090 167.815 ;
        RECT 42.375 167.770 42.545 168.570 ;
        RECT 42.715 168.555 43.925 169.645 ;
        RECT 44.095 168.885 44.610 169.295 ;
        RECT 44.845 168.885 45.015 169.645 ;
        RECT 45.185 169.305 47.215 169.475 ;
        RECT 42.715 168.015 43.235 168.555 ;
        RECT 43.405 167.845 43.925 168.385 ;
        RECT 44.095 168.075 44.435 168.885 ;
        RECT 45.185 168.640 45.355 169.305 ;
        RECT 45.750 168.965 46.875 169.135 ;
        RECT 44.605 168.450 45.355 168.640 ;
        RECT 45.525 168.625 46.535 168.795 ;
        RECT 44.095 167.905 45.325 168.075 ;
        RECT 41.425 167.265 41.595 167.645 ;
        RECT 41.775 167.095 42.105 167.475 ;
        RECT 42.285 167.265 42.545 167.770 ;
        RECT 42.715 167.095 43.925 167.845 ;
        RECT 44.370 167.300 44.615 167.905 ;
        RECT 44.835 167.095 45.345 167.630 ;
        RECT 45.525 167.265 45.715 168.625 ;
        RECT 45.885 168.285 46.160 168.425 ;
        RECT 45.885 168.115 46.165 168.285 ;
        RECT 45.885 167.265 46.160 168.115 ;
        RECT 46.365 167.825 46.535 168.625 ;
        RECT 46.705 167.835 46.875 168.965 ;
        RECT 47.045 168.335 47.215 169.305 ;
        RECT 47.385 168.505 47.555 169.645 ;
        RECT 47.725 168.505 48.060 169.475 ;
        RECT 47.045 168.005 47.240 168.335 ;
        RECT 47.465 168.005 47.720 168.335 ;
        RECT 47.465 167.835 47.635 168.005 ;
        RECT 47.890 167.835 48.060 168.505 ;
        RECT 48.235 168.480 48.525 169.645 ;
        RECT 49.155 168.555 50.825 169.645 ;
        RECT 51.085 168.715 51.255 169.475 ;
        RECT 51.435 168.885 51.765 169.645 ;
        RECT 49.155 168.035 49.905 168.555 ;
        RECT 51.085 168.545 51.750 168.715 ;
        RECT 51.935 168.570 52.205 169.475 ;
        RECT 51.580 168.400 51.750 168.545 ;
        RECT 50.075 167.865 50.825 168.385 ;
        RECT 51.015 167.995 51.345 168.365 ;
        RECT 51.580 168.070 51.865 168.400 ;
        RECT 46.705 167.665 47.635 167.835 ;
        RECT 46.705 167.630 46.880 167.665 ;
        RECT 46.350 167.265 46.880 167.630 ;
        RECT 47.305 167.095 47.635 167.495 ;
        RECT 47.805 167.265 48.060 167.835 ;
        RECT 48.235 167.095 48.525 167.820 ;
        RECT 49.155 167.095 50.825 167.865 ;
        RECT 51.580 167.815 51.750 168.070 ;
        RECT 51.085 167.645 51.750 167.815 ;
        RECT 52.035 167.770 52.205 168.570 ;
        RECT 52.835 168.555 54.505 169.645 ;
        RECT 52.835 168.035 53.585 168.555 ;
        RECT 54.715 168.505 54.945 169.645 ;
        RECT 55.115 168.495 55.445 169.475 ;
        RECT 55.615 168.505 55.825 169.645 ;
        RECT 56.205 168.495 56.535 169.645 ;
        RECT 56.705 168.625 56.875 169.475 ;
        RECT 57.045 168.845 57.375 169.645 ;
        RECT 57.545 168.625 57.715 169.475 ;
        RECT 57.895 168.845 58.135 169.645 ;
        RECT 58.305 168.665 58.635 169.475 ;
        RECT 53.755 167.865 54.505 168.385 ;
        RECT 54.695 168.085 55.025 168.335 ;
        RECT 51.085 167.265 51.255 167.645 ;
        RECT 51.435 167.095 51.765 167.475 ;
        RECT 51.945 167.265 52.205 167.770 ;
        RECT 52.835 167.095 54.505 167.865 ;
        RECT 54.715 167.095 54.945 167.915 ;
        RECT 55.195 167.895 55.445 168.495 ;
        RECT 56.705 168.455 57.715 168.625 ;
        RECT 57.920 168.495 58.635 168.665 ;
        RECT 58.965 168.495 59.295 169.645 ;
        RECT 59.465 168.625 59.635 169.475 ;
        RECT 59.805 168.845 60.135 169.645 ;
        RECT 60.305 168.625 60.475 169.475 ;
        RECT 60.655 168.845 60.895 169.645 ;
        RECT 61.065 168.665 61.395 169.475 ;
        RECT 61.580 169.210 66.925 169.645 ;
        RECT 56.705 167.915 57.200 168.455 ;
        RECT 57.920 168.255 58.090 168.495 ;
        RECT 59.465 168.455 60.475 168.625 ;
        RECT 60.680 168.495 61.395 168.665 ;
        RECT 57.590 168.085 58.090 168.255 ;
        RECT 58.260 168.085 58.640 168.325 ;
        RECT 57.920 167.915 58.090 168.085 ;
        RECT 59.465 167.945 59.960 168.455 ;
        RECT 60.680 168.255 60.850 168.495 ;
        RECT 60.350 168.085 60.850 168.255 ;
        RECT 61.020 168.085 61.400 168.325 ;
        RECT 59.465 167.915 59.965 167.945 ;
        RECT 60.680 167.915 60.850 168.085 ;
        RECT 63.170 167.960 63.520 169.210 ;
        RECT 67.150 168.775 67.435 169.645 ;
        RECT 67.605 169.015 67.865 169.475 ;
        RECT 68.040 169.185 68.295 169.645 ;
        RECT 68.465 169.015 68.725 169.475 ;
        RECT 67.605 168.845 68.725 169.015 ;
        RECT 68.895 168.845 69.205 169.645 ;
        RECT 67.605 168.595 67.865 168.845 ;
        RECT 69.375 168.675 69.685 169.475 ;
        RECT 55.115 167.265 55.445 167.895 ;
        RECT 55.615 167.095 55.825 167.915 ;
        RECT 56.205 167.095 56.535 167.895 ;
        RECT 56.705 167.745 57.715 167.915 ;
        RECT 57.920 167.745 58.555 167.915 ;
        RECT 56.705 167.265 56.875 167.745 ;
        RECT 57.045 167.095 57.375 167.575 ;
        RECT 57.545 167.265 57.715 167.745 ;
        RECT 57.965 167.095 58.205 167.575 ;
        RECT 58.385 167.265 58.555 167.745 ;
        RECT 58.965 167.095 59.295 167.895 ;
        RECT 59.465 167.745 60.475 167.915 ;
        RECT 60.680 167.745 61.315 167.915 ;
        RECT 59.465 167.265 59.635 167.745 ;
        RECT 59.805 167.095 60.135 167.575 ;
        RECT 60.305 167.265 60.475 167.745 ;
        RECT 60.725 167.095 60.965 167.575 ;
        RECT 61.145 167.265 61.315 167.745 ;
        RECT 65.000 167.640 65.340 168.470 ;
        RECT 67.110 168.425 67.865 168.595 ;
        RECT 68.655 168.505 69.685 168.675 ;
        RECT 67.110 167.915 67.515 168.425 ;
        RECT 68.655 168.255 68.825 168.505 ;
        RECT 67.685 168.085 68.825 168.255 ;
        RECT 67.110 167.745 68.760 167.915 ;
        RECT 68.995 167.765 69.345 168.335 ;
        RECT 61.580 167.095 66.925 167.640 ;
        RECT 67.155 167.095 67.435 167.575 ;
        RECT 67.605 167.355 67.865 167.745 ;
        RECT 68.040 167.095 68.295 167.575 ;
        RECT 68.465 167.355 68.760 167.745 ;
        RECT 69.515 167.595 69.685 168.505 ;
        RECT 68.940 167.095 69.215 167.575 ;
        RECT 69.385 167.265 69.685 167.595 ;
        RECT 69.855 168.570 70.125 169.475 ;
        RECT 70.295 168.885 70.625 169.645 ;
        RECT 70.805 168.715 70.975 169.475 ;
        RECT 69.855 167.770 70.025 168.570 ;
        RECT 70.310 168.545 70.975 168.715 ;
        RECT 70.310 168.400 70.480 168.545 ;
        RECT 71.240 168.495 71.500 169.645 ;
        RECT 71.675 168.570 71.930 169.475 ;
        RECT 72.100 168.885 72.430 169.645 ;
        RECT 72.645 168.715 72.815 169.475 ;
        RECT 70.195 168.070 70.480 168.400 ;
        RECT 70.310 167.815 70.480 168.070 ;
        RECT 70.715 167.995 71.045 168.365 ;
        RECT 69.855 167.265 70.115 167.770 ;
        RECT 70.310 167.645 70.975 167.815 ;
        RECT 70.295 167.095 70.625 167.475 ;
        RECT 70.805 167.265 70.975 167.645 ;
        RECT 71.240 167.095 71.500 167.935 ;
        RECT 71.675 167.840 71.845 168.570 ;
        RECT 72.100 168.545 72.815 168.715 ;
        RECT 72.100 168.335 72.270 168.545 ;
        RECT 73.995 168.480 74.285 169.645 ;
        RECT 74.455 168.555 77.965 169.645 ;
        RECT 78.140 169.210 83.485 169.645 ;
        RECT 72.015 168.005 72.270 168.335 ;
        RECT 71.675 167.265 71.930 167.840 ;
        RECT 72.100 167.815 72.270 168.005 ;
        RECT 72.550 167.995 72.905 168.365 ;
        RECT 74.455 168.035 76.145 168.555 ;
        RECT 76.315 167.865 77.965 168.385 ;
        RECT 79.730 167.960 80.080 169.210 ;
        RECT 83.665 168.835 83.960 169.645 ;
        RECT 72.100 167.645 72.815 167.815 ;
        RECT 72.100 167.095 72.430 167.475 ;
        RECT 72.645 167.265 72.815 167.645 ;
        RECT 73.995 167.095 74.285 167.820 ;
        RECT 74.455 167.095 77.965 167.865 ;
        RECT 81.560 167.640 81.900 168.470 ;
        RECT 84.140 168.335 84.385 169.475 ;
        RECT 84.560 168.835 84.820 169.645 ;
        RECT 85.420 169.640 91.695 169.645 ;
        RECT 85.000 168.335 85.250 169.470 ;
        RECT 85.420 168.845 85.680 169.640 ;
        RECT 85.850 168.745 86.110 169.470 ;
        RECT 86.280 168.915 86.540 169.640 ;
        RECT 86.710 168.745 86.970 169.470 ;
        RECT 87.140 168.915 87.400 169.640 ;
        RECT 87.570 168.745 87.830 169.470 ;
        RECT 88.000 168.915 88.260 169.640 ;
        RECT 88.430 168.745 88.690 169.470 ;
        RECT 88.860 168.915 89.105 169.640 ;
        RECT 89.275 168.745 89.535 169.470 ;
        RECT 89.720 168.915 89.965 169.640 ;
        RECT 90.135 168.745 90.395 169.470 ;
        RECT 90.580 168.915 90.825 169.640 ;
        RECT 90.995 168.745 91.255 169.470 ;
        RECT 91.440 168.915 91.695 169.640 ;
        RECT 85.850 168.730 91.255 168.745 ;
        RECT 91.865 168.730 92.155 169.470 ;
        RECT 92.325 168.900 92.595 169.645 ;
        RECT 85.850 168.505 92.595 168.730 ;
        RECT 93.835 168.505 94.045 169.645 ;
        RECT 83.655 167.775 83.970 168.335 ;
        RECT 84.140 168.085 91.260 168.335 ;
        RECT 78.140 167.095 83.485 167.640 ;
        RECT 83.655 167.095 83.960 167.605 ;
        RECT 84.140 167.275 84.390 168.085 ;
        RECT 84.560 167.095 84.820 167.620 ;
        RECT 85.000 167.275 85.250 168.085 ;
        RECT 91.430 167.915 92.595 168.505 ;
        RECT 94.215 168.495 94.545 169.475 ;
        RECT 94.715 168.505 94.945 169.645 ;
        RECT 95.155 168.885 95.670 169.295 ;
        RECT 95.905 168.885 96.075 169.645 ;
        RECT 96.245 169.305 98.275 169.475 ;
        RECT 85.850 167.745 92.595 167.915 ;
        RECT 85.420 167.095 85.680 167.655 ;
        RECT 85.850 167.290 86.110 167.745 ;
        RECT 86.280 167.095 86.540 167.575 ;
        RECT 86.710 167.290 86.970 167.745 ;
        RECT 87.140 167.095 87.400 167.575 ;
        RECT 87.570 167.290 87.830 167.745 ;
        RECT 88.000 167.095 88.245 167.575 ;
        RECT 88.415 167.290 88.690 167.745 ;
        RECT 88.860 167.095 89.105 167.575 ;
        RECT 89.275 167.290 89.535 167.745 ;
        RECT 89.715 167.095 89.965 167.575 ;
        RECT 90.135 167.290 90.395 167.745 ;
        RECT 90.575 167.095 90.825 167.575 ;
        RECT 90.995 167.290 91.255 167.745 ;
        RECT 91.435 167.095 91.695 167.575 ;
        RECT 91.865 167.290 92.125 167.745 ;
        RECT 92.295 167.095 92.595 167.575 ;
        RECT 93.835 167.095 94.045 167.915 ;
        RECT 94.215 167.895 94.465 168.495 ;
        RECT 94.635 168.085 94.965 168.335 ;
        RECT 95.155 168.075 95.495 168.885 ;
        RECT 96.245 168.640 96.415 169.305 ;
        RECT 96.810 168.965 97.935 169.135 ;
        RECT 95.665 168.450 96.415 168.640 ;
        RECT 96.585 168.625 97.595 168.795 ;
        RECT 94.215 167.265 94.545 167.895 ;
        RECT 94.715 167.095 94.945 167.915 ;
        RECT 95.155 167.905 96.385 168.075 ;
        RECT 95.430 167.300 95.675 167.905 ;
        RECT 95.895 167.095 96.405 167.630 ;
        RECT 96.585 167.265 96.775 168.625 ;
        RECT 96.945 167.945 97.220 168.425 ;
        RECT 96.945 167.775 97.225 167.945 ;
        RECT 97.425 167.825 97.595 168.625 ;
        RECT 97.765 167.835 97.935 168.965 ;
        RECT 98.105 168.335 98.275 169.305 ;
        RECT 98.445 168.505 98.615 169.645 ;
        RECT 98.785 168.505 99.120 169.475 ;
        RECT 98.105 168.005 98.300 168.335 ;
        RECT 98.525 168.005 98.780 168.335 ;
        RECT 98.525 167.835 98.695 168.005 ;
        RECT 98.950 167.835 99.120 168.505 ;
        RECT 99.755 168.480 100.045 169.645 ;
        RECT 101.340 168.675 101.670 169.475 ;
        RECT 101.840 168.845 102.170 169.645 ;
        RECT 102.470 168.675 102.800 169.475 ;
        RECT 103.445 168.845 103.695 169.645 ;
        RECT 101.340 168.505 103.775 168.675 ;
        RECT 103.965 168.505 104.135 169.645 ;
        RECT 104.305 168.505 104.645 169.475 ;
        RECT 101.135 168.085 101.485 168.335 ;
        RECT 101.670 167.875 101.840 168.505 ;
        RECT 102.010 168.085 102.340 168.285 ;
        RECT 102.510 168.085 102.840 168.285 ;
        RECT 103.010 168.085 103.430 168.285 ;
        RECT 103.605 168.255 103.775 168.505 ;
        RECT 103.605 168.085 104.300 168.255 ;
        RECT 96.945 167.265 97.220 167.775 ;
        RECT 97.765 167.665 98.695 167.835 ;
        RECT 97.765 167.630 97.940 167.665 ;
        RECT 97.410 167.265 97.940 167.630 ;
        RECT 98.365 167.095 98.695 167.495 ;
        RECT 98.865 167.265 99.120 167.835 ;
        RECT 99.755 167.095 100.045 167.820 ;
        RECT 101.340 167.265 101.840 167.875 ;
        RECT 102.470 167.745 103.695 167.915 ;
        RECT 104.470 167.895 104.645 168.505 ;
        RECT 104.815 168.555 106.485 169.645 ;
        RECT 104.815 168.035 105.565 168.555 ;
        RECT 106.695 168.505 106.925 169.645 ;
        RECT 107.095 168.495 107.425 169.475 ;
        RECT 107.595 168.505 107.805 169.645 ;
        RECT 102.470 167.265 102.800 167.745 ;
        RECT 102.970 167.095 103.195 167.555 ;
        RECT 103.365 167.265 103.695 167.745 ;
        RECT 103.885 167.095 104.135 167.895 ;
        RECT 104.305 167.265 104.645 167.895 ;
        RECT 105.735 167.865 106.485 168.385 ;
        RECT 106.675 168.085 107.005 168.335 ;
        RECT 104.815 167.095 106.485 167.865 ;
        RECT 106.695 167.095 106.925 167.915 ;
        RECT 107.175 167.895 107.425 168.495 ;
        RECT 108.040 168.455 108.295 169.335 ;
        RECT 108.465 168.505 108.770 169.645 ;
        RECT 109.110 169.265 109.440 169.645 ;
        RECT 109.620 169.095 109.790 169.385 ;
        RECT 109.960 169.185 110.210 169.645 ;
        RECT 108.990 168.925 109.790 169.095 ;
        RECT 110.380 169.135 111.250 169.475 ;
        RECT 107.095 167.265 107.425 167.895 ;
        RECT 107.595 167.095 107.805 167.915 ;
        RECT 108.040 167.805 108.250 168.455 ;
        RECT 108.990 168.335 109.160 168.925 ;
        RECT 110.380 168.755 110.550 169.135 ;
        RECT 111.485 169.015 111.655 169.475 ;
        RECT 111.825 169.185 112.195 169.645 ;
        RECT 112.490 169.045 112.660 169.385 ;
        RECT 112.830 169.215 113.160 169.645 ;
        RECT 113.395 169.045 113.565 169.385 ;
        RECT 109.330 168.585 110.550 168.755 ;
        RECT 110.720 168.675 111.180 168.965 ;
        RECT 111.485 168.845 112.045 169.015 ;
        RECT 112.490 168.875 113.565 169.045 ;
        RECT 113.735 169.145 114.415 169.475 ;
        RECT 114.630 169.145 114.880 169.475 ;
        RECT 115.050 169.185 115.300 169.645 ;
        RECT 111.875 168.705 112.045 168.845 ;
        RECT 110.720 168.665 111.685 168.675 ;
        RECT 110.380 168.495 110.550 168.585 ;
        RECT 111.010 168.505 111.685 168.665 ;
        RECT 108.420 168.305 109.160 168.335 ;
        RECT 108.420 168.005 109.335 168.305 ;
        RECT 109.010 167.830 109.335 168.005 ;
        RECT 108.040 167.275 108.295 167.805 ;
        RECT 108.465 167.095 108.770 167.555 ;
        RECT 109.015 167.475 109.335 167.830 ;
        RECT 109.505 168.045 110.045 168.415 ;
        RECT 110.380 168.325 110.785 168.495 ;
        RECT 109.505 167.645 109.745 168.045 ;
        RECT 110.225 167.875 110.445 168.155 ;
        RECT 109.915 167.705 110.445 167.875 ;
        RECT 109.915 167.475 110.085 167.705 ;
        RECT 110.615 167.545 110.785 168.325 ;
        RECT 110.955 167.715 111.305 168.335 ;
        RECT 111.475 167.715 111.685 168.505 ;
        RECT 111.875 168.535 113.375 168.705 ;
        RECT 111.875 167.845 112.045 168.535 ;
        RECT 113.735 168.365 113.905 169.145 ;
        RECT 114.710 169.015 114.880 169.145 ;
        RECT 112.215 168.195 113.905 168.365 ;
        RECT 114.075 168.585 114.540 168.975 ;
        RECT 114.710 168.845 115.105 169.015 ;
        RECT 112.215 168.015 112.385 168.195 ;
        RECT 109.015 167.305 110.085 167.475 ;
        RECT 110.255 167.095 110.445 167.535 ;
        RECT 110.615 167.265 111.565 167.545 ;
        RECT 111.875 167.455 112.135 167.845 ;
        RECT 112.555 167.775 113.345 168.025 ;
        RECT 111.785 167.285 112.135 167.455 ;
        RECT 112.345 167.095 112.675 167.555 ;
        RECT 113.550 167.485 113.720 168.195 ;
        RECT 114.075 167.995 114.245 168.585 ;
        RECT 113.890 167.775 114.245 167.995 ;
        RECT 114.415 167.775 114.765 168.395 ;
        RECT 114.935 167.485 115.105 168.845 ;
        RECT 115.470 168.675 115.795 169.460 ;
        RECT 115.275 167.625 115.735 168.675 ;
        RECT 113.550 167.315 114.405 167.485 ;
        RECT 114.610 167.315 115.105 167.485 ;
        RECT 115.275 167.095 115.605 167.455 ;
        RECT 115.965 167.355 116.135 169.475 ;
        RECT 116.305 169.145 116.635 169.645 ;
        RECT 116.805 168.975 117.060 169.475 ;
        RECT 116.310 168.805 117.060 168.975 ;
        RECT 116.310 167.815 116.540 168.805 ;
        RECT 116.710 167.985 117.060 168.635 ;
        RECT 117.235 168.570 117.505 169.475 ;
        RECT 117.675 168.885 118.005 169.645 ;
        RECT 118.185 168.715 118.355 169.475 ;
        RECT 119.080 169.210 124.425 169.645 ;
        RECT 116.310 167.645 117.060 167.815 ;
        RECT 116.305 167.095 116.635 167.475 ;
        RECT 116.805 167.355 117.060 167.645 ;
        RECT 117.235 167.770 117.405 168.570 ;
        RECT 117.690 168.545 118.355 168.715 ;
        RECT 117.690 168.400 117.860 168.545 ;
        RECT 117.575 168.070 117.860 168.400 ;
        RECT 117.690 167.815 117.860 168.070 ;
        RECT 118.095 167.995 118.425 168.365 ;
        RECT 120.670 167.960 121.020 169.210 ;
        RECT 124.595 168.555 125.805 169.645 ;
        RECT 117.235 167.265 117.495 167.770 ;
        RECT 117.690 167.645 118.355 167.815 ;
        RECT 117.675 167.095 118.005 167.475 ;
        RECT 118.185 167.265 118.355 167.645 ;
        RECT 122.500 167.640 122.840 168.470 ;
        RECT 124.595 168.015 125.115 168.555 ;
        RECT 125.285 167.845 125.805 168.385 ;
        RECT 119.080 167.095 124.425 167.640 ;
        RECT 124.595 167.095 125.805 167.845 ;
        RECT 11.810 166.925 125.890 167.095 ;
        RECT 11.895 166.175 13.105 166.925 ;
        RECT 13.275 166.175 14.485 166.925 ;
        RECT 14.660 166.380 20.005 166.925 ;
        RECT 11.895 165.635 12.415 166.175 ;
        RECT 12.585 165.465 13.105 166.005 ;
        RECT 11.895 164.375 13.105 165.465 ;
        RECT 13.275 165.465 13.795 166.005 ;
        RECT 13.965 165.635 14.485 166.175 ;
        RECT 13.275 164.375 14.485 165.465 ;
        RECT 16.250 164.810 16.600 166.060 ;
        RECT 18.080 165.550 18.420 166.380 ;
        RECT 20.265 166.375 20.435 166.755 ;
        RECT 20.615 166.545 20.945 166.925 ;
        RECT 20.265 166.205 20.930 166.375 ;
        RECT 21.125 166.250 21.385 166.755 ;
        RECT 20.195 165.655 20.525 166.025 ;
        RECT 20.760 165.950 20.930 166.205 ;
        RECT 20.760 165.620 21.045 165.950 ;
        RECT 20.760 165.475 20.930 165.620 ;
        RECT 20.265 165.305 20.930 165.475 ;
        RECT 21.215 165.450 21.385 166.250 ;
        RECT 14.660 164.375 20.005 164.810 ;
        RECT 20.265 164.545 20.435 165.305 ;
        RECT 20.615 164.375 20.945 165.135 ;
        RECT 21.115 164.545 21.385 165.450 ;
        RECT 21.560 166.185 21.815 166.755 ;
        RECT 21.985 166.525 22.315 166.925 ;
        RECT 22.740 166.390 23.270 166.755 ;
        RECT 22.740 166.355 22.915 166.390 ;
        RECT 21.985 166.185 22.915 166.355 ;
        RECT 21.560 165.515 21.730 166.185 ;
        RECT 21.985 166.015 22.155 166.185 ;
        RECT 21.900 165.685 22.155 166.015 ;
        RECT 22.380 165.685 22.575 166.015 ;
        RECT 21.560 164.545 21.895 165.515 ;
        RECT 22.065 164.375 22.235 165.515 ;
        RECT 22.405 164.715 22.575 165.685 ;
        RECT 22.745 165.055 22.915 166.185 ;
        RECT 23.085 165.395 23.255 166.195 ;
        RECT 23.460 165.905 23.735 166.755 ;
        RECT 23.455 165.735 23.735 165.905 ;
        RECT 23.460 165.595 23.735 165.735 ;
        RECT 23.905 165.395 24.095 166.755 ;
        RECT 24.275 166.390 24.785 166.925 ;
        RECT 25.005 166.115 25.250 166.720 ;
        RECT 25.700 166.215 25.955 166.745 ;
        RECT 26.125 166.465 26.430 166.925 ;
        RECT 26.675 166.545 27.745 166.715 ;
        RECT 24.295 165.945 25.525 166.115 ;
        RECT 23.085 165.225 24.095 165.395 ;
        RECT 24.265 165.380 25.015 165.570 ;
        RECT 22.745 164.885 23.870 165.055 ;
        RECT 24.265 164.715 24.435 165.380 ;
        RECT 25.185 165.135 25.525 165.945 ;
        RECT 22.405 164.545 24.435 164.715 ;
        RECT 24.605 164.375 24.775 165.135 ;
        RECT 25.010 164.725 25.525 165.135 ;
        RECT 25.700 165.565 25.910 166.215 ;
        RECT 26.675 166.190 26.995 166.545 ;
        RECT 26.670 166.015 26.995 166.190 ;
        RECT 26.080 165.715 26.995 166.015 ;
        RECT 27.165 165.975 27.405 166.375 ;
        RECT 27.575 166.315 27.745 166.545 ;
        RECT 27.915 166.485 28.105 166.925 ;
        RECT 28.275 166.475 29.225 166.755 ;
        RECT 29.445 166.565 29.795 166.735 ;
        RECT 27.575 166.145 28.105 166.315 ;
        RECT 26.080 165.685 26.820 165.715 ;
        RECT 25.700 164.685 25.955 165.565 ;
        RECT 26.125 164.375 26.430 165.515 ;
        RECT 26.650 165.095 26.820 165.685 ;
        RECT 27.165 165.605 27.705 165.975 ;
        RECT 27.885 165.865 28.105 166.145 ;
        RECT 28.275 165.695 28.445 166.475 ;
        RECT 28.040 165.525 28.445 165.695 ;
        RECT 28.615 165.685 28.965 166.305 ;
        RECT 28.040 165.435 28.210 165.525 ;
        RECT 29.135 165.515 29.345 166.305 ;
        RECT 26.990 165.265 28.210 165.435 ;
        RECT 28.670 165.355 29.345 165.515 ;
        RECT 26.650 164.925 27.450 165.095 ;
        RECT 26.770 164.375 27.100 164.755 ;
        RECT 27.280 164.635 27.450 164.925 ;
        RECT 28.040 164.885 28.210 165.265 ;
        RECT 28.380 165.345 29.345 165.355 ;
        RECT 29.535 166.175 29.795 166.565 ;
        RECT 30.005 166.465 30.335 166.925 ;
        RECT 31.210 166.535 32.065 166.705 ;
        RECT 32.270 166.535 32.765 166.705 ;
        RECT 32.935 166.565 33.265 166.925 ;
        RECT 29.535 165.485 29.705 166.175 ;
        RECT 29.875 165.825 30.045 166.005 ;
        RECT 30.215 165.995 31.005 166.245 ;
        RECT 31.210 165.825 31.380 166.535 ;
        RECT 31.550 166.025 31.905 166.245 ;
        RECT 29.875 165.655 31.565 165.825 ;
        RECT 28.380 165.055 28.840 165.345 ;
        RECT 29.535 165.315 31.035 165.485 ;
        RECT 29.535 165.175 29.705 165.315 ;
        RECT 29.145 165.005 29.705 165.175 ;
        RECT 27.620 164.375 27.870 164.835 ;
        RECT 28.040 164.545 28.910 164.885 ;
        RECT 29.145 164.545 29.315 165.005 ;
        RECT 30.150 164.975 31.225 165.145 ;
        RECT 29.485 164.375 29.855 164.835 ;
        RECT 30.150 164.635 30.320 164.975 ;
        RECT 30.490 164.375 30.820 164.805 ;
        RECT 31.055 164.635 31.225 164.975 ;
        RECT 31.395 164.875 31.565 165.655 ;
        RECT 31.735 165.435 31.905 166.025 ;
        RECT 32.075 165.625 32.425 166.245 ;
        RECT 31.735 165.045 32.200 165.435 ;
        RECT 32.595 165.175 32.765 166.535 ;
        RECT 32.935 165.345 33.395 166.395 ;
        RECT 32.370 165.005 32.765 165.175 ;
        RECT 32.370 164.875 32.540 165.005 ;
        RECT 31.395 164.545 32.075 164.875 ;
        RECT 32.290 164.545 32.540 164.875 ;
        RECT 32.710 164.375 32.960 164.835 ;
        RECT 33.130 164.560 33.455 165.345 ;
        RECT 33.625 164.545 33.795 166.665 ;
        RECT 33.965 166.545 34.295 166.925 ;
        RECT 34.465 166.375 34.720 166.665 ;
        RECT 33.970 166.205 34.720 166.375 ;
        RECT 33.970 165.215 34.200 166.205 ;
        RECT 35.355 166.200 35.645 166.925 ;
        RECT 35.815 166.155 37.485 166.925 ;
        RECT 34.370 165.385 34.720 166.035 ;
        RECT 33.970 165.045 34.720 165.215 ;
        RECT 33.965 164.375 34.295 164.875 ;
        RECT 34.465 164.545 34.720 165.045 ;
        RECT 35.355 164.375 35.645 165.540 ;
        RECT 35.815 165.465 36.565 165.985 ;
        RECT 36.735 165.635 37.485 166.155 ;
        RECT 37.655 166.125 37.995 166.755 ;
        RECT 38.165 166.125 38.415 166.925 ;
        RECT 38.605 166.275 38.935 166.755 ;
        RECT 39.105 166.465 39.330 166.925 ;
        RECT 39.500 166.275 39.830 166.755 ;
        RECT 37.655 165.515 37.830 166.125 ;
        RECT 38.605 166.105 39.830 166.275 ;
        RECT 40.460 166.145 40.960 166.755 ;
        RECT 38.000 165.765 38.695 165.935 ;
        RECT 38.525 165.515 38.695 165.765 ;
        RECT 38.870 165.735 39.290 165.935 ;
        RECT 39.460 165.735 39.790 165.935 ;
        RECT 39.960 165.735 40.290 165.935 ;
        RECT 40.460 165.515 40.630 166.145 ;
        RECT 42.255 166.125 42.595 166.755 ;
        RECT 42.765 166.125 43.015 166.925 ;
        RECT 43.205 166.275 43.535 166.755 ;
        RECT 43.705 166.465 43.930 166.925 ;
        RECT 44.100 166.275 44.430 166.755 ;
        RECT 40.815 165.685 41.165 165.935 ;
        RECT 42.255 165.515 42.430 166.125 ;
        RECT 43.205 166.105 44.430 166.275 ;
        RECT 45.060 166.145 45.560 166.755 ;
        RECT 42.600 165.765 43.295 165.935 ;
        RECT 43.125 165.515 43.295 165.765 ;
        RECT 43.470 165.735 43.890 165.935 ;
        RECT 44.060 165.735 44.390 165.935 ;
        RECT 44.560 165.735 44.890 165.935 ;
        RECT 45.060 165.515 45.230 166.145 ;
        RECT 45.935 166.125 46.275 166.755 ;
        RECT 46.445 166.125 46.695 166.925 ;
        RECT 46.885 166.275 47.215 166.755 ;
        RECT 47.385 166.465 47.610 166.925 ;
        RECT 47.780 166.275 48.110 166.755 ;
        RECT 45.415 165.685 45.765 165.935 ;
        RECT 45.935 165.515 46.110 166.125 ;
        RECT 46.885 166.105 48.110 166.275 ;
        RECT 48.740 166.145 49.240 166.755 ;
        RECT 49.615 166.155 51.285 166.925 ;
        RECT 51.830 166.585 52.085 166.745 ;
        RECT 51.745 166.415 52.085 166.585 ;
        RECT 52.265 166.465 52.550 166.925 ;
        RECT 46.280 165.765 46.975 165.935 ;
        RECT 46.805 165.515 46.975 165.765 ;
        RECT 47.150 165.735 47.570 165.935 ;
        RECT 47.740 165.735 48.070 165.935 ;
        RECT 48.240 165.735 48.570 165.935 ;
        RECT 48.740 165.515 48.910 166.145 ;
        RECT 49.095 165.685 49.445 165.935 ;
        RECT 35.815 164.375 37.485 165.465 ;
        RECT 37.655 164.545 37.995 165.515 ;
        RECT 38.165 164.375 38.335 165.515 ;
        RECT 38.525 165.345 40.960 165.515 ;
        RECT 38.605 164.375 38.855 165.175 ;
        RECT 39.500 164.545 39.830 165.345 ;
        RECT 40.130 164.375 40.460 165.175 ;
        RECT 40.630 164.545 40.960 165.345 ;
        RECT 42.255 164.545 42.595 165.515 ;
        RECT 42.765 164.375 42.935 165.515 ;
        RECT 43.125 165.345 45.560 165.515 ;
        RECT 43.205 164.375 43.455 165.175 ;
        RECT 44.100 164.545 44.430 165.345 ;
        RECT 44.730 164.375 45.060 165.175 ;
        RECT 45.230 164.545 45.560 165.345 ;
        RECT 45.935 164.545 46.275 165.515 ;
        RECT 46.445 164.375 46.615 165.515 ;
        RECT 46.805 165.345 49.240 165.515 ;
        RECT 46.885 164.375 47.135 165.175 ;
        RECT 47.780 164.545 48.110 165.345 ;
        RECT 48.410 164.375 48.740 165.175 ;
        RECT 48.910 164.545 49.240 165.345 ;
        RECT 49.615 165.465 50.365 165.985 ;
        RECT 50.535 165.635 51.285 166.155 ;
        RECT 51.830 166.215 52.085 166.415 ;
        RECT 49.615 164.375 51.285 165.465 ;
        RECT 51.830 165.355 52.010 166.215 ;
        RECT 52.730 166.015 52.980 166.665 ;
        RECT 52.180 165.685 52.980 166.015 ;
        RECT 51.830 164.685 52.085 165.355 ;
        RECT 52.265 164.375 52.550 165.175 ;
        RECT 52.730 165.095 52.980 165.685 ;
        RECT 53.180 166.330 53.500 166.660 ;
        RECT 53.680 166.445 54.340 166.925 ;
        RECT 54.540 166.535 55.390 166.705 ;
        RECT 53.180 165.435 53.370 166.330 ;
        RECT 53.690 166.005 54.350 166.275 ;
        RECT 54.020 165.945 54.350 166.005 ;
        RECT 53.540 165.775 53.870 165.835 ;
        RECT 54.540 165.775 54.710 166.535 ;
        RECT 55.950 166.465 56.270 166.925 ;
        RECT 56.470 166.285 56.720 166.715 ;
        RECT 57.010 166.485 57.420 166.925 ;
        RECT 57.590 166.545 58.605 166.745 ;
        RECT 54.880 166.115 56.130 166.285 ;
        RECT 54.880 165.995 55.210 166.115 ;
        RECT 53.540 165.605 55.440 165.775 ;
        RECT 53.180 165.265 55.100 165.435 ;
        RECT 53.180 165.245 53.500 165.265 ;
        RECT 52.730 164.585 53.060 165.095 ;
        RECT 53.330 164.635 53.500 165.245 ;
        RECT 55.270 165.095 55.440 165.605 ;
        RECT 55.610 165.535 55.790 165.945 ;
        RECT 55.960 165.355 56.130 166.115 ;
        RECT 53.670 164.375 54.000 165.065 ;
        RECT 54.230 164.925 55.440 165.095 ;
        RECT 55.610 165.045 56.130 165.355 ;
        RECT 56.300 165.945 56.720 166.285 ;
        RECT 57.010 165.945 57.420 166.275 ;
        RECT 56.300 165.175 56.490 165.945 ;
        RECT 57.590 165.815 57.760 166.545 ;
        RECT 58.905 166.375 59.075 166.705 ;
        RECT 59.245 166.545 59.575 166.925 ;
        RECT 57.930 165.995 58.280 166.365 ;
        RECT 57.590 165.775 58.010 165.815 ;
        RECT 56.660 165.605 58.010 165.775 ;
        RECT 56.660 165.445 56.910 165.605 ;
        RECT 57.420 165.175 57.670 165.435 ;
        RECT 56.300 164.925 57.670 165.175 ;
        RECT 54.230 164.635 54.470 164.925 ;
        RECT 55.270 164.845 55.440 164.925 ;
        RECT 54.670 164.375 55.090 164.755 ;
        RECT 55.270 164.595 55.900 164.845 ;
        RECT 56.370 164.375 56.700 164.755 ;
        RECT 56.870 164.635 57.040 164.925 ;
        RECT 57.840 164.760 58.010 165.605 ;
        RECT 58.460 165.435 58.680 166.305 ;
        RECT 58.905 166.185 59.600 166.375 ;
        RECT 58.180 165.055 58.680 165.435 ;
        RECT 58.850 165.385 59.260 166.005 ;
        RECT 59.430 165.215 59.600 166.185 ;
        RECT 58.905 165.045 59.600 165.215 ;
        RECT 57.220 164.375 57.600 164.755 ;
        RECT 57.840 164.590 58.670 164.760 ;
        RECT 58.905 164.545 59.075 165.045 ;
        RECT 59.245 164.375 59.575 164.875 ;
        RECT 59.790 164.545 60.015 166.665 ;
        RECT 60.185 166.545 60.515 166.925 ;
        RECT 60.685 166.375 60.855 166.665 ;
        RECT 60.190 166.205 60.855 166.375 ;
        RECT 60.190 165.215 60.420 166.205 ;
        RECT 61.115 166.200 61.405 166.925 ;
        RECT 61.575 166.250 61.835 166.755 ;
        RECT 62.015 166.545 62.345 166.925 ;
        RECT 62.525 166.375 62.695 166.755 ;
        RECT 63.015 166.445 63.295 166.925 ;
        RECT 60.590 165.385 60.940 166.035 ;
        RECT 60.190 165.045 60.855 165.215 ;
        RECT 60.185 164.375 60.515 164.875 ;
        RECT 60.685 164.545 60.855 165.045 ;
        RECT 61.115 164.375 61.405 165.540 ;
        RECT 61.575 165.450 61.745 166.250 ;
        RECT 62.030 166.205 62.695 166.375 ;
        RECT 63.465 166.275 63.725 166.665 ;
        RECT 63.900 166.445 64.155 166.925 ;
        RECT 64.325 166.275 64.620 166.665 ;
        RECT 64.800 166.445 65.075 166.925 ;
        RECT 65.245 166.425 65.545 166.755 ;
        RECT 62.030 165.950 62.200 166.205 ;
        RECT 62.970 166.105 64.620 166.275 ;
        RECT 61.915 165.620 62.200 165.950 ;
        RECT 62.435 165.655 62.765 166.025 ;
        RECT 62.030 165.475 62.200 165.620 ;
        RECT 62.970 165.595 63.375 166.105 ;
        RECT 63.545 165.765 64.685 165.935 ;
        RECT 61.575 164.545 61.845 165.450 ;
        RECT 62.030 165.305 62.695 165.475 ;
        RECT 62.970 165.425 63.725 165.595 ;
        RECT 62.015 164.375 62.345 165.135 ;
        RECT 62.525 164.545 62.695 165.305 ;
        RECT 63.010 164.375 63.295 165.245 ;
        RECT 63.465 165.175 63.725 165.425 ;
        RECT 64.515 165.515 64.685 165.765 ;
        RECT 64.855 165.685 65.205 166.255 ;
        RECT 65.375 165.515 65.545 166.425 ;
        RECT 66.175 166.155 67.845 166.925 ;
        RECT 64.515 165.345 65.545 165.515 ;
        RECT 63.465 165.005 64.585 165.175 ;
        RECT 63.465 164.545 63.725 165.005 ;
        RECT 63.900 164.375 64.155 164.835 ;
        RECT 64.325 164.545 64.585 165.005 ;
        RECT 64.755 164.375 65.065 165.175 ;
        RECT 65.235 164.545 65.545 165.345 ;
        RECT 66.175 165.465 66.925 165.985 ;
        RECT 67.095 165.635 67.845 166.155 ;
        RECT 68.020 166.085 68.280 166.925 ;
        RECT 68.455 166.180 68.710 166.755 ;
        RECT 68.880 166.545 69.210 166.925 ;
        RECT 69.425 166.375 69.595 166.755 ;
        RECT 68.880 166.205 69.595 166.375 ;
        RECT 69.945 166.375 70.115 166.755 ;
        RECT 70.330 166.545 70.660 166.925 ;
        RECT 69.945 166.205 70.660 166.375 ;
        RECT 66.175 164.375 67.845 165.465 ;
        RECT 68.020 164.375 68.280 165.525 ;
        RECT 68.455 165.450 68.625 166.180 ;
        RECT 68.880 166.015 69.050 166.205 ;
        RECT 68.795 165.685 69.050 166.015 ;
        RECT 68.880 165.475 69.050 165.685 ;
        RECT 69.330 165.655 69.685 166.025 ;
        RECT 69.855 165.655 70.210 166.025 ;
        RECT 70.490 166.015 70.660 166.205 ;
        RECT 70.830 166.180 71.085 166.755 ;
        RECT 70.490 165.685 70.745 166.015 ;
        RECT 70.490 165.475 70.660 165.685 ;
        RECT 68.455 164.545 68.710 165.450 ;
        RECT 68.880 165.305 69.595 165.475 ;
        RECT 68.880 164.375 69.210 165.135 ;
        RECT 69.425 164.545 69.595 165.305 ;
        RECT 69.945 165.305 70.660 165.475 ;
        RECT 70.915 165.450 71.085 166.180 ;
        RECT 71.260 166.085 71.520 166.925 ;
        RECT 71.695 166.165 72.405 166.755 ;
        RECT 72.915 166.395 73.245 166.755 ;
        RECT 73.445 166.565 73.775 166.925 ;
        RECT 73.945 166.395 74.275 166.755 ;
        RECT 72.915 166.185 74.275 166.395 ;
        RECT 74.455 166.250 74.715 166.755 ;
        RECT 74.895 166.545 75.225 166.925 ;
        RECT 75.405 166.375 75.575 166.755 ;
        RECT 69.945 164.545 70.115 165.305 ;
        RECT 70.330 164.375 70.660 165.135 ;
        RECT 70.830 164.545 71.085 165.450 ;
        RECT 71.260 164.375 71.520 165.525 ;
        RECT 71.695 165.195 71.900 166.165 ;
        RECT 72.070 165.395 72.400 165.935 ;
        RECT 72.575 165.685 73.070 166.015 ;
        RECT 73.390 165.685 73.765 166.015 ;
        RECT 73.975 165.685 74.285 166.015 ;
        RECT 72.575 165.395 72.900 165.685 ;
        RECT 73.095 165.195 73.425 165.415 ;
        RECT 71.695 164.965 73.425 165.195 ;
        RECT 71.695 164.545 72.395 164.965 ;
        RECT 72.595 164.375 72.925 164.735 ;
        RECT 73.095 164.565 73.425 164.965 ;
        RECT 73.595 164.760 73.765 165.685 ;
        RECT 74.455 165.450 74.625 166.250 ;
        RECT 74.910 166.205 75.575 166.375 ;
        RECT 74.910 165.950 75.080 166.205 ;
        RECT 75.835 166.175 77.045 166.925 ;
        RECT 74.795 165.620 75.080 165.950 ;
        RECT 75.315 165.655 75.645 166.025 ;
        RECT 74.910 165.475 75.080 165.620 ;
        RECT 73.945 164.375 74.275 165.435 ;
        RECT 74.455 164.545 74.725 165.450 ;
        RECT 74.910 165.305 75.575 165.475 ;
        RECT 74.895 164.375 75.225 165.135 ;
        RECT 75.405 164.545 75.575 165.305 ;
        RECT 75.835 165.465 76.355 166.005 ;
        RECT 76.525 165.635 77.045 166.175 ;
        RECT 77.590 166.215 77.845 166.745 ;
        RECT 78.025 166.465 78.310 166.925 ;
        RECT 75.835 164.375 77.045 165.465 ;
        RECT 77.590 165.355 77.770 166.215 ;
        RECT 78.490 166.015 78.740 166.665 ;
        RECT 77.940 165.685 78.740 166.015 ;
        RECT 77.590 164.885 77.845 165.355 ;
        RECT 77.505 164.715 77.845 164.885 ;
        RECT 77.590 164.685 77.845 164.715 ;
        RECT 78.025 164.375 78.310 165.175 ;
        RECT 78.490 165.095 78.740 165.685 ;
        RECT 78.940 166.330 79.260 166.660 ;
        RECT 79.440 166.445 80.100 166.925 ;
        RECT 80.300 166.535 81.150 166.705 ;
        RECT 78.940 165.435 79.130 166.330 ;
        RECT 79.450 166.005 80.110 166.275 ;
        RECT 79.780 165.945 80.110 166.005 ;
        RECT 79.300 165.775 79.630 165.835 ;
        RECT 80.300 165.775 80.470 166.535 ;
        RECT 81.710 166.465 82.030 166.925 ;
        RECT 82.230 166.285 82.480 166.715 ;
        RECT 82.770 166.485 83.180 166.925 ;
        RECT 83.350 166.545 84.365 166.745 ;
        RECT 80.640 166.115 81.890 166.285 ;
        RECT 80.640 165.995 80.970 166.115 ;
        RECT 79.300 165.605 81.200 165.775 ;
        RECT 78.940 165.265 80.860 165.435 ;
        RECT 78.940 165.245 79.260 165.265 ;
        RECT 78.490 164.585 78.820 165.095 ;
        RECT 79.090 164.635 79.260 165.245 ;
        RECT 81.030 165.095 81.200 165.605 ;
        RECT 81.370 165.535 81.550 165.945 ;
        RECT 81.720 165.355 81.890 166.115 ;
        RECT 79.430 164.375 79.760 165.065 ;
        RECT 79.990 164.925 81.200 165.095 ;
        RECT 81.370 165.045 81.890 165.355 ;
        RECT 82.060 165.945 82.480 166.285 ;
        RECT 82.770 165.945 83.180 166.275 ;
        RECT 82.060 165.175 82.250 165.945 ;
        RECT 83.350 165.815 83.520 166.545 ;
        RECT 84.665 166.375 84.835 166.705 ;
        RECT 85.005 166.545 85.335 166.925 ;
        RECT 83.690 165.995 84.040 166.365 ;
        RECT 83.350 165.775 83.770 165.815 ;
        RECT 82.420 165.605 83.770 165.775 ;
        RECT 82.420 165.445 82.670 165.605 ;
        RECT 83.180 165.175 83.430 165.435 ;
        RECT 82.060 164.925 83.430 165.175 ;
        RECT 79.990 164.635 80.230 164.925 ;
        RECT 81.030 164.845 81.200 164.925 ;
        RECT 80.430 164.375 80.850 164.755 ;
        RECT 81.030 164.595 81.660 164.845 ;
        RECT 82.130 164.375 82.460 164.755 ;
        RECT 82.630 164.635 82.800 164.925 ;
        RECT 83.600 164.760 83.770 165.605 ;
        RECT 84.220 165.435 84.440 166.305 ;
        RECT 84.665 166.185 85.360 166.375 ;
        RECT 83.940 165.055 84.440 165.435 ;
        RECT 84.610 165.385 85.020 166.005 ;
        RECT 85.190 165.215 85.360 166.185 ;
        RECT 84.665 165.045 85.360 165.215 ;
        RECT 82.980 164.375 83.360 164.755 ;
        RECT 83.600 164.590 84.430 164.760 ;
        RECT 84.665 164.545 84.835 165.045 ;
        RECT 85.005 164.375 85.335 164.875 ;
        RECT 85.550 164.545 85.775 166.665 ;
        RECT 85.945 166.545 86.275 166.925 ;
        RECT 86.445 166.375 86.615 166.665 ;
        RECT 85.950 166.205 86.615 166.375 ;
        RECT 85.950 165.215 86.180 166.205 ;
        RECT 86.875 166.200 87.165 166.925 ;
        RECT 88.040 166.445 88.340 166.925 ;
        RECT 88.510 166.275 88.770 166.730 ;
        RECT 88.940 166.445 89.200 166.925 ;
        RECT 89.370 166.275 89.630 166.730 ;
        RECT 89.800 166.445 90.060 166.925 ;
        RECT 90.230 166.275 90.490 166.730 ;
        RECT 90.660 166.445 90.920 166.925 ;
        RECT 91.090 166.275 91.350 166.730 ;
        RECT 91.520 166.400 91.780 166.925 ;
        RECT 88.040 166.105 91.350 166.275 ;
        RECT 86.350 165.385 86.700 166.035 ;
        RECT 85.950 165.045 86.615 165.215 ;
        RECT 85.945 164.375 86.275 164.875 ;
        RECT 86.445 164.545 86.615 165.045 ;
        RECT 86.875 164.375 87.165 165.540 ;
        RECT 88.040 165.515 89.010 166.105 ;
        RECT 91.950 165.935 92.200 166.745 ;
        RECT 92.380 166.465 92.625 166.925 ;
        RECT 89.180 165.685 92.200 165.935 ;
        RECT 92.370 165.685 92.685 166.295 ;
        RECT 92.855 166.250 93.115 166.755 ;
        RECT 93.295 166.545 93.625 166.925 ;
        RECT 93.805 166.375 93.975 166.755 ;
        RECT 88.040 165.275 91.350 165.515 ;
        RECT 88.045 164.375 88.340 165.105 ;
        RECT 88.510 164.550 88.770 165.275 ;
        RECT 88.940 164.375 89.200 165.105 ;
        RECT 89.370 164.550 89.630 165.275 ;
        RECT 89.800 164.375 90.060 165.105 ;
        RECT 90.230 164.550 90.490 165.275 ;
        RECT 90.660 164.375 90.920 165.105 ;
        RECT 91.090 164.550 91.350 165.275 ;
        RECT 91.520 164.375 91.780 165.485 ;
        RECT 91.950 164.550 92.200 165.685 ;
        RECT 92.380 164.375 92.675 165.485 ;
        RECT 92.855 165.450 93.025 166.250 ;
        RECT 93.310 166.205 93.975 166.375 ;
        RECT 93.310 165.950 93.480 166.205 ;
        RECT 94.235 166.175 95.445 166.925 ;
        RECT 95.615 166.415 95.920 166.925 ;
        RECT 93.195 165.620 93.480 165.950 ;
        RECT 93.715 165.655 94.045 166.025 ;
        RECT 93.310 165.475 93.480 165.620 ;
        RECT 92.855 164.545 93.125 165.450 ;
        RECT 93.310 165.305 93.975 165.475 ;
        RECT 93.295 164.375 93.625 165.135 ;
        RECT 93.805 164.545 93.975 165.305 ;
        RECT 94.235 165.465 94.755 166.005 ;
        RECT 94.925 165.635 95.445 166.175 ;
        RECT 95.615 165.685 95.930 166.245 ;
        RECT 96.100 165.935 96.350 166.745 ;
        RECT 96.520 166.400 96.780 166.925 ;
        RECT 96.960 165.935 97.210 166.745 ;
        RECT 97.380 166.365 97.640 166.925 ;
        RECT 97.810 166.275 98.070 166.730 ;
        RECT 98.240 166.445 98.500 166.925 ;
        RECT 98.670 166.275 98.930 166.730 ;
        RECT 99.100 166.445 99.360 166.925 ;
        RECT 99.530 166.275 99.790 166.730 ;
        RECT 99.960 166.445 100.205 166.925 ;
        RECT 100.375 166.275 100.650 166.730 ;
        RECT 100.820 166.445 101.065 166.925 ;
        RECT 101.235 166.275 101.495 166.730 ;
        RECT 101.675 166.445 101.925 166.925 ;
        RECT 102.095 166.275 102.355 166.730 ;
        RECT 102.535 166.445 102.785 166.925 ;
        RECT 102.955 166.275 103.215 166.730 ;
        RECT 103.395 166.445 103.655 166.925 ;
        RECT 103.825 166.275 104.085 166.730 ;
        RECT 104.255 166.445 104.555 166.925 ;
        RECT 97.810 166.105 104.555 166.275 ;
        RECT 104.815 166.155 107.405 166.925 ;
        RECT 96.100 165.685 103.220 165.935 ;
        RECT 94.235 164.375 95.445 165.465 ;
        RECT 95.625 164.375 95.920 165.185 ;
        RECT 96.100 164.545 96.345 165.685 ;
        RECT 96.520 164.375 96.780 165.185 ;
        RECT 96.960 164.550 97.210 165.685 ;
        RECT 103.390 165.515 104.555 166.105 ;
        RECT 97.810 165.290 104.555 165.515 ;
        RECT 104.815 165.465 106.025 165.985 ;
        RECT 106.195 165.635 107.405 166.155 ;
        RECT 107.850 166.115 108.095 166.720 ;
        RECT 108.315 166.390 108.825 166.925 ;
        RECT 107.575 165.945 108.805 166.115 ;
        RECT 97.810 165.275 103.215 165.290 ;
        RECT 97.380 164.380 97.640 165.175 ;
        RECT 97.810 164.550 98.070 165.275 ;
        RECT 98.240 164.380 98.500 165.105 ;
        RECT 98.670 164.550 98.930 165.275 ;
        RECT 99.100 164.380 99.360 165.105 ;
        RECT 99.530 164.550 99.790 165.275 ;
        RECT 99.960 164.380 100.220 165.105 ;
        RECT 100.390 164.550 100.650 165.275 ;
        RECT 100.820 164.380 101.065 165.105 ;
        RECT 101.235 164.550 101.495 165.275 ;
        RECT 101.680 164.380 101.925 165.105 ;
        RECT 102.095 164.550 102.355 165.275 ;
        RECT 102.540 164.380 102.785 165.105 ;
        RECT 102.955 164.550 103.215 165.275 ;
        RECT 103.400 164.380 103.655 165.105 ;
        RECT 103.825 164.550 104.115 165.290 ;
        RECT 97.380 164.375 103.655 164.380 ;
        RECT 104.285 164.375 104.555 165.120 ;
        RECT 104.815 164.375 107.405 165.465 ;
        RECT 107.575 165.135 107.915 165.945 ;
        RECT 108.085 165.380 108.835 165.570 ;
        RECT 107.575 164.725 108.090 165.135 ;
        RECT 108.325 164.375 108.495 165.135 ;
        RECT 108.665 164.715 108.835 165.380 ;
        RECT 109.005 165.395 109.195 166.755 ;
        RECT 109.365 166.585 109.640 166.755 ;
        RECT 109.365 166.415 109.645 166.585 ;
        RECT 109.365 165.595 109.640 166.415 ;
        RECT 109.830 166.390 110.360 166.755 ;
        RECT 110.785 166.525 111.115 166.925 ;
        RECT 110.185 166.355 110.360 166.390 ;
        RECT 109.845 165.395 110.015 166.195 ;
        RECT 109.005 165.225 110.015 165.395 ;
        RECT 110.185 166.185 111.115 166.355 ;
        RECT 111.285 166.185 111.540 166.755 ;
        RECT 112.635 166.200 112.925 166.925 ;
        RECT 110.185 165.055 110.355 166.185 ;
        RECT 110.945 166.015 111.115 166.185 ;
        RECT 109.230 164.885 110.355 165.055 ;
        RECT 110.525 165.685 110.720 166.015 ;
        RECT 110.945 165.685 111.200 166.015 ;
        RECT 110.525 164.715 110.695 165.685 ;
        RECT 111.370 165.515 111.540 166.185 ;
        RECT 113.095 166.155 115.685 166.925 ;
        RECT 108.665 164.545 110.695 164.715 ;
        RECT 110.865 164.375 111.035 165.515 ;
        RECT 111.205 164.545 111.540 165.515 ;
        RECT 112.635 164.375 112.925 165.540 ;
        RECT 113.095 165.465 114.305 165.985 ;
        RECT 114.475 165.635 115.685 166.155 ;
        RECT 115.895 166.105 116.125 166.925 ;
        RECT 116.295 166.125 116.625 166.755 ;
        RECT 115.875 165.685 116.205 165.935 ;
        RECT 116.375 165.525 116.625 166.125 ;
        RECT 116.795 166.105 117.005 166.925 ;
        RECT 117.235 166.175 118.445 166.925 ;
        RECT 118.705 166.375 118.875 166.755 ;
        RECT 119.055 166.545 119.385 166.925 ;
        RECT 118.705 166.205 119.370 166.375 ;
        RECT 119.565 166.250 119.825 166.755 ;
        RECT 113.095 164.375 115.685 165.465 ;
        RECT 115.895 164.375 116.125 165.515 ;
        RECT 116.295 164.545 116.625 165.525 ;
        RECT 116.795 164.375 117.005 165.515 ;
        RECT 117.235 165.465 117.755 166.005 ;
        RECT 117.925 165.635 118.445 166.175 ;
        RECT 118.635 165.655 118.965 166.025 ;
        RECT 119.200 165.950 119.370 166.205 ;
        RECT 119.200 165.620 119.485 165.950 ;
        RECT 119.200 165.475 119.370 165.620 ;
        RECT 117.235 164.375 118.445 165.465 ;
        RECT 118.705 165.305 119.370 165.475 ;
        RECT 119.655 165.450 119.825 166.250 ;
        RECT 120.915 166.155 124.425 166.925 ;
        RECT 124.595 166.175 125.805 166.925 ;
        RECT 118.705 164.545 118.875 165.305 ;
        RECT 119.055 164.375 119.385 165.135 ;
        RECT 119.555 164.545 119.825 165.450 ;
        RECT 120.915 165.465 122.605 165.985 ;
        RECT 122.775 165.635 124.425 166.155 ;
        RECT 124.595 165.465 125.115 166.005 ;
        RECT 125.285 165.635 125.805 166.175 ;
        RECT 120.915 164.375 124.425 165.465 ;
        RECT 124.595 164.375 125.805 165.465 ;
        RECT 11.810 164.205 125.890 164.375 ;
        RECT 11.895 163.115 13.105 164.205 ;
        RECT 11.895 162.405 12.415 162.945 ;
        RECT 12.585 162.575 13.105 163.115 ;
        RECT 13.275 163.115 16.785 164.205 ;
        RECT 16.960 163.770 22.305 164.205 ;
        RECT 13.275 162.595 14.965 163.115 ;
        RECT 15.135 162.425 16.785 162.945 ;
        RECT 18.550 162.520 18.900 163.770 ;
        RECT 22.475 163.040 22.765 164.205 ;
        RECT 23.400 163.770 28.745 164.205 ;
        RECT 11.895 161.655 13.105 162.405 ;
        RECT 13.275 161.655 16.785 162.425 ;
        RECT 20.380 162.200 20.720 163.030 ;
        RECT 24.990 162.520 25.340 163.770 ;
        RECT 29.030 163.575 29.315 164.035 ;
        RECT 29.485 163.745 29.755 164.205 ;
        RECT 29.030 163.355 29.985 163.575 ;
        RECT 16.960 161.655 22.305 162.200 ;
        RECT 22.475 161.655 22.765 162.380 ;
        RECT 26.820 162.200 27.160 163.030 ;
        RECT 28.915 162.625 29.605 163.185 ;
        RECT 29.775 162.455 29.985 163.355 ;
        RECT 29.030 162.285 29.985 162.455 ;
        RECT 30.155 163.185 30.555 164.035 ;
        RECT 30.745 163.575 31.025 164.035 ;
        RECT 31.545 163.745 31.870 164.205 ;
        RECT 30.745 163.355 31.870 163.575 ;
        RECT 30.155 162.625 31.250 163.185 ;
        RECT 31.420 162.895 31.870 163.355 ;
        RECT 32.040 163.065 32.425 164.035 ;
        RECT 23.400 161.655 28.745 162.200 ;
        RECT 29.030 161.825 29.315 162.285 ;
        RECT 29.485 161.655 29.755 162.115 ;
        RECT 30.155 161.825 30.555 162.625 ;
        RECT 31.420 162.565 31.975 162.895 ;
        RECT 31.420 162.455 31.870 162.565 ;
        RECT 30.745 162.285 31.870 162.455 ;
        RECT 32.145 162.395 32.425 163.065 ;
        RECT 32.595 163.115 33.805 164.205 ;
        RECT 33.975 163.130 34.245 164.035 ;
        RECT 34.415 163.445 34.745 164.205 ;
        RECT 34.925 163.275 35.095 164.035 ;
        RECT 32.595 162.575 33.115 163.115 ;
        RECT 33.285 162.405 33.805 162.945 ;
        RECT 30.745 161.825 31.025 162.285 ;
        RECT 31.545 161.655 31.870 162.115 ;
        RECT 32.040 161.825 32.425 162.395 ;
        RECT 32.595 161.655 33.805 162.405 ;
        RECT 33.975 162.330 34.145 163.130 ;
        RECT 34.430 163.105 35.095 163.275 ;
        RECT 35.560 163.235 35.890 164.035 ;
        RECT 36.060 163.405 36.390 164.205 ;
        RECT 36.690 163.235 37.020 164.035 ;
        RECT 37.665 163.405 37.915 164.205 ;
        RECT 34.430 162.960 34.600 163.105 ;
        RECT 35.560 163.065 37.995 163.235 ;
        RECT 38.185 163.065 38.355 164.205 ;
        RECT 38.525 163.065 38.865 164.035 ;
        RECT 39.045 163.395 39.340 164.205 ;
        RECT 34.315 162.630 34.600 162.960 ;
        RECT 34.430 162.375 34.600 162.630 ;
        RECT 34.835 162.555 35.165 162.925 ;
        RECT 35.355 162.645 35.705 162.895 ;
        RECT 35.890 162.435 36.060 163.065 ;
        RECT 36.230 162.645 36.560 162.845 ;
        RECT 36.730 162.645 37.060 162.845 ;
        RECT 37.230 162.645 37.650 162.845 ;
        RECT 37.825 162.815 37.995 163.065 ;
        RECT 37.825 162.645 38.520 162.815 ;
        RECT 33.975 161.825 34.235 162.330 ;
        RECT 34.430 162.205 35.095 162.375 ;
        RECT 34.415 161.655 34.745 162.035 ;
        RECT 34.925 161.825 35.095 162.205 ;
        RECT 35.560 161.825 36.060 162.435 ;
        RECT 36.690 162.305 37.915 162.475 ;
        RECT 38.690 162.455 38.865 163.065 ;
        RECT 39.520 162.895 39.765 164.035 ;
        RECT 39.940 163.395 40.200 164.205 ;
        RECT 40.800 164.200 47.075 164.205 ;
        RECT 40.380 162.895 40.630 164.030 ;
        RECT 40.800 163.405 41.060 164.200 ;
        RECT 41.230 163.305 41.490 164.030 ;
        RECT 41.660 163.475 41.920 164.200 ;
        RECT 42.090 163.305 42.350 164.030 ;
        RECT 42.520 163.475 42.780 164.200 ;
        RECT 42.950 163.305 43.210 164.030 ;
        RECT 43.380 163.475 43.640 164.200 ;
        RECT 43.810 163.305 44.070 164.030 ;
        RECT 44.240 163.475 44.485 164.200 ;
        RECT 44.655 163.305 44.915 164.030 ;
        RECT 45.100 163.475 45.345 164.200 ;
        RECT 45.515 163.305 45.775 164.030 ;
        RECT 45.960 163.475 46.205 164.200 ;
        RECT 46.375 163.305 46.635 164.030 ;
        RECT 46.820 163.475 47.075 164.200 ;
        RECT 41.230 163.290 46.635 163.305 ;
        RECT 47.245 163.290 47.535 164.030 ;
        RECT 47.705 163.460 47.975 164.205 ;
        RECT 41.230 163.065 47.975 163.290 ;
        RECT 36.690 161.825 37.020 162.305 ;
        RECT 37.190 161.655 37.415 162.115 ;
        RECT 37.585 161.825 37.915 162.305 ;
        RECT 38.105 161.655 38.355 162.455 ;
        RECT 38.525 161.825 38.865 162.455 ;
        RECT 39.035 162.335 39.350 162.895 ;
        RECT 39.520 162.645 46.640 162.895 ;
        RECT 39.035 161.655 39.340 162.165 ;
        RECT 39.520 161.835 39.770 162.645 ;
        RECT 39.940 161.655 40.200 162.180 ;
        RECT 40.380 161.835 40.630 162.645 ;
        RECT 46.810 162.505 47.975 163.065 ;
        RECT 48.235 163.040 48.525 164.205 ;
        RECT 49.155 163.115 51.745 164.205 ;
        RECT 51.915 163.445 52.430 163.855 ;
        RECT 52.665 163.445 52.835 164.205 ;
        RECT 53.005 163.865 55.035 164.035 ;
        RECT 49.155 162.595 50.365 163.115 ;
        RECT 46.810 162.475 48.005 162.505 ;
        RECT 41.230 162.335 48.005 162.475 ;
        RECT 50.535 162.425 51.745 162.945 ;
        RECT 51.915 162.635 52.255 163.445 ;
        RECT 53.005 163.200 53.175 163.865 ;
        RECT 53.570 163.525 54.695 163.695 ;
        RECT 52.425 163.010 53.175 163.200 ;
        RECT 53.345 163.185 54.355 163.355 ;
        RECT 51.915 162.465 53.145 162.635 ;
        RECT 41.230 162.305 47.975 162.335 ;
        RECT 40.800 161.655 41.060 162.215 ;
        RECT 41.230 161.850 41.490 162.305 ;
        RECT 41.660 161.655 41.920 162.135 ;
        RECT 42.090 161.850 42.350 162.305 ;
        RECT 42.520 161.655 42.780 162.135 ;
        RECT 42.950 161.850 43.210 162.305 ;
        RECT 43.380 161.655 43.625 162.135 ;
        RECT 43.795 161.850 44.070 162.305 ;
        RECT 44.240 161.655 44.485 162.135 ;
        RECT 44.655 161.850 44.915 162.305 ;
        RECT 45.095 161.655 45.345 162.135 ;
        RECT 45.515 161.850 45.775 162.305 ;
        RECT 45.955 161.655 46.205 162.135 ;
        RECT 46.375 161.850 46.635 162.305 ;
        RECT 46.815 161.655 47.075 162.135 ;
        RECT 47.245 161.850 47.505 162.305 ;
        RECT 47.675 161.655 47.975 162.135 ;
        RECT 48.235 161.655 48.525 162.380 ;
        RECT 49.155 161.655 51.745 162.425 ;
        RECT 52.190 161.860 52.435 162.465 ;
        RECT 52.655 161.655 53.165 162.190 ;
        RECT 53.345 161.825 53.535 163.185 ;
        RECT 53.705 162.165 53.980 162.985 ;
        RECT 54.185 162.385 54.355 163.185 ;
        RECT 54.525 162.395 54.695 163.525 ;
        RECT 54.865 162.895 55.035 163.865 ;
        RECT 55.205 163.065 55.375 164.205 ;
        RECT 55.545 163.065 55.880 164.035 ;
        RECT 54.865 162.565 55.060 162.895 ;
        RECT 55.285 162.565 55.540 162.895 ;
        RECT 55.285 162.395 55.455 162.565 ;
        RECT 55.710 162.395 55.880 163.065 ;
        RECT 56.430 163.225 56.685 163.895 ;
        RECT 56.865 163.405 57.150 164.205 ;
        RECT 57.330 163.485 57.660 163.995 ;
        RECT 56.430 162.505 56.610 163.225 ;
        RECT 57.330 162.895 57.580 163.485 ;
        RECT 57.930 163.335 58.100 163.945 ;
        RECT 58.270 163.515 58.600 164.205 ;
        RECT 58.830 163.655 59.070 163.945 ;
        RECT 59.270 163.825 59.690 164.205 ;
        RECT 59.870 163.735 60.500 163.985 ;
        RECT 60.970 163.825 61.300 164.205 ;
        RECT 59.870 163.655 60.040 163.735 ;
        RECT 61.470 163.655 61.640 163.945 ;
        RECT 61.820 163.825 62.200 164.205 ;
        RECT 62.440 163.820 63.270 163.990 ;
        RECT 58.830 163.485 60.040 163.655 ;
        RECT 56.780 162.565 57.580 162.895 ;
        RECT 54.525 162.225 55.455 162.395 ;
        RECT 54.525 162.190 54.700 162.225 ;
        RECT 53.705 161.995 53.985 162.165 ;
        RECT 53.705 161.825 53.980 161.995 ;
        RECT 54.170 161.825 54.700 162.190 ;
        RECT 55.125 161.655 55.455 162.055 ;
        RECT 55.625 161.825 55.880 162.395 ;
        RECT 56.345 162.365 56.610 162.505 ;
        RECT 56.345 162.335 56.685 162.365 ;
        RECT 56.430 161.835 56.685 162.335 ;
        RECT 56.865 161.655 57.150 162.115 ;
        RECT 57.330 161.915 57.580 162.565 ;
        RECT 57.780 163.315 58.100 163.335 ;
        RECT 57.780 163.145 59.700 163.315 ;
        RECT 57.780 162.250 57.970 163.145 ;
        RECT 59.870 162.975 60.040 163.485 ;
        RECT 60.210 163.225 60.730 163.535 ;
        RECT 58.140 162.805 60.040 162.975 ;
        RECT 58.140 162.745 58.470 162.805 ;
        RECT 58.620 162.575 58.950 162.635 ;
        RECT 58.290 162.305 58.950 162.575 ;
        RECT 57.780 161.920 58.100 162.250 ;
        RECT 58.280 161.655 58.940 162.135 ;
        RECT 59.140 162.045 59.310 162.805 ;
        RECT 60.210 162.635 60.390 163.045 ;
        RECT 59.480 162.465 59.810 162.585 ;
        RECT 60.560 162.465 60.730 163.225 ;
        RECT 59.480 162.295 60.730 162.465 ;
        RECT 60.900 163.405 62.270 163.655 ;
        RECT 60.900 162.635 61.090 163.405 ;
        RECT 62.020 163.145 62.270 163.405 ;
        RECT 61.260 162.975 61.510 163.135 ;
        RECT 62.440 162.975 62.610 163.820 ;
        RECT 63.505 163.535 63.675 164.035 ;
        RECT 63.845 163.705 64.175 164.205 ;
        RECT 62.780 163.145 63.280 163.525 ;
        RECT 63.505 163.365 64.200 163.535 ;
        RECT 61.260 162.805 62.610 162.975 ;
        RECT 62.190 162.765 62.610 162.805 ;
        RECT 60.900 162.295 61.320 162.635 ;
        RECT 61.610 162.305 62.020 162.635 ;
        RECT 59.140 161.875 59.990 162.045 ;
        RECT 60.550 161.655 60.870 162.115 ;
        RECT 61.070 161.865 61.320 162.295 ;
        RECT 61.610 161.655 62.020 162.095 ;
        RECT 62.190 162.035 62.360 162.765 ;
        RECT 62.530 162.215 62.880 162.585 ;
        RECT 63.060 162.275 63.280 163.145 ;
        RECT 63.450 162.575 63.860 163.195 ;
        RECT 64.030 162.395 64.200 163.365 ;
        RECT 63.505 162.205 64.200 162.395 ;
        RECT 62.190 161.835 63.205 162.035 ;
        RECT 63.505 161.875 63.675 162.205 ;
        RECT 63.845 161.655 64.175 162.035 ;
        RECT 64.390 161.915 64.615 164.035 ;
        RECT 64.785 163.705 65.115 164.205 ;
        RECT 65.285 163.535 65.455 164.035 ;
        RECT 64.790 163.365 65.455 163.535 ;
        RECT 64.790 162.375 65.020 163.365 ;
        RECT 65.190 162.545 65.540 163.195 ;
        RECT 66.175 163.115 67.845 164.205 ;
        RECT 68.015 163.130 68.285 164.035 ;
        RECT 68.455 163.445 68.785 164.205 ;
        RECT 68.965 163.275 69.135 164.035 ;
        RECT 66.175 162.595 66.925 163.115 ;
        RECT 67.095 162.425 67.845 162.945 ;
        RECT 64.790 162.205 65.455 162.375 ;
        RECT 64.785 161.655 65.115 162.035 ;
        RECT 65.285 161.915 65.455 162.205 ;
        RECT 66.175 161.655 67.845 162.425 ;
        RECT 68.015 162.330 68.185 163.130 ;
        RECT 68.470 163.105 69.135 163.275 ;
        RECT 69.485 163.275 69.655 164.035 ;
        RECT 69.870 163.445 70.200 164.205 ;
        RECT 69.485 163.105 70.200 163.275 ;
        RECT 70.370 163.130 70.625 164.035 ;
        RECT 68.470 162.960 68.640 163.105 ;
        RECT 68.355 162.630 68.640 162.960 ;
        RECT 68.470 162.375 68.640 162.630 ;
        RECT 68.875 162.555 69.205 162.925 ;
        RECT 69.395 162.555 69.750 162.925 ;
        RECT 70.030 162.895 70.200 163.105 ;
        RECT 70.030 162.565 70.285 162.895 ;
        RECT 70.030 162.375 70.200 162.565 ;
        RECT 70.455 162.400 70.625 163.130 ;
        RECT 70.800 163.055 71.060 164.205 ;
        RECT 71.245 163.145 71.575 164.205 ;
        RECT 71.755 162.895 71.925 163.865 ;
        RECT 72.095 163.615 72.425 164.015 ;
        RECT 72.595 163.845 72.925 164.205 ;
        RECT 73.125 163.615 73.825 164.035 ;
        RECT 72.095 163.385 73.825 163.615 ;
        RECT 72.095 163.165 72.425 163.385 ;
        RECT 72.620 162.895 72.945 163.185 ;
        RECT 71.235 162.565 71.545 162.895 ;
        RECT 71.755 162.565 72.130 162.895 ;
        RECT 72.450 162.565 72.945 162.895 ;
        RECT 73.120 162.645 73.450 163.185 ;
        RECT 68.015 161.825 68.275 162.330 ;
        RECT 68.470 162.205 69.135 162.375 ;
        RECT 68.455 161.655 68.785 162.035 ;
        RECT 68.965 161.825 69.135 162.205 ;
        RECT 69.485 162.205 70.200 162.375 ;
        RECT 69.485 161.825 69.655 162.205 ;
        RECT 69.870 161.655 70.200 162.035 ;
        RECT 70.370 161.825 70.625 162.400 ;
        RECT 70.800 161.655 71.060 162.495 ;
        RECT 73.620 162.415 73.825 163.385 ;
        RECT 73.995 163.040 74.285 164.205 ;
        RECT 74.915 163.115 76.585 164.205 ;
        RECT 76.755 163.445 77.270 163.855 ;
        RECT 77.505 163.445 77.675 164.205 ;
        RECT 77.845 163.865 79.875 164.035 ;
        RECT 74.915 162.595 75.665 163.115 ;
        RECT 75.835 162.425 76.585 162.945 ;
        RECT 76.755 162.635 77.095 163.445 ;
        RECT 77.845 163.200 78.015 163.865 ;
        RECT 78.410 163.525 79.535 163.695 ;
        RECT 77.265 163.010 78.015 163.200 ;
        RECT 78.185 163.185 79.195 163.355 ;
        RECT 76.755 162.465 77.985 162.635 ;
        RECT 71.245 162.185 72.605 162.395 ;
        RECT 71.245 161.825 71.575 162.185 ;
        RECT 71.745 161.655 72.075 162.015 ;
        RECT 72.275 161.825 72.605 162.185 ;
        RECT 73.115 161.825 73.825 162.415 ;
        RECT 73.995 161.655 74.285 162.380 ;
        RECT 74.915 161.655 76.585 162.425 ;
        RECT 77.030 161.860 77.275 162.465 ;
        RECT 77.495 161.655 78.005 162.190 ;
        RECT 78.185 161.825 78.375 163.185 ;
        RECT 78.545 162.165 78.820 162.985 ;
        RECT 79.025 162.385 79.195 163.185 ;
        RECT 79.365 162.395 79.535 163.525 ;
        RECT 79.705 162.895 79.875 163.865 ;
        RECT 80.045 163.065 80.215 164.205 ;
        RECT 80.385 163.065 80.720 164.035 ;
        RECT 79.705 162.565 79.900 162.895 ;
        RECT 80.125 162.565 80.380 162.895 ;
        RECT 80.125 162.395 80.295 162.565 ;
        RECT 80.550 162.395 80.720 163.065 ;
        RECT 79.365 162.225 80.295 162.395 ;
        RECT 79.365 162.190 79.540 162.225 ;
        RECT 78.545 161.995 78.825 162.165 ;
        RECT 78.545 161.825 78.820 161.995 ;
        RECT 79.010 161.825 79.540 162.190 ;
        RECT 79.965 161.655 80.295 162.055 ;
        RECT 80.465 161.825 80.720 162.395 ;
        RECT 81.270 163.225 81.525 163.895 ;
        RECT 81.705 163.405 81.990 164.205 ;
        RECT 82.170 163.485 82.500 163.995 ;
        RECT 81.270 162.365 81.450 163.225 ;
        RECT 82.170 162.895 82.420 163.485 ;
        RECT 82.770 163.335 82.940 163.945 ;
        RECT 83.110 163.515 83.440 164.205 ;
        RECT 83.670 163.655 83.910 163.945 ;
        RECT 84.110 163.825 84.530 164.205 ;
        RECT 84.710 163.735 85.340 163.985 ;
        RECT 85.810 163.825 86.140 164.205 ;
        RECT 84.710 163.655 84.880 163.735 ;
        RECT 86.310 163.655 86.480 163.945 ;
        RECT 86.660 163.825 87.040 164.205 ;
        RECT 87.280 163.820 88.110 163.990 ;
        RECT 83.670 163.485 84.880 163.655 ;
        RECT 81.620 162.565 82.420 162.895 ;
        RECT 81.270 162.165 81.525 162.365 ;
        RECT 81.185 161.995 81.525 162.165 ;
        RECT 81.270 161.835 81.525 161.995 ;
        RECT 81.705 161.655 81.990 162.115 ;
        RECT 82.170 161.915 82.420 162.565 ;
        RECT 82.620 163.315 82.940 163.335 ;
        RECT 82.620 163.145 84.540 163.315 ;
        RECT 82.620 162.250 82.810 163.145 ;
        RECT 84.710 162.975 84.880 163.485 ;
        RECT 85.050 163.225 85.570 163.535 ;
        RECT 82.980 162.805 84.880 162.975 ;
        RECT 82.980 162.745 83.310 162.805 ;
        RECT 83.460 162.575 83.790 162.635 ;
        RECT 83.130 162.305 83.790 162.575 ;
        RECT 82.620 161.920 82.940 162.250 ;
        RECT 83.120 161.655 83.780 162.135 ;
        RECT 83.980 162.045 84.150 162.805 ;
        RECT 85.050 162.635 85.230 163.045 ;
        RECT 84.320 162.465 84.650 162.585 ;
        RECT 85.400 162.465 85.570 163.225 ;
        RECT 84.320 162.295 85.570 162.465 ;
        RECT 85.740 163.405 87.110 163.655 ;
        RECT 85.740 162.635 85.930 163.405 ;
        RECT 86.860 163.145 87.110 163.405 ;
        RECT 86.100 162.975 86.350 163.135 ;
        RECT 87.280 162.975 87.450 163.820 ;
        RECT 88.345 163.535 88.515 164.035 ;
        RECT 88.685 163.705 89.015 164.205 ;
        RECT 87.620 163.145 88.120 163.525 ;
        RECT 88.345 163.365 89.040 163.535 ;
        RECT 86.100 162.805 87.450 162.975 ;
        RECT 87.030 162.765 87.450 162.805 ;
        RECT 85.740 162.295 86.160 162.635 ;
        RECT 86.450 162.305 86.860 162.635 ;
        RECT 83.980 161.875 84.830 162.045 ;
        RECT 85.390 161.655 85.710 162.115 ;
        RECT 85.910 161.865 86.160 162.295 ;
        RECT 86.450 161.655 86.860 162.095 ;
        RECT 87.030 162.035 87.200 162.765 ;
        RECT 87.370 162.215 87.720 162.585 ;
        RECT 87.900 162.275 88.120 163.145 ;
        RECT 88.290 162.575 88.700 163.195 ;
        RECT 88.870 162.395 89.040 163.365 ;
        RECT 88.345 162.205 89.040 162.395 ;
        RECT 87.030 161.835 88.045 162.035 ;
        RECT 88.345 161.875 88.515 162.205 ;
        RECT 88.685 161.655 89.015 162.035 ;
        RECT 89.230 161.915 89.455 164.035 ;
        RECT 89.625 163.705 89.955 164.205 ;
        RECT 90.125 163.535 90.295 164.035 ;
        RECT 89.630 163.365 90.295 163.535 ;
        RECT 89.630 162.375 89.860 163.365 ;
        RECT 90.030 162.545 90.380 163.195 ;
        RECT 90.560 163.015 90.815 163.895 ;
        RECT 90.985 163.065 91.290 164.205 ;
        RECT 91.630 163.825 91.960 164.205 ;
        RECT 92.140 163.655 92.310 163.945 ;
        RECT 92.480 163.745 92.730 164.205 ;
        RECT 91.510 163.485 92.310 163.655 ;
        RECT 92.900 163.695 93.770 164.035 ;
        RECT 89.630 162.205 90.295 162.375 ;
        RECT 89.625 161.655 89.955 162.035 ;
        RECT 90.125 161.915 90.295 162.205 ;
        RECT 90.560 162.365 90.770 163.015 ;
        RECT 91.510 162.895 91.680 163.485 ;
        RECT 92.900 163.315 93.070 163.695 ;
        RECT 94.005 163.575 94.175 164.035 ;
        RECT 94.345 163.745 94.715 164.205 ;
        RECT 95.010 163.605 95.180 163.945 ;
        RECT 95.350 163.775 95.680 164.205 ;
        RECT 95.915 163.605 96.085 163.945 ;
        RECT 91.850 163.145 93.070 163.315 ;
        RECT 93.240 163.235 93.700 163.525 ;
        RECT 94.005 163.405 94.565 163.575 ;
        RECT 95.010 163.435 96.085 163.605 ;
        RECT 96.255 163.705 96.935 164.035 ;
        RECT 97.150 163.705 97.400 164.035 ;
        RECT 97.570 163.745 97.820 164.205 ;
        RECT 94.395 163.265 94.565 163.405 ;
        RECT 93.240 163.225 94.205 163.235 ;
        RECT 92.900 163.055 93.070 163.145 ;
        RECT 93.530 163.065 94.205 163.225 ;
        RECT 90.940 162.865 91.680 162.895 ;
        RECT 90.940 162.565 91.855 162.865 ;
        RECT 91.530 162.390 91.855 162.565 ;
        RECT 90.560 161.835 90.815 162.365 ;
        RECT 90.985 161.655 91.290 162.115 ;
        RECT 91.535 162.035 91.855 162.390 ;
        RECT 92.025 162.605 92.565 162.975 ;
        RECT 92.900 162.885 93.305 163.055 ;
        RECT 92.025 162.205 92.265 162.605 ;
        RECT 92.745 162.435 92.965 162.715 ;
        RECT 92.435 162.265 92.965 162.435 ;
        RECT 92.435 162.035 92.605 162.265 ;
        RECT 93.135 162.105 93.305 162.885 ;
        RECT 93.475 162.275 93.825 162.895 ;
        RECT 93.995 162.275 94.205 163.065 ;
        RECT 94.395 163.095 95.895 163.265 ;
        RECT 94.395 162.405 94.565 163.095 ;
        RECT 96.255 162.925 96.425 163.705 ;
        RECT 97.230 163.575 97.400 163.705 ;
        RECT 94.735 162.755 96.425 162.925 ;
        RECT 96.595 163.145 97.060 163.535 ;
        RECT 97.230 163.405 97.625 163.575 ;
        RECT 94.735 162.575 94.905 162.755 ;
        RECT 91.535 161.865 92.605 162.035 ;
        RECT 92.775 161.655 92.965 162.095 ;
        RECT 93.135 161.825 94.085 162.105 ;
        RECT 94.395 162.015 94.655 162.405 ;
        RECT 95.075 162.335 95.865 162.585 ;
        RECT 94.305 161.845 94.655 162.015 ;
        RECT 94.865 161.655 95.195 162.115 ;
        RECT 96.070 162.045 96.240 162.755 ;
        RECT 96.595 162.555 96.765 163.145 ;
        RECT 96.410 162.335 96.765 162.555 ;
        RECT 96.935 162.335 97.285 162.955 ;
        RECT 97.455 162.045 97.625 163.405 ;
        RECT 97.990 163.235 98.315 164.020 ;
        RECT 97.795 162.185 98.255 163.235 ;
        RECT 96.070 161.875 96.925 162.045 ;
        RECT 97.130 161.875 97.625 162.045 ;
        RECT 97.795 161.655 98.125 162.015 ;
        RECT 98.485 161.915 98.655 164.035 ;
        RECT 98.825 163.705 99.155 164.205 ;
        RECT 99.325 163.535 99.580 164.035 ;
        RECT 98.830 163.365 99.580 163.535 ;
        RECT 98.830 162.375 99.060 163.365 ;
        RECT 99.230 162.545 99.580 163.195 ;
        RECT 99.755 163.040 100.045 164.205 ;
        RECT 100.215 163.065 100.555 164.035 ;
        RECT 100.725 163.065 100.895 164.205 ;
        RECT 101.165 163.405 101.415 164.205 ;
        RECT 102.060 163.235 102.390 164.035 ;
        RECT 102.690 163.405 103.020 164.205 ;
        RECT 103.190 163.235 103.520 164.035 ;
        RECT 101.085 163.065 103.520 163.235 ;
        RECT 103.895 163.065 104.235 164.035 ;
        RECT 104.405 163.065 104.575 164.205 ;
        RECT 104.845 163.405 105.095 164.205 ;
        RECT 105.740 163.235 106.070 164.035 ;
        RECT 106.370 163.405 106.700 164.205 ;
        RECT 106.870 163.235 107.200 164.035 ;
        RECT 108.040 163.770 113.385 164.205 ;
        RECT 104.765 163.065 107.200 163.235 ;
        RECT 100.215 162.455 100.390 163.065 ;
        RECT 101.085 162.815 101.255 163.065 ;
        RECT 100.560 162.645 101.255 162.815 ;
        RECT 101.430 162.645 101.850 162.845 ;
        RECT 102.020 162.645 102.350 162.845 ;
        RECT 102.520 162.645 102.850 162.845 ;
        RECT 98.830 162.205 99.580 162.375 ;
        RECT 98.825 161.655 99.155 162.035 ;
        RECT 99.325 161.915 99.580 162.205 ;
        RECT 99.755 161.655 100.045 162.380 ;
        RECT 100.215 161.825 100.555 162.455 ;
        RECT 100.725 161.655 100.975 162.455 ;
        RECT 101.165 162.305 102.390 162.475 ;
        RECT 101.165 161.825 101.495 162.305 ;
        RECT 101.665 161.655 101.890 162.115 ;
        RECT 102.060 161.825 102.390 162.305 ;
        RECT 103.020 162.435 103.190 163.065 ;
        RECT 103.375 162.645 103.725 162.895 ;
        RECT 103.895 162.455 104.070 163.065 ;
        RECT 104.765 162.815 104.935 163.065 ;
        RECT 104.240 162.645 104.935 162.815 ;
        RECT 105.110 162.645 105.530 162.845 ;
        RECT 105.700 162.645 106.030 162.845 ;
        RECT 106.200 162.645 106.530 162.845 ;
        RECT 103.020 161.825 103.520 162.435 ;
        RECT 103.895 161.825 104.235 162.455 ;
        RECT 104.405 161.655 104.655 162.455 ;
        RECT 104.845 162.305 106.070 162.475 ;
        RECT 104.845 161.825 105.175 162.305 ;
        RECT 105.345 161.655 105.570 162.115 ;
        RECT 105.740 161.825 106.070 162.305 ;
        RECT 106.700 162.435 106.870 163.065 ;
        RECT 107.055 162.645 107.405 162.895 ;
        RECT 109.630 162.520 109.980 163.770 ;
        RECT 106.700 161.825 107.200 162.435 ;
        RECT 111.460 162.200 111.800 163.030 ;
        RECT 113.560 163.015 113.815 163.895 ;
        RECT 113.985 163.065 114.290 164.205 ;
        RECT 114.630 163.825 114.960 164.205 ;
        RECT 115.140 163.655 115.310 163.945 ;
        RECT 115.480 163.745 115.730 164.205 ;
        RECT 114.510 163.485 115.310 163.655 ;
        RECT 115.900 163.695 116.770 164.035 ;
        RECT 113.560 162.365 113.770 163.015 ;
        RECT 114.510 162.895 114.680 163.485 ;
        RECT 115.900 163.315 116.070 163.695 ;
        RECT 117.005 163.575 117.175 164.035 ;
        RECT 117.345 163.745 117.715 164.205 ;
        RECT 118.010 163.605 118.180 163.945 ;
        RECT 118.350 163.775 118.680 164.205 ;
        RECT 118.915 163.605 119.085 163.945 ;
        RECT 114.850 163.145 116.070 163.315 ;
        RECT 116.240 163.235 116.700 163.525 ;
        RECT 117.005 163.405 117.565 163.575 ;
        RECT 118.010 163.435 119.085 163.605 ;
        RECT 119.255 163.705 119.935 164.035 ;
        RECT 120.150 163.705 120.400 164.035 ;
        RECT 120.570 163.745 120.820 164.205 ;
        RECT 117.395 163.265 117.565 163.405 ;
        RECT 116.240 163.225 117.205 163.235 ;
        RECT 115.900 163.055 116.070 163.145 ;
        RECT 116.530 163.065 117.205 163.225 ;
        RECT 113.940 162.865 114.680 162.895 ;
        RECT 113.940 162.565 114.855 162.865 ;
        RECT 114.530 162.390 114.855 162.565 ;
        RECT 108.040 161.655 113.385 162.200 ;
        RECT 113.560 161.835 113.815 162.365 ;
        RECT 113.985 161.655 114.290 162.115 ;
        RECT 114.535 162.035 114.855 162.390 ;
        RECT 115.025 162.605 115.565 162.975 ;
        RECT 115.900 162.885 116.305 163.055 ;
        RECT 115.025 162.205 115.265 162.605 ;
        RECT 115.745 162.435 115.965 162.715 ;
        RECT 115.435 162.265 115.965 162.435 ;
        RECT 115.435 162.035 115.605 162.265 ;
        RECT 116.135 162.105 116.305 162.885 ;
        RECT 116.475 162.275 116.825 162.895 ;
        RECT 116.995 162.275 117.205 163.065 ;
        RECT 117.395 163.095 118.895 163.265 ;
        RECT 117.395 162.405 117.565 163.095 ;
        RECT 119.255 162.925 119.425 163.705 ;
        RECT 120.230 163.575 120.400 163.705 ;
        RECT 117.735 162.755 119.425 162.925 ;
        RECT 119.595 163.145 120.060 163.535 ;
        RECT 120.230 163.405 120.625 163.575 ;
        RECT 117.735 162.575 117.905 162.755 ;
        RECT 114.535 161.865 115.605 162.035 ;
        RECT 115.775 161.655 115.965 162.095 ;
        RECT 116.135 161.825 117.085 162.105 ;
        RECT 117.395 162.015 117.655 162.405 ;
        RECT 118.075 162.335 118.865 162.585 ;
        RECT 117.305 161.845 117.655 162.015 ;
        RECT 117.865 161.655 118.195 162.115 ;
        RECT 119.070 162.045 119.240 162.755 ;
        RECT 119.595 162.555 119.765 163.145 ;
        RECT 119.410 162.335 119.765 162.555 ;
        RECT 119.935 162.335 120.285 162.955 ;
        RECT 120.455 162.045 120.625 163.405 ;
        RECT 120.990 163.235 121.315 164.020 ;
        RECT 120.795 162.185 121.255 163.235 ;
        RECT 119.070 161.875 119.925 162.045 ;
        RECT 120.130 161.875 120.625 162.045 ;
        RECT 120.795 161.655 121.125 162.015 ;
        RECT 121.485 161.915 121.655 164.035 ;
        RECT 121.825 163.705 122.155 164.205 ;
        RECT 122.325 163.535 122.580 164.035 ;
        RECT 121.830 163.365 122.580 163.535 ;
        RECT 121.830 162.375 122.060 163.365 ;
        RECT 122.230 162.545 122.580 163.195 ;
        RECT 122.755 163.115 124.425 164.205 ;
        RECT 124.595 163.115 125.805 164.205 ;
        RECT 122.755 162.595 123.505 163.115 ;
        RECT 123.675 162.425 124.425 162.945 ;
        RECT 124.595 162.575 125.115 163.115 ;
        RECT 121.830 162.205 122.580 162.375 ;
        RECT 121.825 161.655 122.155 162.035 ;
        RECT 122.325 161.915 122.580 162.205 ;
        RECT 122.755 161.655 124.425 162.425 ;
        RECT 125.285 162.405 125.805 162.945 ;
        RECT 124.595 161.655 125.805 162.405 ;
        RECT 11.810 161.485 125.890 161.655 ;
        RECT 11.895 160.735 13.105 161.485 ;
        RECT 14.200 160.940 19.545 161.485 ;
        RECT 11.895 160.195 12.415 160.735 ;
        RECT 12.585 160.025 13.105 160.565 ;
        RECT 11.895 158.935 13.105 160.025 ;
        RECT 15.790 159.370 16.140 160.620 ;
        RECT 17.620 160.110 17.960 160.940 ;
        RECT 19.990 160.675 20.235 161.280 ;
        RECT 20.455 160.950 20.965 161.485 ;
        RECT 19.715 160.505 20.945 160.675 ;
        RECT 19.715 159.695 20.055 160.505 ;
        RECT 20.225 159.940 20.975 160.130 ;
        RECT 14.200 158.935 19.545 159.370 ;
        RECT 19.715 159.285 20.230 159.695 ;
        RECT 20.465 158.935 20.635 159.695 ;
        RECT 20.805 159.275 20.975 159.940 ;
        RECT 21.145 159.955 21.335 161.315 ;
        RECT 21.505 161.145 21.780 161.315 ;
        RECT 21.505 160.975 21.785 161.145 ;
        RECT 21.505 160.155 21.780 160.975 ;
        RECT 21.970 160.950 22.500 161.315 ;
        RECT 22.925 161.085 23.255 161.485 ;
        RECT 22.325 160.915 22.500 160.950 ;
        RECT 21.985 159.955 22.155 160.755 ;
        RECT 21.145 159.785 22.155 159.955 ;
        RECT 22.325 160.745 23.255 160.915 ;
        RECT 23.425 160.745 23.680 161.315 ;
        RECT 23.860 160.940 29.205 161.485 ;
        RECT 22.325 159.615 22.495 160.745 ;
        RECT 23.085 160.575 23.255 160.745 ;
        RECT 21.370 159.445 22.495 159.615 ;
        RECT 22.665 160.245 22.860 160.575 ;
        RECT 23.085 160.245 23.340 160.575 ;
        RECT 22.665 159.275 22.835 160.245 ;
        RECT 23.510 160.075 23.680 160.745 ;
        RECT 20.805 159.105 22.835 159.275 ;
        RECT 23.005 158.935 23.175 160.075 ;
        RECT 23.345 159.105 23.680 160.075 ;
        RECT 25.450 159.370 25.800 160.620 ;
        RECT 27.280 160.110 27.620 160.940 ;
        RECT 29.650 160.675 29.895 161.280 ;
        RECT 30.115 160.950 30.625 161.485 ;
        RECT 29.375 160.505 30.605 160.675 ;
        RECT 29.375 159.695 29.715 160.505 ;
        RECT 29.885 159.940 30.635 160.130 ;
        RECT 23.860 158.935 29.205 159.370 ;
        RECT 29.375 159.285 29.890 159.695 ;
        RECT 30.125 158.935 30.295 159.695 ;
        RECT 30.465 159.275 30.635 159.940 ;
        RECT 30.805 159.955 30.995 161.315 ;
        RECT 31.165 160.465 31.440 161.315 ;
        RECT 31.630 160.950 32.160 161.315 ;
        RECT 32.585 161.085 32.915 161.485 ;
        RECT 31.985 160.915 32.160 160.950 ;
        RECT 31.165 160.295 31.445 160.465 ;
        RECT 31.165 160.155 31.440 160.295 ;
        RECT 31.645 159.955 31.815 160.755 ;
        RECT 30.805 159.785 31.815 159.955 ;
        RECT 31.985 160.745 32.915 160.915 ;
        RECT 33.085 160.745 33.340 161.315 ;
        RECT 31.985 159.615 32.155 160.745 ;
        RECT 32.745 160.575 32.915 160.745 ;
        RECT 31.030 159.445 32.155 159.615 ;
        RECT 32.325 160.245 32.520 160.575 ;
        RECT 32.745 160.245 33.000 160.575 ;
        RECT 32.325 159.275 32.495 160.245 ;
        RECT 33.170 160.075 33.340 160.745 ;
        RECT 33.515 160.715 35.185 161.485 ;
        RECT 35.355 160.760 35.645 161.485 ;
        RECT 30.465 159.105 32.495 159.275 ;
        RECT 32.665 158.935 32.835 160.075 ;
        RECT 33.005 159.105 33.340 160.075 ;
        RECT 33.515 160.025 34.265 160.545 ;
        RECT 34.435 160.195 35.185 160.715 ;
        RECT 36.940 160.705 37.440 161.315 ;
        RECT 36.735 160.245 37.085 160.495 ;
        RECT 33.515 158.935 35.185 160.025 ;
        RECT 35.355 158.935 35.645 160.100 ;
        RECT 37.270 160.075 37.440 160.705 ;
        RECT 38.070 160.835 38.400 161.315 ;
        RECT 38.570 161.025 38.795 161.485 ;
        RECT 38.965 160.835 39.295 161.315 ;
        RECT 38.070 160.665 39.295 160.835 ;
        RECT 39.485 160.685 39.735 161.485 ;
        RECT 39.905 160.685 40.245 161.315 ;
        RECT 40.525 161.005 40.695 161.485 ;
        RECT 40.865 160.835 41.195 161.310 ;
        RECT 41.365 161.005 41.535 161.485 ;
        RECT 41.705 160.835 42.035 161.310 ;
        RECT 42.205 161.005 42.375 161.485 ;
        RECT 42.545 160.835 42.875 161.310 ;
        RECT 43.045 161.005 43.215 161.485 ;
        RECT 43.385 160.835 43.715 161.310 ;
        RECT 43.885 161.005 44.055 161.485 ;
        RECT 44.225 160.835 44.555 161.310 ;
        RECT 44.725 161.005 44.895 161.485 ;
        RECT 45.145 161.310 45.315 161.315 ;
        RECT 45.065 160.835 45.395 161.310 ;
        RECT 45.565 161.005 45.735 161.485 ;
        RECT 45.985 161.310 46.155 161.315 ;
        RECT 45.905 160.835 46.235 161.310 ;
        RECT 46.405 161.005 46.575 161.485 ;
        RECT 46.825 161.310 47.075 161.315 ;
        RECT 46.745 160.835 47.075 161.310 ;
        RECT 47.245 161.005 47.415 161.485 ;
        RECT 47.585 160.835 47.915 161.310 ;
        RECT 48.085 161.005 48.255 161.485 ;
        RECT 48.425 160.835 48.755 161.310 ;
        RECT 48.925 161.005 49.095 161.485 ;
        RECT 49.265 160.835 49.595 161.310 ;
        RECT 49.765 161.005 49.935 161.485 ;
        RECT 50.105 160.835 50.435 161.310 ;
        RECT 50.605 161.005 50.775 161.485 ;
        RECT 50.945 160.835 51.275 161.310 ;
        RECT 37.610 160.295 37.940 160.495 ;
        RECT 38.110 160.295 38.440 160.495 ;
        RECT 38.610 160.295 39.030 160.495 ;
        RECT 39.205 160.325 39.900 160.495 ;
        RECT 39.205 160.075 39.375 160.325 ;
        RECT 40.070 160.075 40.245 160.685 ;
        RECT 36.940 159.905 39.375 160.075 ;
        RECT 36.940 159.105 37.270 159.905 ;
        RECT 37.440 158.935 37.770 159.735 ;
        RECT 38.070 159.105 38.400 159.905 ;
        RECT 39.045 158.935 39.295 159.735 ;
        RECT 39.565 158.935 39.735 160.075 ;
        RECT 39.905 159.105 40.245 160.075 ;
        RECT 40.415 160.665 47.075 160.835 ;
        RECT 47.245 160.665 49.595 160.835 ;
        RECT 49.765 160.665 51.275 160.835 ;
        RECT 51.455 160.685 51.795 161.315 ;
        RECT 51.965 160.685 52.215 161.485 ;
        RECT 52.405 160.835 52.735 161.315 ;
        RECT 52.905 161.025 53.130 161.485 ;
        RECT 53.300 160.835 53.630 161.315 ;
        RECT 40.415 160.125 40.690 160.665 ;
        RECT 47.245 160.495 47.420 160.665 ;
        RECT 49.765 160.495 49.935 160.665 ;
        RECT 40.860 160.295 47.420 160.495 ;
        RECT 47.625 160.295 49.935 160.495 ;
        RECT 50.105 160.295 51.280 160.495 ;
        RECT 47.245 160.125 47.420 160.295 ;
        RECT 49.765 160.125 49.935 160.295 ;
        RECT 40.415 159.955 47.075 160.125 ;
        RECT 47.245 159.955 49.595 160.125 ;
        RECT 49.765 159.955 51.275 160.125 ;
        RECT 40.525 158.935 40.695 159.735 ;
        RECT 40.865 159.105 41.195 159.955 ;
        RECT 41.365 158.935 41.535 159.735 ;
        RECT 41.705 159.105 42.035 159.955 ;
        RECT 42.205 158.935 42.375 159.735 ;
        RECT 42.545 159.105 42.875 159.955 ;
        RECT 43.045 158.935 43.215 159.735 ;
        RECT 43.385 159.105 43.715 159.955 ;
        RECT 43.885 158.935 44.055 159.735 ;
        RECT 44.225 159.105 44.555 159.955 ;
        RECT 44.725 158.935 44.895 159.735 ;
        RECT 45.065 159.105 45.395 159.955 ;
        RECT 45.565 158.935 45.735 159.735 ;
        RECT 45.905 159.105 46.235 159.955 ;
        RECT 46.405 158.935 46.575 159.735 ;
        RECT 46.745 159.105 47.075 159.955 ;
        RECT 47.245 158.935 47.415 159.735 ;
        RECT 47.585 159.105 47.915 159.955 ;
        RECT 48.085 158.935 48.255 159.735 ;
        RECT 48.425 159.105 48.755 159.955 ;
        RECT 48.925 158.935 49.095 159.735 ;
        RECT 49.265 159.105 49.595 159.955 ;
        RECT 49.765 158.935 49.935 159.785 ;
        RECT 50.105 159.105 50.435 159.955 ;
        RECT 50.605 158.935 50.775 159.785 ;
        RECT 50.945 159.105 51.275 159.955 ;
        RECT 51.455 160.075 51.630 160.685 ;
        RECT 52.405 160.665 53.630 160.835 ;
        RECT 54.260 160.705 54.760 161.315 ;
        RECT 55.135 160.735 56.345 161.485 ;
        RECT 51.800 160.325 52.495 160.495 ;
        RECT 52.325 160.075 52.495 160.325 ;
        RECT 52.670 160.295 53.090 160.495 ;
        RECT 53.260 160.295 53.590 160.495 ;
        RECT 53.760 160.295 54.090 160.495 ;
        RECT 54.260 160.075 54.430 160.705 ;
        RECT 54.615 160.245 54.965 160.495 ;
        RECT 51.455 159.105 51.795 160.075 ;
        RECT 51.965 158.935 52.135 160.075 ;
        RECT 52.325 159.905 54.760 160.075 ;
        RECT 52.405 158.935 52.655 159.735 ;
        RECT 53.300 159.105 53.630 159.905 ;
        RECT 53.930 158.935 54.260 159.735 ;
        RECT 54.430 159.105 54.760 159.905 ;
        RECT 55.135 160.025 55.655 160.565 ;
        RECT 55.825 160.195 56.345 160.735 ;
        RECT 56.790 160.675 57.035 161.280 ;
        RECT 57.255 160.950 57.765 161.485 ;
        RECT 56.515 160.505 57.745 160.675 ;
        RECT 55.135 158.935 56.345 160.025 ;
        RECT 56.515 159.695 56.855 160.505 ;
        RECT 57.025 159.940 57.775 160.130 ;
        RECT 56.515 159.285 57.030 159.695 ;
        RECT 57.265 158.935 57.435 159.695 ;
        RECT 57.605 159.275 57.775 159.940 ;
        RECT 57.945 159.955 58.135 161.315 ;
        RECT 58.305 161.145 58.580 161.315 ;
        RECT 58.305 160.975 58.585 161.145 ;
        RECT 58.305 160.155 58.580 160.975 ;
        RECT 58.770 160.950 59.300 161.315 ;
        RECT 59.725 161.085 60.055 161.485 ;
        RECT 59.125 160.915 59.300 160.950 ;
        RECT 58.785 159.955 58.955 160.755 ;
        RECT 57.945 159.785 58.955 159.955 ;
        RECT 59.125 160.745 60.055 160.915 ;
        RECT 60.225 160.745 60.480 161.315 ;
        RECT 61.115 160.760 61.405 161.485 ;
        RECT 61.665 160.935 61.835 161.315 ;
        RECT 62.015 161.105 62.345 161.485 ;
        RECT 61.665 160.765 62.330 160.935 ;
        RECT 62.525 160.810 62.785 161.315 ;
        RECT 59.125 159.615 59.295 160.745 ;
        RECT 59.885 160.575 60.055 160.745 ;
        RECT 58.170 159.445 59.295 159.615 ;
        RECT 59.465 160.245 59.660 160.575 ;
        RECT 59.885 160.245 60.140 160.575 ;
        RECT 59.465 159.275 59.635 160.245 ;
        RECT 60.310 160.075 60.480 160.745 ;
        RECT 61.595 160.215 61.925 160.585 ;
        RECT 62.160 160.510 62.330 160.765 ;
        RECT 62.160 160.180 62.445 160.510 ;
        RECT 57.605 159.105 59.635 159.275 ;
        RECT 59.805 158.935 59.975 160.075 ;
        RECT 60.145 159.105 60.480 160.075 ;
        RECT 61.115 158.935 61.405 160.100 ;
        RECT 62.160 160.035 62.330 160.180 ;
        RECT 61.665 159.865 62.330 160.035 ;
        RECT 62.615 160.010 62.785 160.810 ;
        RECT 62.955 160.715 64.625 161.485 ;
        RECT 61.665 159.105 61.835 159.865 ;
        RECT 62.015 158.935 62.345 159.695 ;
        RECT 62.515 159.105 62.785 160.010 ;
        RECT 62.955 160.025 63.705 160.545 ;
        RECT 63.875 160.195 64.625 160.715 ;
        RECT 64.800 160.645 65.060 161.485 ;
        RECT 65.235 160.740 65.490 161.315 ;
        RECT 65.660 161.105 65.990 161.485 ;
        RECT 66.205 160.935 66.375 161.315 ;
        RECT 65.660 160.765 66.375 160.935 ;
        RECT 62.955 158.935 64.625 160.025 ;
        RECT 64.800 158.935 65.060 160.085 ;
        RECT 65.235 160.010 65.405 160.740 ;
        RECT 65.660 160.575 65.830 160.765 ;
        RECT 66.640 160.645 66.900 161.485 ;
        RECT 67.075 160.740 67.330 161.315 ;
        RECT 67.500 161.105 67.830 161.485 ;
        RECT 68.045 160.935 68.215 161.315 ;
        RECT 67.500 160.765 68.215 160.935 ;
        RECT 65.575 160.245 65.830 160.575 ;
        RECT 65.660 160.035 65.830 160.245 ;
        RECT 66.110 160.215 66.465 160.585 ;
        RECT 65.235 159.105 65.490 160.010 ;
        RECT 65.660 159.865 66.375 160.035 ;
        RECT 65.660 158.935 65.990 159.695 ;
        RECT 66.205 159.105 66.375 159.865 ;
        RECT 66.640 158.935 66.900 160.085 ;
        RECT 67.075 160.010 67.245 160.740 ;
        RECT 67.500 160.575 67.670 160.765 ;
        RECT 68.480 160.645 68.740 161.485 ;
        RECT 68.915 160.740 69.170 161.315 ;
        RECT 69.340 161.105 69.670 161.485 ;
        RECT 69.885 160.935 70.055 161.315 ;
        RECT 69.340 160.765 70.055 160.935 ;
        RECT 67.415 160.245 67.670 160.575 ;
        RECT 67.500 160.035 67.670 160.245 ;
        RECT 67.950 160.215 68.305 160.585 ;
        RECT 67.075 159.105 67.330 160.010 ;
        RECT 67.500 159.865 68.215 160.035 ;
        RECT 67.500 158.935 67.830 159.695 ;
        RECT 68.045 159.105 68.215 159.865 ;
        RECT 68.480 158.935 68.740 160.085 ;
        RECT 68.915 160.010 69.085 160.740 ;
        RECT 69.340 160.575 69.510 160.765 ;
        RECT 70.780 160.645 71.040 161.485 ;
        RECT 71.215 160.740 71.470 161.315 ;
        RECT 71.640 161.105 71.970 161.485 ;
        RECT 72.185 160.935 72.355 161.315 ;
        RECT 71.640 160.765 72.355 160.935 ;
        RECT 69.255 160.245 69.510 160.575 ;
        RECT 69.340 160.035 69.510 160.245 ;
        RECT 69.790 160.215 70.145 160.585 ;
        RECT 68.915 159.105 69.170 160.010 ;
        RECT 69.340 159.865 70.055 160.035 ;
        RECT 69.340 158.935 69.670 159.695 ;
        RECT 69.885 159.105 70.055 159.865 ;
        RECT 70.780 158.935 71.040 160.085 ;
        RECT 71.215 160.010 71.385 160.740 ;
        RECT 71.640 160.575 71.810 160.765 ;
        RECT 72.615 160.735 73.825 161.485 ;
        RECT 71.555 160.245 71.810 160.575 ;
        RECT 71.640 160.035 71.810 160.245 ;
        RECT 72.090 160.215 72.445 160.585 ;
        RECT 71.215 159.105 71.470 160.010 ;
        RECT 71.640 159.865 72.355 160.035 ;
        RECT 71.640 158.935 71.970 159.695 ;
        RECT 72.185 159.105 72.355 159.865 ;
        RECT 72.615 160.025 73.135 160.565 ;
        RECT 73.305 160.195 73.825 160.735 ;
        RECT 73.995 160.985 74.295 161.315 ;
        RECT 74.465 161.005 74.740 161.485 ;
        RECT 73.995 160.075 74.165 160.985 ;
        RECT 74.920 160.835 75.215 161.225 ;
        RECT 75.385 161.005 75.640 161.485 ;
        RECT 75.815 160.835 76.075 161.225 ;
        RECT 76.245 161.005 76.525 161.485 ;
        RECT 74.335 160.245 74.685 160.815 ;
        RECT 74.920 160.665 76.570 160.835 ;
        RECT 76.960 160.705 77.460 161.315 ;
        RECT 74.855 160.325 75.995 160.495 ;
        RECT 74.855 160.075 75.025 160.325 ;
        RECT 76.165 160.155 76.570 160.665 ;
        RECT 76.755 160.245 77.105 160.495 ;
        RECT 72.615 158.935 73.825 160.025 ;
        RECT 73.995 159.905 75.025 160.075 ;
        RECT 75.815 159.985 76.570 160.155 ;
        RECT 77.290 160.075 77.460 160.705 ;
        RECT 78.090 160.835 78.420 161.315 ;
        RECT 78.590 161.025 78.815 161.485 ;
        RECT 78.985 160.835 79.315 161.315 ;
        RECT 78.090 160.665 79.315 160.835 ;
        RECT 79.505 160.685 79.755 161.485 ;
        RECT 79.925 160.685 80.265 161.315 ;
        RECT 80.435 160.715 82.105 161.485 ;
        RECT 77.630 160.295 77.960 160.495 ;
        RECT 78.130 160.295 78.460 160.495 ;
        RECT 78.630 160.295 79.050 160.495 ;
        RECT 79.225 160.325 79.920 160.495 ;
        RECT 79.225 160.075 79.395 160.325 ;
        RECT 80.090 160.075 80.265 160.685 ;
        RECT 73.995 159.105 74.305 159.905 ;
        RECT 75.815 159.735 76.075 159.985 ;
        RECT 76.960 159.905 79.395 160.075 ;
        RECT 74.475 158.935 74.785 159.735 ;
        RECT 74.955 159.565 76.075 159.735 ;
        RECT 74.955 159.105 75.215 159.565 ;
        RECT 75.385 158.935 75.640 159.395 ;
        RECT 75.815 159.105 76.075 159.565 ;
        RECT 76.245 158.935 76.530 159.805 ;
        RECT 76.960 159.105 77.290 159.905 ;
        RECT 77.460 158.935 77.790 159.735 ;
        RECT 78.090 159.105 78.420 159.905 ;
        RECT 79.065 158.935 79.315 159.735 ;
        RECT 79.585 158.935 79.755 160.075 ;
        RECT 79.925 159.105 80.265 160.075 ;
        RECT 80.435 160.025 81.185 160.545 ;
        RECT 81.355 160.195 82.105 160.715 ;
        RECT 82.550 160.675 82.795 161.280 ;
        RECT 83.015 160.950 83.525 161.485 ;
        RECT 82.275 160.505 83.505 160.675 ;
        RECT 80.435 158.935 82.105 160.025 ;
        RECT 82.275 159.695 82.615 160.505 ;
        RECT 82.785 159.940 83.535 160.130 ;
        RECT 82.275 159.285 82.790 159.695 ;
        RECT 83.025 158.935 83.195 159.695 ;
        RECT 83.365 159.275 83.535 159.940 ;
        RECT 83.705 159.955 83.895 161.315 ;
        RECT 84.065 161.145 84.340 161.315 ;
        RECT 84.065 160.975 84.345 161.145 ;
        RECT 84.065 160.155 84.340 160.975 ;
        RECT 84.530 160.950 85.060 161.315 ;
        RECT 85.485 161.085 85.815 161.485 ;
        RECT 84.885 160.915 85.060 160.950 ;
        RECT 84.545 159.955 84.715 160.755 ;
        RECT 83.705 159.785 84.715 159.955 ;
        RECT 84.885 160.745 85.815 160.915 ;
        RECT 85.985 160.745 86.240 161.315 ;
        RECT 86.875 160.760 87.165 161.485 ;
        RECT 87.425 160.935 87.595 161.315 ;
        RECT 87.775 161.105 88.105 161.485 ;
        RECT 87.425 160.765 88.090 160.935 ;
        RECT 88.285 160.810 88.545 161.315 ;
        RECT 84.885 159.615 85.055 160.745 ;
        RECT 85.645 160.575 85.815 160.745 ;
        RECT 83.930 159.445 85.055 159.615 ;
        RECT 85.225 160.245 85.420 160.575 ;
        RECT 85.645 160.245 85.900 160.575 ;
        RECT 85.225 159.275 85.395 160.245 ;
        RECT 86.070 160.075 86.240 160.745 ;
        RECT 87.355 160.215 87.685 160.585 ;
        RECT 87.920 160.510 88.090 160.765 ;
        RECT 87.920 160.180 88.205 160.510 ;
        RECT 83.365 159.105 85.395 159.275 ;
        RECT 85.565 158.935 85.735 160.075 ;
        RECT 85.905 159.105 86.240 160.075 ;
        RECT 86.875 158.935 87.165 160.100 ;
        RECT 87.920 160.035 88.090 160.180 ;
        RECT 87.425 159.865 88.090 160.035 ;
        RECT 88.375 160.010 88.545 160.810 ;
        RECT 88.775 160.665 88.985 161.485 ;
        RECT 89.155 160.685 89.485 161.315 ;
        RECT 89.155 160.085 89.405 160.685 ;
        RECT 89.655 160.665 89.885 161.485 ;
        RECT 90.645 160.935 90.815 161.315 ;
        RECT 90.995 161.105 91.325 161.485 ;
        RECT 90.645 160.765 91.310 160.935 ;
        RECT 91.505 160.810 91.765 161.315 ;
        RECT 89.575 160.245 89.905 160.495 ;
        RECT 90.575 160.215 90.905 160.585 ;
        RECT 91.140 160.510 91.310 160.765 ;
        RECT 91.140 160.180 91.425 160.510 ;
        RECT 87.425 159.105 87.595 159.865 ;
        RECT 87.775 158.935 88.105 159.695 ;
        RECT 88.275 159.105 88.545 160.010 ;
        RECT 88.775 158.935 88.985 160.075 ;
        RECT 89.155 159.105 89.485 160.085 ;
        RECT 89.655 158.935 89.885 160.075 ;
        RECT 91.140 160.035 91.310 160.180 ;
        RECT 90.645 159.865 91.310 160.035 ;
        RECT 91.595 160.010 91.765 160.810 ;
        RECT 91.995 160.665 92.205 161.485 ;
        RECT 92.375 160.685 92.705 161.315 ;
        RECT 92.375 160.085 92.625 160.685 ;
        RECT 92.875 160.665 93.105 161.485 ;
        RECT 93.690 160.775 93.945 161.305 ;
        RECT 94.125 161.025 94.410 161.485 ;
        RECT 92.795 160.245 93.125 160.495 ;
        RECT 90.645 159.105 90.815 159.865 ;
        RECT 90.995 158.935 91.325 159.695 ;
        RECT 91.495 159.105 91.765 160.010 ;
        RECT 91.995 158.935 92.205 160.075 ;
        RECT 92.375 159.105 92.705 160.085 ;
        RECT 92.875 158.935 93.105 160.075 ;
        RECT 93.690 159.915 93.870 160.775 ;
        RECT 94.590 160.575 94.840 161.225 ;
        RECT 94.040 160.245 94.840 160.575 ;
        RECT 93.690 159.445 93.945 159.915 ;
        RECT 93.605 159.275 93.945 159.445 ;
        RECT 93.690 159.245 93.945 159.275 ;
        RECT 94.125 158.935 94.410 159.735 ;
        RECT 94.590 159.655 94.840 160.245 ;
        RECT 95.040 160.890 95.360 161.220 ;
        RECT 95.540 161.005 96.200 161.485 ;
        RECT 96.400 161.095 97.250 161.265 ;
        RECT 95.040 159.995 95.230 160.890 ;
        RECT 95.550 160.565 96.210 160.835 ;
        RECT 95.880 160.505 96.210 160.565 ;
        RECT 95.400 160.335 95.730 160.395 ;
        RECT 96.400 160.335 96.570 161.095 ;
        RECT 97.810 161.025 98.130 161.485 ;
        RECT 98.330 160.845 98.580 161.275 ;
        RECT 98.870 161.045 99.280 161.485 ;
        RECT 99.450 161.105 100.465 161.305 ;
        RECT 96.740 160.675 97.990 160.845 ;
        RECT 96.740 160.555 97.070 160.675 ;
        RECT 95.400 160.165 97.300 160.335 ;
        RECT 95.040 159.825 96.960 159.995 ;
        RECT 95.040 159.805 95.360 159.825 ;
        RECT 94.590 159.145 94.920 159.655 ;
        RECT 95.190 159.195 95.360 159.805 ;
        RECT 97.130 159.655 97.300 160.165 ;
        RECT 97.470 160.095 97.650 160.505 ;
        RECT 97.820 159.915 97.990 160.675 ;
        RECT 95.530 158.935 95.860 159.625 ;
        RECT 96.090 159.485 97.300 159.655 ;
        RECT 97.470 159.605 97.990 159.915 ;
        RECT 98.160 160.505 98.580 160.845 ;
        RECT 98.870 160.505 99.280 160.835 ;
        RECT 98.160 159.735 98.350 160.505 ;
        RECT 99.450 160.375 99.620 161.105 ;
        RECT 100.765 160.935 100.935 161.265 ;
        RECT 101.105 161.105 101.435 161.485 ;
        RECT 99.790 160.555 100.140 160.925 ;
        RECT 99.450 160.335 99.870 160.375 ;
        RECT 98.520 160.165 99.870 160.335 ;
        RECT 98.520 160.005 98.770 160.165 ;
        RECT 99.280 159.735 99.530 159.995 ;
        RECT 98.160 159.485 99.530 159.735 ;
        RECT 96.090 159.195 96.330 159.485 ;
        RECT 97.130 159.405 97.300 159.485 ;
        RECT 96.530 158.935 96.950 159.315 ;
        RECT 97.130 159.155 97.760 159.405 ;
        RECT 98.230 158.935 98.560 159.315 ;
        RECT 98.730 159.195 98.900 159.485 ;
        RECT 99.700 159.320 99.870 160.165 ;
        RECT 100.320 159.995 100.540 160.865 ;
        RECT 100.765 160.745 101.460 160.935 ;
        RECT 100.040 159.615 100.540 159.995 ;
        RECT 100.710 159.945 101.120 160.565 ;
        RECT 101.290 159.775 101.460 160.745 ;
        RECT 100.765 159.605 101.460 159.775 ;
        RECT 99.080 158.935 99.460 159.315 ;
        RECT 99.700 159.150 100.530 159.320 ;
        RECT 100.765 159.105 100.935 159.605 ;
        RECT 101.105 158.935 101.435 159.435 ;
        RECT 101.650 159.105 101.875 161.225 ;
        RECT 102.045 161.105 102.375 161.485 ;
        RECT 102.545 160.935 102.715 161.225 ;
        RECT 102.050 160.765 102.715 160.935 ;
        RECT 102.050 159.775 102.280 160.765 ;
        RECT 102.975 160.715 104.645 161.485 ;
        RECT 102.450 159.945 102.800 160.595 ;
        RECT 102.975 160.025 103.725 160.545 ;
        RECT 103.895 160.195 104.645 160.715 ;
        RECT 104.815 160.685 105.155 161.315 ;
        RECT 105.325 160.685 105.575 161.485 ;
        RECT 105.765 160.835 106.095 161.315 ;
        RECT 106.265 161.025 106.490 161.485 ;
        RECT 106.660 160.835 106.990 161.315 ;
        RECT 104.815 160.075 104.990 160.685 ;
        RECT 105.765 160.665 106.990 160.835 ;
        RECT 107.620 160.705 108.120 161.315 ;
        RECT 108.955 160.715 112.465 161.485 ;
        RECT 112.635 160.760 112.925 161.485 ;
        RECT 105.160 160.325 105.855 160.495 ;
        RECT 105.685 160.075 105.855 160.325 ;
        RECT 106.030 160.295 106.450 160.495 ;
        RECT 106.620 160.295 106.950 160.495 ;
        RECT 107.120 160.295 107.450 160.495 ;
        RECT 107.620 160.075 107.790 160.705 ;
        RECT 107.975 160.245 108.325 160.495 ;
        RECT 102.050 159.605 102.715 159.775 ;
        RECT 102.045 158.935 102.375 159.435 ;
        RECT 102.545 159.105 102.715 159.605 ;
        RECT 102.975 158.935 104.645 160.025 ;
        RECT 104.815 159.105 105.155 160.075 ;
        RECT 105.325 158.935 105.495 160.075 ;
        RECT 105.685 159.905 108.120 160.075 ;
        RECT 105.765 158.935 106.015 159.735 ;
        RECT 106.660 159.105 106.990 159.905 ;
        RECT 107.290 158.935 107.620 159.735 ;
        RECT 107.790 159.105 108.120 159.905 ;
        RECT 108.955 160.025 110.645 160.545 ;
        RECT 110.815 160.195 112.465 160.715 ;
        RECT 113.370 160.675 113.615 161.280 ;
        RECT 113.835 160.950 114.345 161.485 ;
        RECT 113.095 160.505 114.325 160.675 ;
        RECT 108.955 158.935 112.465 160.025 ;
        RECT 112.635 158.935 112.925 160.100 ;
        RECT 113.095 159.695 113.435 160.505 ;
        RECT 113.605 159.940 114.355 160.130 ;
        RECT 113.095 159.285 113.610 159.695 ;
        RECT 113.845 158.935 114.015 159.695 ;
        RECT 114.185 159.275 114.355 159.940 ;
        RECT 114.525 159.955 114.715 161.315 ;
        RECT 114.885 161.145 115.160 161.315 ;
        RECT 114.885 160.975 115.165 161.145 ;
        RECT 114.885 160.155 115.160 160.975 ;
        RECT 115.350 160.950 115.880 161.315 ;
        RECT 116.305 161.085 116.635 161.485 ;
        RECT 115.705 160.915 115.880 160.950 ;
        RECT 115.365 159.955 115.535 160.755 ;
        RECT 114.525 159.785 115.535 159.955 ;
        RECT 115.705 160.745 116.635 160.915 ;
        RECT 116.805 160.745 117.060 161.315 ;
        RECT 115.705 159.615 115.875 160.745 ;
        RECT 116.465 160.575 116.635 160.745 ;
        RECT 114.750 159.445 115.875 159.615 ;
        RECT 116.045 160.245 116.240 160.575 ;
        RECT 116.465 160.245 116.720 160.575 ;
        RECT 116.045 159.275 116.215 160.245 ;
        RECT 116.890 160.075 117.060 160.745 ;
        RECT 117.735 160.665 117.965 161.485 ;
        RECT 118.135 160.685 118.465 161.315 ;
        RECT 117.715 160.245 118.045 160.495 ;
        RECT 118.215 160.085 118.465 160.685 ;
        RECT 118.635 160.665 118.845 161.485 ;
        RECT 119.625 160.935 119.795 161.315 ;
        RECT 119.975 161.105 120.305 161.485 ;
        RECT 119.625 160.765 120.290 160.935 ;
        RECT 120.485 160.810 120.745 161.315 ;
        RECT 119.555 160.215 119.885 160.585 ;
        RECT 120.120 160.510 120.290 160.765 ;
        RECT 114.185 159.105 116.215 159.275 ;
        RECT 116.385 158.935 116.555 160.075 ;
        RECT 116.725 159.105 117.060 160.075 ;
        RECT 117.735 158.935 117.965 160.075 ;
        RECT 118.135 159.105 118.465 160.085 ;
        RECT 120.120 160.180 120.405 160.510 ;
        RECT 118.635 158.935 118.845 160.075 ;
        RECT 120.120 160.035 120.290 160.180 ;
        RECT 119.625 159.865 120.290 160.035 ;
        RECT 120.575 160.010 120.745 160.810 ;
        RECT 120.915 160.715 124.425 161.485 ;
        RECT 124.595 160.735 125.805 161.485 ;
        RECT 119.625 159.105 119.795 159.865 ;
        RECT 119.975 158.935 120.305 159.695 ;
        RECT 120.475 159.105 120.745 160.010 ;
        RECT 120.915 160.025 122.605 160.545 ;
        RECT 122.775 160.195 124.425 160.715 ;
        RECT 124.595 160.025 125.115 160.565 ;
        RECT 125.285 160.195 125.805 160.735 ;
        RECT 120.915 158.935 124.425 160.025 ;
        RECT 124.595 158.935 125.805 160.025 ;
        RECT 11.810 158.765 125.890 158.935 ;
        RECT 11.895 157.675 13.105 158.765 ;
        RECT 11.895 156.965 12.415 157.505 ;
        RECT 12.585 157.135 13.105 157.675 ;
        RECT 13.280 157.575 13.535 158.455 ;
        RECT 13.705 157.625 14.010 158.765 ;
        RECT 14.350 158.385 14.680 158.765 ;
        RECT 14.860 158.215 15.030 158.505 ;
        RECT 15.200 158.305 15.450 158.765 ;
        RECT 14.230 158.045 15.030 158.215 ;
        RECT 15.620 158.255 16.490 158.595 ;
        RECT 11.895 156.215 13.105 156.965 ;
        RECT 13.280 156.925 13.490 157.575 ;
        RECT 14.230 157.455 14.400 158.045 ;
        RECT 15.620 157.875 15.790 158.255 ;
        RECT 16.725 158.135 16.895 158.595 ;
        RECT 17.065 158.305 17.435 158.765 ;
        RECT 17.730 158.165 17.900 158.505 ;
        RECT 18.070 158.335 18.400 158.765 ;
        RECT 18.635 158.165 18.805 158.505 ;
        RECT 14.570 157.705 15.790 157.875 ;
        RECT 15.960 157.795 16.420 158.085 ;
        RECT 16.725 157.965 17.285 158.135 ;
        RECT 17.730 157.995 18.805 158.165 ;
        RECT 18.975 158.265 19.655 158.595 ;
        RECT 19.870 158.265 20.120 158.595 ;
        RECT 20.290 158.305 20.540 158.765 ;
        RECT 17.115 157.825 17.285 157.965 ;
        RECT 15.960 157.785 16.925 157.795 ;
        RECT 15.620 157.615 15.790 157.705 ;
        RECT 16.250 157.625 16.925 157.785 ;
        RECT 13.660 157.425 14.400 157.455 ;
        RECT 13.660 157.125 14.575 157.425 ;
        RECT 14.250 156.950 14.575 157.125 ;
        RECT 13.280 156.395 13.535 156.925 ;
        RECT 13.705 156.215 14.010 156.675 ;
        RECT 14.255 156.595 14.575 156.950 ;
        RECT 14.745 157.165 15.285 157.535 ;
        RECT 15.620 157.445 16.025 157.615 ;
        RECT 14.745 156.765 14.985 157.165 ;
        RECT 15.465 156.995 15.685 157.275 ;
        RECT 15.155 156.825 15.685 156.995 ;
        RECT 15.155 156.595 15.325 156.825 ;
        RECT 15.855 156.665 16.025 157.445 ;
        RECT 16.195 156.835 16.545 157.455 ;
        RECT 16.715 156.835 16.925 157.625 ;
        RECT 17.115 157.655 18.615 157.825 ;
        RECT 17.115 156.965 17.285 157.655 ;
        RECT 18.975 157.485 19.145 158.265 ;
        RECT 19.950 158.135 20.120 158.265 ;
        RECT 17.455 157.315 19.145 157.485 ;
        RECT 19.315 157.705 19.780 158.095 ;
        RECT 19.950 157.965 20.345 158.135 ;
        RECT 17.455 157.135 17.625 157.315 ;
        RECT 14.255 156.425 15.325 156.595 ;
        RECT 15.495 156.215 15.685 156.655 ;
        RECT 15.855 156.385 16.805 156.665 ;
        RECT 17.115 156.575 17.375 156.965 ;
        RECT 17.795 156.895 18.585 157.145 ;
        RECT 17.025 156.405 17.375 156.575 ;
        RECT 17.585 156.215 17.915 156.675 ;
        RECT 18.790 156.605 18.960 157.315 ;
        RECT 19.315 157.115 19.485 157.705 ;
        RECT 19.130 156.895 19.485 157.115 ;
        RECT 19.655 156.895 20.005 157.515 ;
        RECT 20.175 156.605 20.345 157.965 ;
        RECT 20.710 157.795 21.035 158.580 ;
        RECT 20.515 156.745 20.975 157.795 ;
        RECT 18.790 156.435 19.645 156.605 ;
        RECT 19.850 156.435 20.345 156.605 ;
        RECT 20.515 156.215 20.845 156.575 ;
        RECT 21.205 156.475 21.375 158.595 ;
        RECT 21.545 158.265 21.875 158.765 ;
        RECT 22.045 158.095 22.300 158.595 ;
        RECT 21.550 157.925 22.300 158.095 ;
        RECT 21.550 156.935 21.780 157.925 ;
        RECT 21.950 157.105 22.300 157.755 ;
        RECT 22.475 157.600 22.765 158.765 ;
        RECT 22.935 157.690 23.205 158.595 ;
        RECT 23.375 158.005 23.705 158.765 ;
        RECT 23.885 157.835 24.055 158.595 ;
        RECT 21.550 156.765 22.300 156.935 ;
        RECT 21.545 156.215 21.875 156.595 ;
        RECT 22.045 156.475 22.300 156.765 ;
        RECT 22.475 156.215 22.765 156.940 ;
        RECT 22.935 156.890 23.105 157.690 ;
        RECT 23.390 157.665 24.055 157.835 ;
        RECT 24.315 157.675 25.985 158.765 ;
        RECT 23.390 157.520 23.560 157.665 ;
        RECT 23.275 157.190 23.560 157.520 ;
        RECT 23.390 156.935 23.560 157.190 ;
        RECT 23.795 157.115 24.125 157.485 ;
        RECT 24.315 157.155 25.065 157.675 ;
        RECT 26.195 157.625 26.425 158.765 ;
        RECT 26.595 157.615 26.925 158.595 ;
        RECT 27.095 157.625 27.305 158.765 ;
        RECT 27.625 158.020 27.895 158.765 ;
        RECT 28.525 158.760 34.800 158.765 ;
        RECT 28.065 157.850 28.355 158.590 ;
        RECT 28.525 158.035 28.780 158.760 ;
        RECT 28.965 157.865 29.225 158.590 ;
        RECT 29.395 158.035 29.640 158.760 ;
        RECT 29.825 157.865 30.085 158.590 ;
        RECT 30.255 158.035 30.500 158.760 ;
        RECT 30.685 157.865 30.945 158.590 ;
        RECT 31.115 158.035 31.360 158.760 ;
        RECT 31.530 157.865 31.790 158.590 ;
        RECT 31.960 158.035 32.220 158.760 ;
        RECT 32.390 157.865 32.650 158.590 ;
        RECT 32.820 158.035 33.080 158.760 ;
        RECT 33.250 157.865 33.510 158.590 ;
        RECT 33.680 158.035 33.940 158.760 ;
        RECT 34.110 157.865 34.370 158.590 ;
        RECT 34.540 157.965 34.800 158.760 ;
        RECT 28.965 157.850 34.370 157.865 ;
        RECT 27.625 157.625 34.370 157.850 ;
        RECT 25.235 156.985 25.985 157.505 ;
        RECT 26.175 157.205 26.505 157.455 ;
        RECT 22.935 156.385 23.195 156.890 ;
        RECT 23.390 156.765 24.055 156.935 ;
        RECT 23.375 156.215 23.705 156.595 ;
        RECT 23.885 156.385 24.055 156.765 ;
        RECT 24.315 156.215 25.985 156.985 ;
        RECT 26.195 156.215 26.425 157.035 ;
        RECT 26.675 157.015 26.925 157.615 ;
        RECT 27.625 157.035 28.790 157.625 ;
        RECT 34.970 157.455 35.220 158.590 ;
        RECT 35.400 157.955 35.660 158.765 ;
        RECT 35.835 157.455 36.080 158.595 ;
        RECT 36.260 157.955 36.555 158.765 ;
        RECT 37.400 157.795 37.730 158.595 ;
        RECT 37.900 157.965 38.230 158.765 ;
        RECT 38.530 157.795 38.860 158.595 ;
        RECT 39.505 157.965 39.755 158.765 ;
        RECT 37.400 157.625 39.835 157.795 ;
        RECT 40.025 157.625 40.195 158.765 ;
        RECT 40.365 157.625 40.705 158.595 ;
        RECT 28.960 157.205 36.080 157.455 ;
        RECT 26.595 156.385 26.925 157.015 ;
        RECT 27.095 156.215 27.305 157.035 ;
        RECT 27.625 156.865 34.370 157.035 ;
        RECT 27.625 156.215 27.925 156.695 ;
        RECT 28.095 156.410 28.355 156.865 ;
        RECT 28.525 156.215 28.785 156.695 ;
        RECT 28.965 156.410 29.225 156.865 ;
        RECT 29.395 156.215 29.645 156.695 ;
        RECT 29.825 156.410 30.085 156.865 ;
        RECT 30.255 156.215 30.505 156.695 ;
        RECT 30.685 156.410 30.945 156.865 ;
        RECT 31.115 156.215 31.360 156.695 ;
        RECT 31.530 156.410 31.805 156.865 ;
        RECT 31.975 156.215 32.220 156.695 ;
        RECT 32.390 156.410 32.650 156.865 ;
        RECT 32.820 156.215 33.080 156.695 ;
        RECT 33.250 156.410 33.510 156.865 ;
        RECT 33.680 156.215 33.940 156.695 ;
        RECT 34.110 156.410 34.370 156.865 ;
        RECT 34.540 156.215 34.800 156.775 ;
        RECT 34.970 156.395 35.220 157.205 ;
        RECT 35.400 156.215 35.660 156.740 ;
        RECT 35.830 156.395 36.080 157.205 ;
        RECT 36.250 156.895 36.565 157.455 ;
        RECT 37.195 157.205 37.545 157.455 ;
        RECT 37.730 156.995 37.900 157.625 ;
        RECT 38.070 157.205 38.400 157.405 ;
        RECT 38.570 157.205 38.900 157.405 ;
        RECT 39.070 157.205 39.490 157.405 ;
        RECT 39.665 157.375 39.835 157.625 ;
        RECT 39.665 157.205 40.360 157.375 ;
        RECT 36.260 156.215 36.565 156.725 ;
        RECT 37.400 156.385 37.900 156.995 ;
        RECT 38.530 156.865 39.755 157.035 ;
        RECT 40.530 157.015 40.705 157.625 ;
        RECT 38.530 156.385 38.860 156.865 ;
        RECT 39.030 156.215 39.255 156.675 ;
        RECT 39.425 156.385 39.755 156.865 ;
        RECT 39.945 156.215 40.195 157.015 ;
        RECT 40.365 156.385 40.705 157.015 ;
        RECT 40.875 157.625 41.215 158.595 ;
        RECT 41.385 157.625 41.555 158.765 ;
        RECT 41.825 157.965 42.075 158.765 ;
        RECT 42.720 157.795 43.050 158.595 ;
        RECT 43.350 157.965 43.680 158.765 ;
        RECT 43.850 157.795 44.180 158.595 ;
        RECT 41.745 157.625 44.180 157.795 ;
        RECT 44.555 157.625 44.895 158.595 ;
        RECT 45.065 157.625 45.235 158.765 ;
        RECT 45.505 157.965 45.755 158.765 ;
        RECT 46.400 157.795 46.730 158.595 ;
        RECT 47.030 157.965 47.360 158.765 ;
        RECT 47.530 157.795 47.860 158.595 ;
        RECT 45.425 157.625 47.860 157.795 ;
        RECT 40.875 157.015 41.050 157.625 ;
        RECT 41.745 157.375 41.915 157.625 ;
        RECT 41.220 157.205 41.915 157.375 ;
        RECT 42.090 157.205 42.510 157.405 ;
        RECT 42.680 157.205 43.010 157.405 ;
        RECT 43.180 157.205 43.510 157.405 ;
        RECT 40.875 156.385 41.215 157.015 ;
        RECT 41.385 156.215 41.635 157.015 ;
        RECT 41.825 156.865 43.050 157.035 ;
        RECT 41.825 156.385 42.155 156.865 ;
        RECT 42.325 156.215 42.550 156.675 ;
        RECT 42.720 156.385 43.050 156.865 ;
        RECT 43.680 156.995 43.850 157.625 ;
        RECT 44.035 157.205 44.385 157.455 ;
        RECT 44.555 157.015 44.730 157.625 ;
        RECT 45.425 157.375 45.595 157.625 ;
        RECT 44.900 157.205 45.595 157.375 ;
        RECT 45.770 157.205 46.190 157.405 ;
        RECT 46.360 157.205 46.690 157.405 ;
        RECT 46.860 157.205 47.190 157.405 ;
        RECT 43.680 156.385 44.180 156.995 ;
        RECT 44.555 156.385 44.895 157.015 ;
        RECT 45.065 156.215 45.315 157.015 ;
        RECT 45.505 156.865 46.730 157.035 ;
        RECT 45.505 156.385 45.835 156.865 ;
        RECT 46.005 156.215 46.230 156.675 ;
        RECT 46.400 156.385 46.730 156.865 ;
        RECT 47.360 156.995 47.530 157.625 ;
        RECT 48.235 157.600 48.525 158.765 ;
        RECT 49.155 157.675 51.745 158.765 ;
        RECT 51.915 158.005 52.430 158.415 ;
        RECT 52.665 158.005 52.835 158.765 ;
        RECT 53.005 158.425 55.035 158.595 ;
        RECT 47.715 157.205 48.065 157.455 ;
        RECT 49.155 157.155 50.365 157.675 ;
        RECT 47.360 156.385 47.860 156.995 ;
        RECT 50.535 156.985 51.745 157.505 ;
        RECT 51.915 157.195 52.255 158.005 ;
        RECT 53.005 157.760 53.175 158.425 ;
        RECT 53.570 158.085 54.695 158.255 ;
        RECT 52.425 157.570 53.175 157.760 ;
        RECT 53.345 157.745 54.355 157.915 ;
        RECT 51.915 157.025 53.145 157.195 ;
        RECT 48.235 156.215 48.525 156.940 ;
        RECT 49.155 156.215 51.745 156.985 ;
        RECT 52.190 156.420 52.435 157.025 ;
        RECT 52.655 156.215 53.165 156.750 ;
        RECT 53.345 156.385 53.535 157.745 ;
        RECT 53.705 156.725 53.980 157.545 ;
        RECT 54.185 156.945 54.355 157.745 ;
        RECT 54.525 156.955 54.695 158.085 ;
        RECT 54.865 157.455 55.035 158.425 ;
        RECT 55.205 157.625 55.375 158.765 ;
        RECT 55.545 157.625 55.880 158.595 ;
        RECT 54.865 157.125 55.060 157.455 ;
        RECT 55.285 157.125 55.540 157.455 ;
        RECT 55.285 156.955 55.455 157.125 ;
        RECT 55.710 156.955 55.880 157.625 ;
        RECT 56.430 157.785 56.685 158.455 ;
        RECT 56.865 157.965 57.150 158.765 ;
        RECT 57.330 158.045 57.660 158.555 ;
        RECT 56.430 157.065 56.610 157.785 ;
        RECT 57.330 157.455 57.580 158.045 ;
        RECT 57.930 157.895 58.100 158.505 ;
        RECT 58.270 158.075 58.600 158.765 ;
        RECT 58.830 158.215 59.070 158.505 ;
        RECT 59.270 158.385 59.690 158.765 ;
        RECT 59.870 158.295 60.500 158.545 ;
        RECT 60.970 158.385 61.300 158.765 ;
        RECT 59.870 158.215 60.040 158.295 ;
        RECT 61.470 158.215 61.640 158.505 ;
        RECT 61.820 158.385 62.200 158.765 ;
        RECT 62.440 158.380 63.270 158.550 ;
        RECT 58.830 158.045 60.040 158.215 ;
        RECT 56.780 157.125 57.580 157.455 ;
        RECT 54.525 156.785 55.455 156.955 ;
        RECT 54.525 156.750 54.700 156.785 ;
        RECT 53.705 156.555 53.985 156.725 ;
        RECT 53.705 156.385 53.980 156.555 ;
        RECT 54.170 156.385 54.700 156.750 ;
        RECT 55.125 156.215 55.455 156.615 ;
        RECT 55.625 156.385 55.880 156.955 ;
        RECT 56.345 156.925 56.610 157.065 ;
        RECT 56.345 156.895 56.685 156.925 ;
        RECT 56.430 156.395 56.685 156.895 ;
        RECT 56.865 156.215 57.150 156.675 ;
        RECT 57.330 156.475 57.580 157.125 ;
        RECT 57.780 157.875 58.100 157.895 ;
        RECT 57.780 157.705 59.700 157.875 ;
        RECT 57.780 156.810 57.970 157.705 ;
        RECT 59.870 157.535 60.040 158.045 ;
        RECT 60.210 157.785 60.730 158.095 ;
        RECT 58.140 157.365 60.040 157.535 ;
        RECT 58.140 157.305 58.470 157.365 ;
        RECT 58.620 157.135 58.950 157.195 ;
        RECT 58.290 156.865 58.950 157.135 ;
        RECT 57.780 156.480 58.100 156.810 ;
        RECT 58.280 156.215 58.940 156.695 ;
        RECT 59.140 156.605 59.310 157.365 ;
        RECT 60.210 157.195 60.390 157.605 ;
        RECT 59.480 157.025 59.810 157.145 ;
        RECT 60.560 157.025 60.730 157.785 ;
        RECT 59.480 156.855 60.730 157.025 ;
        RECT 60.900 157.965 62.270 158.215 ;
        RECT 60.900 157.195 61.090 157.965 ;
        RECT 62.020 157.705 62.270 157.965 ;
        RECT 61.260 157.535 61.510 157.695 ;
        RECT 62.440 157.535 62.610 158.380 ;
        RECT 63.505 158.095 63.675 158.595 ;
        RECT 63.845 158.265 64.175 158.765 ;
        RECT 62.780 157.705 63.280 158.085 ;
        RECT 63.505 157.925 64.200 158.095 ;
        RECT 61.260 157.365 62.610 157.535 ;
        RECT 62.190 157.325 62.610 157.365 ;
        RECT 60.900 156.855 61.320 157.195 ;
        RECT 61.610 156.865 62.020 157.195 ;
        RECT 59.140 156.435 59.990 156.605 ;
        RECT 60.550 156.215 60.870 156.675 ;
        RECT 61.070 156.425 61.320 156.855 ;
        RECT 61.610 156.215 62.020 156.655 ;
        RECT 62.190 156.595 62.360 157.325 ;
        RECT 62.530 156.775 62.880 157.145 ;
        RECT 63.060 156.835 63.280 157.705 ;
        RECT 63.450 157.135 63.860 157.755 ;
        RECT 64.030 156.955 64.200 157.925 ;
        RECT 63.505 156.765 64.200 156.955 ;
        RECT 62.190 156.395 63.205 156.595 ;
        RECT 63.505 156.435 63.675 156.765 ;
        RECT 63.845 156.215 64.175 156.595 ;
        RECT 64.390 156.475 64.615 158.595 ;
        RECT 64.785 158.265 65.115 158.765 ;
        RECT 65.285 158.095 65.455 158.595 ;
        RECT 64.790 157.925 65.455 158.095 ;
        RECT 64.790 156.935 65.020 157.925 ;
        RECT 66.725 157.835 66.895 158.595 ;
        RECT 67.110 158.005 67.440 158.765 ;
        RECT 65.190 157.105 65.540 157.755 ;
        RECT 66.725 157.665 67.440 157.835 ;
        RECT 67.610 157.690 67.865 158.595 ;
        RECT 66.635 157.115 66.990 157.485 ;
        RECT 67.270 157.455 67.440 157.665 ;
        RECT 67.270 157.125 67.525 157.455 ;
        RECT 67.270 156.935 67.440 157.125 ;
        RECT 67.695 156.960 67.865 157.690 ;
        RECT 68.040 157.615 68.300 158.765 ;
        RECT 68.565 157.835 68.735 158.595 ;
        RECT 68.950 158.005 69.280 158.765 ;
        RECT 68.565 157.665 69.280 157.835 ;
        RECT 69.450 157.690 69.705 158.595 ;
        RECT 68.475 157.115 68.830 157.485 ;
        RECT 69.110 157.455 69.280 157.665 ;
        RECT 69.110 157.125 69.365 157.455 ;
        RECT 64.790 156.765 65.455 156.935 ;
        RECT 64.785 156.215 65.115 156.595 ;
        RECT 65.285 156.475 65.455 156.765 ;
        RECT 66.725 156.765 67.440 156.935 ;
        RECT 66.725 156.385 66.895 156.765 ;
        RECT 67.110 156.215 67.440 156.595 ;
        RECT 67.610 156.385 67.865 156.960 ;
        RECT 68.040 156.215 68.300 157.055 ;
        RECT 69.110 156.935 69.280 157.125 ;
        RECT 69.535 156.960 69.705 157.690 ;
        RECT 69.880 157.615 70.140 158.765 ;
        RECT 71.240 157.615 71.500 158.765 ;
        RECT 71.675 157.690 71.930 158.595 ;
        RECT 72.100 158.005 72.430 158.765 ;
        RECT 72.645 157.835 72.815 158.595 ;
        RECT 68.565 156.765 69.280 156.935 ;
        RECT 68.565 156.385 68.735 156.765 ;
        RECT 68.950 156.215 69.280 156.595 ;
        RECT 69.450 156.385 69.705 156.960 ;
        RECT 69.880 156.215 70.140 157.055 ;
        RECT 71.240 156.215 71.500 157.055 ;
        RECT 71.675 156.960 71.845 157.690 ;
        RECT 72.100 157.665 72.815 157.835 ;
        RECT 72.100 157.455 72.270 157.665 ;
        RECT 73.995 157.600 74.285 158.765 ;
        RECT 74.455 157.675 76.125 158.765 ;
        RECT 72.015 157.125 72.270 157.455 ;
        RECT 71.675 156.385 71.930 156.960 ;
        RECT 72.100 156.935 72.270 157.125 ;
        RECT 72.550 157.115 72.905 157.485 ;
        RECT 74.455 157.155 75.205 157.675 ;
        RECT 76.295 157.625 76.635 158.595 ;
        RECT 76.805 157.625 76.975 158.765 ;
        RECT 77.245 157.965 77.495 158.765 ;
        RECT 78.140 157.795 78.470 158.595 ;
        RECT 78.770 157.965 79.100 158.765 ;
        RECT 79.270 157.795 79.600 158.595 ;
        RECT 77.165 157.625 79.600 157.795 ;
        RECT 80.435 158.005 80.950 158.415 ;
        RECT 81.185 158.005 81.355 158.765 ;
        RECT 81.525 158.425 83.555 158.595 ;
        RECT 75.375 156.985 76.125 157.505 ;
        RECT 72.100 156.765 72.815 156.935 ;
        RECT 72.100 156.215 72.430 156.595 ;
        RECT 72.645 156.385 72.815 156.765 ;
        RECT 73.995 156.215 74.285 156.940 ;
        RECT 74.455 156.215 76.125 156.985 ;
        RECT 76.295 157.065 76.470 157.625 ;
        RECT 77.165 157.375 77.335 157.625 ;
        RECT 76.640 157.205 77.335 157.375 ;
        RECT 77.510 157.205 77.930 157.405 ;
        RECT 78.100 157.205 78.430 157.405 ;
        RECT 78.600 157.205 78.930 157.405 ;
        RECT 76.295 157.015 76.525 157.065 ;
        RECT 76.295 156.385 76.635 157.015 ;
        RECT 76.805 156.215 77.055 157.015 ;
        RECT 77.245 156.865 78.470 157.035 ;
        RECT 77.245 156.385 77.575 156.865 ;
        RECT 77.745 156.215 77.970 156.675 ;
        RECT 78.140 156.385 78.470 156.865 ;
        RECT 79.100 156.995 79.270 157.625 ;
        RECT 79.455 157.205 79.805 157.455 ;
        RECT 80.435 157.195 80.775 158.005 ;
        RECT 81.525 157.760 81.695 158.425 ;
        RECT 82.090 158.085 83.215 158.255 ;
        RECT 80.945 157.570 81.695 157.760 ;
        RECT 81.865 157.745 82.875 157.915 ;
        RECT 80.435 157.025 81.665 157.195 ;
        RECT 79.100 156.385 79.600 156.995 ;
        RECT 80.710 156.420 80.955 157.025 ;
        RECT 81.175 156.215 81.685 156.750 ;
        RECT 81.865 156.385 82.055 157.745 ;
        RECT 82.225 157.065 82.500 157.545 ;
        RECT 82.225 156.895 82.505 157.065 ;
        RECT 82.705 156.945 82.875 157.745 ;
        RECT 83.045 156.955 83.215 158.085 ;
        RECT 83.385 157.455 83.555 158.425 ;
        RECT 83.725 157.625 83.895 158.765 ;
        RECT 84.065 157.625 84.400 158.595 ;
        RECT 83.385 157.125 83.580 157.455 ;
        RECT 83.805 157.125 84.060 157.455 ;
        RECT 83.805 156.955 83.975 157.125 ;
        RECT 84.230 156.955 84.400 157.625 ;
        RECT 82.225 156.385 82.500 156.895 ;
        RECT 83.045 156.785 83.975 156.955 ;
        RECT 83.045 156.750 83.220 156.785 ;
        RECT 82.690 156.385 83.220 156.750 ;
        RECT 83.645 156.215 83.975 156.615 ;
        RECT 84.145 156.385 84.400 156.955 ;
        RECT 84.950 157.785 85.205 158.455 ;
        RECT 85.385 157.965 85.670 158.765 ;
        RECT 85.850 158.045 86.180 158.555 ;
        RECT 84.950 156.925 85.130 157.785 ;
        RECT 85.850 157.455 86.100 158.045 ;
        RECT 86.450 157.895 86.620 158.505 ;
        RECT 86.790 158.075 87.120 158.765 ;
        RECT 87.350 158.215 87.590 158.505 ;
        RECT 87.790 158.385 88.210 158.765 ;
        RECT 88.390 158.295 89.020 158.545 ;
        RECT 89.490 158.385 89.820 158.765 ;
        RECT 88.390 158.215 88.560 158.295 ;
        RECT 89.990 158.215 90.160 158.505 ;
        RECT 90.340 158.385 90.720 158.765 ;
        RECT 90.960 158.380 91.790 158.550 ;
        RECT 87.350 158.045 88.560 158.215 ;
        RECT 85.300 157.125 86.100 157.455 ;
        RECT 84.950 156.725 85.205 156.925 ;
        RECT 84.865 156.555 85.205 156.725 ;
        RECT 84.950 156.395 85.205 156.555 ;
        RECT 85.385 156.215 85.670 156.675 ;
        RECT 85.850 156.475 86.100 157.125 ;
        RECT 86.300 157.875 86.620 157.895 ;
        RECT 86.300 157.705 88.220 157.875 ;
        RECT 86.300 156.810 86.490 157.705 ;
        RECT 88.390 157.535 88.560 158.045 ;
        RECT 88.730 157.785 89.250 158.095 ;
        RECT 86.660 157.365 88.560 157.535 ;
        RECT 86.660 157.305 86.990 157.365 ;
        RECT 87.140 157.135 87.470 157.195 ;
        RECT 86.810 156.865 87.470 157.135 ;
        RECT 86.300 156.480 86.620 156.810 ;
        RECT 86.800 156.215 87.460 156.695 ;
        RECT 87.660 156.605 87.830 157.365 ;
        RECT 88.730 157.195 88.910 157.605 ;
        RECT 88.000 157.025 88.330 157.145 ;
        RECT 89.080 157.025 89.250 157.785 ;
        RECT 88.000 156.855 89.250 157.025 ;
        RECT 89.420 157.965 90.790 158.215 ;
        RECT 89.420 157.195 89.610 157.965 ;
        RECT 90.540 157.705 90.790 157.965 ;
        RECT 89.780 157.535 90.030 157.695 ;
        RECT 90.960 157.535 91.130 158.380 ;
        RECT 92.025 158.095 92.195 158.595 ;
        RECT 92.365 158.265 92.695 158.765 ;
        RECT 91.300 157.705 91.800 158.085 ;
        RECT 92.025 157.925 92.720 158.095 ;
        RECT 89.780 157.365 91.130 157.535 ;
        RECT 90.710 157.325 91.130 157.365 ;
        RECT 89.420 156.855 89.840 157.195 ;
        RECT 90.130 156.865 90.540 157.195 ;
        RECT 87.660 156.435 88.510 156.605 ;
        RECT 89.070 156.215 89.390 156.675 ;
        RECT 89.590 156.425 89.840 156.855 ;
        RECT 90.130 156.215 90.540 156.655 ;
        RECT 90.710 156.595 90.880 157.325 ;
        RECT 91.050 156.775 91.400 157.145 ;
        RECT 91.580 156.835 91.800 157.705 ;
        RECT 91.970 157.135 92.380 157.755 ;
        RECT 92.550 156.955 92.720 157.925 ;
        RECT 92.025 156.765 92.720 156.955 ;
        RECT 90.710 156.395 91.725 156.595 ;
        RECT 92.025 156.435 92.195 156.765 ;
        RECT 92.365 156.215 92.695 156.595 ;
        RECT 92.910 156.475 93.135 158.595 ;
        RECT 93.305 158.265 93.635 158.765 ;
        RECT 93.805 158.095 93.975 158.595 ;
        RECT 93.310 157.925 93.975 158.095 ;
        RECT 93.310 156.935 93.540 157.925 ;
        RECT 93.710 157.105 94.060 157.755 ;
        RECT 94.275 157.625 94.505 158.765 ;
        RECT 94.675 157.615 95.005 158.595 ;
        RECT 95.175 157.625 95.385 158.765 ;
        RECT 95.615 158.005 96.130 158.415 ;
        RECT 96.365 158.005 96.535 158.765 ;
        RECT 96.705 158.425 98.735 158.595 ;
        RECT 94.255 157.205 94.585 157.455 ;
        RECT 93.310 156.765 93.975 156.935 ;
        RECT 93.305 156.215 93.635 156.595 ;
        RECT 93.805 156.475 93.975 156.765 ;
        RECT 94.275 156.215 94.505 157.035 ;
        RECT 94.755 157.015 95.005 157.615 ;
        RECT 95.615 157.195 95.955 158.005 ;
        RECT 96.705 157.760 96.875 158.425 ;
        RECT 97.270 158.085 98.395 158.255 ;
        RECT 96.125 157.570 96.875 157.760 ;
        RECT 97.045 157.745 98.055 157.915 ;
        RECT 94.675 156.385 95.005 157.015 ;
        RECT 95.175 156.215 95.385 157.035 ;
        RECT 95.615 157.025 96.845 157.195 ;
        RECT 95.890 156.420 96.135 157.025 ;
        RECT 96.355 156.215 96.865 156.750 ;
        RECT 97.045 156.385 97.235 157.745 ;
        RECT 97.405 156.725 97.680 157.545 ;
        RECT 97.885 156.945 98.055 157.745 ;
        RECT 98.225 156.955 98.395 158.085 ;
        RECT 98.565 157.455 98.735 158.425 ;
        RECT 98.905 157.625 99.075 158.765 ;
        RECT 99.245 157.625 99.580 158.595 ;
        RECT 98.565 157.125 98.760 157.455 ;
        RECT 98.985 157.125 99.240 157.455 ;
        RECT 98.985 156.955 99.155 157.125 ;
        RECT 99.410 156.955 99.580 157.625 ;
        RECT 99.755 157.600 100.045 158.765 ;
        RECT 100.305 157.835 100.475 158.595 ;
        RECT 100.655 158.005 100.985 158.765 ;
        RECT 100.305 157.665 100.970 157.835 ;
        RECT 101.155 157.690 101.425 158.595 ;
        RECT 100.800 157.520 100.970 157.665 ;
        RECT 100.235 157.115 100.565 157.485 ;
        RECT 100.800 157.190 101.085 157.520 ;
        RECT 98.225 156.785 99.155 156.955 ;
        RECT 98.225 156.750 98.400 156.785 ;
        RECT 97.405 156.555 97.685 156.725 ;
        RECT 97.405 156.385 97.680 156.555 ;
        RECT 97.870 156.385 98.400 156.750 ;
        RECT 98.825 156.215 99.155 156.615 ;
        RECT 99.325 156.385 99.580 156.955 ;
        RECT 99.755 156.215 100.045 156.940 ;
        RECT 100.800 156.935 100.970 157.190 ;
        RECT 100.305 156.765 100.970 156.935 ;
        RECT 101.255 156.890 101.425 157.690 ;
        RECT 102.185 157.595 102.515 158.765 ;
        RECT 102.715 157.425 103.045 158.595 ;
        RECT 103.245 157.595 103.575 158.765 ;
        RECT 103.775 157.425 104.135 158.595 ;
        RECT 104.305 157.625 104.635 158.765 ;
        RECT 105.735 157.625 106.075 158.595 ;
        RECT 106.245 157.625 106.415 158.765 ;
        RECT 106.685 157.965 106.935 158.765 ;
        RECT 107.580 157.795 107.910 158.595 ;
        RECT 108.210 157.965 108.540 158.765 ;
        RECT 108.710 157.795 109.040 158.595 ;
        RECT 106.605 157.625 109.040 157.795 ;
        RECT 110.335 158.005 110.850 158.415 ;
        RECT 111.085 158.005 111.255 158.765 ;
        RECT 111.425 158.425 113.455 158.595 ;
        RECT 105.735 157.575 105.965 157.625 ;
        RECT 102.715 157.145 104.135 157.425 ;
        RECT 100.305 156.385 100.475 156.765 ;
        RECT 100.655 156.215 100.985 156.595 ;
        RECT 101.165 156.385 101.425 156.890 ;
        RECT 102.725 156.215 103.055 156.905 ;
        RECT 103.775 156.810 104.135 157.145 ;
        RECT 104.305 156.875 104.645 157.455 ;
        RECT 105.735 157.015 105.910 157.575 ;
        RECT 106.605 157.375 106.775 157.625 ;
        RECT 106.080 157.205 106.775 157.375 ;
        RECT 106.950 157.205 107.370 157.405 ;
        RECT 107.540 157.205 107.870 157.405 ;
        RECT 108.040 157.205 108.370 157.405 ;
        RECT 103.515 156.385 104.135 156.810 ;
        RECT 104.305 156.215 104.635 156.705 ;
        RECT 105.735 156.385 106.075 157.015 ;
        RECT 106.245 156.215 106.495 157.015 ;
        RECT 106.685 156.865 107.910 157.035 ;
        RECT 106.685 156.385 107.015 156.865 ;
        RECT 107.185 156.215 107.410 156.675 ;
        RECT 107.580 156.385 107.910 156.865 ;
        RECT 108.540 156.995 108.710 157.625 ;
        RECT 108.895 157.205 109.245 157.455 ;
        RECT 110.335 157.195 110.675 158.005 ;
        RECT 111.425 157.760 111.595 158.425 ;
        RECT 111.990 158.085 113.115 158.255 ;
        RECT 110.845 157.570 111.595 157.760 ;
        RECT 111.765 157.745 112.775 157.915 ;
        RECT 110.335 157.025 111.565 157.195 ;
        RECT 108.540 156.385 109.040 156.995 ;
        RECT 110.610 156.420 110.855 157.025 ;
        RECT 111.075 156.215 111.585 156.750 ;
        RECT 111.765 156.385 111.955 157.745 ;
        RECT 112.125 157.065 112.400 157.545 ;
        RECT 112.125 156.895 112.405 157.065 ;
        RECT 112.605 156.945 112.775 157.745 ;
        RECT 112.945 156.955 113.115 158.085 ;
        RECT 113.285 157.455 113.455 158.425 ;
        RECT 113.625 157.625 113.795 158.765 ;
        RECT 113.965 157.625 114.300 158.595 ;
        RECT 113.285 157.125 113.480 157.455 ;
        RECT 113.705 157.125 113.960 157.455 ;
        RECT 113.705 156.955 113.875 157.125 ;
        RECT 114.130 156.955 114.300 157.625 ;
        RECT 114.850 157.785 115.105 158.455 ;
        RECT 115.285 157.965 115.570 158.765 ;
        RECT 115.750 158.045 116.080 158.555 ;
        RECT 114.850 157.405 115.030 157.785 ;
        RECT 115.750 157.455 116.000 158.045 ;
        RECT 116.350 157.895 116.520 158.505 ;
        RECT 116.690 158.075 117.020 158.765 ;
        RECT 117.250 158.215 117.490 158.505 ;
        RECT 117.690 158.385 118.110 158.765 ;
        RECT 118.290 158.295 118.920 158.545 ;
        RECT 119.390 158.385 119.720 158.765 ;
        RECT 118.290 158.215 118.460 158.295 ;
        RECT 119.890 158.215 120.060 158.505 ;
        RECT 120.240 158.385 120.620 158.765 ;
        RECT 120.860 158.380 121.690 158.550 ;
        RECT 117.250 158.045 118.460 158.215 ;
        RECT 114.765 157.235 115.030 157.405 ;
        RECT 112.125 156.385 112.400 156.895 ;
        RECT 112.945 156.785 113.875 156.955 ;
        RECT 112.945 156.750 113.120 156.785 ;
        RECT 112.590 156.385 113.120 156.750 ;
        RECT 113.545 156.215 113.875 156.615 ;
        RECT 114.045 156.385 114.300 156.955 ;
        RECT 114.850 156.925 115.030 157.235 ;
        RECT 115.200 157.125 116.000 157.455 ;
        RECT 114.850 156.395 115.105 156.925 ;
        RECT 115.285 156.215 115.570 156.675 ;
        RECT 115.750 156.475 116.000 157.125 ;
        RECT 116.200 157.875 116.520 157.895 ;
        RECT 116.200 157.705 118.120 157.875 ;
        RECT 116.200 156.810 116.390 157.705 ;
        RECT 118.290 157.535 118.460 158.045 ;
        RECT 118.630 157.785 119.150 158.095 ;
        RECT 116.560 157.365 118.460 157.535 ;
        RECT 116.560 157.305 116.890 157.365 ;
        RECT 117.040 157.135 117.370 157.195 ;
        RECT 116.710 156.865 117.370 157.135 ;
        RECT 116.200 156.480 116.520 156.810 ;
        RECT 116.700 156.215 117.360 156.695 ;
        RECT 117.560 156.605 117.730 157.365 ;
        RECT 118.630 157.195 118.810 157.605 ;
        RECT 117.900 157.025 118.230 157.145 ;
        RECT 118.980 157.025 119.150 157.785 ;
        RECT 117.900 156.855 119.150 157.025 ;
        RECT 119.320 157.965 120.690 158.215 ;
        RECT 119.320 157.195 119.510 157.965 ;
        RECT 120.440 157.705 120.690 157.965 ;
        RECT 119.680 157.535 119.930 157.695 ;
        RECT 120.860 157.535 121.030 158.380 ;
        RECT 121.925 158.095 122.095 158.595 ;
        RECT 122.265 158.265 122.595 158.765 ;
        RECT 121.200 157.705 121.700 158.085 ;
        RECT 121.925 157.925 122.620 158.095 ;
        RECT 119.680 157.365 121.030 157.535 ;
        RECT 120.610 157.325 121.030 157.365 ;
        RECT 119.320 156.855 119.740 157.195 ;
        RECT 120.030 156.865 120.440 157.195 ;
        RECT 117.560 156.435 118.410 156.605 ;
        RECT 118.970 156.215 119.290 156.675 ;
        RECT 119.490 156.425 119.740 156.855 ;
        RECT 120.030 156.215 120.440 156.655 ;
        RECT 120.610 156.595 120.780 157.325 ;
        RECT 120.950 156.775 121.300 157.145 ;
        RECT 121.480 156.835 121.700 157.705 ;
        RECT 121.870 157.135 122.280 157.755 ;
        RECT 122.450 156.955 122.620 157.925 ;
        RECT 121.925 156.765 122.620 156.955 ;
        RECT 120.610 156.395 121.625 156.595 ;
        RECT 121.925 156.435 122.095 156.765 ;
        RECT 122.265 156.215 122.595 156.595 ;
        RECT 122.810 156.475 123.035 158.595 ;
        RECT 123.205 158.265 123.535 158.765 ;
        RECT 123.705 158.095 123.875 158.595 ;
        RECT 123.210 157.925 123.875 158.095 ;
        RECT 123.210 156.935 123.440 157.925 ;
        RECT 123.610 157.105 123.960 157.755 ;
        RECT 124.595 157.675 125.805 158.765 ;
        RECT 124.595 157.135 125.115 157.675 ;
        RECT 125.285 156.965 125.805 157.505 ;
        RECT 123.210 156.765 123.875 156.935 ;
        RECT 123.205 156.215 123.535 156.595 ;
        RECT 123.705 156.475 123.875 156.765 ;
        RECT 124.595 156.215 125.805 156.965 ;
        RECT 11.810 156.045 125.890 156.215 ;
        RECT 11.895 155.295 13.105 156.045 ;
        RECT 11.895 154.755 12.415 155.295 ;
        RECT 13.335 155.225 13.545 156.045 ;
        RECT 13.715 155.245 14.045 155.875 ;
        RECT 12.585 154.585 13.105 155.125 ;
        RECT 13.715 154.645 13.965 155.245 ;
        RECT 14.215 155.225 14.445 156.045 ;
        RECT 14.660 155.335 14.915 155.865 ;
        RECT 15.085 155.585 15.390 156.045 ;
        RECT 15.635 155.665 16.705 155.835 ;
        RECT 14.135 154.805 14.465 155.055 ;
        RECT 14.660 154.685 14.870 155.335 ;
        RECT 15.635 155.310 15.955 155.665 ;
        RECT 15.630 155.135 15.955 155.310 ;
        RECT 15.040 154.835 15.955 155.135 ;
        RECT 16.125 155.095 16.365 155.495 ;
        RECT 16.535 155.435 16.705 155.665 ;
        RECT 16.875 155.605 17.065 156.045 ;
        RECT 17.235 155.595 18.185 155.875 ;
        RECT 18.405 155.685 18.755 155.855 ;
        RECT 16.535 155.265 17.065 155.435 ;
        RECT 15.040 154.805 15.780 154.835 ;
        RECT 11.895 153.495 13.105 154.585 ;
        RECT 13.335 153.495 13.545 154.635 ;
        RECT 13.715 153.665 14.045 154.645 ;
        RECT 14.215 153.495 14.445 154.635 ;
        RECT 14.660 153.805 14.915 154.685 ;
        RECT 15.085 153.495 15.390 154.635 ;
        RECT 15.610 154.215 15.780 154.805 ;
        RECT 16.125 154.725 16.665 155.095 ;
        RECT 16.845 154.985 17.065 155.265 ;
        RECT 17.235 154.815 17.405 155.595 ;
        RECT 17.000 154.645 17.405 154.815 ;
        RECT 17.575 154.805 17.925 155.425 ;
        RECT 17.000 154.555 17.170 154.645 ;
        RECT 18.095 154.635 18.305 155.425 ;
        RECT 15.950 154.385 17.170 154.555 ;
        RECT 17.630 154.475 18.305 154.635 ;
        RECT 15.610 154.045 16.410 154.215 ;
        RECT 15.730 153.495 16.060 153.875 ;
        RECT 16.240 153.755 16.410 154.045 ;
        RECT 17.000 154.005 17.170 154.385 ;
        RECT 17.340 154.465 18.305 154.475 ;
        RECT 18.495 155.295 18.755 155.685 ;
        RECT 18.965 155.585 19.295 156.045 ;
        RECT 20.170 155.655 21.025 155.825 ;
        RECT 21.230 155.655 21.725 155.825 ;
        RECT 21.895 155.685 22.225 156.045 ;
        RECT 18.495 154.605 18.665 155.295 ;
        RECT 18.835 154.945 19.005 155.125 ;
        RECT 19.175 155.115 19.965 155.365 ;
        RECT 20.170 154.945 20.340 155.655 ;
        RECT 20.510 155.145 20.865 155.365 ;
        RECT 18.835 154.775 20.525 154.945 ;
        RECT 17.340 154.175 17.800 154.465 ;
        RECT 18.495 154.435 19.995 154.605 ;
        RECT 18.495 154.295 18.665 154.435 ;
        RECT 18.105 154.125 18.665 154.295 ;
        RECT 16.580 153.495 16.830 153.955 ;
        RECT 17.000 153.665 17.870 154.005 ;
        RECT 18.105 153.665 18.275 154.125 ;
        RECT 19.110 154.095 20.185 154.265 ;
        RECT 18.445 153.495 18.815 153.955 ;
        RECT 19.110 153.755 19.280 154.095 ;
        RECT 19.450 153.495 19.780 153.925 ;
        RECT 20.015 153.755 20.185 154.095 ;
        RECT 20.355 153.995 20.525 154.775 ;
        RECT 20.695 154.555 20.865 155.145 ;
        RECT 21.035 154.745 21.385 155.365 ;
        RECT 20.695 154.165 21.160 154.555 ;
        RECT 21.555 154.295 21.725 155.655 ;
        RECT 21.895 154.465 22.355 155.515 ;
        RECT 21.330 154.125 21.725 154.295 ;
        RECT 21.330 153.995 21.500 154.125 ;
        RECT 20.355 153.665 21.035 153.995 ;
        RECT 21.250 153.665 21.500 153.995 ;
        RECT 21.670 153.495 21.920 153.955 ;
        RECT 22.090 153.680 22.415 154.465 ;
        RECT 22.585 153.665 22.755 155.785 ;
        RECT 22.925 155.665 23.255 156.045 ;
        RECT 23.425 155.495 23.680 155.785 ;
        RECT 22.930 155.325 23.680 155.495 ;
        RECT 24.775 155.370 25.035 155.875 ;
        RECT 25.215 155.665 25.545 156.045 ;
        RECT 25.725 155.495 25.895 155.875 ;
        RECT 22.930 154.335 23.160 155.325 ;
        RECT 23.330 154.505 23.680 155.155 ;
        RECT 24.775 154.570 24.945 155.370 ;
        RECT 25.230 155.325 25.895 155.495 ;
        RECT 26.160 155.335 26.415 155.865 ;
        RECT 26.585 155.585 26.890 156.045 ;
        RECT 27.135 155.665 28.205 155.835 ;
        RECT 25.230 155.070 25.400 155.325 ;
        RECT 25.115 154.740 25.400 155.070 ;
        RECT 25.635 154.775 25.965 155.145 ;
        RECT 25.230 154.595 25.400 154.740 ;
        RECT 26.160 154.685 26.370 155.335 ;
        RECT 27.135 155.310 27.455 155.665 ;
        RECT 27.130 155.135 27.455 155.310 ;
        RECT 26.540 154.835 27.455 155.135 ;
        RECT 27.625 155.095 27.865 155.495 ;
        RECT 28.035 155.435 28.205 155.665 ;
        RECT 28.375 155.605 28.565 156.045 ;
        RECT 28.735 155.595 29.685 155.875 ;
        RECT 29.905 155.685 30.255 155.855 ;
        RECT 28.035 155.265 28.565 155.435 ;
        RECT 26.540 154.805 27.280 154.835 ;
        RECT 22.930 154.165 23.680 154.335 ;
        RECT 22.925 153.495 23.255 153.995 ;
        RECT 23.425 153.665 23.680 154.165 ;
        RECT 24.775 153.665 25.045 154.570 ;
        RECT 25.230 154.425 25.895 154.595 ;
        RECT 25.215 153.495 25.545 154.255 ;
        RECT 25.725 153.665 25.895 154.425 ;
        RECT 26.160 153.805 26.415 154.685 ;
        RECT 26.585 153.495 26.890 154.635 ;
        RECT 27.110 154.215 27.280 154.805 ;
        RECT 27.625 154.725 28.165 155.095 ;
        RECT 28.345 154.985 28.565 155.265 ;
        RECT 28.735 154.815 28.905 155.595 ;
        RECT 28.500 154.645 28.905 154.815 ;
        RECT 29.075 154.805 29.425 155.425 ;
        RECT 28.500 154.555 28.670 154.645 ;
        RECT 29.595 154.635 29.805 155.425 ;
        RECT 27.450 154.385 28.670 154.555 ;
        RECT 29.130 154.475 29.805 154.635 ;
        RECT 27.110 154.045 27.910 154.215 ;
        RECT 27.230 153.495 27.560 153.875 ;
        RECT 27.740 153.755 27.910 154.045 ;
        RECT 28.500 154.005 28.670 154.385 ;
        RECT 28.840 154.465 29.805 154.475 ;
        RECT 29.995 155.295 30.255 155.685 ;
        RECT 30.465 155.585 30.795 156.045 ;
        RECT 31.670 155.655 32.525 155.825 ;
        RECT 32.730 155.655 33.225 155.825 ;
        RECT 33.395 155.685 33.725 156.045 ;
        RECT 29.995 154.605 30.165 155.295 ;
        RECT 30.335 154.945 30.505 155.125 ;
        RECT 30.675 155.115 31.465 155.365 ;
        RECT 31.670 154.945 31.840 155.655 ;
        RECT 32.010 155.145 32.365 155.365 ;
        RECT 30.335 154.775 32.025 154.945 ;
        RECT 28.840 154.175 29.300 154.465 ;
        RECT 29.995 154.435 31.495 154.605 ;
        RECT 29.995 154.295 30.165 154.435 ;
        RECT 29.605 154.125 30.165 154.295 ;
        RECT 28.080 153.495 28.330 153.955 ;
        RECT 28.500 153.665 29.370 154.005 ;
        RECT 29.605 153.665 29.775 154.125 ;
        RECT 30.610 154.095 31.685 154.265 ;
        RECT 29.945 153.495 30.315 153.955 ;
        RECT 30.610 153.755 30.780 154.095 ;
        RECT 30.950 153.495 31.280 153.925 ;
        RECT 31.515 153.755 31.685 154.095 ;
        RECT 31.855 153.995 32.025 154.775 ;
        RECT 32.195 154.555 32.365 155.145 ;
        RECT 32.535 154.745 32.885 155.365 ;
        RECT 32.195 154.165 32.660 154.555 ;
        RECT 33.055 154.295 33.225 155.655 ;
        RECT 33.395 154.465 33.855 155.515 ;
        RECT 32.830 154.125 33.225 154.295 ;
        RECT 32.830 153.995 33.000 154.125 ;
        RECT 31.855 153.665 32.535 153.995 ;
        RECT 32.750 153.665 33.000 153.995 ;
        RECT 33.170 153.495 33.420 153.955 ;
        RECT 33.590 153.680 33.915 154.465 ;
        RECT 34.085 153.665 34.255 155.785 ;
        RECT 34.425 155.665 34.755 156.045 ;
        RECT 34.925 155.495 35.180 155.785 ;
        RECT 34.430 155.325 35.180 155.495 ;
        RECT 34.430 154.335 34.660 155.325 ;
        RECT 35.355 155.320 35.645 156.045 ;
        RECT 36.485 155.355 36.815 156.045 ;
        RECT 37.275 155.450 37.895 155.875 ;
        RECT 38.065 155.555 38.395 156.045 ;
        RECT 34.830 154.505 35.180 155.155 ;
        RECT 37.535 155.115 37.895 155.450 ;
        RECT 36.475 154.835 37.895 155.115 ;
        RECT 34.430 154.165 35.180 154.335 ;
        RECT 34.425 153.495 34.755 153.995 ;
        RECT 34.925 153.665 35.180 154.165 ;
        RECT 35.355 153.495 35.645 154.660 ;
        RECT 35.945 153.495 36.275 154.665 ;
        RECT 36.475 153.665 36.805 154.835 ;
        RECT 37.005 153.495 37.335 154.665 ;
        RECT 37.535 153.665 37.895 154.835 ;
        RECT 38.065 154.805 38.405 155.385 ;
        RECT 38.575 155.295 39.785 156.045 ;
        RECT 38.065 153.495 38.395 154.635 ;
        RECT 38.575 154.585 39.095 155.125 ;
        RECT 39.265 154.755 39.785 155.295 ;
        RECT 39.955 155.275 43.465 156.045 ;
        RECT 39.955 154.585 41.645 155.105 ;
        RECT 41.815 154.755 43.465 155.275 ;
        RECT 43.635 155.245 43.975 155.875 ;
        RECT 44.145 155.245 44.395 156.045 ;
        RECT 44.585 155.395 44.915 155.875 ;
        RECT 45.085 155.585 45.310 156.045 ;
        RECT 45.480 155.395 45.810 155.875 ;
        RECT 43.635 154.635 43.810 155.245 ;
        RECT 44.585 155.225 45.810 155.395 ;
        RECT 46.440 155.265 46.940 155.875 ;
        RECT 43.980 154.885 44.675 155.055 ;
        RECT 44.505 154.635 44.675 154.885 ;
        RECT 44.850 154.855 45.270 155.055 ;
        RECT 45.440 154.855 45.770 155.055 ;
        RECT 45.940 154.855 46.270 155.055 ;
        RECT 46.440 154.635 46.610 155.265 ;
        RECT 47.315 155.245 47.655 155.875 ;
        RECT 47.825 155.245 48.075 156.045 ;
        RECT 48.265 155.395 48.595 155.875 ;
        RECT 48.765 155.585 48.990 156.045 ;
        RECT 49.160 155.395 49.490 155.875 ;
        RECT 46.795 154.805 47.145 155.055 ;
        RECT 47.315 154.635 47.490 155.245 ;
        RECT 48.265 155.225 49.490 155.395 ;
        RECT 50.120 155.265 50.620 155.875 ;
        RECT 47.660 154.885 48.355 155.055 ;
        RECT 48.185 154.635 48.355 154.885 ;
        RECT 48.530 154.855 48.950 155.055 ;
        RECT 49.120 154.855 49.450 155.055 ;
        RECT 49.620 154.855 49.950 155.055 ;
        RECT 50.120 154.635 50.290 155.265 ;
        RECT 50.995 155.245 51.335 155.875 ;
        RECT 51.505 155.245 51.755 156.045 ;
        RECT 51.945 155.395 52.275 155.875 ;
        RECT 52.445 155.585 52.670 156.045 ;
        RECT 52.840 155.395 53.170 155.875 ;
        RECT 50.475 154.805 50.825 155.055 ;
        RECT 50.995 154.635 51.170 155.245 ;
        RECT 51.945 155.225 53.170 155.395 ;
        RECT 53.800 155.265 54.300 155.875 ;
        RECT 55.135 155.275 56.805 156.045 ;
        RECT 51.340 154.885 52.035 155.055 ;
        RECT 51.865 154.635 52.035 154.885 ;
        RECT 52.210 154.855 52.630 155.055 ;
        RECT 52.800 154.855 53.130 155.055 ;
        RECT 53.300 154.855 53.630 155.055 ;
        RECT 53.800 154.635 53.970 155.265 ;
        RECT 54.155 154.805 54.505 155.055 ;
        RECT 38.575 153.495 39.785 154.585 ;
        RECT 39.955 153.495 43.465 154.585 ;
        RECT 43.635 153.665 43.975 154.635 ;
        RECT 44.145 153.495 44.315 154.635 ;
        RECT 44.505 154.465 46.940 154.635 ;
        RECT 44.585 153.495 44.835 154.295 ;
        RECT 45.480 153.665 45.810 154.465 ;
        RECT 46.110 153.495 46.440 154.295 ;
        RECT 46.610 153.665 46.940 154.465 ;
        RECT 47.315 153.665 47.655 154.635 ;
        RECT 47.825 153.495 47.995 154.635 ;
        RECT 48.185 154.465 50.620 154.635 ;
        RECT 48.265 153.495 48.515 154.295 ;
        RECT 49.160 153.665 49.490 154.465 ;
        RECT 49.790 153.495 50.120 154.295 ;
        RECT 50.290 153.665 50.620 154.465 ;
        RECT 50.995 153.665 51.335 154.635 ;
        RECT 51.505 153.495 51.675 154.635 ;
        RECT 51.865 154.465 54.300 154.635 ;
        RECT 51.945 153.495 52.195 154.295 ;
        RECT 52.840 153.665 53.170 154.465 ;
        RECT 53.470 153.495 53.800 154.295 ;
        RECT 53.970 153.665 54.300 154.465 ;
        RECT 55.135 154.585 55.885 155.105 ;
        RECT 56.055 154.755 56.805 155.275 ;
        RECT 57.015 155.225 57.245 156.045 ;
        RECT 57.415 155.245 57.745 155.875 ;
        RECT 56.995 154.805 57.325 155.055 ;
        RECT 57.495 154.645 57.745 155.245 ;
        RECT 57.915 155.225 58.125 156.045 ;
        RECT 58.395 155.225 58.625 156.045 ;
        RECT 58.795 155.245 59.125 155.875 ;
        RECT 58.375 154.805 58.705 155.055 ;
        RECT 58.875 154.645 59.125 155.245 ;
        RECT 59.295 155.225 59.505 156.045 ;
        RECT 59.825 155.495 59.995 155.875 ;
        RECT 60.175 155.665 60.505 156.045 ;
        RECT 59.825 155.325 60.490 155.495 ;
        RECT 60.685 155.370 60.945 155.875 ;
        RECT 59.755 154.775 60.085 155.145 ;
        RECT 60.320 155.070 60.490 155.325 ;
        RECT 55.135 153.495 56.805 154.585 ;
        RECT 57.015 153.495 57.245 154.635 ;
        RECT 57.415 153.665 57.745 154.645 ;
        RECT 57.915 153.495 58.125 154.635 ;
        RECT 58.395 153.495 58.625 154.635 ;
        RECT 58.795 153.665 59.125 154.645 ;
        RECT 60.320 154.740 60.605 155.070 ;
        RECT 59.295 153.495 59.505 154.635 ;
        RECT 60.320 154.595 60.490 154.740 ;
        RECT 59.825 154.425 60.490 154.595 ;
        RECT 60.775 154.570 60.945 155.370 ;
        RECT 61.115 155.320 61.405 156.045 ;
        RECT 61.575 155.295 62.785 156.045 ;
        RECT 59.825 153.665 59.995 154.425 ;
        RECT 60.175 153.495 60.505 154.255 ;
        RECT 60.675 153.665 60.945 154.570 ;
        RECT 61.115 153.495 61.405 154.660 ;
        RECT 61.575 154.585 62.095 155.125 ;
        RECT 62.265 154.755 62.785 155.295 ;
        RECT 62.955 155.275 66.465 156.045 ;
        RECT 62.955 154.585 64.645 155.105 ;
        RECT 64.815 154.755 66.465 155.275 ;
        RECT 66.785 155.245 67.115 156.045 ;
        RECT 67.285 155.395 67.455 155.875 ;
        RECT 67.625 155.565 67.955 156.045 ;
        RECT 68.125 155.395 68.295 155.875 ;
        RECT 68.545 155.565 68.785 156.045 ;
        RECT 68.965 155.395 69.135 155.875 ;
        RECT 67.285 155.225 68.295 155.395 ;
        RECT 68.500 155.225 69.135 155.395 ;
        RECT 69.395 155.275 72.905 156.045 ;
        RECT 67.285 154.685 67.780 155.225 ;
        RECT 68.500 155.055 68.670 155.225 ;
        RECT 68.170 154.885 68.670 155.055 ;
        RECT 61.575 153.495 62.785 154.585 ;
        RECT 62.955 153.495 66.465 154.585 ;
        RECT 66.785 153.495 67.115 154.645 ;
        RECT 67.285 154.515 68.295 154.685 ;
        RECT 67.285 153.665 67.455 154.515 ;
        RECT 67.625 153.495 67.955 154.295 ;
        RECT 68.125 153.665 68.295 154.515 ;
        RECT 68.500 154.645 68.670 154.885 ;
        RECT 68.840 154.815 69.220 155.055 ;
        RECT 68.500 154.475 69.215 154.645 ;
        RECT 68.475 153.495 68.715 154.295 ;
        RECT 68.885 153.665 69.215 154.475 ;
        RECT 69.395 154.585 71.085 155.105 ;
        RECT 71.255 154.755 72.905 155.275 ;
        RECT 73.280 155.265 73.780 155.875 ;
        RECT 73.075 154.805 73.425 155.055 ;
        RECT 73.610 154.635 73.780 155.265 ;
        RECT 74.410 155.395 74.740 155.875 ;
        RECT 74.910 155.585 75.135 156.045 ;
        RECT 75.305 155.395 75.635 155.875 ;
        RECT 74.410 155.225 75.635 155.395 ;
        RECT 75.825 155.245 76.075 156.045 ;
        RECT 76.245 155.245 76.585 155.875 ;
        RECT 73.950 154.855 74.280 155.055 ;
        RECT 74.450 154.855 74.780 155.055 ;
        RECT 74.950 154.855 75.370 155.055 ;
        RECT 75.545 154.885 76.240 155.055 ;
        RECT 75.545 154.635 75.715 154.885 ;
        RECT 76.410 154.635 76.585 155.245 ;
        RECT 69.395 153.495 72.905 154.585 ;
        RECT 73.280 154.465 75.715 154.635 ;
        RECT 73.280 153.665 73.610 154.465 ;
        RECT 73.780 153.495 74.110 154.295 ;
        RECT 74.410 153.665 74.740 154.465 ;
        RECT 75.385 153.495 75.635 154.295 ;
        RECT 75.905 153.495 76.075 154.635 ;
        RECT 76.245 153.665 76.585 154.635 ;
        RECT 76.755 155.245 77.095 155.875 ;
        RECT 77.265 155.245 77.515 156.045 ;
        RECT 77.705 155.395 78.035 155.875 ;
        RECT 78.205 155.585 78.430 156.045 ;
        RECT 78.600 155.395 78.930 155.875 ;
        RECT 76.755 154.635 76.930 155.245 ;
        RECT 77.705 155.225 78.930 155.395 ;
        RECT 79.560 155.265 80.060 155.875 ;
        RECT 81.360 155.500 86.705 156.045 ;
        RECT 77.100 154.885 77.795 155.055 ;
        RECT 77.625 154.635 77.795 154.885 ;
        RECT 77.970 154.855 78.390 155.055 ;
        RECT 78.560 154.855 78.890 155.055 ;
        RECT 79.060 154.855 79.390 155.055 ;
        RECT 79.560 154.635 79.730 155.265 ;
        RECT 79.915 154.805 80.265 155.055 ;
        RECT 76.755 153.665 77.095 154.635 ;
        RECT 77.265 153.495 77.435 154.635 ;
        RECT 77.625 154.465 80.060 154.635 ;
        RECT 77.705 153.495 77.955 154.295 ;
        RECT 78.600 153.665 78.930 154.465 ;
        RECT 79.230 153.495 79.560 154.295 ;
        RECT 79.730 153.665 80.060 154.465 ;
        RECT 82.950 153.930 83.300 155.180 ;
        RECT 84.780 154.670 85.120 155.500 ;
        RECT 86.875 155.320 87.165 156.045 ;
        RECT 87.795 155.275 90.385 156.045 ;
        RECT 90.560 155.500 95.905 156.045 ;
        RECT 96.080 155.500 101.425 156.045 ;
        RECT 81.360 153.495 86.705 153.930 ;
        RECT 86.875 153.495 87.165 154.660 ;
        RECT 87.795 154.585 89.005 155.105 ;
        RECT 89.175 154.755 90.385 155.275 ;
        RECT 87.795 153.495 90.385 154.585 ;
        RECT 92.150 153.930 92.500 155.180 ;
        RECT 93.980 154.670 94.320 155.500 ;
        RECT 97.670 153.930 98.020 155.180 ;
        RECT 99.500 154.670 99.840 155.500 ;
        RECT 101.800 155.265 102.300 155.875 ;
        RECT 101.595 154.805 101.945 155.055 ;
        RECT 102.130 154.635 102.300 155.265 ;
        RECT 102.930 155.395 103.260 155.875 ;
        RECT 103.430 155.585 103.655 156.045 ;
        RECT 103.825 155.395 104.155 155.875 ;
        RECT 102.930 155.225 104.155 155.395 ;
        RECT 104.345 155.245 104.595 156.045 ;
        RECT 104.765 155.245 105.105 155.875 ;
        RECT 102.470 154.855 102.800 155.055 ;
        RECT 102.970 154.855 103.300 155.055 ;
        RECT 103.470 154.855 103.890 155.055 ;
        RECT 104.065 154.885 104.760 155.055 ;
        RECT 104.065 154.635 104.235 154.885 ;
        RECT 104.930 154.635 105.105 155.245 ;
        RECT 101.800 154.465 104.235 154.635 ;
        RECT 90.560 153.495 95.905 153.930 ;
        RECT 96.080 153.495 101.425 153.930 ;
        RECT 101.800 153.665 102.130 154.465 ;
        RECT 102.300 153.495 102.630 154.295 ;
        RECT 102.930 153.665 103.260 154.465 ;
        RECT 103.905 153.495 104.155 154.295 ;
        RECT 104.425 153.495 104.595 154.635 ;
        RECT 104.765 153.665 105.105 154.635 ;
        RECT 105.275 155.245 105.615 155.875 ;
        RECT 105.785 155.245 106.035 156.045 ;
        RECT 106.225 155.395 106.555 155.875 ;
        RECT 106.725 155.585 106.950 156.045 ;
        RECT 107.120 155.395 107.450 155.875 ;
        RECT 105.275 154.635 105.450 155.245 ;
        RECT 106.225 155.225 107.450 155.395 ;
        RECT 108.080 155.265 108.580 155.875 ;
        RECT 108.955 155.275 112.465 156.045 ;
        RECT 112.635 155.320 112.925 156.045 ;
        RECT 113.095 155.295 114.305 156.045 ;
        RECT 105.620 154.885 106.315 155.055 ;
        RECT 106.145 154.635 106.315 154.885 ;
        RECT 106.490 154.855 106.910 155.055 ;
        RECT 107.080 154.855 107.410 155.055 ;
        RECT 107.580 154.855 107.910 155.055 ;
        RECT 108.080 154.635 108.250 155.265 ;
        RECT 108.435 154.805 108.785 155.055 ;
        RECT 105.275 153.665 105.615 154.635 ;
        RECT 105.785 153.495 105.955 154.635 ;
        RECT 106.145 154.465 108.580 154.635 ;
        RECT 106.225 153.495 106.475 154.295 ;
        RECT 107.120 153.665 107.450 154.465 ;
        RECT 107.750 153.495 108.080 154.295 ;
        RECT 108.250 153.665 108.580 154.465 ;
        RECT 108.955 154.585 110.645 155.105 ;
        RECT 110.815 154.755 112.465 155.275 ;
        RECT 108.955 153.495 112.465 154.585 ;
        RECT 112.635 153.495 112.925 154.660 ;
        RECT 113.095 154.585 113.615 155.125 ;
        RECT 113.785 154.755 114.305 155.295 ;
        RECT 114.625 155.245 114.955 156.045 ;
        RECT 115.125 155.395 115.295 155.875 ;
        RECT 115.465 155.565 115.795 156.045 ;
        RECT 115.965 155.395 116.135 155.875 ;
        RECT 116.385 155.565 116.625 156.045 ;
        RECT 116.805 155.395 116.975 155.875 ;
        RECT 115.125 155.225 116.135 155.395 ;
        RECT 116.340 155.225 116.975 155.395 ;
        RECT 117.235 155.275 118.905 156.045 ;
        RECT 119.080 155.500 124.425 156.045 ;
        RECT 115.125 155.195 115.625 155.225 ;
        RECT 115.125 154.685 115.620 155.195 ;
        RECT 116.340 155.055 116.510 155.225 ;
        RECT 116.010 154.885 116.510 155.055 ;
        RECT 113.095 153.495 114.305 154.585 ;
        RECT 114.625 153.495 114.955 154.645 ;
        RECT 115.125 154.515 116.135 154.685 ;
        RECT 115.125 153.665 115.295 154.515 ;
        RECT 115.465 153.495 115.795 154.295 ;
        RECT 115.965 153.665 116.135 154.515 ;
        RECT 116.340 154.645 116.510 154.885 ;
        RECT 116.680 154.815 117.060 155.055 ;
        RECT 116.340 154.475 117.055 154.645 ;
        RECT 116.315 153.495 116.555 154.295 ;
        RECT 116.725 153.665 117.055 154.475 ;
        RECT 117.235 154.585 117.985 155.105 ;
        RECT 118.155 154.755 118.905 155.275 ;
        RECT 117.235 153.495 118.905 154.585 ;
        RECT 120.670 153.930 121.020 155.180 ;
        RECT 122.500 154.670 122.840 155.500 ;
        RECT 124.595 155.295 125.805 156.045 ;
        RECT 124.595 154.585 125.115 155.125 ;
        RECT 125.285 154.755 125.805 155.295 ;
        RECT 119.080 153.495 124.425 153.930 ;
        RECT 124.595 153.495 125.805 154.585 ;
        RECT 11.810 153.325 125.890 153.495 ;
        RECT 11.895 152.235 13.105 153.325 ;
        RECT 11.895 151.525 12.415 152.065 ;
        RECT 12.585 151.695 13.105 152.235 ;
        RECT 13.280 152.135 13.535 153.015 ;
        RECT 13.705 152.185 14.010 153.325 ;
        RECT 14.350 152.945 14.680 153.325 ;
        RECT 14.860 152.775 15.030 153.065 ;
        RECT 15.200 152.865 15.450 153.325 ;
        RECT 14.230 152.605 15.030 152.775 ;
        RECT 15.620 152.815 16.490 153.155 ;
        RECT 11.895 150.775 13.105 151.525 ;
        RECT 13.280 151.485 13.490 152.135 ;
        RECT 14.230 152.015 14.400 152.605 ;
        RECT 15.620 152.435 15.790 152.815 ;
        RECT 16.725 152.695 16.895 153.155 ;
        RECT 17.065 152.865 17.435 153.325 ;
        RECT 17.730 152.725 17.900 153.065 ;
        RECT 18.070 152.895 18.400 153.325 ;
        RECT 18.635 152.725 18.805 153.065 ;
        RECT 14.570 152.265 15.790 152.435 ;
        RECT 15.960 152.355 16.420 152.645 ;
        RECT 16.725 152.525 17.285 152.695 ;
        RECT 17.730 152.555 18.805 152.725 ;
        RECT 18.975 152.825 19.655 153.155 ;
        RECT 19.870 152.825 20.120 153.155 ;
        RECT 20.290 152.865 20.540 153.325 ;
        RECT 17.115 152.385 17.285 152.525 ;
        RECT 15.960 152.345 16.925 152.355 ;
        RECT 15.620 152.175 15.790 152.265 ;
        RECT 16.250 152.185 16.925 152.345 ;
        RECT 13.660 151.985 14.400 152.015 ;
        RECT 13.660 151.685 14.575 151.985 ;
        RECT 14.250 151.510 14.575 151.685 ;
        RECT 13.280 150.955 13.535 151.485 ;
        RECT 13.705 150.775 14.010 151.235 ;
        RECT 14.255 151.155 14.575 151.510 ;
        RECT 14.745 151.725 15.285 152.095 ;
        RECT 15.620 152.005 16.025 152.175 ;
        RECT 14.745 151.325 14.985 151.725 ;
        RECT 15.465 151.555 15.685 151.835 ;
        RECT 15.155 151.385 15.685 151.555 ;
        RECT 15.155 151.155 15.325 151.385 ;
        RECT 15.855 151.225 16.025 152.005 ;
        RECT 16.195 151.395 16.545 152.015 ;
        RECT 16.715 151.395 16.925 152.185 ;
        RECT 17.115 152.215 18.615 152.385 ;
        RECT 17.115 151.525 17.285 152.215 ;
        RECT 18.975 152.045 19.145 152.825 ;
        RECT 19.950 152.695 20.120 152.825 ;
        RECT 17.455 151.875 19.145 152.045 ;
        RECT 19.315 152.265 19.780 152.655 ;
        RECT 19.950 152.525 20.345 152.695 ;
        RECT 17.455 151.695 17.625 151.875 ;
        RECT 14.255 150.985 15.325 151.155 ;
        RECT 15.495 150.775 15.685 151.215 ;
        RECT 15.855 150.945 16.805 151.225 ;
        RECT 17.115 151.135 17.375 151.525 ;
        RECT 17.795 151.455 18.585 151.705 ;
        RECT 17.025 150.965 17.375 151.135 ;
        RECT 17.585 150.775 17.915 151.235 ;
        RECT 18.790 151.165 18.960 151.875 ;
        RECT 19.315 151.675 19.485 152.265 ;
        RECT 19.130 151.455 19.485 151.675 ;
        RECT 19.655 151.455 20.005 152.075 ;
        RECT 20.175 151.165 20.345 152.525 ;
        RECT 20.710 152.355 21.035 153.140 ;
        RECT 20.515 151.305 20.975 152.355 ;
        RECT 18.790 150.995 19.645 151.165 ;
        RECT 19.850 150.995 20.345 151.165 ;
        RECT 20.515 150.775 20.845 151.135 ;
        RECT 21.205 151.035 21.375 153.155 ;
        RECT 21.545 152.825 21.875 153.325 ;
        RECT 22.045 152.655 22.300 153.155 ;
        RECT 21.550 152.485 22.300 152.655 ;
        RECT 21.550 151.495 21.780 152.485 ;
        RECT 21.950 151.665 22.300 152.315 ;
        RECT 22.475 152.160 22.765 153.325 ;
        RECT 22.940 152.185 23.275 153.155 ;
        RECT 23.445 152.185 23.615 153.325 ;
        RECT 23.785 152.985 25.815 153.155 ;
        RECT 22.940 151.515 23.110 152.185 ;
        RECT 23.785 152.015 23.955 152.985 ;
        RECT 23.280 151.685 23.535 152.015 ;
        RECT 23.760 151.685 23.955 152.015 ;
        RECT 24.125 152.645 25.250 152.815 ;
        RECT 23.365 151.515 23.535 151.685 ;
        RECT 24.125 151.515 24.295 152.645 ;
        RECT 21.550 151.325 22.300 151.495 ;
        RECT 21.545 150.775 21.875 151.155 ;
        RECT 22.045 151.035 22.300 151.325 ;
        RECT 22.475 150.775 22.765 151.500 ;
        RECT 22.940 150.945 23.195 151.515 ;
        RECT 23.365 151.345 24.295 151.515 ;
        RECT 24.465 152.305 25.475 152.475 ;
        RECT 24.465 151.505 24.635 152.305 ;
        RECT 24.840 151.625 25.115 152.105 ;
        RECT 24.835 151.455 25.115 151.625 ;
        RECT 24.120 151.310 24.295 151.345 ;
        RECT 23.365 150.775 23.695 151.175 ;
        RECT 24.120 150.945 24.650 151.310 ;
        RECT 24.840 150.945 25.115 151.455 ;
        RECT 25.285 150.945 25.475 152.305 ;
        RECT 25.645 152.320 25.815 152.985 ;
        RECT 25.985 152.565 26.155 153.325 ;
        RECT 26.390 152.565 26.905 152.975 ;
        RECT 25.645 152.130 26.395 152.320 ;
        RECT 26.565 151.755 26.905 152.565 ;
        RECT 25.675 151.585 26.905 151.755 ;
        RECT 28.000 152.135 28.255 153.015 ;
        RECT 28.425 152.185 28.730 153.325 ;
        RECT 29.070 152.945 29.400 153.325 ;
        RECT 29.580 152.775 29.750 153.065 ;
        RECT 29.920 152.865 30.170 153.325 ;
        RECT 28.950 152.605 29.750 152.775 ;
        RECT 30.340 152.815 31.210 153.155 ;
        RECT 25.655 150.775 26.165 151.310 ;
        RECT 26.385 150.980 26.630 151.585 ;
        RECT 28.000 151.485 28.210 152.135 ;
        RECT 28.950 152.015 29.120 152.605 ;
        RECT 30.340 152.435 30.510 152.815 ;
        RECT 31.445 152.695 31.615 153.155 ;
        RECT 31.785 152.865 32.155 153.325 ;
        RECT 32.450 152.725 32.620 153.065 ;
        RECT 32.790 152.895 33.120 153.325 ;
        RECT 33.355 152.725 33.525 153.065 ;
        RECT 29.290 152.265 30.510 152.435 ;
        RECT 30.680 152.355 31.140 152.645 ;
        RECT 31.445 152.525 32.005 152.695 ;
        RECT 32.450 152.555 33.525 152.725 ;
        RECT 33.695 152.825 34.375 153.155 ;
        RECT 34.590 152.825 34.840 153.155 ;
        RECT 35.010 152.865 35.260 153.325 ;
        RECT 31.835 152.385 32.005 152.525 ;
        RECT 30.680 152.345 31.645 152.355 ;
        RECT 30.340 152.175 30.510 152.265 ;
        RECT 30.970 152.185 31.645 152.345 ;
        RECT 28.380 151.985 29.120 152.015 ;
        RECT 28.380 151.685 29.295 151.985 ;
        RECT 28.970 151.510 29.295 151.685 ;
        RECT 28.000 150.955 28.255 151.485 ;
        RECT 28.425 150.775 28.730 151.235 ;
        RECT 28.975 151.155 29.295 151.510 ;
        RECT 29.465 151.725 30.005 152.095 ;
        RECT 30.340 152.005 30.745 152.175 ;
        RECT 29.465 151.325 29.705 151.725 ;
        RECT 30.185 151.555 30.405 151.835 ;
        RECT 29.875 151.385 30.405 151.555 ;
        RECT 29.875 151.155 30.045 151.385 ;
        RECT 30.575 151.225 30.745 152.005 ;
        RECT 30.915 151.395 31.265 152.015 ;
        RECT 31.435 151.395 31.645 152.185 ;
        RECT 31.835 152.215 33.335 152.385 ;
        RECT 31.835 151.525 32.005 152.215 ;
        RECT 33.695 152.045 33.865 152.825 ;
        RECT 34.670 152.695 34.840 152.825 ;
        RECT 32.175 151.875 33.865 152.045 ;
        RECT 34.035 152.265 34.500 152.655 ;
        RECT 34.670 152.525 35.065 152.695 ;
        RECT 32.175 151.695 32.345 151.875 ;
        RECT 28.975 150.985 30.045 151.155 ;
        RECT 30.215 150.775 30.405 151.215 ;
        RECT 30.575 150.945 31.525 151.225 ;
        RECT 31.835 151.135 32.095 151.525 ;
        RECT 32.515 151.455 33.305 151.705 ;
        RECT 31.745 150.965 32.095 151.135 ;
        RECT 32.305 150.775 32.635 151.235 ;
        RECT 33.510 151.165 33.680 151.875 ;
        RECT 34.035 151.675 34.205 152.265 ;
        RECT 33.850 151.455 34.205 151.675 ;
        RECT 34.375 151.455 34.725 152.075 ;
        RECT 34.895 151.165 35.065 152.525 ;
        RECT 35.430 152.355 35.755 153.140 ;
        RECT 35.235 151.305 35.695 152.355 ;
        RECT 33.510 150.995 34.365 151.165 ;
        RECT 34.570 150.995 35.065 151.165 ;
        RECT 35.235 150.775 35.565 151.135 ;
        RECT 35.925 151.035 36.095 153.155 ;
        RECT 36.265 152.825 36.595 153.325 ;
        RECT 36.765 152.655 37.020 153.155 ;
        RECT 36.270 152.485 37.020 152.655 ;
        RECT 36.270 151.495 36.500 152.485 ;
        RECT 36.670 151.665 37.020 152.315 ;
        RECT 37.195 152.250 37.465 153.155 ;
        RECT 37.635 152.565 37.965 153.325 ;
        RECT 38.145 152.395 38.315 153.155 ;
        RECT 36.270 151.325 37.020 151.495 ;
        RECT 36.265 150.775 36.595 151.155 ;
        RECT 36.765 151.035 37.020 151.325 ;
        RECT 37.195 151.450 37.365 152.250 ;
        RECT 37.650 152.225 38.315 152.395 ;
        RECT 39.035 152.235 41.625 153.325 ;
        RECT 42.000 152.355 42.330 153.155 ;
        RECT 42.500 152.525 42.830 153.325 ;
        RECT 43.130 152.355 43.460 153.155 ;
        RECT 44.105 152.525 44.355 153.325 ;
        RECT 37.650 152.080 37.820 152.225 ;
        RECT 37.535 151.750 37.820 152.080 ;
        RECT 37.650 151.495 37.820 151.750 ;
        RECT 38.055 151.675 38.385 152.045 ;
        RECT 39.035 151.715 40.245 152.235 ;
        RECT 42.000 152.185 44.435 152.355 ;
        RECT 44.625 152.185 44.795 153.325 ;
        RECT 44.965 152.185 45.305 153.155 ;
        RECT 40.415 151.545 41.625 152.065 ;
        RECT 41.795 151.765 42.145 152.015 ;
        RECT 42.330 151.555 42.500 152.185 ;
        RECT 42.670 151.765 43.000 151.965 ;
        RECT 43.170 151.765 43.500 151.965 ;
        RECT 43.670 151.765 44.090 151.965 ;
        RECT 44.265 151.935 44.435 152.185 ;
        RECT 44.265 151.765 44.960 151.935 ;
        RECT 37.195 150.945 37.455 151.450 ;
        RECT 37.650 151.325 38.315 151.495 ;
        RECT 37.635 150.775 37.965 151.155 ;
        RECT 38.145 150.945 38.315 151.325 ;
        RECT 39.035 150.775 41.625 151.545 ;
        RECT 42.000 150.945 42.500 151.555 ;
        RECT 43.130 151.425 44.355 151.595 ;
        RECT 45.130 151.575 45.305 152.185 ;
        RECT 45.475 152.235 48.065 153.325 ;
        RECT 45.475 151.715 46.685 152.235 ;
        RECT 48.235 152.160 48.525 153.325 ;
        RECT 49.155 152.235 50.825 153.325 ;
        RECT 43.130 150.945 43.460 151.425 ;
        RECT 43.630 150.775 43.855 151.235 ;
        RECT 44.025 150.945 44.355 151.425 ;
        RECT 44.545 150.775 44.795 151.575 ;
        RECT 44.965 150.945 45.305 151.575 ;
        RECT 46.855 151.545 48.065 152.065 ;
        RECT 49.155 151.715 49.905 152.235 ;
        RECT 50.995 152.185 51.335 153.155 ;
        RECT 51.505 152.185 51.675 153.325 ;
        RECT 51.945 152.525 52.195 153.325 ;
        RECT 52.840 152.355 53.170 153.155 ;
        RECT 53.470 152.525 53.800 153.325 ;
        RECT 53.970 152.355 54.300 153.155 ;
        RECT 51.865 152.185 54.300 152.355 ;
        RECT 55.595 152.235 59.105 153.325 ;
        RECT 59.280 152.890 64.625 153.325 ;
        RECT 64.800 152.890 70.145 153.325 ;
        RECT 50.075 151.545 50.825 152.065 ;
        RECT 45.475 150.775 48.065 151.545 ;
        RECT 48.235 150.775 48.525 151.500 ;
        RECT 49.155 150.775 50.825 151.545 ;
        RECT 50.995 151.625 51.170 152.185 ;
        RECT 51.865 151.935 52.035 152.185 ;
        RECT 51.340 151.765 52.035 151.935 ;
        RECT 52.210 151.765 52.630 151.965 ;
        RECT 52.800 151.765 53.130 151.965 ;
        RECT 53.300 151.765 53.630 151.965 ;
        RECT 50.995 151.575 51.225 151.625 ;
        RECT 50.995 150.945 51.335 151.575 ;
        RECT 51.505 150.775 51.755 151.575 ;
        RECT 51.945 151.425 53.170 151.595 ;
        RECT 51.945 150.945 52.275 151.425 ;
        RECT 52.445 150.775 52.670 151.235 ;
        RECT 52.840 150.945 53.170 151.425 ;
        RECT 53.800 151.555 53.970 152.185 ;
        RECT 54.155 151.765 54.505 152.015 ;
        RECT 55.595 151.715 57.285 152.235 ;
        RECT 53.800 150.945 54.300 151.555 ;
        RECT 57.455 151.545 59.105 152.065 ;
        RECT 60.870 151.640 61.220 152.890 ;
        RECT 55.595 150.775 59.105 151.545 ;
        RECT 62.700 151.320 63.040 152.150 ;
        RECT 66.390 151.640 66.740 152.890 ;
        RECT 70.520 152.355 70.850 153.155 ;
        RECT 71.020 152.525 71.350 153.325 ;
        RECT 71.650 152.355 71.980 153.155 ;
        RECT 72.625 152.525 72.875 153.325 ;
        RECT 70.520 152.185 72.955 152.355 ;
        RECT 73.145 152.185 73.315 153.325 ;
        RECT 73.485 152.185 73.825 153.155 ;
        RECT 68.220 151.320 68.560 152.150 ;
        RECT 70.315 151.765 70.665 152.015 ;
        RECT 70.850 151.555 71.020 152.185 ;
        RECT 71.190 151.765 71.520 151.965 ;
        RECT 71.690 151.765 72.020 151.965 ;
        RECT 72.190 151.765 72.610 151.965 ;
        RECT 72.785 151.935 72.955 152.185 ;
        RECT 72.785 151.765 73.480 151.935 ;
        RECT 59.280 150.775 64.625 151.320 ;
        RECT 64.800 150.775 70.145 151.320 ;
        RECT 70.520 150.945 71.020 151.555 ;
        RECT 71.650 151.425 72.875 151.595 ;
        RECT 73.650 151.575 73.825 152.185 ;
        RECT 73.995 152.160 74.285 153.325 ;
        RECT 74.455 152.235 76.125 153.325 ;
        RECT 74.455 151.715 75.205 152.235 ;
        RECT 76.295 152.185 76.635 153.155 ;
        RECT 76.805 152.185 76.975 153.325 ;
        RECT 77.245 152.525 77.495 153.325 ;
        RECT 78.140 152.355 78.470 153.155 ;
        RECT 78.770 152.525 79.100 153.325 ;
        RECT 79.270 152.355 79.600 153.155 ;
        RECT 77.165 152.185 79.600 152.355 ;
        RECT 79.975 152.185 80.315 153.155 ;
        RECT 80.485 152.185 80.655 153.325 ;
        RECT 80.925 152.525 81.175 153.325 ;
        RECT 81.820 152.355 82.150 153.155 ;
        RECT 82.450 152.525 82.780 153.325 ;
        RECT 82.950 152.355 83.280 153.155 ;
        RECT 80.845 152.185 83.280 152.355 ;
        RECT 83.655 152.235 84.865 153.325 ;
        RECT 85.040 152.890 90.385 153.325 ;
        RECT 90.560 152.890 95.905 153.325 ;
        RECT 71.650 150.945 71.980 151.425 ;
        RECT 72.150 150.775 72.375 151.235 ;
        RECT 72.545 150.945 72.875 151.425 ;
        RECT 73.065 150.775 73.315 151.575 ;
        RECT 73.485 150.945 73.825 151.575 ;
        RECT 75.375 151.545 76.125 152.065 ;
        RECT 73.995 150.775 74.285 151.500 ;
        RECT 74.455 150.775 76.125 151.545 ;
        RECT 76.295 151.575 76.470 152.185 ;
        RECT 77.165 151.935 77.335 152.185 ;
        RECT 76.640 151.765 77.335 151.935 ;
        RECT 77.510 151.765 77.930 151.965 ;
        RECT 78.100 151.765 78.430 151.965 ;
        RECT 78.600 151.765 78.930 151.965 ;
        RECT 76.295 150.945 76.635 151.575 ;
        RECT 76.805 150.775 77.055 151.575 ;
        RECT 77.245 151.425 78.470 151.595 ;
        RECT 77.245 150.945 77.575 151.425 ;
        RECT 77.745 150.775 77.970 151.235 ;
        RECT 78.140 150.945 78.470 151.425 ;
        RECT 79.100 151.555 79.270 152.185 ;
        RECT 79.455 151.765 79.805 152.015 ;
        RECT 79.975 151.575 80.150 152.185 ;
        RECT 80.845 151.935 81.015 152.185 ;
        RECT 80.320 151.765 81.015 151.935 ;
        RECT 81.190 151.765 81.610 151.965 ;
        RECT 81.780 151.765 82.110 151.965 ;
        RECT 82.280 151.765 82.610 151.965 ;
        RECT 79.100 150.945 79.600 151.555 ;
        RECT 79.975 150.945 80.315 151.575 ;
        RECT 80.485 150.775 80.735 151.575 ;
        RECT 80.925 151.425 82.150 151.595 ;
        RECT 80.925 150.945 81.255 151.425 ;
        RECT 81.425 150.775 81.650 151.235 ;
        RECT 81.820 150.945 82.150 151.425 ;
        RECT 82.780 151.555 82.950 152.185 ;
        RECT 83.135 151.765 83.485 152.015 ;
        RECT 83.655 151.695 84.175 152.235 ;
        RECT 82.780 150.945 83.280 151.555 ;
        RECT 84.345 151.525 84.865 152.065 ;
        RECT 86.630 151.640 86.980 152.890 ;
        RECT 83.655 150.775 84.865 151.525 ;
        RECT 88.460 151.320 88.800 152.150 ;
        RECT 92.150 151.640 92.500 152.890 ;
        RECT 96.075 152.185 96.415 153.155 ;
        RECT 96.585 152.185 96.755 153.325 ;
        RECT 97.025 152.525 97.275 153.325 ;
        RECT 97.920 152.355 98.250 153.155 ;
        RECT 98.550 152.525 98.880 153.325 ;
        RECT 99.050 152.355 99.380 153.155 ;
        RECT 96.945 152.185 99.380 152.355 ;
        RECT 93.980 151.320 94.320 152.150 ;
        RECT 96.075 151.575 96.250 152.185 ;
        RECT 96.945 151.935 97.115 152.185 ;
        RECT 96.420 151.765 97.115 151.935 ;
        RECT 97.290 151.765 97.710 151.965 ;
        RECT 97.880 151.765 98.210 151.965 ;
        RECT 98.380 151.765 98.710 151.965 ;
        RECT 85.040 150.775 90.385 151.320 ;
        RECT 90.560 150.775 95.905 151.320 ;
        RECT 96.075 150.945 96.415 151.575 ;
        RECT 96.585 150.775 96.835 151.575 ;
        RECT 97.025 151.425 98.250 151.595 ;
        RECT 97.025 150.945 97.355 151.425 ;
        RECT 97.525 150.775 97.750 151.235 ;
        RECT 97.920 150.945 98.250 151.425 ;
        RECT 98.880 151.555 99.050 152.185 ;
        RECT 99.755 152.160 100.045 153.325 ;
        RECT 100.215 152.235 101.425 153.325 ;
        RECT 99.235 151.765 99.585 152.015 ;
        RECT 100.215 151.695 100.735 152.235 ;
        RECT 101.595 152.185 101.935 153.155 ;
        RECT 102.105 152.185 102.275 153.325 ;
        RECT 102.545 152.525 102.795 153.325 ;
        RECT 103.440 152.355 103.770 153.155 ;
        RECT 104.070 152.525 104.400 153.325 ;
        RECT 104.570 152.355 104.900 153.155 ;
        RECT 102.465 152.185 104.900 152.355 ;
        RECT 106.195 152.185 106.535 153.155 ;
        RECT 106.705 152.185 106.875 153.325 ;
        RECT 107.145 152.525 107.395 153.325 ;
        RECT 108.040 152.355 108.370 153.155 ;
        RECT 108.670 152.525 109.000 153.325 ;
        RECT 109.170 152.355 109.500 153.155 ;
        RECT 107.065 152.185 109.500 152.355 ;
        RECT 110.345 152.345 110.675 153.155 ;
        RECT 110.845 152.525 111.085 153.325 ;
        RECT 98.880 150.945 99.380 151.555 ;
        RECT 100.905 151.525 101.425 152.065 ;
        RECT 99.755 150.775 100.045 151.500 ;
        RECT 100.215 150.775 101.425 151.525 ;
        RECT 101.595 151.575 101.770 152.185 ;
        RECT 102.465 151.935 102.635 152.185 ;
        RECT 101.940 151.765 102.635 151.935 ;
        RECT 102.810 151.765 103.230 151.965 ;
        RECT 103.400 151.765 103.730 151.965 ;
        RECT 103.900 151.765 104.230 151.965 ;
        RECT 101.595 150.945 101.935 151.575 ;
        RECT 102.105 150.775 102.355 151.575 ;
        RECT 102.545 151.425 103.770 151.595 ;
        RECT 102.545 150.945 102.875 151.425 ;
        RECT 103.045 150.775 103.270 151.235 ;
        RECT 103.440 150.945 103.770 151.425 ;
        RECT 104.400 151.555 104.570 152.185 ;
        RECT 104.755 151.765 105.105 152.015 ;
        RECT 106.195 151.575 106.370 152.185 ;
        RECT 107.065 151.935 107.235 152.185 ;
        RECT 106.540 151.765 107.235 151.935 ;
        RECT 107.410 151.765 107.830 151.965 ;
        RECT 108.000 151.765 108.330 151.965 ;
        RECT 108.500 151.765 108.830 151.965 ;
        RECT 104.400 150.945 104.900 151.555 ;
        RECT 106.195 150.945 106.535 151.575 ;
        RECT 106.705 150.775 106.955 151.575 ;
        RECT 107.145 151.425 108.370 151.595 ;
        RECT 107.145 150.945 107.475 151.425 ;
        RECT 107.645 150.775 107.870 151.235 ;
        RECT 108.040 150.945 108.370 151.425 ;
        RECT 109.000 151.555 109.170 152.185 ;
        RECT 110.345 152.175 111.060 152.345 ;
        RECT 109.355 151.765 109.705 152.015 ;
        RECT 110.340 151.765 110.720 152.005 ;
        RECT 110.890 151.935 111.060 152.175 ;
        RECT 111.265 152.305 111.435 153.155 ;
        RECT 111.605 152.525 111.935 153.325 ;
        RECT 112.105 152.305 112.275 153.155 ;
        RECT 111.265 152.135 112.275 152.305 ;
        RECT 112.445 152.175 112.775 153.325 ;
        RECT 110.890 151.765 111.390 151.935 ;
        RECT 110.890 151.595 111.060 151.765 ;
        RECT 111.780 151.595 112.275 152.135 ;
        RECT 109.000 150.945 109.500 151.555 ;
        RECT 110.425 151.425 111.060 151.595 ;
        RECT 111.265 151.425 112.275 151.595 ;
        RECT 113.100 152.135 113.355 153.015 ;
        RECT 113.525 152.185 113.830 153.325 ;
        RECT 114.170 152.945 114.500 153.325 ;
        RECT 114.680 152.775 114.850 153.065 ;
        RECT 115.020 152.865 115.270 153.325 ;
        RECT 114.050 152.605 114.850 152.775 ;
        RECT 115.440 152.815 116.310 153.155 ;
        RECT 110.425 150.945 110.595 151.425 ;
        RECT 110.775 150.775 111.015 151.255 ;
        RECT 111.265 150.945 111.435 151.425 ;
        RECT 111.605 150.775 111.935 151.255 ;
        RECT 112.105 150.945 112.275 151.425 ;
        RECT 112.445 150.775 112.775 151.575 ;
        RECT 113.100 151.485 113.310 152.135 ;
        RECT 114.050 152.015 114.220 152.605 ;
        RECT 115.440 152.435 115.610 152.815 ;
        RECT 116.545 152.695 116.715 153.155 ;
        RECT 116.885 152.865 117.255 153.325 ;
        RECT 117.550 152.725 117.720 153.065 ;
        RECT 117.890 152.895 118.220 153.325 ;
        RECT 118.455 152.725 118.625 153.065 ;
        RECT 114.390 152.265 115.610 152.435 ;
        RECT 115.780 152.355 116.240 152.645 ;
        RECT 116.545 152.525 117.105 152.695 ;
        RECT 117.550 152.555 118.625 152.725 ;
        RECT 118.795 152.825 119.475 153.155 ;
        RECT 119.690 152.825 119.940 153.155 ;
        RECT 120.110 152.865 120.360 153.325 ;
        RECT 116.935 152.385 117.105 152.525 ;
        RECT 115.780 152.345 116.745 152.355 ;
        RECT 115.440 152.175 115.610 152.265 ;
        RECT 116.070 152.185 116.745 152.345 ;
        RECT 113.480 151.985 114.220 152.015 ;
        RECT 113.480 151.685 114.395 151.985 ;
        RECT 114.070 151.510 114.395 151.685 ;
        RECT 113.100 150.955 113.355 151.485 ;
        RECT 113.525 150.775 113.830 151.235 ;
        RECT 114.075 151.155 114.395 151.510 ;
        RECT 114.565 151.725 115.105 152.095 ;
        RECT 115.440 152.005 115.845 152.175 ;
        RECT 114.565 151.325 114.805 151.725 ;
        RECT 115.285 151.555 115.505 151.835 ;
        RECT 114.975 151.385 115.505 151.555 ;
        RECT 114.975 151.155 115.145 151.385 ;
        RECT 115.675 151.225 115.845 152.005 ;
        RECT 116.015 151.395 116.365 152.015 ;
        RECT 116.535 151.395 116.745 152.185 ;
        RECT 116.935 152.215 118.435 152.385 ;
        RECT 116.935 151.525 117.105 152.215 ;
        RECT 118.795 152.045 118.965 152.825 ;
        RECT 119.770 152.695 119.940 152.825 ;
        RECT 117.275 151.875 118.965 152.045 ;
        RECT 119.135 152.265 119.600 152.655 ;
        RECT 119.770 152.525 120.165 152.695 ;
        RECT 117.275 151.695 117.445 151.875 ;
        RECT 114.075 150.985 115.145 151.155 ;
        RECT 115.315 150.775 115.505 151.215 ;
        RECT 115.675 150.945 116.625 151.225 ;
        RECT 116.935 151.135 117.195 151.525 ;
        RECT 117.615 151.455 118.405 151.705 ;
        RECT 116.845 150.965 117.195 151.135 ;
        RECT 117.405 150.775 117.735 151.235 ;
        RECT 118.610 151.165 118.780 151.875 ;
        RECT 119.135 151.675 119.305 152.265 ;
        RECT 118.950 151.455 119.305 151.675 ;
        RECT 119.475 151.455 119.825 152.075 ;
        RECT 119.995 151.165 120.165 152.525 ;
        RECT 120.530 152.355 120.855 153.140 ;
        RECT 120.335 151.305 120.795 152.355 ;
        RECT 118.610 150.995 119.465 151.165 ;
        RECT 119.670 150.995 120.165 151.165 ;
        RECT 120.335 150.775 120.665 151.135 ;
        RECT 121.025 151.035 121.195 153.155 ;
        RECT 121.365 152.825 121.695 153.325 ;
        RECT 121.865 152.655 122.120 153.155 ;
        RECT 121.370 152.485 122.120 152.655 ;
        RECT 121.370 151.495 121.600 152.485 ;
        RECT 121.770 151.665 122.120 152.315 ;
        RECT 122.755 152.235 124.425 153.325 ;
        RECT 124.595 152.235 125.805 153.325 ;
        RECT 122.755 151.715 123.505 152.235 ;
        RECT 123.675 151.545 124.425 152.065 ;
        RECT 124.595 151.695 125.115 152.235 ;
        RECT 121.370 151.325 122.120 151.495 ;
        RECT 121.365 150.775 121.695 151.155 ;
        RECT 121.865 151.035 122.120 151.325 ;
        RECT 122.755 150.775 124.425 151.545 ;
        RECT 125.285 151.525 125.805 152.065 ;
        RECT 124.595 150.775 125.805 151.525 ;
        RECT 11.810 150.605 125.890 150.775 ;
        RECT 11.895 149.855 13.105 150.605 ;
        RECT 11.895 149.315 12.415 149.855 ;
        RECT 13.735 149.835 15.405 150.605 ;
        RECT 12.585 149.145 13.105 149.685 ;
        RECT 11.895 148.055 13.105 149.145 ;
        RECT 13.735 149.145 14.485 149.665 ;
        RECT 14.655 149.315 15.405 149.835 ;
        RECT 15.615 149.785 15.845 150.605 ;
        RECT 16.015 149.805 16.345 150.435 ;
        RECT 15.595 149.365 15.925 149.615 ;
        RECT 16.095 149.205 16.345 149.805 ;
        RECT 16.515 149.785 16.725 150.605 ;
        RECT 17.015 149.785 17.225 150.605 ;
        RECT 17.395 149.805 17.725 150.435 ;
        RECT 13.735 148.055 15.405 149.145 ;
        RECT 15.615 148.055 15.845 149.195 ;
        RECT 16.015 148.225 16.345 149.205 ;
        RECT 17.395 149.205 17.645 149.805 ;
        RECT 17.895 149.785 18.125 150.605 ;
        RECT 18.425 150.055 18.595 150.435 ;
        RECT 18.775 150.225 19.105 150.605 ;
        RECT 18.425 149.885 19.090 150.055 ;
        RECT 19.285 149.930 19.545 150.435 ;
        RECT 17.815 149.365 18.145 149.615 ;
        RECT 18.355 149.335 18.685 149.705 ;
        RECT 18.920 149.630 19.090 149.885 ;
        RECT 18.920 149.300 19.205 149.630 ;
        RECT 16.515 148.055 16.725 149.195 ;
        RECT 17.015 148.055 17.225 149.195 ;
        RECT 17.395 148.225 17.725 149.205 ;
        RECT 17.895 148.055 18.125 149.195 ;
        RECT 18.920 149.155 19.090 149.300 ;
        RECT 18.425 148.985 19.090 149.155 ;
        RECT 19.375 149.130 19.545 149.930 ;
        RECT 18.425 148.225 18.595 148.985 ;
        RECT 18.775 148.055 19.105 148.815 ;
        RECT 19.275 148.225 19.545 149.130 ;
        RECT 19.720 149.865 19.975 150.435 ;
        RECT 20.145 150.205 20.475 150.605 ;
        RECT 20.900 150.070 21.430 150.435 ;
        RECT 21.620 150.265 21.895 150.435 ;
        RECT 21.615 150.095 21.895 150.265 ;
        RECT 20.900 150.035 21.075 150.070 ;
        RECT 20.145 149.865 21.075 150.035 ;
        RECT 19.720 149.195 19.890 149.865 ;
        RECT 20.145 149.695 20.315 149.865 ;
        RECT 20.060 149.365 20.315 149.695 ;
        RECT 20.540 149.365 20.735 149.695 ;
        RECT 19.720 148.225 20.055 149.195 ;
        RECT 20.225 148.055 20.395 149.195 ;
        RECT 20.565 148.395 20.735 149.365 ;
        RECT 20.905 148.735 21.075 149.865 ;
        RECT 21.245 149.075 21.415 149.875 ;
        RECT 21.620 149.275 21.895 150.095 ;
        RECT 22.065 149.075 22.255 150.435 ;
        RECT 22.435 150.070 22.945 150.605 ;
        RECT 23.165 149.795 23.410 150.400 ;
        RECT 23.855 149.835 25.525 150.605 ;
        RECT 22.455 149.625 23.685 149.795 ;
        RECT 21.245 148.905 22.255 149.075 ;
        RECT 22.425 149.060 23.175 149.250 ;
        RECT 20.905 148.565 22.030 148.735 ;
        RECT 22.425 148.395 22.595 149.060 ;
        RECT 23.345 148.815 23.685 149.625 ;
        RECT 20.565 148.225 22.595 148.395 ;
        RECT 22.765 148.055 22.935 148.815 ;
        RECT 23.170 148.405 23.685 148.815 ;
        RECT 23.855 149.145 24.605 149.665 ;
        RECT 24.775 149.315 25.525 149.835 ;
        RECT 25.735 149.785 25.965 150.605 ;
        RECT 26.135 149.805 26.465 150.435 ;
        RECT 25.715 149.365 26.045 149.615 ;
        RECT 26.215 149.205 26.465 149.805 ;
        RECT 26.635 149.785 26.845 150.605 ;
        RECT 27.350 149.795 27.595 150.400 ;
        RECT 27.815 150.070 28.325 150.605 ;
        RECT 23.855 148.055 25.525 149.145 ;
        RECT 25.735 148.055 25.965 149.195 ;
        RECT 26.135 148.225 26.465 149.205 ;
        RECT 27.075 149.625 28.305 149.795 ;
        RECT 26.635 148.055 26.845 149.195 ;
        RECT 27.075 148.815 27.415 149.625 ;
        RECT 27.585 149.060 28.335 149.250 ;
        RECT 27.075 148.405 27.590 148.815 ;
        RECT 27.825 148.055 27.995 148.815 ;
        RECT 28.165 148.395 28.335 149.060 ;
        RECT 28.505 149.075 28.695 150.435 ;
        RECT 28.865 150.265 29.140 150.435 ;
        RECT 28.865 150.095 29.145 150.265 ;
        RECT 28.865 149.275 29.140 150.095 ;
        RECT 29.330 150.070 29.860 150.435 ;
        RECT 30.285 150.205 30.615 150.605 ;
        RECT 29.685 150.035 29.860 150.070 ;
        RECT 29.345 149.075 29.515 149.875 ;
        RECT 28.505 148.905 29.515 149.075 ;
        RECT 29.685 149.865 30.615 150.035 ;
        RECT 30.785 149.865 31.040 150.435 ;
        RECT 29.685 148.735 29.855 149.865 ;
        RECT 30.445 149.695 30.615 149.865 ;
        RECT 28.730 148.565 29.855 148.735 ;
        RECT 30.025 149.365 30.220 149.695 ;
        RECT 30.445 149.365 30.700 149.695 ;
        RECT 30.025 148.395 30.195 149.365 ;
        RECT 30.870 149.195 31.040 149.865 ;
        RECT 31.490 149.795 31.735 150.400 ;
        RECT 31.955 150.070 32.465 150.605 ;
        RECT 28.165 148.225 30.195 148.395 ;
        RECT 30.365 148.055 30.535 149.195 ;
        RECT 30.705 148.225 31.040 149.195 ;
        RECT 31.215 149.625 32.445 149.795 ;
        RECT 31.215 148.815 31.555 149.625 ;
        RECT 31.725 149.060 32.475 149.250 ;
        RECT 31.215 148.405 31.730 148.815 ;
        RECT 31.965 148.055 32.135 148.815 ;
        RECT 32.305 148.395 32.475 149.060 ;
        RECT 32.645 149.075 32.835 150.435 ;
        RECT 33.005 150.265 33.280 150.435 ;
        RECT 33.005 150.095 33.285 150.265 ;
        RECT 33.005 149.275 33.280 150.095 ;
        RECT 33.470 150.070 34.000 150.435 ;
        RECT 34.425 150.205 34.755 150.605 ;
        RECT 33.825 150.035 34.000 150.070 ;
        RECT 33.485 149.075 33.655 149.875 ;
        RECT 32.645 148.905 33.655 149.075 ;
        RECT 33.825 149.865 34.755 150.035 ;
        RECT 34.925 149.865 35.180 150.435 ;
        RECT 35.355 149.880 35.645 150.605 ;
        RECT 35.815 149.930 36.075 150.435 ;
        RECT 36.255 150.225 36.585 150.605 ;
        RECT 36.765 150.055 36.935 150.435 ;
        RECT 33.825 148.735 33.995 149.865 ;
        RECT 34.585 149.695 34.755 149.865 ;
        RECT 32.870 148.565 33.995 148.735 ;
        RECT 34.165 149.365 34.360 149.695 ;
        RECT 34.585 149.365 34.840 149.695 ;
        RECT 34.165 148.395 34.335 149.365 ;
        RECT 35.010 149.195 35.180 149.865 ;
        RECT 32.305 148.225 34.335 148.395 ;
        RECT 34.505 148.055 34.675 149.195 ;
        RECT 34.845 148.225 35.180 149.195 ;
        RECT 35.355 148.055 35.645 149.220 ;
        RECT 35.815 149.130 35.985 149.930 ;
        RECT 36.270 149.885 36.935 150.055 ;
        RECT 36.270 149.630 36.440 149.885 ;
        RECT 37.195 149.835 38.865 150.605 ;
        RECT 36.155 149.300 36.440 149.630 ;
        RECT 36.675 149.335 37.005 149.705 ;
        RECT 36.270 149.155 36.440 149.300 ;
        RECT 35.815 148.225 36.085 149.130 ;
        RECT 36.270 148.985 36.935 149.155 ;
        RECT 36.255 148.055 36.585 148.815 ;
        RECT 36.765 148.225 36.935 148.985 ;
        RECT 37.195 149.145 37.945 149.665 ;
        RECT 38.115 149.315 38.865 149.835 ;
        RECT 39.035 149.805 39.375 150.435 ;
        RECT 39.545 149.805 39.795 150.605 ;
        RECT 39.985 149.955 40.315 150.435 ;
        RECT 40.485 150.145 40.710 150.605 ;
        RECT 40.880 149.955 41.210 150.435 ;
        RECT 39.035 149.195 39.210 149.805 ;
        RECT 39.985 149.785 41.210 149.955 ;
        RECT 41.840 149.825 42.340 150.435 ;
        RECT 42.920 149.825 43.420 150.435 ;
        RECT 39.380 149.445 40.075 149.615 ;
        RECT 39.905 149.195 40.075 149.445 ;
        RECT 40.250 149.415 40.670 149.615 ;
        RECT 40.840 149.415 41.170 149.615 ;
        RECT 41.340 149.415 41.670 149.615 ;
        RECT 41.840 149.195 42.010 149.825 ;
        RECT 42.195 149.365 42.545 149.615 ;
        RECT 42.715 149.365 43.065 149.615 ;
        RECT 43.250 149.195 43.420 149.825 ;
        RECT 44.050 149.955 44.380 150.435 ;
        RECT 44.550 150.145 44.775 150.605 ;
        RECT 44.945 149.955 45.275 150.435 ;
        RECT 44.050 149.785 45.275 149.955 ;
        RECT 45.465 149.805 45.715 150.605 ;
        RECT 45.885 149.805 46.225 150.435 ;
        RECT 46.855 149.835 49.445 150.605 ;
        RECT 43.590 149.415 43.920 149.615 ;
        RECT 44.090 149.415 44.420 149.615 ;
        RECT 44.590 149.415 45.010 149.615 ;
        RECT 45.185 149.445 45.880 149.615 ;
        RECT 45.185 149.195 45.355 149.445 ;
        RECT 46.050 149.195 46.225 149.805 ;
        RECT 37.195 148.055 38.865 149.145 ;
        RECT 39.035 148.225 39.375 149.195 ;
        RECT 39.545 148.055 39.715 149.195 ;
        RECT 39.905 149.025 42.340 149.195 ;
        RECT 39.985 148.055 40.235 148.855 ;
        RECT 40.880 148.225 41.210 149.025 ;
        RECT 41.510 148.055 41.840 148.855 ;
        RECT 42.010 148.225 42.340 149.025 ;
        RECT 42.920 149.025 45.355 149.195 ;
        RECT 42.920 148.225 43.250 149.025 ;
        RECT 43.420 148.055 43.750 148.855 ;
        RECT 44.050 148.225 44.380 149.025 ;
        RECT 45.025 148.055 45.275 148.855 ;
        RECT 45.545 148.055 45.715 149.195 ;
        RECT 45.885 148.225 46.225 149.195 ;
        RECT 46.855 149.145 48.065 149.665 ;
        RECT 48.235 149.315 49.445 149.835 ;
        RECT 49.615 149.805 49.955 150.435 ;
        RECT 50.125 149.805 50.375 150.605 ;
        RECT 50.565 149.955 50.895 150.435 ;
        RECT 51.065 150.145 51.290 150.605 ;
        RECT 51.460 149.955 51.790 150.435 ;
        RECT 49.615 149.195 49.790 149.805 ;
        RECT 50.565 149.785 51.790 149.955 ;
        RECT 52.420 149.825 52.920 150.435 ;
        RECT 53.755 149.835 55.425 150.605 ;
        RECT 55.600 150.060 60.945 150.605 ;
        RECT 49.960 149.445 50.655 149.615 ;
        RECT 50.485 149.195 50.655 149.445 ;
        RECT 50.830 149.415 51.250 149.615 ;
        RECT 51.420 149.415 51.750 149.615 ;
        RECT 51.920 149.415 52.250 149.615 ;
        RECT 52.420 149.195 52.590 149.825 ;
        RECT 52.775 149.365 53.125 149.615 ;
        RECT 46.855 148.055 49.445 149.145 ;
        RECT 49.615 148.225 49.955 149.195 ;
        RECT 50.125 148.055 50.295 149.195 ;
        RECT 50.485 149.025 52.920 149.195 ;
        RECT 50.565 148.055 50.815 148.855 ;
        RECT 51.460 148.225 51.790 149.025 ;
        RECT 52.090 148.055 52.420 148.855 ;
        RECT 52.590 148.225 52.920 149.025 ;
        RECT 53.755 149.145 54.505 149.665 ;
        RECT 54.675 149.315 55.425 149.835 ;
        RECT 53.755 148.055 55.425 149.145 ;
        RECT 57.190 148.490 57.540 149.740 ;
        RECT 59.020 149.230 59.360 150.060 ;
        RECT 61.115 149.880 61.405 150.605 ;
        RECT 61.575 149.835 63.245 150.605 ;
        RECT 55.600 148.055 60.945 148.490 ;
        RECT 61.115 148.055 61.405 149.220 ;
        RECT 61.575 149.145 62.325 149.665 ;
        RECT 62.495 149.315 63.245 149.835 ;
        RECT 63.455 149.785 63.685 150.605 ;
        RECT 63.855 149.805 64.185 150.435 ;
        RECT 63.435 149.365 63.765 149.615 ;
        RECT 63.935 149.205 64.185 149.805 ;
        RECT 64.355 149.785 64.565 150.605 ;
        RECT 65.345 150.055 65.515 150.435 ;
        RECT 65.695 150.225 66.025 150.605 ;
        RECT 65.345 149.885 66.010 150.055 ;
        RECT 66.205 149.930 66.465 150.435 ;
        RECT 65.275 149.335 65.605 149.705 ;
        RECT 65.840 149.630 66.010 149.885 ;
        RECT 61.575 148.055 63.245 149.145 ;
        RECT 63.455 148.055 63.685 149.195 ;
        RECT 63.855 148.225 64.185 149.205 ;
        RECT 65.840 149.300 66.125 149.630 ;
        RECT 64.355 148.055 64.565 149.195 ;
        RECT 65.840 149.155 66.010 149.300 ;
        RECT 65.345 148.985 66.010 149.155 ;
        RECT 66.295 149.130 66.465 149.930 ;
        RECT 66.635 149.835 69.225 150.605 ;
        RECT 69.485 150.055 69.655 150.435 ;
        RECT 69.870 150.225 70.200 150.605 ;
        RECT 69.485 149.885 70.200 150.055 ;
        RECT 65.345 148.225 65.515 148.985 ;
        RECT 65.695 148.055 66.025 148.815 ;
        RECT 66.195 148.225 66.465 149.130 ;
        RECT 66.635 149.145 67.845 149.665 ;
        RECT 68.015 149.315 69.225 149.835 ;
        RECT 69.395 149.335 69.750 149.705 ;
        RECT 70.030 149.695 70.200 149.885 ;
        RECT 70.370 149.860 70.625 150.435 ;
        RECT 70.030 149.365 70.285 149.695 ;
        RECT 70.030 149.155 70.200 149.365 ;
        RECT 66.635 148.055 69.225 149.145 ;
        RECT 69.485 148.985 70.200 149.155 ;
        RECT 70.455 149.130 70.625 149.860 ;
        RECT 70.800 149.765 71.060 150.605 ;
        RECT 71.240 149.765 71.500 150.605 ;
        RECT 71.675 149.860 71.930 150.435 ;
        RECT 72.100 150.225 72.430 150.605 ;
        RECT 72.645 150.055 72.815 150.435 ;
        RECT 72.100 149.885 72.815 150.055 ;
        RECT 69.485 148.225 69.655 148.985 ;
        RECT 69.870 148.055 70.200 148.815 ;
        RECT 70.370 148.225 70.625 149.130 ;
        RECT 70.800 148.055 71.060 149.205 ;
        RECT 71.240 148.055 71.500 149.205 ;
        RECT 71.675 149.130 71.845 149.860 ;
        RECT 72.100 149.695 72.270 149.885 ;
        RECT 73.535 149.835 76.125 150.605 ;
        RECT 72.015 149.365 72.270 149.695 ;
        RECT 72.100 149.155 72.270 149.365 ;
        RECT 72.550 149.335 72.905 149.705 ;
        RECT 71.675 148.225 71.930 149.130 ;
        RECT 72.100 148.985 72.815 149.155 ;
        RECT 72.100 148.055 72.430 148.815 ;
        RECT 72.645 148.225 72.815 148.985 ;
        RECT 73.535 149.145 74.745 149.665 ;
        RECT 74.915 149.315 76.125 149.835 ;
        RECT 76.295 149.805 76.635 150.435 ;
        RECT 76.805 149.805 77.055 150.605 ;
        RECT 77.245 149.955 77.575 150.435 ;
        RECT 77.745 150.145 77.970 150.605 ;
        RECT 78.140 149.955 78.470 150.435 ;
        RECT 76.295 149.195 76.470 149.805 ;
        RECT 77.245 149.785 78.470 149.955 ;
        RECT 79.100 149.825 79.600 150.435 ;
        RECT 79.975 149.855 81.185 150.605 ;
        RECT 81.360 150.060 86.705 150.605 ;
        RECT 76.640 149.445 77.335 149.615 ;
        RECT 77.165 149.195 77.335 149.445 ;
        RECT 77.510 149.415 77.930 149.615 ;
        RECT 78.100 149.415 78.430 149.615 ;
        RECT 78.600 149.415 78.930 149.615 ;
        RECT 79.100 149.195 79.270 149.825 ;
        RECT 79.455 149.365 79.805 149.615 ;
        RECT 73.535 148.055 76.125 149.145 ;
        RECT 76.295 148.225 76.635 149.195 ;
        RECT 76.805 148.055 76.975 149.195 ;
        RECT 77.165 149.025 79.600 149.195 ;
        RECT 77.245 148.055 77.495 148.855 ;
        RECT 78.140 148.225 78.470 149.025 ;
        RECT 78.770 148.055 79.100 148.855 ;
        RECT 79.270 148.225 79.600 149.025 ;
        RECT 79.975 149.145 80.495 149.685 ;
        RECT 80.665 149.315 81.185 149.855 ;
        RECT 79.975 148.055 81.185 149.145 ;
        RECT 82.950 148.490 83.300 149.740 ;
        RECT 84.780 149.230 85.120 150.060 ;
        RECT 86.875 149.880 87.165 150.605 ;
        RECT 87.395 149.785 87.605 150.605 ;
        RECT 87.775 149.805 88.105 150.435 ;
        RECT 81.360 148.055 86.705 148.490 ;
        RECT 86.875 148.055 87.165 149.220 ;
        RECT 87.775 149.205 88.025 149.805 ;
        RECT 88.275 149.785 88.505 150.605 ;
        RECT 89.180 149.895 89.435 150.425 ;
        RECT 89.605 150.145 89.910 150.605 ;
        RECT 90.155 150.225 91.225 150.395 ;
        RECT 88.195 149.365 88.525 149.615 ;
        RECT 89.180 149.245 89.390 149.895 ;
        RECT 90.155 149.870 90.475 150.225 ;
        RECT 90.150 149.695 90.475 149.870 ;
        RECT 89.560 149.395 90.475 149.695 ;
        RECT 90.645 149.655 90.885 150.055 ;
        RECT 91.055 149.995 91.225 150.225 ;
        RECT 91.395 150.165 91.585 150.605 ;
        RECT 91.755 150.155 92.705 150.435 ;
        RECT 92.925 150.245 93.275 150.415 ;
        RECT 91.055 149.825 91.585 149.995 ;
        RECT 89.560 149.365 90.300 149.395 ;
        RECT 87.395 148.055 87.605 149.195 ;
        RECT 87.775 148.225 88.105 149.205 ;
        RECT 88.275 148.055 88.505 149.195 ;
        RECT 89.180 148.365 89.435 149.245 ;
        RECT 89.605 148.055 89.910 149.195 ;
        RECT 90.130 148.775 90.300 149.365 ;
        RECT 90.645 149.285 91.185 149.655 ;
        RECT 91.365 149.545 91.585 149.825 ;
        RECT 91.755 149.375 91.925 150.155 ;
        RECT 91.520 149.205 91.925 149.375 ;
        RECT 92.095 149.365 92.445 149.985 ;
        RECT 91.520 149.115 91.690 149.205 ;
        RECT 92.615 149.195 92.825 149.985 ;
        RECT 90.470 148.945 91.690 149.115 ;
        RECT 92.150 149.035 92.825 149.195 ;
        RECT 90.130 148.605 90.930 148.775 ;
        RECT 90.250 148.055 90.580 148.435 ;
        RECT 90.760 148.315 90.930 148.605 ;
        RECT 91.520 148.565 91.690 148.945 ;
        RECT 91.860 149.025 92.825 149.035 ;
        RECT 93.015 149.855 93.275 150.245 ;
        RECT 93.485 150.145 93.815 150.605 ;
        RECT 94.690 150.215 95.545 150.385 ;
        RECT 95.750 150.215 96.245 150.385 ;
        RECT 96.415 150.245 96.745 150.605 ;
        RECT 93.015 149.165 93.185 149.855 ;
        RECT 93.355 149.505 93.525 149.685 ;
        RECT 93.695 149.675 94.485 149.925 ;
        RECT 94.690 149.505 94.860 150.215 ;
        RECT 95.030 149.705 95.385 149.925 ;
        RECT 93.355 149.335 95.045 149.505 ;
        RECT 91.860 148.735 92.320 149.025 ;
        RECT 93.015 148.995 94.515 149.165 ;
        RECT 93.015 148.855 93.185 148.995 ;
        RECT 92.625 148.685 93.185 148.855 ;
        RECT 91.100 148.055 91.350 148.515 ;
        RECT 91.520 148.225 92.390 148.565 ;
        RECT 92.625 148.225 92.795 148.685 ;
        RECT 93.630 148.655 94.705 148.825 ;
        RECT 92.965 148.055 93.335 148.515 ;
        RECT 93.630 148.315 93.800 148.655 ;
        RECT 93.970 148.055 94.300 148.485 ;
        RECT 94.535 148.315 94.705 148.655 ;
        RECT 94.875 148.555 95.045 149.335 ;
        RECT 95.215 149.115 95.385 149.705 ;
        RECT 95.555 149.305 95.905 149.925 ;
        RECT 95.215 148.725 95.680 149.115 ;
        RECT 96.075 148.855 96.245 150.215 ;
        RECT 96.415 149.025 96.875 150.075 ;
        RECT 95.850 148.685 96.245 148.855 ;
        RECT 95.850 148.555 96.020 148.685 ;
        RECT 94.875 148.225 95.555 148.555 ;
        RECT 95.770 148.225 96.020 148.555 ;
        RECT 96.190 148.055 96.440 148.515 ;
        RECT 96.610 148.240 96.935 149.025 ;
        RECT 97.105 148.225 97.275 150.345 ;
        RECT 97.445 150.225 97.775 150.605 ;
        RECT 97.945 150.055 98.200 150.345 ;
        RECT 99.300 150.060 104.645 150.605 ;
        RECT 97.450 149.885 98.200 150.055 ;
        RECT 97.450 148.895 97.680 149.885 ;
        RECT 97.850 149.065 98.200 149.715 ;
        RECT 97.450 148.725 98.200 148.895 ;
        RECT 97.445 148.055 97.775 148.555 ;
        RECT 97.945 148.225 98.200 148.725 ;
        RECT 100.890 148.490 101.240 149.740 ;
        RECT 102.720 149.230 103.060 150.060 ;
        RECT 104.815 149.930 105.085 150.275 ;
        RECT 105.275 150.205 105.655 150.605 ;
        RECT 105.825 150.035 105.995 150.385 ;
        RECT 106.165 150.205 106.495 150.605 ;
        RECT 106.695 150.035 106.865 150.385 ;
        RECT 107.065 150.105 107.395 150.605 ;
        RECT 104.815 149.195 104.985 149.930 ;
        RECT 105.255 149.865 106.865 150.035 ;
        RECT 105.255 149.695 105.425 149.865 ;
        RECT 105.155 149.365 105.425 149.695 ;
        RECT 105.595 149.365 106.000 149.695 ;
        RECT 105.255 149.195 105.425 149.365 ;
        RECT 99.300 148.055 104.645 148.490 ;
        RECT 104.815 148.225 105.085 149.195 ;
        RECT 105.255 149.025 105.980 149.195 ;
        RECT 106.170 149.075 106.880 149.695 ;
        RECT 107.050 149.365 107.400 149.935 ;
        RECT 107.575 149.855 108.785 150.605 ;
        RECT 105.810 148.905 105.980 149.025 ;
        RECT 107.080 148.905 107.400 149.195 ;
        RECT 105.295 148.055 105.575 148.855 ;
        RECT 105.810 148.735 107.400 148.905 ;
        RECT 107.575 149.145 108.095 149.685 ;
        RECT 108.265 149.315 108.785 149.855 ;
        RECT 108.955 149.835 112.465 150.605 ;
        RECT 112.635 149.880 112.925 150.605 ;
        RECT 113.555 149.835 116.145 150.605 ;
        RECT 108.955 149.145 110.645 149.665 ;
        RECT 110.815 149.315 112.465 149.835 ;
        RECT 105.745 148.275 107.400 148.565 ;
        RECT 107.575 148.055 108.785 149.145 ;
        RECT 108.955 148.055 112.465 149.145 ;
        RECT 112.635 148.055 112.925 149.220 ;
        RECT 113.555 149.145 114.765 149.665 ;
        RECT 114.935 149.315 116.145 149.835 ;
        RECT 116.375 149.785 116.585 150.605 ;
        RECT 116.755 149.805 117.085 150.435 ;
        RECT 116.755 149.205 117.005 149.805 ;
        RECT 117.255 149.785 117.485 150.605 ;
        RECT 117.785 150.055 117.955 150.435 ;
        RECT 118.135 150.225 118.465 150.605 ;
        RECT 117.785 149.885 118.450 150.055 ;
        RECT 118.645 149.930 118.905 150.435 ;
        RECT 119.080 150.060 124.425 150.605 ;
        RECT 117.175 149.365 117.505 149.615 ;
        RECT 117.715 149.335 118.045 149.705 ;
        RECT 118.280 149.630 118.450 149.885 ;
        RECT 118.280 149.300 118.565 149.630 ;
        RECT 113.555 148.055 116.145 149.145 ;
        RECT 116.375 148.055 116.585 149.195 ;
        RECT 116.755 148.225 117.085 149.205 ;
        RECT 117.255 148.055 117.485 149.195 ;
        RECT 118.280 149.155 118.450 149.300 ;
        RECT 117.785 148.985 118.450 149.155 ;
        RECT 118.735 149.130 118.905 149.930 ;
        RECT 117.785 148.225 117.955 148.985 ;
        RECT 118.135 148.055 118.465 148.815 ;
        RECT 118.635 148.225 118.905 149.130 ;
        RECT 120.670 148.490 121.020 149.740 ;
        RECT 122.500 149.230 122.840 150.060 ;
        RECT 124.595 149.855 125.805 150.605 ;
        RECT 124.595 149.145 125.115 149.685 ;
        RECT 125.285 149.315 125.805 149.855 ;
        RECT 119.080 148.055 124.425 148.490 ;
        RECT 124.595 148.055 125.805 149.145 ;
        RECT 11.810 147.885 125.890 148.055 ;
        RECT 11.895 146.795 13.105 147.885 ;
        RECT 11.895 146.085 12.415 146.625 ;
        RECT 12.585 146.255 13.105 146.795 ;
        RECT 13.275 146.795 16.785 147.885 ;
        RECT 16.960 147.450 22.305 147.885 ;
        RECT 13.275 146.275 14.965 146.795 ;
        RECT 15.135 146.105 16.785 146.625 ;
        RECT 18.550 146.200 18.900 147.450 ;
        RECT 22.475 146.720 22.765 147.885 ;
        RECT 23.855 146.795 27.365 147.885 ;
        RECT 27.540 147.450 32.885 147.885 ;
        RECT 33.060 147.450 38.405 147.885 ;
        RECT 11.895 145.335 13.105 146.085 ;
        RECT 13.275 145.335 16.785 146.105 ;
        RECT 20.380 145.880 20.720 146.710 ;
        RECT 23.855 146.275 25.545 146.795 ;
        RECT 25.715 146.105 27.365 146.625 ;
        RECT 29.130 146.200 29.480 147.450 ;
        RECT 16.960 145.335 22.305 145.880 ;
        RECT 22.475 145.335 22.765 146.060 ;
        RECT 23.855 145.335 27.365 146.105 ;
        RECT 30.960 145.880 31.300 146.710 ;
        RECT 34.650 146.200 35.000 147.450 ;
        RECT 38.780 146.915 39.110 147.715 ;
        RECT 39.280 147.085 39.610 147.885 ;
        RECT 39.910 146.915 40.240 147.715 ;
        RECT 40.885 147.085 41.135 147.885 ;
        RECT 38.780 146.745 41.215 146.915 ;
        RECT 41.405 146.745 41.575 147.885 ;
        RECT 41.745 146.745 42.085 147.715 ;
        RECT 42.460 146.915 42.790 147.715 ;
        RECT 42.960 147.085 43.290 147.885 ;
        RECT 43.590 146.915 43.920 147.715 ;
        RECT 44.565 147.085 44.815 147.885 ;
        RECT 42.460 146.745 44.895 146.915 ;
        RECT 45.085 146.745 45.255 147.885 ;
        RECT 45.425 146.745 45.765 147.715 ;
        RECT 36.480 145.880 36.820 146.710 ;
        RECT 38.575 146.325 38.925 146.575 ;
        RECT 39.110 146.115 39.280 146.745 ;
        RECT 39.450 146.325 39.780 146.525 ;
        RECT 39.950 146.325 40.280 146.525 ;
        RECT 40.450 146.325 40.870 146.525 ;
        RECT 41.045 146.495 41.215 146.745 ;
        RECT 41.045 146.325 41.740 146.495 ;
        RECT 27.540 145.335 32.885 145.880 ;
        RECT 33.060 145.335 38.405 145.880 ;
        RECT 38.780 145.505 39.280 146.115 ;
        RECT 39.910 145.985 41.135 146.155 ;
        RECT 41.910 146.135 42.085 146.745 ;
        RECT 42.255 146.325 42.605 146.575 ;
        RECT 39.910 145.505 40.240 145.985 ;
        RECT 40.410 145.335 40.635 145.795 ;
        RECT 40.805 145.505 41.135 145.985 ;
        RECT 41.325 145.335 41.575 146.135 ;
        RECT 41.745 145.505 42.085 146.135 ;
        RECT 42.790 146.115 42.960 146.745 ;
        RECT 43.130 146.325 43.460 146.525 ;
        RECT 43.630 146.325 43.960 146.525 ;
        RECT 44.130 146.325 44.550 146.525 ;
        RECT 44.725 146.495 44.895 146.745 ;
        RECT 44.725 146.325 45.420 146.495 ;
        RECT 42.460 145.505 42.960 146.115 ;
        RECT 43.590 145.985 44.815 146.155 ;
        RECT 45.590 146.135 45.765 146.745 ;
        RECT 46.395 146.795 48.065 147.885 ;
        RECT 46.395 146.275 47.145 146.795 ;
        RECT 48.235 146.720 48.525 147.885 ;
        RECT 48.695 146.795 52.205 147.885 ;
        RECT 43.590 145.505 43.920 145.985 ;
        RECT 44.090 145.335 44.315 145.795 ;
        RECT 44.485 145.505 44.815 145.985 ;
        RECT 45.005 145.335 45.255 146.135 ;
        RECT 45.425 145.505 45.765 146.135 ;
        RECT 47.315 146.105 48.065 146.625 ;
        RECT 48.695 146.275 50.385 146.795 ;
        RECT 52.375 146.745 52.715 147.715 ;
        RECT 52.885 146.745 53.055 147.885 ;
        RECT 53.325 147.085 53.575 147.885 ;
        RECT 54.220 146.915 54.550 147.715 ;
        RECT 54.850 147.085 55.180 147.885 ;
        RECT 55.350 146.915 55.680 147.715 ;
        RECT 53.245 146.745 55.680 146.915 ;
        RECT 56.055 146.745 56.395 147.715 ;
        RECT 56.565 146.745 56.735 147.885 ;
        RECT 57.005 147.085 57.255 147.885 ;
        RECT 57.900 146.915 58.230 147.715 ;
        RECT 58.530 147.085 58.860 147.885 ;
        RECT 59.030 146.915 59.360 147.715 ;
        RECT 59.825 147.140 60.095 147.885 ;
        RECT 60.725 147.880 67.000 147.885 ;
        RECT 60.265 146.970 60.555 147.710 ;
        RECT 60.725 147.155 60.980 147.880 ;
        RECT 61.165 146.985 61.425 147.710 ;
        RECT 61.595 147.155 61.840 147.880 ;
        RECT 62.025 146.985 62.285 147.710 ;
        RECT 62.455 147.155 62.700 147.880 ;
        RECT 62.885 146.985 63.145 147.710 ;
        RECT 63.315 147.155 63.560 147.880 ;
        RECT 63.730 146.985 63.990 147.710 ;
        RECT 64.160 147.155 64.420 147.880 ;
        RECT 64.590 146.985 64.850 147.710 ;
        RECT 65.020 147.155 65.280 147.880 ;
        RECT 65.450 146.985 65.710 147.710 ;
        RECT 65.880 147.155 66.140 147.880 ;
        RECT 66.310 146.985 66.570 147.710 ;
        RECT 66.740 147.085 67.000 147.880 ;
        RECT 61.165 146.970 66.570 146.985 ;
        RECT 56.925 146.745 59.360 146.915 ;
        RECT 59.825 146.745 66.570 146.970 ;
        RECT 50.555 146.105 52.205 146.625 ;
        RECT 46.395 145.335 48.065 146.105 ;
        RECT 48.235 145.335 48.525 146.060 ;
        RECT 48.695 145.335 52.205 146.105 ;
        RECT 52.375 146.135 52.550 146.745 ;
        RECT 53.245 146.495 53.415 146.745 ;
        RECT 52.720 146.325 53.415 146.495 ;
        RECT 53.590 146.325 54.010 146.525 ;
        RECT 54.180 146.325 54.510 146.525 ;
        RECT 54.680 146.325 55.010 146.525 ;
        RECT 52.375 145.505 52.715 146.135 ;
        RECT 52.885 145.335 53.135 146.135 ;
        RECT 53.325 145.985 54.550 146.155 ;
        RECT 53.325 145.505 53.655 145.985 ;
        RECT 53.825 145.335 54.050 145.795 ;
        RECT 54.220 145.505 54.550 145.985 ;
        RECT 55.180 146.115 55.350 146.745 ;
        RECT 55.535 146.325 55.885 146.575 ;
        RECT 56.055 146.135 56.230 146.745 ;
        RECT 56.925 146.495 57.095 146.745 ;
        RECT 56.400 146.325 57.095 146.495 ;
        RECT 57.270 146.325 57.690 146.525 ;
        RECT 57.860 146.325 58.190 146.525 ;
        RECT 58.360 146.325 58.690 146.525 ;
        RECT 55.180 145.505 55.680 146.115 ;
        RECT 56.055 145.505 56.395 146.135 ;
        RECT 56.565 145.335 56.815 146.135 ;
        RECT 57.005 145.985 58.230 146.155 ;
        RECT 57.005 145.505 57.335 145.985 ;
        RECT 57.505 145.335 57.730 145.795 ;
        RECT 57.900 145.505 58.230 145.985 ;
        RECT 58.860 146.115 59.030 146.745 ;
        RECT 59.215 146.325 59.565 146.575 ;
        RECT 59.825 146.155 60.990 146.745 ;
        RECT 67.170 146.575 67.420 147.710 ;
        RECT 67.600 147.075 67.860 147.885 ;
        RECT 68.035 146.575 68.280 147.715 ;
        RECT 68.460 147.075 68.755 147.885 ;
        RECT 68.940 146.735 69.200 147.885 ;
        RECT 69.375 146.810 69.630 147.715 ;
        RECT 69.800 147.125 70.130 147.885 ;
        RECT 70.345 146.955 70.515 147.715 ;
        RECT 61.160 146.325 68.280 146.575 ;
        RECT 58.860 145.505 59.360 146.115 ;
        RECT 59.825 145.985 66.570 146.155 ;
        RECT 59.825 145.335 60.125 145.815 ;
        RECT 60.295 145.530 60.555 145.985 ;
        RECT 60.725 145.335 60.985 145.815 ;
        RECT 61.165 145.530 61.425 145.985 ;
        RECT 61.595 145.335 61.845 145.815 ;
        RECT 62.025 145.530 62.285 145.985 ;
        RECT 62.455 145.335 62.705 145.815 ;
        RECT 62.885 145.530 63.145 145.985 ;
        RECT 63.315 145.335 63.560 145.815 ;
        RECT 63.730 145.530 64.005 145.985 ;
        RECT 64.175 145.335 64.420 145.815 ;
        RECT 64.590 145.530 64.850 145.985 ;
        RECT 65.020 145.335 65.280 145.815 ;
        RECT 65.450 145.530 65.710 145.985 ;
        RECT 65.880 145.335 66.140 145.815 ;
        RECT 66.310 145.530 66.570 145.985 ;
        RECT 66.740 145.335 67.000 145.895 ;
        RECT 67.170 145.515 67.420 146.325 ;
        RECT 67.600 145.335 67.860 145.860 ;
        RECT 68.030 145.515 68.280 146.325 ;
        RECT 68.450 146.015 68.765 146.575 ;
        RECT 68.460 145.335 68.765 145.845 ;
        RECT 68.940 145.335 69.200 146.175 ;
        RECT 69.375 146.080 69.545 146.810 ;
        RECT 69.800 146.785 70.515 146.955 ;
        RECT 71.245 146.825 71.575 147.885 ;
        RECT 69.800 146.575 69.970 146.785 ;
        RECT 69.715 146.245 69.970 146.575 ;
        RECT 69.375 145.505 69.630 146.080 ;
        RECT 69.800 146.055 69.970 146.245 ;
        RECT 70.250 146.235 70.605 146.605 ;
        RECT 71.755 146.575 71.925 147.545 ;
        RECT 72.095 147.295 72.425 147.695 ;
        RECT 72.595 147.525 72.925 147.885 ;
        RECT 73.125 147.295 73.825 147.715 ;
        RECT 72.095 147.065 73.825 147.295 ;
        RECT 72.095 146.845 72.425 147.065 ;
        RECT 72.620 146.575 72.945 146.865 ;
        RECT 71.235 146.245 71.545 146.575 ;
        RECT 71.755 146.245 72.130 146.575 ;
        RECT 72.450 146.245 72.945 146.575 ;
        RECT 73.120 146.325 73.450 146.865 ;
        RECT 73.620 146.095 73.825 147.065 ;
        RECT 73.995 146.720 74.285 147.885 ;
        RECT 74.545 146.955 74.715 147.715 ;
        RECT 74.930 147.125 75.260 147.885 ;
        RECT 74.545 146.785 75.260 146.955 ;
        RECT 75.430 146.810 75.685 147.715 ;
        RECT 74.455 146.235 74.810 146.605 ;
        RECT 75.090 146.575 75.260 146.785 ;
        RECT 75.090 146.245 75.345 146.575 ;
        RECT 69.800 145.885 70.515 146.055 ;
        RECT 69.800 145.335 70.130 145.715 ;
        RECT 70.345 145.505 70.515 145.885 ;
        RECT 71.245 145.865 72.605 146.075 ;
        RECT 71.245 145.505 71.575 145.865 ;
        RECT 71.745 145.335 72.075 145.695 ;
        RECT 72.275 145.505 72.605 145.865 ;
        RECT 73.115 145.505 73.825 146.095 ;
        RECT 73.995 145.335 74.285 146.060 ;
        RECT 75.090 146.055 75.260 146.245 ;
        RECT 75.515 146.080 75.685 146.810 ;
        RECT 75.860 146.735 76.120 147.885 ;
        RECT 76.385 146.955 76.555 147.715 ;
        RECT 76.770 147.125 77.100 147.885 ;
        RECT 76.385 146.785 77.100 146.955 ;
        RECT 77.270 146.810 77.525 147.715 ;
        RECT 76.295 146.235 76.650 146.605 ;
        RECT 76.930 146.575 77.100 146.785 ;
        RECT 76.930 146.245 77.185 146.575 ;
        RECT 74.545 145.885 75.260 146.055 ;
        RECT 74.545 145.505 74.715 145.885 ;
        RECT 74.930 145.335 75.260 145.715 ;
        RECT 75.430 145.505 75.685 146.080 ;
        RECT 75.860 145.335 76.120 146.175 ;
        RECT 76.930 146.055 77.100 146.245 ;
        RECT 77.355 146.080 77.525 146.810 ;
        RECT 77.700 146.735 77.960 147.885 ;
        RECT 79.055 146.795 82.565 147.885 ;
        RECT 83.110 146.905 83.365 147.575 ;
        RECT 83.545 147.085 83.830 147.885 ;
        RECT 84.010 147.165 84.340 147.675 ;
        RECT 79.055 146.275 80.745 146.795 ;
        RECT 76.385 145.885 77.100 146.055 ;
        RECT 76.385 145.505 76.555 145.885 ;
        RECT 76.770 145.335 77.100 145.715 ;
        RECT 77.270 145.505 77.525 146.080 ;
        RECT 77.700 145.335 77.960 146.175 ;
        RECT 80.915 146.105 82.565 146.625 ;
        RECT 79.055 145.335 82.565 146.105 ;
        RECT 83.110 146.045 83.290 146.905 ;
        RECT 84.010 146.575 84.260 147.165 ;
        RECT 84.610 147.015 84.780 147.625 ;
        RECT 84.950 147.195 85.280 147.885 ;
        RECT 85.510 147.335 85.750 147.625 ;
        RECT 85.950 147.505 86.370 147.885 ;
        RECT 86.550 147.415 87.180 147.665 ;
        RECT 87.650 147.505 87.980 147.885 ;
        RECT 86.550 147.335 86.720 147.415 ;
        RECT 88.150 147.335 88.320 147.625 ;
        RECT 88.500 147.505 88.880 147.885 ;
        RECT 89.120 147.500 89.950 147.670 ;
        RECT 85.510 147.165 86.720 147.335 ;
        RECT 83.460 146.245 84.260 146.575 ;
        RECT 83.110 145.845 83.365 146.045 ;
        RECT 83.025 145.675 83.365 145.845 ;
        RECT 83.110 145.515 83.365 145.675 ;
        RECT 83.545 145.335 83.830 145.795 ;
        RECT 84.010 145.595 84.260 146.245 ;
        RECT 84.460 146.995 84.780 147.015 ;
        RECT 84.460 146.825 86.380 146.995 ;
        RECT 84.460 145.930 84.650 146.825 ;
        RECT 86.550 146.655 86.720 147.165 ;
        RECT 86.890 146.905 87.410 147.215 ;
        RECT 84.820 146.485 86.720 146.655 ;
        RECT 84.820 146.425 85.150 146.485 ;
        RECT 85.300 146.255 85.630 146.315 ;
        RECT 84.970 145.985 85.630 146.255 ;
        RECT 84.460 145.600 84.780 145.930 ;
        RECT 84.960 145.335 85.620 145.815 ;
        RECT 85.820 145.725 85.990 146.485 ;
        RECT 86.890 146.315 87.070 146.725 ;
        RECT 86.160 146.145 86.490 146.265 ;
        RECT 87.240 146.145 87.410 146.905 ;
        RECT 86.160 145.975 87.410 146.145 ;
        RECT 87.580 147.085 88.950 147.335 ;
        RECT 87.580 146.315 87.770 147.085 ;
        RECT 88.700 146.825 88.950 147.085 ;
        RECT 87.940 146.655 88.190 146.815 ;
        RECT 89.120 146.655 89.290 147.500 ;
        RECT 90.185 147.215 90.355 147.715 ;
        RECT 90.525 147.385 90.855 147.885 ;
        RECT 89.460 146.825 89.960 147.205 ;
        RECT 90.185 147.045 90.880 147.215 ;
        RECT 87.940 146.485 89.290 146.655 ;
        RECT 88.870 146.445 89.290 146.485 ;
        RECT 87.580 145.975 88.000 146.315 ;
        RECT 88.290 145.985 88.700 146.315 ;
        RECT 85.820 145.555 86.670 145.725 ;
        RECT 87.230 145.335 87.550 145.795 ;
        RECT 87.750 145.545 88.000 145.975 ;
        RECT 88.290 145.335 88.700 145.775 ;
        RECT 88.870 145.715 89.040 146.445 ;
        RECT 89.210 145.895 89.560 146.265 ;
        RECT 89.740 145.955 89.960 146.825 ;
        RECT 90.130 146.255 90.540 146.875 ;
        RECT 90.710 146.075 90.880 147.045 ;
        RECT 90.185 145.885 90.880 146.075 ;
        RECT 88.870 145.515 89.885 145.715 ;
        RECT 90.185 145.555 90.355 145.885 ;
        RECT 90.525 145.335 90.855 145.715 ;
        RECT 91.070 145.595 91.295 147.715 ;
        RECT 91.465 147.385 91.795 147.885 ;
        RECT 91.965 147.215 92.135 147.715 ;
        RECT 91.470 147.045 92.135 147.215 ;
        RECT 91.470 146.055 91.700 147.045 ;
        RECT 91.870 146.225 92.220 146.875 ;
        RECT 92.455 146.745 92.665 147.885 ;
        RECT 92.835 146.735 93.165 147.715 ;
        RECT 93.335 146.745 93.565 147.885 ;
        RECT 94.325 146.955 94.495 147.715 ;
        RECT 94.675 147.125 95.005 147.885 ;
        RECT 94.325 146.785 94.990 146.955 ;
        RECT 95.175 146.810 95.445 147.715 ;
        RECT 91.470 145.885 92.135 146.055 ;
        RECT 91.465 145.335 91.795 145.715 ;
        RECT 91.965 145.595 92.135 145.885 ;
        RECT 92.455 145.335 92.665 146.155 ;
        RECT 92.835 146.135 93.085 146.735 ;
        RECT 94.820 146.640 94.990 146.785 ;
        RECT 93.255 146.325 93.585 146.575 ;
        RECT 94.255 146.235 94.585 146.605 ;
        RECT 94.820 146.310 95.105 146.640 ;
        RECT 92.835 145.505 93.165 146.135 ;
        RECT 93.335 145.335 93.565 146.155 ;
        RECT 94.820 146.055 94.990 146.310 ;
        RECT 94.325 145.885 94.990 146.055 ;
        RECT 95.275 146.010 95.445 146.810 ;
        RECT 95.615 146.795 96.825 147.885 ;
        RECT 97.000 147.375 98.655 147.665 ;
        RECT 97.000 147.035 98.590 147.205 ;
        RECT 98.825 147.085 99.105 147.885 ;
        RECT 95.615 146.255 96.135 146.795 ;
        RECT 97.000 146.745 97.320 147.035 ;
        RECT 98.420 146.915 98.590 147.035 ;
        RECT 97.515 146.695 98.230 146.865 ;
        RECT 98.420 146.745 99.145 146.915 ;
        RECT 99.315 146.745 99.585 147.715 ;
        RECT 96.305 146.085 96.825 146.625 ;
        RECT 94.325 145.505 94.495 145.885 ;
        RECT 94.675 145.335 95.005 145.715 ;
        RECT 95.185 145.505 95.445 146.010 ;
        RECT 95.615 145.335 96.825 146.085 ;
        RECT 97.000 146.005 97.350 146.575 ;
        RECT 97.520 146.245 98.230 146.695 ;
        RECT 98.975 146.575 99.145 146.745 ;
        RECT 98.400 146.245 98.805 146.575 ;
        RECT 98.975 146.245 99.245 146.575 ;
        RECT 98.975 146.075 99.145 146.245 ;
        RECT 97.535 145.905 99.145 146.075 ;
        RECT 99.415 146.010 99.585 146.745 ;
        RECT 99.755 146.720 100.045 147.885 ;
        RECT 100.675 146.795 102.345 147.885 ;
        RECT 100.675 146.275 101.425 146.795 ;
        RECT 102.515 146.745 102.855 147.715 ;
        RECT 103.025 146.745 103.195 147.885 ;
        RECT 103.465 147.085 103.715 147.885 ;
        RECT 104.360 146.915 104.690 147.715 ;
        RECT 104.990 147.085 105.320 147.885 ;
        RECT 105.490 146.915 105.820 147.715 ;
        RECT 103.385 146.745 105.820 146.915 ;
        RECT 106.655 146.745 106.995 147.715 ;
        RECT 107.165 146.745 107.335 147.885 ;
        RECT 107.605 147.085 107.855 147.885 ;
        RECT 108.500 146.915 108.830 147.715 ;
        RECT 109.130 147.085 109.460 147.885 ;
        RECT 109.630 146.915 109.960 147.715 ;
        RECT 107.525 146.745 109.960 146.915 ;
        RECT 111.255 147.125 111.770 147.535 ;
        RECT 112.005 147.125 112.175 147.885 ;
        RECT 112.345 147.545 114.375 147.715 ;
        RECT 101.595 146.105 102.345 146.625 ;
        RECT 97.005 145.335 97.335 145.835 ;
        RECT 97.535 145.555 97.705 145.905 ;
        RECT 97.905 145.335 98.235 145.735 ;
        RECT 98.405 145.555 98.575 145.905 ;
        RECT 98.745 145.335 99.125 145.735 ;
        RECT 99.315 145.665 99.585 146.010 ;
        RECT 99.755 145.335 100.045 146.060 ;
        RECT 100.675 145.335 102.345 146.105 ;
        RECT 102.515 146.185 102.690 146.745 ;
        RECT 103.385 146.495 103.555 146.745 ;
        RECT 102.860 146.325 103.555 146.495 ;
        RECT 103.730 146.325 104.150 146.525 ;
        RECT 104.320 146.325 104.650 146.525 ;
        RECT 104.820 146.325 105.150 146.525 ;
        RECT 102.515 146.135 102.745 146.185 ;
        RECT 102.515 145.505 102.855 146.135 ;
        RECT 103.025 145.335 103.275 146.135 ;
        RECT 103.465 145.985 104.690 146.155 ;
        RECT 103.465 145.505 103.795 145.985 ;
        RECT 103.965 145.335 104.190 145.795 ;
        RECT 104.360 145.505 104.690 145.985 ;
        RECT 105.320 146.115 105.490 146.745 ;
        RECT 105.675 146.325 106.025 146.575 ;
        RECT 106.655 146.135 106.830 146.745 ;
        RECT 107.525 146.495 107.695 146.745 ;
        RECT 107.000 146.325 107.695 146.495 ;
        RECT 107.870 146.325 108.290 146.525 ;
        RECT 108.460 146.325 108.790 146.525 ;
        RECT 108.960 146.325 109.290 146.525 ;
        RECT 105.320 145.505 105.820 146.115 ;
        RECT 106.655 145.505 106.995 146.135 ;
        RECT 107.165 145.335 107.415 146.135 ;
        RECT 107.605 145.985 108.830 146.155 ;
        RECT 107.605 145.505 107.935 145.985 ;
        RECT 108.105 145.335 108.330 145.795 ;
        RECT 108.500 145.505 108.830 145.985 ;
        RECT 109.460 146.115 109.630 146.745 ;
        RECT 109.815 146.325 110.165 146.575 ;
        RECT 111.255 146.315 111.595 147.125 ;
        RECT 112.345 146.880 112.515 147.545 ;
        RECT 112.910 147.205 114.035 147.375 ;
        RECT 111.765 146.690 112.515 146.880 ;
        RECT 112.685 146.865 113.695 147.035 ;
        RECT 111.255 146.145 112.485 146.315 ;
        RECT 109.460 145.505 109.960 146.115 ;
        RECT 111.530 145.540 111.775 146.145 ;
        RECT 111.995 145.335 112.505 145.870 ;
        RECT 112.685 145.505 112.875 146.865 ;
        RECT 113.045 145.845 113.320 146.665 ;
        RECT 113.525 146.065 113.695 146.865 ;
        RECT 113.865 146.075 114.035 147.205 ;
        RECT 114.205 146.575 114.375 147.545 ;
        RECT 114.545 146.745 114.715 147.885 ;
        RECT 114.885 146.745 115.220 147.715 ;
        RECT 114.205 146.245 114.400 146.575 ;
        RECT 114.625 146.245 114.880 146.575 ;
        RECT 114.625 146.075 114.795 146.245 ;
        RECT 115.050 146.075 115.220 146.745 ;
        RECT 115.855 146.795 117.525 147.885 ;
        RECT 115.855 146.275 116.605 146.795 ;
        RECT 117.735 146.745 117.965 147.885 ;
        RECT 118.135 146.735 118.465 147.715 ;
        RECT 118.635 146.745 118.845 147.885 ;
        RECT 119.625 146.955 119.795 147.715 ;
        RECT 119.975 147.125 120.305 147.885 ;
        RECT 119.625 146.785 120.290 146.955 ;
        RECT 120.475 146.810 120.745 147.715 ;
        RECT 116.775 146.105 117.525 146.625 ;
        RECT 117.715 146.325 118.045 146.575 ;
        RECT 113.865 145.905 114.795 146.075 ;
        RECT 113.865 145.870 114.040 145.905 ;
        RECT 113.045 145.675 113.325 145.845 ;
        RECT 113.045 145.505 113.320 145.675 ;
        RECT 113.510 145.505 114.040 145.870 ;
        RECT 114.465 145.335 114.795 145.735 ;
        RECT 114.965 145.505 115.220 146.075 ;
        RECT 115.855 145.335 117.525 146.105 ;
        RECT 117.735 145.335 117.965 146.155 ;
        RECT 118.215 146.135 118.465 146.735 ;
        RECT 120.120 146.640 120.290 146.785 ;
        RECT 119.555 146.235 119.885 146.605 ;
        RECT 120.120 146.310 120.405 146.640 ;
        RECT 118.135 145.505 118.465 146.135 ;
        RECT 118.635 145.335 118.845 146.155 ;
        RECT 120.120 146.055 120.290 146.310 ;
        RECT 119.625 145.885 120.290 146.055 ;
        RECT 120.575 146.010 120.745 146.810 ;
        RECT 120.915 146.795 124.425 147.885 ;
        RECT 124.595 146.795 125.805 147.885 ;
        RECT 120.915 146.275 122.605 146.795 ;
        RECT 122.775 146.105 124.425 146.625 ;
        RECT 124.595 146.255 125.115 146.795 ;
        RECT 119.625 145.505 119.795 145.885 ;
        RECT 119.975 145.335 120.305 145.715 ;
        RECT 120.485 145.505 120.745 146.010 ;
        RECT 120.915 145.335 124.425 146.105 ;
        RECT 125.285 146.085 125.805 146.625 ;
        RECT 124.595 145.335 125.805 146.085 ;
        RECT 11.810 145.165 125.890 145.335 ;
        RECT 11.895 144.415 13.105 145.165 ;
        RECT 14.110 144.455 14.365 144.985 ;
        RECT 14.545 144.705 14.830 145.165 ;
        RECT 11.895 143.875 12.415 144.415 ;
        RECT 12.585 143.705 13.105 144.245 ;
        RECT 11.895 142.615 13.105 143.705 ;
        RECT 14.110 143.595 14.290 144.455 ;
        RECT 15.010 144.255 15.260 144.905 ;
        RECT 14.460 143.925 15.260 144.255 ;
        RECT 14.110 143.125 14.365 143.595 ;
        RECT 14.025 142.955 14.365 143.125 ;
        RECT 14.110 142.925 14.365 142.955 ;
        RECT 14.545 142.615 14.830 143.415 ;
        RECT 15.010 143.335 15.260 143.925 ;
        RECT 15.460 144.570 15.780 144.900 ;
        RECT 15.960 144.685 16.620 145.165 ;
        RECT 16.820 144.775 17.670 144.945 ;
        RECT 15.460 143.675 15.650 144.570 ;
        RECT 15.970 144.245 16.630 144.515 ;
        RECT 16.300 144.185 16.630 144.245 ;
        RECT 15.820 144.015 16.150 144.075 ;
        RECT 16.820 144.015 16.990 144.775 ;
        RECT 18.230 144.705 18.550 145.165 ;
        RECT 18.750 144.525 19.000 144.955 ;
        RECT 19.290 144.725 19.700 145.165 ;
        RECT 19.870 144.785 20.885 144.985 ;
        RECT 17.160 144.355 18.410 144.525 ;
        RECT 17.160 144.235 17.490 144.355 ;
        RECT 15.820 143.845 17.720 144.015 ;
        RECT 15.460 143.505 17.380 143.675 ;
        RECT 15.460 143.485 15.780 143.505 ;
        RECT 15.010 142.825 15.340 143.335 ;
        RECT 15.610 142.875 15.780 143.485 ;
        RECT 17.550 143.335 17.720 143.845 ;
        RECT 17.890 143.775 18.070 144.185 ;
        RECT 18.240 143.595 18.410 144.355 ;
        RECT 15.950 142.615 16.280 143.305 ;
        RECT 16.510 143.165 17.720 143.335 ;
        RECT 17.890 143.285 18.410 143.595 ;
        RECT 18.580 144.185 19.000 144.525 ;
        RECT 19.290 144.185 19.700 144.515 ;
        RECT 18.580 143.415 18.770 144.185 ;
        RECT 19.870 144.055 20.040 144.785 ;
        RECT 21.185 144.615 21.355 144.945 ;
        RECT 21.525 144.785 21.855 145.165 ;
        RECT 20.210 144.235 20.560 144.605 ;
        RECT 19.870 144.015 20.290 144.055 ;
        RECT 18.940 143.845 20.290 144.015 ;
        RECT 18.940 143.685 19.190 143.845 ;
        RECT 19.700 143.415 19.950 143.675 ;
        RECT 18.580 143.165 19.950 143.415 ;
        RECT 16.510 142.875 16.750 143.165 ;
        RECT 17.550 143.085 17.720 143.165 ;
        RECT 16.950 142.615 17.370 142.995 ;
        RECT 17.550 142.835 18.180 143.085 ;
        RECT 18.650 142.615 18.980 142.995 ;
        RECT 19.150 142.875 19.320 143.165 ;
        RECT 20.120 143.000 20.290 143.845 ;
        RECT 20.740 143.675 20.960 144.545 ;
        RECT 21.185 144.425 21.880 144.615 ;
        RECT 20.460 143.295 20.960 143.675 ;
        RECT 21.130 143.625 21.540 144.245 ;
        RECT 21.710 143.455 21.880 144.425 ;
        RECT 21.185 143.285 21.880 143.455 ;
        RECT 19.500 142.615 19.880 142.995 ;
        RECT 20.120 142.830 20.950 143.000 ;
        RECT 21.185 142.785 21.355 143.285 ;
        RECT 21.525 142.615 21.855 143.115 ;
        RECT 22.070 142.785 22.295 144.905 ;
        RECT 22.465 144.785 22.795 145.165 ;
        RECT 22.965 144.615 23.135 144.905 ;
        RECT 24.320 144.620 29.665 145.165 ;
        RECT 29.840 144.620 35.185 145.165 ;
        RECT 22.470 144.445 23.135 144.615 ;
        RECT 22.470 143.455 22.700 144.445 ;
        RECT 22.870 143.625 23.220 144.275 ;
        RECT 22.470 143.285 23.135 143.455 ;
        RECT 22.465 142.615 22.795 143.115 ;
        RECT 22.965 142.785 23.135 143.285 ;
        RECT 25.910 143.050 26.260 144.300 ;
        RECT 27.740 143.790 28.080 144.620 ;
        RECT 31.430 143.050 31.780 144.300 ;
        RECT 33.260 143.790 33.600 144.620 ;
        RECT 35.355 144.440 35.645 145.165 ;
        RECT 36.735 144.490 37.005 144.835 ;
        RECT 37.195 144.765 37.575 145.165 ;
        RECT 37.745 144.595 37.915 144.945 ;
        RECT 38.085 144.765 38.415 145.165 ;
        RECT 38.615 144.595 38.785 144.945 ;
        RECT 38.985 144.665 39.315 145.165 ;
        RECT 24.320 142.615 29.665 143.050 ;
        RECT 29.840 142.615 35.185 143.050 ;
        RECT 35.355 142.615 35.645 143.780 ;
        RECT 36.735 143.755 36.905 144.490 ;
        RECT 37.175 144.425 38.785 144.595 ;
        RECT 37.175 144.255 37.345 144.425 ;
        RECT 37.075 143.925 37.345 144.255 ;
        RECT 37.515 143.925 37.920 144.255 ;
        RECT 37.175 143.755 37.345 143.925 ;
        RECT 36.735 142.785 37.005 143.755 ;
        RECT 37.175 143.585 37.900 143.755 ;
        RECT 38.090 143.635 38.800 144.255 ;
        RECT 38.970 143.925 39.320 144.495 ;
        RECT 39.955 144.490 40.225 144.835 ;
        RECT 40.415 144.765 40.795 145.165 ;
        RECT 40.965 144.595 41.135 144.945 ;
        RECT 41.305 144.765 41.635 145.165 ;
        RECT 41.835 144.595 42.005 144.945 ;
        RECT 42.205 144.665 42.535 145.165 ;
        RECT 39.955 143.755 40.125 144.490 ;
        RECT 40.395 144.425 42.005 144.595 ;
        RECT 40.395 144.255 40.565 144.425 ;
        RECT 40.295 143.925 40.565 144.255 ;
        RECT 40.735 143.925 41.140 144.255 ;
        RECT 40.395 143.755 40.565 143.925 ;
        RECT 41.310 143.805 42.020 144.255 ;
        RECT 42.190 143.925 42.540 144.495 ;
        RECT 42.715 144.365 43.055 144.995 ;
        RECT 43.225 144.365 43.475 145.165 ;
        RECT 43.665 144.515 43.995 144.995 ;
        RECT 44.165 144.705 44.390 145.165 ;
        RECT 44.560 144.515 44.890 144.995 ;
        RECT 42.715 144.315 42.945 144.365 ;
        RECT 43.665 144.345 44.890 144.515 ;
        RECT 45.520 144.385 46.020 144.995 ;
        RECT 46.400 144.620 51.745 145.165 ;
        RECT 37.730 143.465 37.900 143.585 ;
        RECT 39.000 143.465 39.320 143.755 ;
        RECT 37.215 142.615 37.495 143.415 ;
        RECT 37.730 143.295 39.320 143.465 ;
        RECT 37.665 142.835 39.320 143.125 ;
        RECT 39.955 142.785 40.225 143.755 ;
        RECT 40.395 143.585 41.120 143.755 ;
        RECT 41.310 143.635 42.025 143.805 ;
        RECT 42.715 143.755 42.890 144.315 ;
        RECT 43.060 144.005 43.755 144.175 ;
        RECT 43.930 144.145 44.350 144.175 ;
        RECT 43.585 143.755 43.755 144.005 ;
        RECT 43.925 143.975 44.350 144.145 ;
        RECT 44.520 143.975 44.850 144.175 ;
        RECT 45.020 143.975 45.350 144.175 ;
        RECT 45.520 143.755 45.690 144.385 ;
        RECT 45.875 143.925 46.225 144.175 ;
        RECT 40.950 143.465 41.120 143.585 ;
        RECT 42.220 143.465 42.540 143.755 ;
        RECT 40.435 142.615 40.715 143.415 ;
        RECT 40.950 143.295 42.540 143.465 ;
        RECT 40.885 142.835 42.540 143.125 ;
        RECT 42.715 142.785 43.055 143.755 ;
        RECT 43.225 142.615 43.395 143.755 ;
        RECT 43.585 143.585 46.020 143.755 ;
        RECT 43.665 142.615 43.915 143.415 ;
        RECT 44.560 142.785 44.890 143.585 ;
        RECT 45.190 142.615 45.520 143.415 ;
        RECT 45.690 142.785 46.020 143.585 ;
        RECT 47.990 143.050 48.340 144.300 ;
        RECT 49.820 143.790 50.160 144.620 ;
        RECT 52.005 144.615 52.175 144.995 ;
        RECT 52.355 144.785 52.685 145.165 ;
        RECT 52.005 144.445 52.670 144.615 ;
        RECT 52.865 144.490 53.125 144.995 ;
        RECT 51.935 143.895 52.265 144.265 ;
        RECT 52.500 144.190 52.670 144.445 ;
        RECT 52.500 143.860 52.785 144.190 ;
        RECT 52.500 143.715 52.670 143.860 ;
        RECT 52.005 143.545 52.670 143.715 ;
        RECT 52.955 143.690 53.125 144.490 ;
        RECT 46.400 142.615 51.745 143.050 ;
        RECT 52.005 142.785 52.175 143.545 ;
        RECT 52.355 142.615 52.685 143.375 ;
        RECT 52.855 142.785 53.125 143.690 ;
        RECT 53.295 144.365 53.635 144.995 ;
        RECT 53.805 144.365 54.055 145.165 ;
        RECT 54.245 144.515 54.575 144.995 ;
        RECT 54.745 144.705 54.970 145.165 ;
        RECT 55.140 144.515 55.470 144.995 ;
        RECT 53.295 143.755 53.470 144.365 ;
        RECT 54.245 144.345 55.470 144.515 ;
        RECT 56.100 144.385 56.600 144.995 ;
        RECT 53.640 144.005 54.335 144.175 ;
        RECT 54.165 143.755 54.335 144.005 ;
        RECT 54.510 143.975 54.930 144.175 ;
        RECT 55.100 143.975 55.430 144.175 ;
        RECT 55.600 143.975 55.930 144.175 ;
        RECT 56.100 143.755 56.270 144.385 ;
        RECT 57.250 144.355 57.495 144.960 ;
        RECT 57.715 144.630 58.225 145.165 ;
        RECT 56.975 144.185 58.205 144.355 ;
        RECT 56.455 143.925 56.805 144.175 ;
        RECT 53.295 142.785 53.635 143.755 ;
        RECT 53.805 142.615 53.975 143.755 ;
        RECT 54.165 143.585 56.600 143.755 ;
        RECT 54.245 142.615 54.495 143.415 ;
        RECT 55.140 142.785 55.470 143.585 ;
        RECT 55.770 142.615 56.100 143.415 ;
        RECT 56.270 142.785 56.600 143.585 ;
        RECT 56.975 143.375 57.315 144.185 ;
        RECT 57.485 143.620 58.235 143.810 ;
        RECT 56.975 142.965 57.490 143.375 ;
        RECT 57.725 142.615 57.895 143.375 ;
        RECT 58.065 142.955 58.235 143.620 ;
        RECT 58.405 143.635 58.595 144.995 ;
        RECT 58.765 144.145 59.040 144.995 ;
        RECT 59.230 144.630 59.760 144.995 ;
        RECT 60.185 144.765 60.515 145.165 ;
        RECT 59.585 144.595 59.760 144.630 ;
        RECT 58.765 143.975 59.045 144.145 ;
        RECT 58.765 143.835 59.040 143.975 ;
        RECT 59.245 143.635 59.415 144.435 ;
        RECT 58.405 143.465 59.415 143.635 ;
        RECT 59.585 144.425 60.515 144.595 ;
        RECT 60.685 144.425 60.940 144.995 ;
        RECT 61.115 144.440 61.405 145.165 ;
        RECT 61.950 144.485 62.205 144.985 ;
        RECT 62.385 144.705 62.670 145.165 ;
        RECT 61.865 144.455 62.205 144.485 ;
        RECT 59.585 143.295 59.755 144.425 ;
        RECT 60.345 144.255 60.515 144.425 ;
        RECT 58.630 143.125 59.755 143.295 ;
        RECT 59.925 143.925 60.120 144.255 ;
        RECT 60.345 143.925 60.600 144.255 ;
        RECT 59.925 142.955 60.095 143.925 ;
        RECT 60.770 143.755 60.940 144.425 ;
        RECT 61.865 144.315 62.130 144.455 ;
        RECT 58.065 142.785 60.095 142.955 ;
        RECT 60.265 142.615 60.435 143.755 ;
        RECT 60.605 142.785 60.940 143.755 ;
        RECT 61.115 142.615 61.405 143.780 ;
        RECT 61.950 143.595 62.130 144.315 ;
        RECT 62.850 144.255 63.100 144.905 ;
        RECT 62.300 143.925 63.100 144.255 ;
        RECT 61.950 142.925 62.205 143.595 ;
        RECT 62.385 142.615 62.670 143.415 ;
        RECT 62.850 143.335 63.100 143.925 ;
        RECT 63.300 144.570 63.620 144.900 ;
        RECT 63.800 144.685 64.460 145.165 ;
        RECT 64.660 144.775 65.510 144.945 ;
        RECT 63.300 143.675 63.490 144.570 ;
        RECT 63.810 144.245 64.470 144.515 ;
        RECT 64.140 144.185 64.470 144.245 ;
        RECT 63.660 144.015 63.990 144.075 ;
        RECT 64.660 144.015 64.830 144.775 ;
        RECT 66.070 144.705 66.390 145.165 ;
        RECT 66.590 144.525 66.840 144.955 ;
        RECT 67.130 144.725 67.540 145.165 ;
        RECT 67.710 144.785 68.725 144.985 ;
        RECT 65.000 144.355 66.250 144.525 ;
        RECT 65.000 144.235 65.330 144.355 ;
        RECT 63.660 143.845 65.560 144.015 ;
        RECT 63.300 143.505 65.220 143.675 ;
        RECT 63.300 143.485 63.620 143.505 ;
        RECT 62.850 142.825 63.180 143.335 ;
        RECT 63.450 142.875 63.620 143.485 ;
        RECT 65.390 143.335 65.560 143.845 ;
        RECT 65.730 143.775 65.910 144.185 ;
        RECT 66.080 143.595 66.250 144.355 ;
        RECT 63.790 142.615 64.120 143.305 ;
        RECT 64.350 143.165 65.560 143.335 ;
        RECT 65.730 143.285 66.250 143.595 ;
        RECT 66.420 144.185 66.840 144.525 ;
        RECT 67.130 144.185 67.540 144.515 ;
        RECT 66.420 143.415 66.610 144.185 ;
        RECT 67.710 144.055 67.880 144.785 ;
        RECT 69.025 144.615 69.195 144.945 ;
        RECT 69.365 144.785 69.695 145.165 ;
        RECT 68.050 144.235 68.400 144.605 ;
        RECT 67.710 144.015 68.130 144.055 ;
        RECT 66.780 143.845 68.130 144.015 ;
        RECT 66.780 143.685 67.030 143.845 ;
        RECT 67.540 143.415 67.790 143.675 ;
        RECT 66.420 143.165 67.790 143.415 ;
        RECT 64.350 142.875 64.590 143.165 ;
        RECT 65.390 143.085 65.560 143.165 ;
        RECT 64.790 142.615 65.210 142.995 ;
        RECT 65.390 142.835 66.020 143.085 ;
        RECT 66.490 142.615 66.820 142.995 ;
        RECT 66.990 142.875 67.160 143.165 ;
        RECT 67.960 143.000 68.130 143.845 ;
        RECT 68.580 143.675 68.800 144.545 ;
        RECT 69.025 144.425 69.720 144.615 ;
        RECT 68.300 143.295 68.800 143.675 ;
        RECT 68.970 143.625 69.380 144.245 ;
        RECT 69.550 143.455 69.720 144.425 ;
        RECT 69.025 143.285 69.720 143.455 ;
        RECT 67.340 142.615 67.720 142.995 ;
        RECT 67.960 142.830 68.790 143.000 ;
        RECT 69.025 142.785 69.195 143.285 ;
        RECT 69.365 142.615 69.695 143.115 ;
        RECT 69.910 142.785 70.135 144.905 ;
        RECT 70.305 144.785 70.635 145.165 ;
        RECT 70.805 144.615 70.975 144.905 ;
        RECT 71.295 144.685 71.575 145.165 ;
        RECT 70.310 144.445 70.975 144.615 ;
        RECT 71.745 144.515 72.005 144.905 ;
        RECT 72.180 144.685 72.435 145.165 ;
        RECT 72.605 144.515 72.900 144.905 ;
        RECT 73.080 144.685 73.355 145.165 ;
        RECT 73.525 144.665 73.825 144.995 ;
        RECT 70.310 143.455 70.540 144.445 ;
        RECT 71.250 144.345 72.900 144.515 ;
        RECT 70.710 143.625 71.060 144.275 ;
        RECT 71.250 143.835 71.655 144.345 ;
        RECT 71.825 144.005 72.965 144.175 ;
        RECT 71.250 143.665 72.005 143.835 ;
        RECT 70.310 143.285 70.975 143.455 ;
        RECT 70.305 142.615 70.635 143.115 ;
        RECT 70.805 142.785 70.975 143.285 ;
        RECT 71.290 142.615 71.575 143.485 ;
        RECT 71.745 143.415 72.005 143.665 ;
        RECT 72.795 143.755 72.965 144.005 ;
        RECT 73.135 143.925 73.485 144.495 ;
        RECT 73.655 143.755 73.825 144.665 ;
        RECT 74.085 144.615 74.255 144.995 ;
        RECT 74.470 144.785 74.800 145.165 ;
        RECT 74.085 144.445 74.800 144.615 ;
        RECT 73.995 143.895 74.350 144.265 ;
        RECT 74.630 144.255 74.800 144.445 ;
        RECT 74.970 144.420 75.225 144.995 ;
        RECT 74.630 143.925 74.885 144.255 ;
        RECT 72.795 143.585 73.825 143.755 ;
        RECT 74.630 143.715 74.800 143.925 ;
        RECT 71.745 143.245 72.865 143.415 ;
        RECT 71.745 142.785 72.005 143.245 ;
        RECT 72.180 142.615 72.435 143.075 ;
        RECT 72.605 142.785 72.865 143.245 ;
        RECT 73.035 142.615 73.345 143.415 ;
        RECT 73.515 142.785 73.825 143.585 ;
        RECT 74.085 143.545 74.800 143.715 ;
        RECT 75.055 143.690 75.225 144.420 ;
        RECT 75.400 144.325 75.660 145.165 ;
        RECT 76.295 144.665 76.595 144.995 ;
        RECT 76.765 144.685 77.040 145.165 ;
        RECT 74.085 142.785 74.255 143.545 ;
        RECT 74.470 142.615 74.800 143.375 ;
        RECT 74.970 142.785 75.225 143.690 ;
        RECT 75.400 142.615 75.660 143.765 ;
        RECT 76.295 143.755 76.465 144.665 ;
        RECT 77.220 144.515 77.515 144.905 ;
        RECT 77.685 144.685 77.940 145.165 ;
        RECT 78.115 144.515 78.375 144.905 ;
        RECT 78.545 144.685 78.825 145.165 ;
        RECT 76.635 143.925 76.985 144.495 ;
        RECT 77.220 144.345 78.870 144.515 ;
        RECT 79.055 144.395 82.565 145.165 ;
        RECT 77.155 144.005 78.295 144.175 ;
        RECT 77.155 143.755 77.325 144.005 ;
        RECT 78.465 143.835 78.870 144.345 ;
        RECT 76.295 143.585 77.325 143.755 ;
        RECT 78.115 143.665 78.870 143.835 ;
        RECT 79.055 143.705 80.745 144.225 ;
        RECT 80.915 143.875 82.565 144.395 ;
        RECT 83.010 144.355 83.255 144.960 ;
        RECT 83.475 144.630 83.985 145.165 ;
        RECT 82.735 144.185 83.965 144.355 ;
        RECT 76.295 142.785 76.605 143.585 ;
        RECT 78.115 143.415 78.375 143.665 ;
        RECT 76.775 142.615 77.085 143.415 ;
        RECT 77.255 143.245 78.375 143.415 ;
        RECT 77.255 142.785 77.515 143.245 ;
        RECT 77.685 142.615 77.940 143.075 ;
        RECT 78.115 142.785 78.375 143.245 ;
        RECT 78.545 142.615 78.830 143.485 ;
        RECT 79.055 142.615 82.565 143.705 ;
        RECT 82.735 143.375 83.075 144.185 ;
        RECT 83.245 143.620 83.995 143.810 ;
        RECT 82.735 142.965 83.250 143.375 ;
        RECT 83.485 142.615 83.655 143.375 ;
        RECT 83.825 142.955 83.995 143.620 ;
        RECT 84.165 143.635 84.355 144.995 ;
        RECT 84.525 144.145 84.800 144.995 ;
        RECT 84.990 144.630 85.520 144.995 ;
        RECT 85.945 144.765 86.275 145.165 ;
        RECT 85.345 144.595 85.520 144.630 ;
        RECT 84.525 143.975 84.805 144.145 ;
        RECT 84.525 143.835 84.800 143.975 ;
        RECT 85.005 143.635 85.175 144.435 ;
        RECT 84.165 143.465 85.175 143.635 ;
        RECT 85.345 144.425 86.275 144.595 ;
        RECT 86.445 144.425 86.700 144.995 ;
        RECT 86.875 144.440 87.165 145.165 ;
        RECT 87.885 144.615 88.055 144.995 ;
        RECT 88.235 144.785 88.565 145.165 ;
        RECT 87.885 144.445 88.550 144.615 ;
        RECT 88.745 144.490 89.005 144.995 ;
        RECT 85.345 143.295 85.515 144.425 ;
        RECT 86.105 144.255 86.275 144.425 ;
        RECT 84.390 143.125 85.515 143.295 ;
        RECT 85.685 143.925 85.880 144.255 ;
        RECT 86.105 143.925 86.360 144.255 ;
        RECT 85.685 142.955 85.855 143.925 ;
        RECT 86.530 143.755 86.700 144.425 ;
        RECT 87.815 143.895 88.145 144.265 ;
        RECT 88.380 144.190 88.550 144.445 ;
        RECT 88.380 143.860 88.665 144.190 ;
        RECT 83.825 142.785 85.855 142.955 ;
        RECT 86.025 142.615 86.195 143.755 ;
        RECT 86.365 142.785 86.700 143.755 ;
        RECT 86.875 142.615 87.165 143.780 ;
        RECT 88.380 143.715 88.550 143.860 ;
        RECT 87.885 143.545 88.550 143.715 ;
        RECT 88.835 143.690 89.005 144.490 ;
        RECT 89.450 144.355 89.695 144.960 ;
        RECT 89.915 144.630 90.425 145.165 ;
        RECT 87.885 142.785 88.055 143.545 ;
        RECT 88.235 142.615 88.565 143.375 ;
        RECT 88.735 142.785 89.005 143.690 ;
        RECT 89.175 144.185 90.405 144.355 ;
        RECT 89.175 143.375 89.515 144.185 ;
        RECT 89.685 143.620 90.435 143.810 ;
        RECT 89.175 142.965 89.690 143.375 ;
        RECT 89.925 142.615 90.095 143.375 ;
        RECT 90.265 142.955 90.435 143.620 ;
        RECT 90.605 143.635 90.795 144.995 ;
        RECT 90.965 144.145 91.240 144.995 ;
        RECT 91.430 144.630 91.960 144.995 ;
        RECT 92.385 144.765 92.715 145.165 ;
        RECT 91.785 144.595 91.960 144.630 ;
        RECT 90.965 143.975 91.245 144.145 ;
        RECT 90.965 143.835 91.240 143.975 ;
        RECT 91.445 143.635 91.615 144.435 ;
        RECT 90.605 143.465 91.615 143.635 ;
        RECT 91.785 144.425 92.715 144.595 ;
        RECT 92.885 144.425 93.140 144.995 ;
        RECT 91.785 143.295 91.955 144.425 ;
        RECT 92.545 144.255 92.715 144.425 ;
        RECT 90.830 143.125 91.955 143.295 ;
        RECT 92.125 143.925 92.320 144.255 ;
        RECT 92.545 143.925 92.800 144.255 ;
        RECT 92.125 142.955 92.295 143.925 ;
        RECT 92.970 143.755 93.140 144.425 ;
        RECT 93.315 144.395 94.985 145.165 ;
        RECT 95.160 144.620 100.505 145.165 ;
        RECT 90.265 142.785 92.295 142.955 ;
        RECT 92.465 142.615 92.635 143.755 ;
        RECT 92.805 142.785 93.140 143.755 ;
        RECT 93.315 143.705 94.065 144.225 ;
        RECT 94.235 143.875 94.985 144.395 ;
        RECT 93.315 142.615 94.985 143.705 ;
        RECT 96.750 143.050 97.100 144.300 ;
        RECT 98.580 143.790 98.920 144.620 ;
        RECT 100.675 144.490 100.945 144.835 ;
        RECT 101.135 144.765 101.515 145.165 ;
        RECT 101.685 144.595 101.855 144.945 ;
        RECT 102.025 144.765 102.355 145.165 ;
        RECT 102.555 144.595 102.725 144.945 ;
        RECT 102.925 144.665 103.255 145.165 ;
        RECT 100.675 143.755 100.845 144.490 ;
        RECT 101.115 144.425 102.725 144.595 ;
        RECT 103.550 144.535 103.835 144.995 ;
        RECT 104.005 144.705 104.275 145.165 ;
        RECT 101.115 144.255 101.285 144.425 ;
        RECT 101.015 143.925 101.285 144.255 ;
        RECT 101.455 143.925 101.860 144.255 ;
        RECT 101.115 143.755 101.285 143.925 ;
        RECT 102.030 143.805 102.740 144.255 ;
        RECT 102.910 143.925 103.260 144.495 ;
        RECT 103.550 144.365 104.505 144.535 ;
        RECT 95.160 142.615 100.505 143.050 ;
        RECT 100.675 142.785 100.945 143.755 ;
        RECT 101.115 143.585 101.840 143.755 ;
        RECT 102.030 143.635 102.745 143.805 ;
        RECT 101.670 143.465 101.840 143.585 ;
        RECT 102.940 143.465 103.260 143.755 ;
        RECT 103.435 143.635 104.125 144.195 ;
        RECT 104.295 143.465 104.505 144.365 ;
        RECT 101.155 142.615 101.435 143.415 ;
        RECT 101.670 143.295 103.260 143.465 ;
        RECT 103.550 143.245 104.505 143.465 ;
        RECT 104.675 144.195 105.075 144.995 ;
        RECT 105.265 144.535 105.545 144.995 ;
        RECT 106.065 144.705 106.390 145.165 ;
        RECT 105.265 144.365 106.390 144.535 ;
        RECT 106.560 144.425 106.945 144.995 ;
        RECT 105.940 144.255 106.390 144.365 ;
        RECT 104.675 143.635 105.770 144.195 ;
        RECT 105.940 143.925 106.495 144.255 ;
        RECT 101.605 142.835 103.260 143.125 ;
        RECT 103.550 142.785 103.835 143.245 ;
        RECT 104.005 142.615 104.275 143.075 ;
        RECT 104.675 142.785 105.075 143.635 ;
        RECT 105.940 143.465 106.390 143.925 ;
        RECT 106.665 143.755 106.945 144.425 ;
        RECT 105.265 143.245 106.390 143.465 ;
        RECT 105.265 142.785 105.545 143.245 ;
        RECT 106.065 142.615 106.390 143.075 ;
        RECT 106.560 142.785 106.945 143.755 ;
        RECT 107.115 144.365 107.455 144.995 ;
        RECT 107.625 144.365 107.875 145.165 ;
        RECT 108.065 144.515 108.395 144.995 ;
        RECT 108.565 144.705 108.790 145.165 ;
        RECT 108.960 144.515 109.290 144.995 ;
        RECT 107.115 144.315 107.345 144.365 ;
        RECT 108.065 144.345 109.290 144.515 ;
        RECT 109.920 144.385 110.420 144.995 ;
        RECT 110.795 144.395 112.465 145.165 ;
        RECT 112.635 144.440 112.925 145.165 ;
        RECT 113.095 144.415 114.305 145.165 ;
        RECT 107.115 143.755 107.290 144.315 ;
        RECT 107.460 144.005 108.155 144.175 ;
        RECT 107.985 143.755 108.155 144.005 ;
        RECT 108.330 143.975 108.750 144.175 ;
        RECT 108.920 143.975 109.250 144.175 ;
        RECT 109.420 143.975 109.750 144.175 ;
        RECT 109.920 143.755 110.090 144.385 ;
        RECT 110.275 143.925 110.625 144.175 ;
        RECT 107.115 142.785 107.455 143.755 ;
        RECT 107.625 142.615 107.795 143.755 ;
        RECT 107.985 143.585 110.420 143.755 ;
        RECT 108.065 142.615 108.315 143.415 ;
        RECT 108.960 142.785 109.290 143.585 ;
        RECT 109.590 142.615 109.920 143.415 ;
        RECT 110.090 142.785 110.420 143.585 ;
        RECT 110.795 143.705 111.545 144.225 ;
        RECT 111.715 143.875 112.465 144.395 ;
        RECT 110.795 142.615 112.465 143.705 ;
        RECT 112.635 142.615 112.925 143.780 ;
        RECT 113.095 143.705 113.615 144.245 ;
        RECT 113.785 143.875 114.305 144.415 ;
        RECT 114.850 144.455 115.105 144.985 ;
        RECT 115.285 144.705 115.570 145.165 ;
        RECT 114.850 143.805 115.030 144.455 ;
        RECT 115.750 144.255 116.000 144.905 ;
        RECT 115.200 143.925 116.000 144.255 ;
        RECT 113.095 142.615 114.305 143.705 ;
        RECT 114.765 143.635 115.030 143.805 ;
        RECT 114.850 143.595 115.030 143.635 ;
        RECT 114.850 142.925 115.105 143.595 ;
        RECT 115.285 142.615 115.570 143.415 ;
        RECT 115.750 143.335 116.000 143.925 ;
        RECT 116.200 144.570 116.520 144.900 ;
        RECT 116.700 144.685 117.360 145.165 ;
        RECT 117.560 144.775 118.410 144.945 ;
        RECT 116.200 143.675 116.390 144.570 ;
        RECT 116.710 144.245 117.370 144.515 ;
        RECT 117.040 144.185 117.370 144.245 ;
        RECT 116.560 144.015 116.890 144.075 ;
        RECT 117.560 144.015 117.730 144.775 ;
        RECT 118.970 144.705 119.290 145.165 ;
        RECT 119.490 144.525 119.740 144.955 ;
        RECT 120.030 144.725 120.440 145.165 ;
        RECT 120.610 144.785 121.625 144.985 ;
        RECT 117.900 144.355 119.150 144.525 ;
        RECT 117.900 144.235 118.230 144.355 ;
        RECT 116.560 143.845 118.460 144.015 ;
        RECT 116.200 143.505 118.120 143.675 ;
        RECT 116.200 143.485 116.520 143.505 ;
        RECT 115.750 142.825 116.080 143.335 ;
        RECT 116.350 142.875 116.520 143.485 ;
        RECT 118.290 143.335 118.460 143.845 ;
        RECT 118.630 143.775 118.810 144.185 ;
        RECT 118.980 143.595 119.150 144.355 ;
        RECT 116.690 142.615 117.020 143.305 ;
        RECT 117.250 143.165 118.460 143.335 ;
        RECT 118.630 143.285 119.150 143.595 ;
        RECT 119.320 144.185 119.740 144.525 ;
        RECT 120.030 144.185 120.440 144.515 ;
        RECT 119.320 143.415 119.510 144.185 ;
        RECT 120.610 144.055 120.780 144.785 ;
        RECT 121.925 144.615 122.095 144.945 ;
        RECT 122.265 144.785 122.595 145.165 ;
        RECT 120.950 144.235 121.300 144.605 ;
        RECT 120.610 144.015 121.030 144.055 ;
        RECT 119.680 143.845 121.030 144.015 ;
        RECT 119.680 143.685 119.930 143.845 ;
        RECT 120.440 143.415 120.690 143.675 ;
        RECT 119.320 143.165 120.690 143.415 ;
        RECT 117.250 142.875 117.490 143.165 ;
        RECT 118.290 143.085 118.460 143.165 ;
        RECT 117.690 142.615 118.110 142.995 ;
        RECT 118.290 142.835 118.920 143.085 ;
        RECT 119.390 142.615 119.720 142.995 ;
        RECT 119.890 142.875 120.060 143.165 ;
        RECT 120.860 143.000 121.030 143.845 ;
        RECT 121.480 143.675 121.700 144.545 ;
        RECT 121.925 144.425 122.620 144.615 ;
        RECT 121.200 143.295 121.700 143.675 ;
        RECT 121.870 143.625 122.280 144.245 ;
        RECT 122.450 143.455 122.620 144.425 ;
        RECT 121.925 143.285 122.620 143.455 ;
        RECT 120.240 142.615 120.620 142.995 ;
        RECT 120.860 142.830 121.690 143.000 ;
        RECT 121.925 142.785 122.095 143.285 ;
        RECT 122.265 142.615 122.595 143.115 ;
        RECT 122.810 142.785 123.035 144.905 ;
        RECT 123.205 144.785 123.535 145.165 ;
        RECT 123.705 144.615 123.875 144.905 ;
        RECT 123.210 144.445 123.875 144.615 ;
        RECT 123.210 143.455 123.440 144.445 ;
        RECT 124.595 144.415 125.805 145.165 ;
        RECT 123.610 143.625 123.960 144.275 ;
        RECT 124.595 143.705 125.115 144.245 ;
        RECT 125.285 143.875 125.805 144.415 ;
        RECT 123.210 143.285 123.875 143.455 ;
        RECT 123.205 142.615 123.535 143.115 ;
        RECT 123.705 142.785 123.875 143.285 ;
        RECT 124.595 142.615 125.805 143.705 ;
        RECT 11.810 142.445 125.890 142.615 ;
        RECT 11.895 141.355 13.105 142.445 ;
        RECT 11.895 140.645 12.415 141.185 ;
        RECT 12.585 140.815 13.105 141.355 ;
        RECT 13.735 141.355 15.405 142.445 ;
        RECT 15.580 142.010 20.925 142.445 ;
        RECT 13.735 140.835 14.485 141.355 ;
        RECT 14.655 140.665 15.405 141.185 ;
        RECT 17.170 140.760 17.520 142.010 ;
        RECT 21.185 141.515 21.355 142.275 ;
        RECT 21.535 141.685 21.865 142.445 ;
        RECT 21.185 141.345 21.850 141.515 ;
        RECT 22.035 141.370 22.305 142.275 ;
        RECT 11.895 139.895 13.105 140.645 ;
        RECT 13.735 139.895 15.405 140.665 ;
        RECT 19.000 140.440 19.340 141.270 ;
        RECT 21.680 141.200 21.850 141.345 ;
        RECT 21.115 140.795 21.445 141.165 ;
        RECT 21.680 140.870 21.965 141.200 ;
        RECT 21.680 140.615 21.850 140.870 ;
        RECT 21.185 140.445 21.850 140.615 ;
        RECT 22.135 140.570 22.305 141.370 ;
        RECT 22.475 141.280 22.765 142.445 ;
        RECT 22.975 141.305 23.205 142.445 ;
        RECT 23.375 141.295 23.705 142.275 ;
        RECT 23.875 141.305 24.085 142.445 ;
        RECT 24.315 141.355 25.985 142.445 ;
        RECT 26.155 141.685 26.670 142.095 ;
        RECT 26.905 141.685 27.075 142.445 ;
        RECT 27.245 142.105 29.275 142.275 ;
        RECT 22.955 140.885 23.285 141.135 ;
        RECT 15.580 139.895 20.925 140.440 ;
        RECT 21.185 140.065 21.355 140.445 ;
        RECT 21.535 139.895 21.865 140.275 ;
        RECT 22.045 140.065 22.305 140.570 ;
        RECT 22.475 139.895 22.765 140.620 ;
        RECT 22.975 139.895 23.205 140.715 ;
        RECT 23.455 140.695 23.705 141.295 ;
        RECT 24.315 140.835 25.065 141.355 ;
        RECT 23.375 140.065 23.705 140.695 ;
        RECT 23.875 139.895 24.085 140.715 ;
        RECT 25.235 140.665 25.985 141.185 ;
        RECT 26.155 140.875 26.495 141.685 ;
        RECT 27.245 141.440 27.415 142.105 ;
        RECT 27.810 141.765 28.935 141.935 ;
        RECT 26.665 141.250 27.415 141.440 ;
        RECT 27.585 141.425 28.595 141.595 ;
        RECT 26.155 140.705 27.385 140.875 ;
        RECT 24.315 139.895 25.985 140.665 ;
        RECT 26.430 140.100 26.675 140.705 ;
        RECT 26.895 139.895 27.405 140.430 ;
        RECT 27.585 140.065 27.775 141.425 ;
        RECT 27.945 141.085 28.220 141.225 ;
        RECT 27.945 140.915 28.225 141.085 ;
        RECT 27.945 140.065 28.220 140.915 ;
        RECT 28.425 140.625 28.595 141.425 ;
        RECT 28.765 140.635 28.935 141.765 ;
        RECT 29.105 141.135 29.275 142.105 ;
        RECT 29.445 141.305 29.615 142.445 ;
        RECT 29.785 141.305 30.120 142.275 ;
        RECT 29.105 140.805 29.300 141.135 ;
        RECT 29.525 140.805 29.780 141.135 ;
        RECT 29.525 140.635 29.695 140.805 ;
        RECT 29.950 140.635 30.120 141.305 ;
        RECT 30.295 141.355 31.965 142.445 ;
        RECT 32.335 141.775 32.615 142.445 ;
        RECT 32.785 141.555 33.085 142.105 ;
        RECT 33.285 141.725 33.615 142.445 ;
        RECT 33.805 141.725 34.265 142.275 ;
        RECT 30.295 140.835 31.045 141.355 ;
        RECT 31.215 140.665 31.965 141.185 ;
        RECT 32.150 141.135 32.415 141.495 ;
        RECT 32.785 141.385 33.725 141.555 ;
        RECT 33.555 141.135 33.725 141.385 ;
        RECT 32.150 140.885 32.825 141.135 ;
        RECT 33.045 140.885 33.385 141.135 ;
        RECT 33.555 140.805 33.845 141.135 ;
        RECT 33.555 140.715 33.725 140.805 ;
        RECT 28.765 140.465 29.695 140.635 ;
        RECT 28.765 140.430 28.940 140.465 ;
        RECT 28.410 140.065 28.940 140.430 ;
        RECT 29.365 139.895 29.695 140.295 ;
        RECT 29.865 140.065 30.120 140.635 ;
        RECT 30.295 139.895 31.965 140.665 ;
        RECT 32.335 140.525 33.725 140.715 ;
        RECT 32.335 140.165 32.665 140.525 ;
        RECT 34.015 140.355 34.265 141.725 ;
        RECT 33.285 139.895 33.535 140.355 ;
        RECT 33.705 140.065 34.265 140.355 ;
        RECT 34.435 141.305 34.705 142.275 ;
        RECT 34.915 141.645 35.195 142.445 ;
        RECT 35.365 141.935 37.020 142.225 ;
        RECT 35.430 141.595 37.020 141.765 ;
        RECT 35.430 141.475 35.600 141.595 ;
        RECT 34.875 141.305 35.600 141.475 ;
        RECT 34.435 140.570 34.605 141.305 ;
        RECT 34.875 141.135 35.045 141.305 ;
        RECT 35.790 141.255 36.505 141.425 ;
        RECT 36.700 141.305 37.020 141.595 ;
        RECT 37.195 141.305 37.465 142.275 ;
        RECT 37.675 141.645 37.955 142.445 ;
        RECT 38.125 141.935 39.780 142.225 ;
        RECT 40.155 141.775 40.435 142.445 ;
        RECT 38.190 141.595 39.780 141.765 ;
        RECT 38.190 141.475 38.360 141.595 ;
        RECT 37.635 141.305 38.360 141.475 ;
        RECT 34.775 140.805 35.045 141.135 ;
        RECT 35.215 140.805 35.620 141.135 ;
        RECT 35.790 140.805 36.500 141.255 ;
        RECT 34.875 140.635 35.045 140.805 ;
        RECT 34.435 140.225 34.705 140.570 ;
        RECT 34.875 140.465 36.485 140.635 ;
        RECT 36.670 140.565 37.020 141.135 ;
        RECT 37.195 140.570 37.365 141.305 ;
        RECT 37.635 141.135 37.805 141.305 ;
        RECT 37.535 140.805 37.805 141.135 ;
        RECT 37.975 140.805 38.380 141.135 ;
        RECT 38.550 140.805 39.260 141.425 ;
        RECT 39.460 141.305 39.780 141.595 ;
        RECT 40.605 141.555 40.905 142.105 ;
        RECT 41.105 141.725 41.435 142.445 ;
        RECT 41.625 141.725 42.085 142.275 ;
        RECT 42.720 142.010 48.065 142.445 ;
        RECT 39.970 141.135 40.235 141.495 ;
        RECT 40.605 141.385 41.545 141.555 ;
        RECT 41.375 141.135 41.545 141.385 ;
        RECT 37.635 140.635 37.805 140.805 ;
        RECT 34.895 139.895 35.275 140.295 ;
        RECT 35.445 140.115 35.615 140.465 ;
        RECT 35.785 139.895 36.115 140.295 ;
        RECT 36.315 140.115 36.485 140.465 ;
        RECT 36.685 139.895 37.015 140.395 ;
        RECT 37.195 140.225 37.465 140.570 ;
        RECT 37.635 140.465 39.245 140.635 ;
        RECT 39.430 140.565 39.780 141.135 ;
        RECT 39.970 140.885 40.645 141.135 ;
        RECT 40.865 140.885 41.205 141.135 ;
        RECT 41.375 140.805 41.665 141.135 ;
        RECT 41.375 140.715 41.545 140.805 ;
        RECT 37.655 139.895 38.035 140.295 ;
        RECT 38.205 140.115 38.375 140.465 ;
        RECT 38.545 139.895 38.875 140.295 ;
        RECT 39.075 140.115 39.245 140.465 ;
        RECT 40.155 140.525 41.545 140.715 ;
        RECT 39.445 139.895 39.775 140.395 ;
        RECT 40.155 140.165 40.485 140.525 ;
        RECT 41.835 140.355 42.085 141.725 ;
        RECT 44.310 140.760 44.660 142.010 ;
        RECT 48.235 141.280 48.525 142.445 ;
        RECT 46.140 140.440 46.480 141.270 ;
        RECT 48.700 141.255 48.955 142.135 ;
        RECT 49.125 141.305 49.430 142.445 ;
        RECT 49.770 142.065 50.100 142.445 ;
        RECT 50.280 141.895 50.450 142.185 ;
        RECT 50.620 141.985 50.870 142.445 ;
        RECT 49.650 141.725 50.450 141.895 ;
        RECT 51.040 141.935 51.910 142.275 ;
        RECT 41.105 139.895 41.355 140.355 ;
        RECT 41.525 140.065 42.085 140.355 ;
        RECT 42.720 139.895 48.065 140.440 ;
        RECT 48.235 139.895 48.525 140.620 ;
        RECT 48.700 140.605 48.910 141.255 ;
        RECT 49.650 141.135 49.820 141.725 ;
        RECT 51.040 141.555 51.210 141.935 ;
        RECT 52.145 141.815 52.315 142.275 ;
        RECT 52.485 141.985 52.855 142.445 ;
        RECT 53.150 141.845 53.320 142.185 ;
        RECT 53.490 142.015 53.820 142.445 ;
        RECT 54.055 141.845 54.225 142.185 ;
        RECT 49.990 141.385 51.210 141.555 ;
        RECT 51.380 141.475 51.840 141.765 ;
        RECT 52.145 141.645 52.705 141.815 ;
        RECT 53.150 141.675 54.225 141.845 ;
        RECT 54.395 141.945 55.075 142.275 ;
        RECT 55.290 141.945 55.540 142.275 ;
        RECT 55.710 141.985 55.960 142.445 ;
        RECT 52.535 141.505 52.705 141.645 ;
        RECT 51.380 141.465 52.345 141.475 ;
        RECT 51.040 141.295 51.210 141.385 ;
        RECT 51.670 141.305 52.345 141.465 ;
        RECT 49.080 141.105 49.820 141.135 ;
        RECT 49.080 140.805 49.995 141.105 ;
        RECT 49.670 140.630 49.995 140.805 ;
        RECT 48.700 140.075 48.955 140.605 ;
        RECT 49.125 139.895 49.430 140.355 ;
        RECT 49.675 140.275 49.995 140.630 ;
        RECT 50.165 140.845 50.705 141.215 ;
        RECT 51.040 141.125 51.445 141.295 ;
        RECT 50.165 140.445 50.405 140.845 ;
        RECT 50.885 140.675 51.105 140.955 ;
        RECT 50.575 140.505 51.105 140.675 ;
        RECT 50.575 140.275 50.745 140.505 ;
        RECT 51.275 140.345 51.445 141.125 ;
        RECT 51.615 140.515 51.965 141.135 ;
        RECT 52.135 140.515 52.345 141.305 ;
        RECT 52.535 141.335 54.035 141.505 ;
        RECT 52.535 140.645 52.705 141.335 ;
        RECT 54.395 141.165 54.565 141.945 ;
        RECT 55.370 141.815 55.540 141.945 ;
        RECT 52.875 140.995 54.565 141.165 ;
        RECT 54.735 141.385 55.200 141.775 ;
        RECT 55.370 141.645 55.765 141.815 ;
        RECT 52.875 140.815 53.045 140.995 ;
        RECT 49.675 140.105 50.745 140.275 ;
        RECT 50.915 139.895 51.105 140.335 ;
        RECT 51.275 140.065 52.225 140.345 ;
        RECT 52.535 140.255 52.795 140.645 ;
        RECT 53.215 140.575 54.005 140.825 ;
        RECT 52.445 140.085 52.795 140.255 ;
        RECT 53.005 139.895 53.335 140.355 ;
        RECT 54.210 140.285 54.380 140.995 ;
        RECT 54.735 140.795 54.905 141.385 ;
        RECT 54.550 140.575 54.905 140.795 ;
        RECT 55.075 140.575 55.425 141.195 ;
        RECT 55.595 140.285 55.765 141.645 ;
        RECT 56.130 141.475 56.455 142.260 ;
        RECT 55.935 140.425 56.395 141.475 ;
        RECT 54.210 140.115 55.065 140.285 ;
        RECT 55.270 140.115 55.765 140.285 ;
        RECT 55.935 139.895 56.265 140.255 ;
        RECT 56.625 140.155 56.795 142.275 ;
        RECT 56.965 141.945 57.295 142.445 ;
        RECT 57.465 141.775 57.720 142.275 ;
        RECT 56.970 141.605 57.720 141.775 ;
        RECT 56.970 140.615 57.200 141.605 ;
        RECT 57.370 140.785 57.720 141.435 ;
        RECT 57.895 141.305 58.235 142.275 ;
        RECT 58.405 141.305 58.575 142.445 ;
        RECT 58.845 141.645 59.095 142.445 ;
        RECT 59.740 141.475 60.070 142.275 ;
        RECT 60.370 141.645 60.700 142.445 ;
        RECT 60.870 141.475 61.200 142.275 ;
        RECT 58.765 141.305 61.200 141.475 ;
        RECT 62.035 141.355 63.705 142.445 ;
        RECT 64.250 141.465 64.505 142.135 ;
        RECT 64.685 141.645 64.970 142.445 ;
        RECT 65.150 141.725 65.480 142.235 ;
        RECT 57.895 140.695 58.070 141.305 ;
        RECT 58.765 141.055 58.935 141.305 ;
        RECT 58.240 140.885 58.935 141.055 ;
        RECT 59.110 140.885 59.530 141.085 ;
        RECT 59.700 140.885 60.030 141.085 ;
        RECT 60.200 140.885 60.530 141.085 ;
        RECT 56.970 140.445 57.720 140.615 ;
        RECT 56.965 139.895 57.295 140.275 ;
        RECT 57.465 140.155 57.720 140.445 ;
        RECT 57.895 140.065 58.235 140.695 ;
        RECT 58.405 139.895 58.655 140.695 ;
        RECT 58.845 140.545 60.070 140.715 ;
        RECT 58.845 140.065 59.175 140.545 ;
        RECT 59.345 139.895 59.570 140.355 ;
        RECT 59.740 140.065 60.070 140.545 ;
        RECT 60.700 140.675 60.870 141.305 ;
        RECT 61.055 140.885 61.405 141.135 ;
        RECT 62.035 140.835 62.785 141.355 ;
        RECT 60.700 140.065 61.200 140.675 ;
        RECT 62.955 140.665 63.705 141.185 ;
        RECT 62.035 139.895 63.705 140.665 ;
        RECT 64.250 140.605 64.430 141.465 ;
        RECT 65.150 141.135 65.400 141.725 ;
        RECT 65.750 141.575 65.920 142.185 ;
        RECT 66.090 141.755 66.420 142.445 ;
        RECT 66.650 141.895 66.890 142.185 ;
        RECT 67.090 142.065 67.510 142.445 ;
        RECT 67.690 141.975 68.320 142.225 ;
        RECT 68.790 142.065 69.120 142.445 ;
        RECT 67.690 141.895 67.860 141.975 ;
        RECT 69.290 141.895 69.460 142.185 ;
        RECT 69.640 142.065 70.020 142.445 ;
        RECT 70.260 142.060 71.090 142.230 ;
        RECT 66.650 141.725 67.860 141.895 ;
        RECT 64.600 140.805 65.400 141.135 ;
        RECT 64.250 140.405 64.505 140.605 ;
        RECT 64.165 140.235 64.505 140.405 ;
        RECT 64.250 140.075 64.505 140.235 ;
        RECT 64.685 139.895 64.970 140.355 ;
        RECT 65.150 140.155 65.400 140.805 ;
        RECT 65.600 141.555 65.920 141.575 ;
        RECT 65.600 141.385 67.520 141.555 ;
        RECT 65.600 140.490 65.790 141.385 ;
        RECT 67.690 141.215 67.860 141.725 ;
        RECT 68.030 141.465 68.550 141.775 ;
        RECT 65.960 141.045 67.860 141.215 ;
        RECT 65.960 140.985 66.290 141.045 ;
        RECT 66.440 140.815 66.770 140.875 ;
        RECT 66.110 140.545 66.770 140.815 ;
        RECT 65.600 140.160 65.920 140.490 ;
        RECT 66.100 139.895 66.760 140.375 ;
        RECT 66.960 140.285 67.130 141.045 ;
        RECT 68.030 140.875 68.210 141.285 ;
        RECT 67.300 140.705 67.630 140.825 ;
        RECT 68.380 140.705 68.550 141.465 ;
        RECT 67.300 140.535 68.550 140.705 ;
        RECT 68.720 141.645 70.090 141.895 ;
        RECT 68.720 140.875 68.910 141.645 ;
        RECT 69.840 141.385 70.090 141.645 ;
        RECT 69.080 141.215 69.330 141.375 ;
        RECT 70.260 141.215 70.430 142.060 ;
        RECT 71.325 141.775 71.495 142.275 ;
        RECT 71.665 141.945 71.995 142.445 ;
        RECT 70.600 141.385 71.100 141.765 ;
        RECT 71.325 141.605 72.020 141.775 ;
        RECT 69.080 141.045 70.430 141.215 ;
        RECT 70.010 141.005 70.430 141.045 ;
        RECT 68.720 140.535 69.140 140.875 ;
        RECT 69.430 140.545 69.840 140.875 ;
        RECT 66.960 140.115 67.810 140.285 ;
        RECT 68.370 139.895 68.690 140.355 ;
        RECT 68.890 140.105 69.140 140.535 ;
        RECT 69.430 139.895 69.840 140.335 ;
        RECT 70.010 140.275 70.180 141.005 ;
        RECT 70.350 140.455 70.700 140.825 ;
        RECT 70.880 140.515 71.100 141.385 ;
        RECT 71.270 140.815 71.680 141.435 ;
        RECT 71.850 140.635 72.020 141.605 ;
        RECT 71.325 140.445 72.020 140.635 ;
        RECT 70.010 140.075 71.025 140.275 ;
        RECT 71.325 140.115 71.495 140.445 ;
        RECT 71.665 139.895 71.995 140.275 ;
        RECT 72.210 140.155 72.435 142.275 ;
        RECT 72.605 141.945 72.935 142.445 ;
        RECT 73.105 141.775 73.275 142.275 ;
        RECT 72.610 141.605 73.275 141.775 ;
        RECT 72.610 140.615 72.840 141.605 ;
        RECT 73.010 140.785 73.360 141.435 ;
        RECT 73.995 141.280 74.285 142.445 ;
        RECT 75.375 141.305 75.645 142.275 ;
        RECT 75.855 141.645 76.135 142.445 ;
        RECT 76.305 141.935 77.960 142.225 ;
        RECT 76.370 141.595 77.960 141.765 ;
        RECT 76.370 141.475 76.540 141.595 ;
        RECT 75.815 141.305 76.540 141.475 ;
        RECT 72.610 140.445 73.275 140.615 ;
        RECT 72.605 139.895 72.935 140.275 ;
        RECT 73.105 140.155 73.275 140.445 ;
        RECT 73.995 139.895 74.285 140.620 ;
        RECT 75.375 140.570 75.545 141.305 ;
        RECT 75.815 141.135 75.985 141.305 ;
        RECT 76.730 141.255 77.445 141.425 ;
        RECT 77.640 141.305 77.960 141.595 ;
        RECT 78.135 141.305 78.475 142.275 ;
        RECT 78.645 141.305 78.815 142.445 ;
        RECT 79.085 141.645 79.335 142.445 ;
        RECT 79.980 141.475 80.310 142.275 ;
        RECT 80.610 141.645 80.940 142.445 ;
        RECT 81.110 141.475 81.440 142.275 ;
        RECT 79.005 141.305 81.440 141.475 ;
        RECT 82.190 141.465 82.445 142.135 ;
        RECT 82.625 141.645 82.910 142.445 ;
        RECT 83.090 141.725 83.420 142.235 ;
        RECT 75.715 140.805 75.985 141.135 ;
        RECT 76.155 140.805 76.560 141.135 ;
        RECT 76.730 140.805 77.440 141.255 ;
        RECT 75.815 140.635 75.985 140.805 ;
        RECT 75.375 140.225 75.645 140.570 ;
        RECT 75.815 140.465 77.425 140.635 ;
        RECT 77.610 140.565 77.960 141.135 ;
        RECT 78.135 140.745 78.310 141.305 ;
        RECT 79.005 141.055 79.175 141.305 ;
        RECT 78.480 140.885 79.175 141.055 ;
        RECT 79.350 140.885 79.770 141.085 ;
        RECT 79.940 140.885 80.270 141.085 ;
        RECT 80.440 140.885 80.770 141.085 ;
        RECT 78.135 140.695 78.365 140.745 ;
        RECT 75.835 139.895 76.215 140.295 ;
        RECT 76.385 140.115 76.555 140.465 ;
        RECT 76.725 139.895 77.055 140.295 ;
        RECT 77.255 140.115 77.425 140.465 ;
        RECT 77.625 139.895 77.955 140.395 ;
        RECT 78.135 140.065 78.475 140.695 ;
        RECT 78.645 139.895 78.895 140.695 ;
        RECT 79.085 140.545 80.310 140.715 ;
        RECT 79.085 140.065 79.415 140.545 ;
        RECT 79.585 139.895 79.810 140.355 ;
        RECT 79.980 140.065 80.310 140.545 ;
        RECT 80.940 140.675 81.110 141.305 ;
        RECT 81.295 140.885 81.645 141.135 ;
        RECT 80.940 140.065 81.440 140.675 ;
        RECT 82.190 140.605 82.370 141.465 ;
        RECT 83.090 141.135 83.340 141.725 ;
        RECT 83.690 141.575 83.860 142.185 ;
        RECT 84.030 141.755 84.360 142.445 ;
        RECT 84.590 141.895 84.830 142.185 ;
        RECT 85.030 142.065 85.450 142.445 ;
        RECT 85.630 141.975 86.260 142.225 ;
        RECT 86.730 142.065 87.060 142.445 ;
        RECT 85.630 141.895 85.800 141.975 ;
        RECT 87.230 141.895 87.400 142.185 ;
        RECT 87.580 142.065 87.960 142.445 ;
        RECT 88.200 142.060 89.030 142.230 ;
        RECT 84.590 141.725 85.800 141.895 ;
        RECT 82.540 140.805 83.340 141.135 ;
        RECT 82.190 140.405 82.445 140.605 ;
        RECT 82.105 140.235 82.445 140.405 ;
        RECT 82.190 140.075 82.445 140.235 ;
        RECT 82.625 139.895 82.910 140.355 ;
        RECT 83.090 140.155 83.340 140.805 ;
        RECT 83.540 141.555 83.860 141.575 ;
        RECT 83.540 141.385 85.460 141.555 ;
        RECT 83.540 140.490 83.730 141.385 ;
        RECT 85.630 141.215 85.800 141.725 ;
        RECT 85.970 141.465 86.490 141.775 ;
        RECT 83.900 141.045 85.800 141.215 ;
        RECT 83.900 140.985 84.230 141.045 ;
        RECT 84.380 140.815 84.710 140.875 ;
        RECT 84.050 140.545 84.710 140.815 ;
        RECT 83.540 140.160 83.860 140.490 ;
        RECT 84.040 139.895 84.700 140.375 ;
        RECT 84.900 140.285 85.070 141.045 ;
        RECT 85.970 140.875 86.150 141.285 ;
        RECT 85.240 140.705 85.570 140.825 ;
        RECT 86.320 140.705 86.490 141.465 ;
        RECT 85.240 140.535 86.490 140.705 ;
        RECT 86.660 141.645 88.030 141.895 ;
        RECT 86.660 140.875 86.850 141.645 ;
        RECT 87.780 141.385 88.030 141.645 ;
        RECT 87.020 141.215 87.270 141.375 ;
        RECT 88.200 141.215 88.370 142.060 ;
        RECT 89.265 141.775 89.435 142.275 ;
        RECT 89.605 141.945 89.935 142.445 ;
        RECT 88.540 141.385 89.040 141.765 ;
        RECT 89.265 141.605 89.960 141.775 ;
        RECT 87.020 141.045 88.370 141.215 ;
        RECT 87.950 141.005 88.370 141.045 ;
        RECT 86.660 140.535 87.080 140.875 ;
        RECT 87.370 140.545 87.780 140.875 ;
        RECT 84.900 140.115 85.750 140.285 ;
        RECT 86.310 139.895 86.630 140.355 ;
        RECT 86.830 140.105 87.080 140.535 ;
        RECT 87.370 139.895 87.780 140.335 ;
        RECT 87.950 140.275 88.120 141.005 ;
        RECT 88.290 140.455 88.640 140.825 ;
        RECT 88.820 140.515 89.040 141.385 ;
        RECT 89.210 140.815 89.620 141.435 ;
        RECT 89.790 140.635 89.960 141.605 ;
        RECT 89.265 140.445 89.960 140.635 ;
        RECT 87.950 140.075 88.965 140.275 ;
        RECT 89.265 140.115 89.435 140.445 ;
        RECT 89.605 139.895 89.935 140.275 ;
        RECT 90.150 140.155 90.375 142.275 ;
        RECT 90.545 141.945 90.875 142.445 ;
        RECT 91.045 141.775 91.215 142.275 ;
        RECT 90.550 141.605 91.215 141.775 ;
        RECT 90.550 140.615 90.780 141.605 ;
        RECT 90.950 140.785 91.300 141.435 ;
        RECT 91.475 141.355 93.145 142.445 ;
        RECT 93.320 141.935 94.975 142.225 ;
        RECT 93.320 141.595 94.910 141.765 ;
        RECT 95.145 141.645 95.425 142.445 ;
        RECT 91.475 140.835 92.225 141.355 ;
        RECT 93.320 141.305 93.640 141.595 ;
        RECT 94.740 141.475 94.910 141.595 ;
        RECT 92.395 140.665 93.145 141.185 ;
        RECT 90.550 140.445 91.215 140.615 ;
        RECT 90.545 139.895 90.875 140.275 ;
        RECT 91.045 140.155 91.215 140.445 ;
        RECT 91.475 139.895 93.145 140.665 ;
        RECT 93.320 140.565 93.670 141.135 ;
        RECT 93.840 140.805 94.550 141.425 ;
        RECT 94.740 141.305 95.465 141.475 ;
        RECT 95.635 141.305 95.905 142.275 ;
        RECT 95.295 141.135 95.465 141.305 ;
        RECT 94.720 140.805 95.125 141.135 ;
        RECT 95.295 140.805 95.565 141.135 ;
        RECT 95.295 140.635 95.465 140.805 ;
        RECT 93.855 140.465 95.465 140.635 ;
        RECT 95.735 140.570 95.905 141.305 ;
        RECT 93.325 139.895 93.655 140.395 ;
        RECT 93.855 140.115 94.025 140.465 ;
        RECT 94.225 139.895 94.555 140.295 ;
        RECT 94.725 140.115 94.895 140.465 ;
        RECT 95.065 139.895 95.445 140.295 ;
        RECT 95.635 140.225 95.905 140.570 ;
        RECT 96.075 141.305 96.415 142.275 ;
        RECT 96.585 141.305 96.755 142.445 ;
        RECT 97.025 141.645 97.275 142.445 ;
        RECT 97.920 141.475 98.250 142.275 ;
        RECT 98.550 141.645 98.880 142.445 ;
        RECT 99.050 141.475 99.380 142.275 ;
        RECT 96.945 141.305 99.380 141.475 ;
        RECT 96.075 140.745 96.250 141.305 ;
        RECT 96.945 141.055 97.115 141.305 ;
        RECT 96.420 140.885 97.115 141.055 ;
        RECT 97.290 140.885 97.710 141.085 ;
        RECT 97.880 140.885 98.210 141.085 ;
        RECT 98.380 140.885 98.710 141.085 ;
        RECT 96.075 140.695 96.305 140.745 ;
        RECT 96.075 140.065 96.415 140.695 ;
        RECT 96.585 139.895 96.835 140.695 ;
        RECT 97.025 140.545 98.250 140.715 ;
        RECT 97.025 140.065 97.355 140.545 ;
        RECT 97.525 139.895 97.750 140.355 ;
        RECT 97.920 140.065 98.250 140.545 ;
        RECT 98.880 140.675 99.050 141.305 ;
        RECT 99.755 141.280 100.045 142.445 ;
        RECT 100.215 141.355 103.725 142.445 ;
        RECT 99.235 140.885 99.585 141.135 ;
        RECT 100.215 140.835 101.905 141.355 ;
        RECT 103.895 141.305 104.235 142.275 ;
        RECT 104.405 141.305 104.575 142.445 ;
        RECT 104.845 141.645 105.095 142.445 ;
        RECT 105.740 141.475 106.070 142.275 ;
        RECT 106.370 141.645 106.700 142.445 ;
        RECT 106.870 141.475 107.200 142.275 ;
        RECT 104.765 141.305 107.200 141.475 ;
        RECT 107.575 141.355 109.245 142.445 ;
        RECT 109.415 141.685 109.930 142.095 ;
        RECT 110.165 141.685 110.335 142.445 ;
        RECT 110.505 142.105 112.535 142.275 ;
        RECT 98.880 140.065 99.380 140.675 ;
        RECT 102.075 140.665 103.725 141.185 ;
        RECT 99.755 139.895 100.045 140.620 ;
        RECT 100.215 139.895 103.725 140.665 ;
        RECT 103.895 140.695 104.070 141.305 ;
        RECT 104.765 141.055 104.935 141.305 ;
        RECT 104.240 140.885 104.935 141.055 ;
        RECT 105.110 140.885 105.530 141.085 ;
        RECT 105.700 140.885 106.030 141.085 ;
        RECT 106.200 140.885 106.530 141.085 ;
        RECT 103.895 140.065 104.235 140.695 ;
        RECT 104.405 139.895 104.655 140.695 ;
        RECT 104.845 140.545 106.070 140.715 ;
        RECT 104.845 140.065 105.175 140.545 ;
        RECT 105.345 139.895 105.570 140.355 ;
        RECT 105.740 140.065 106.070 140.545 ;
        RECT 106.700 140.675 106.870 141.305 ;
        RECT 107.055 140.885 107.405 141.135 ;
        RECT 107.575 140.835 108.325 141.355 ;
        RECT 106.700 140.065 107.200 140.675 ;
        RECT 108.495 140.665 109.245 141.185 ;
        RECT 109.415 140.875 109.755 141.685 ;
        RECT 110.505 141.440 110.675 142.105 ;
        RECT 111.070 141.765 112.195 141.935 ;
        RECT 109.925 141.250 110.675 141.440 ;
        RECT 110.845 141.425 111.855 141.595 ;
        RECT 109.415 140.705 110.645 140.875 ;
        RECT 107.575 139.895 109.245 140.665 ;
        RECT 109.690 140.100 109.935 140.705 ;
        RECT 110.155 139.895 110.665 140.430 ;
        RECT 110.845 140.065 111.035 141.425 ;
        RECT 111.205 140.405 111.480 141.225 ;
        RECT 111.685 140.625 111.855 141.425 ;
        RECT 112.025 140.635 112.195 141.765 ;
        RECT 112.365 141.135 112.535 142.105 ;
        RECT 112.705 141.305 112.875 142.445 ;
        RECT 113.045 141.305 113.380 142.275 ;
        RECT 112.365 140.805 112.560 141.135 ;
        RECT 112.785 140.805 113.040 141.135 ;
        RECT 112.785 140.635 112.955 140.805 ;
        RECT 113.210 140.635 113.380 141.305 ;
        RECT 113.555 141.685 114.070 142.095 ;
        RECT 114.305 141.685 114.475 142.445 ;
        RECT 114.645 142.105 116.675 142.275 ;
        RECT 113.555 140.875 113.895 141.685 ;
        RECT 114.645 141.440 114.815 142.105 ;
        RECT 115.210 141.765 116.335 141.935 ;
        RECT 114.065 141.250 114.815 141.440 ;
        RECT 114.985 141.425 115.995 141.595 ;
        RECT 113.555 140.705 114.785 140.875 ;
        RECT 112.025 140.465 112.955 140.635 ;
        RECT 112.025 140.430 112.200 140.465 ;
        RECT 111.205 140.235 111.485 140.405 ;
        RECT 111.205 140.065 111.480 140.235 ;
        RECT 111.670 140.065 112.200 140.430 ;
        RECT 112.625 139.895 112.955 140.295 ;
        RECT 113.125 140.065 113.380 140.635 ;
        RECT 113.830 140.100 114.075 140.705 ;
        RECT 114.295 139.895 114.805 140.430 ;
        RECT 114.985 140.065 115.175 141.425 ;
        RECT 115.345 141.085 115.620 141.225 ;
        RECT 115.345 140.915 115.625 141.085 ;
        RECT 115.345 140.065 115.620 140.915 ;
        RECT 115.825 140.625 115.995 141.425 ;
        RECT 116.165 140.635 116.335 141.765 ;
        RECT 116.505 141.135 116.675 142.105 ;
        RECT 116.845 141.305 117.015 142.445 ;
        RECT 117.185 141.305 117.520 142.275 ;
        RECT 117.735 141.305 117.965 142.445 ;
        RECT 116.505 140.805 116.700 141.135 ;
        RECT 116.925 140.805 117.180 141.135 ;
        RECT 116.925 140.635 117.095 140.805 ;
        RECT 117.350 140.635 117.520 141.305 ;
        RECT 118.135 141.295 118.465 142.275 ;
        RECT 118.635 141.305 118.845 142.445 ;
        RECT 119.625 141.515 119.795 142.275 ;
        RECT 119.975 141.685 120.305 142.445 ;
        RECT 119.625 141.345 120.290 141.515 ;
        RECT 120.475 141.370 120.745 142.275 ;
        RECT 117.715 140.885 118.045 141.135 ;
        RECT 116.165 140.465 117.095 140.635 ;
        RECT 116.165 140.430 116.340 140.465 ;
        RECT 115.810 140.065 116.340 140.430 ;
        RECT 116.765 139.895 117.095 140.295 ;
        RECT 117.265 140.065 117.520 140.635 ;
        RECT 117.735 139.895 117.965 140.715 ;
        RECT 118.215 140.695 118.465 141.295 ;
        RECT 120.120 141.200 120.290 141.345 ;
        RECT 119.555 140.795 119.885 141.165 ;
        RECT 120.120 140.870 120.405 141.200 ;
        RECT 118.135 140.065 118.465 140.695 ;
        RECT 118.635 139.895 118.845 140.715 ;
        RECT 120.120 140.615 120.290 140.870 ;
        RECT 119.625 140.445 120.290 140.615 ;
        RECT 120.575 140.570 120.745 141.370 ;
        RECT 120.915 141.355 124.425 142.445 ;
        RECT 124.595 141.355 125.805 142.445 ;
        RECT 120.915 140.835 122.605 141.355 ;
        RECT 122.775 140.665 124.425 141.185 ;
        RECT 124.595 140.815 125.115 141.355 ;
        RECT 119.625 140.065 119.795 140.445 ;
        RECT 119.975 139.895 120.305 140.275 ;
        RECT 120.485 140.065 120.745 140.570 ;
        RECT 120.915 139.895 124.425 140.665 ;
        RECT 125.285 140.645 125.805 141.185 ;
        RECT 124.595 139.895 125.805 140.645 ;
        RECT 11.810 139.725 125.890 139.895 ;
        RECT 11.895 138.975 13.105 139.725 ;
        RECT 11.895 138.435 12.415 138.975 ;
        RECT 14.255 138.905 14.465 139.725 ;
        RECT 14.635 138.925 14.965 139.555 ;
        RECT 12.585 138.265 13.105 138.805 ;
        RECT 14.635 138.325 14.885 138.925 ;
        RECT 15.135 138.905 15.365 139.725 ;
        RECT 15.850 138.915 16.095 139.520 ;
        RECT 16.315 139.190 16.825 139.725 ;
        RECT 15.575 138.745 16.805 138.915 ;
        RECT 15.055 138.485 15.385 138.735 ;
        RECT 11.895 137.175 13.105 138.265 ;
        RECT 14.255 137.175 14.465 138.315 ;
        RECT 14.635 137.345 14.965 138.325 ;
        RECT 15.135 137.175 15.365 138.315 ;
        RECT 15.575 137.935 15.915 138.745 ;
        RECT 16.085 138.180 16.835 138.370 ;
        RECT 15.575 137.525 16.090 137.935 ;
        RECT 16.325 137.175 16.495 137.935 ;
        RECT 16.665 137.515 16.835 138.180 ;
        RECT 17.005 138.195 17.195 139.555 ;
        RECT 17.365 139.385 17.640 139.555 ;
        RECT 17.365 139.215 17.645 139.385 ;
        RECT 17.365 138.395 17.640 139.215 ;
        RECT 17.830 139.190 18.360 139.555 ;
        RECT 18.785 139.325 19.115 139.725 ;
        RECT 18.185 139.155 18.360 139.190 ;
        RECT 17.845 138.195 18.015 138.995 ;
        RECT 17.005 138.025 18.015 138.195 ;
        RECT 18.185 138.985 19.115 139.155 ;
        RECT 19.285 138.985 19.540 139.555 ;
        RECT 20.090 139.045 20.345 139.545 ;
        RECT 20.525 139.265 20.810 139.725 ;
        RECT 18.185 137.855 18.355 138.985 ;
        RECT 18.945 138.815 19.115 138.985 ;
        RECT 17.230 137.685 18.355 137.855 ;
        RECT 18.525 138.485 18.720 138.815 ;
        RECT 18.945 138.485 19.200 138.815 ;
        RECT 18.525 137.515 18.695 138.485 ;
        RECT 19.370 138.315 19.540 138.985 ;
        RECT 20.005 139.015 20.345 139.045 ;
        RECT 20.005 138.875 20.270 139.015 ;
        RECT 16.665 137.345 18.695 137.515 ;
        RECT 18.865 137.175 19.035 138.315 ;
        RECT 19.205 137.345 19.540 138.315 ;
        RECT 20.090 138.155 20.270 138.875 ;
        RECT 20.990 138.815 21.240 139.465 ;
        RECT 20.440 138.485 21.240 138.815 ;
        RECT 20.090 137.485 20.345 138.155 ;
        RECT 20.525 137.175 20.810 137.975 ;
        RECT 20.990 137.895 21.240 138.485 ;
        RECT 21.440 139.130 21.760 139.460 ;
        RECT 21.940 139.245 22.600 139.725 ;
        RECT 22.800 139.335 23.650 139.505 ;
        RECT 21.440 138.235 21.630 139.130 ;
        RECT 21.950 138.805 22.610 139.075 ;
        RECT 22.280 138.745 22.610 138.805 ;
        RECT 21.800 138.575 22.130 138.635 ;
        RECT 22.800 138.575 22.970 139.335 ;
        RECT 24.210 139.265 24.530 139.725 ;
        RECT 24.730 139.085 24.980 139.515 ;
        RECT 25.270 139.285 25.680 139.725 ;
        RECT 25.850 139.345 26.865 139.545 ;
        RECT 23.140 138.915 24.390 139.085 ;
        RECT 23.140 138.795 23.470 138.915 ;
        RECT 21.800 138.405 23.700 138.575 ;
        RECT 21.440 138.065 23.360 138.235 ;
        RECT 21.440 138.045 21.760 138.065 ;
        RECT 20.990 137.385 21.320 137.895 ;
        RECT 21.590 137.435 21.760 138.045 ;
        RECT 23.530 137.895 23.700 138.405 ;
        RECT 23.870 138.335 24.050 138.745 ;
        RECT 24.220 138.155 24.390 138.915 ;
        RECT 21.930 137.175 22.260 137.865 ;
        RECT 22.490 137.725 23.700 137.895 ;
        RECT 23.870 137.845 24.390 138.155 ;
        RECT 24.560 138.745 24.980 139.085 ;
        RECT 25.270 138.745 25.680 139.075 ;
        RECT 24.560 137.975 24.750 138.745 ;
        RECT 25.850 138.615 26.020 139.345 ;
        RECT 27.165 139.175 27.335 139.505 ;
        RECT 27.505 139.345 27.835 139.725 ;
        RECT 26.190 138.795 26.540 139.165 ;
        RECT 25.850 138.575 26.270 138.615 ;
        RECT 24.920 138.405 26.270 138.575 ;
        RECT 24.920 138.245 25.170 138.405 ;
        RECT 25.680 137.975 25.930 138.235 ;
        RECT 24.560 137.725 25.930 137.975 ;
        RECT 22.490 137.435 22.730 137.725 ;
        RECT 23.530 137.645 23.700 137.725 ;
        RECT 22.930 137.175 23.350 137.555 ;
        RECT 23.530 137.395 24.160 137.645 ;
        RECT 24.630 137.175 24.960 137.555 ;
        RECT 25.130 137.435 25.300 137.725 ;
        RECT 26.100 137.560 26.270 138.405 ;
        RECT 26.720 138.235 26.940 139.105 ;
        RECT 27.165 138.985 27.860 139.175 ;
        RECT 26.440 137.855 26.940 138.235 ;
        RECT 27.110 138.185 27.520 138.805 ;
        RECT 27.690 138.015 27.860 138.985 ;
        RECT 27.165 137.845 27.860 138.015 ;
        RECT 25.480 137.175 25.860 137.555 ;
        RECT 26.100 137.390 26.930 137.560 ;
        RECT 27.165 137.345 27.335 137.845 ;
        RECT 27.505 137.175 27.835 137.675 ;
        RECT 28.050 137.345 28.275 139.465 ;
        RECT 28.445 139.345 28.775 139.725 ;
        RECT 28.945 139.175 29.115 139.465 ;
        RECT 28.450 139.005 29.115 139.175 ;
        RECT 29.375 139.050 29.635 139.555 ;
        RECT 29.815 139.345 30.145 139.725 ;
        RECT 30.325 139.175 30.495 139.555 ;
        RECT 28.450 138.015 28.680 139.005 ;
        RECT 28.850 138.185 29.200 138.835 ;
        RECT 29.375 138.250 29.545 139.050 ;
        RECT 29.830 139.005 30.495 139.175 ;
        RECT 29.830 138.750 30.000 139.005 ;
        RECT 31.490 138.915 31.735 139.520 ;
        RECT 31.955 139.190 32.465 139.725 ;
        RECT 29.715 138.420 30.000 138.750 ;
        RECT 30.235 138.455 30.565 138.825 ;
        RECT 31.215 138.745 32.445 138.915 ;
        RECT 29.830 138.275 30.000 138.420 ;
        RECT 28.450 137.845 29.115 138.015 ;
        RECT 28.445 137.175 28.775 137.675 ;
        RECT 28.945 137.345 29.115 137.845 ;
        RECT 29.375 137.345 29.645 138.250 ;
        RECT 29.830 138.105 30.495 138.275 ;
        RECT 29.815 137.175 30.145 137.935 ;
        RECT 30.325 137.345 30.495 138.105 ;
        RECT 31.215 137.935 31.555 138.745 ;
        RECT 31.725 138.180 32.475 138.370 ;
        RECT 31.215 137.525 31.730 137.935 ;
        RECT 31.965 137.175 32.135 137.935 ;
        RECT 32.305 137.515 32.475 138.180 ;
        RECT 32.645 138.195 32.835 139.555 ;
        RECT 33.005 138.705 33.280 139.555 ;
        RECT 33.470 139.190 34.000 139.555 ;
        RECT 34.425 139.325 34.755 139.725 ;
        RECT 33.825 139.155 34.000 139.190 ;
        RECT 33.005 138.535 33.285 138.705 ;
        RECT 33.005 138.395 33.280 138.535 ;
        RECT 33.485 138.195 33.655 138.995 ;
        RECT 32.645 138.025 33.655 138.195 ;
        RECT 33.825 138.985 34.755 139.155 ;
        RECT 34.925 138.985 35.180 139.555 ;
        RECT 35.355 139.000 35.645 139.725 ;
        RECT 36.015 139.095 36.345 139.455 ;
        RECT 36.965 139.265 37.215 139.725 ;
        RECT 37.385 139.265 37.945 139.555 ;
        RECT 33.825 137.855 33.995 138.985 ;
        RECT 34.585 138.815 34.755 138.985 ;
        RECT 32.870 137.685 33.995 137.855 ;
        RECT 34.165 138.485 34.360 138.815 ;
        RECT 34.585 138.485 34.840 138.815 ;
        RECT 34.165 137.515 34.335 138.485 ;
        RECT 35.010 138.315 35.180 138.985 ;
        RECT 36.015 138.905 37.405 139.095 ;
        RECT 37.235 138.815 37.405 138.905 ;
        RECT 35.830 138.485 36.505 138.735 ;
        RECT 36.725 138.485 37.065 138.735 ;
        RECT 37.235 138.485 37.525 138.815 ;
        RECT 32.305 137.345 34.335 137.515 ;
        RECT 34.505 137.175 34.675 138.315 ;
        RECT 34.845 137.345 35.180 138.315 ;
        RECT 35.355 137.175 35.645 138.340 ;
        RECT 35.830 138.125 36.095 138.485 ;
        RECT 37.235 138.235 37.405 138.485 ;
        RECT 36.465 138.065 37.405 138.235 ;
        RECT 36.015 137.175 36.295 137.845 ;
        RECT 36.465 137.515 36.765 138.065 ;
        RECT 37.695 137.895 37.945 139.265 ;
        RECT 36.965 137.175 37.295 137.895 ;
        RECT 37.485 137.345 37.945 137.895 ;
        RECT 38.115 139.265 38.675 139.555 ;
        RECT 38.845 139.265 39.095 139.725 ;
        RECT 38.115 137.895 38.365 139.265 ;
        RECT 39.715 139.095 40.045 139.455 ;
        RECT 38.655 138.905 40.045 139.095 ;
        RECT 40.415 138.955 43.925 139.725 ;
        RECT 44.105 139.225 44.435 139.725 ;
        RECT 44.635 139.155 44.805 139.505 ;
        RECT 45.005 139.325 45.335 139.725 ;
        RECT 45.505 139.155 45.675 139.505 ;
        RECT 45.845 139.325 46.225 139.725 ;
        RECT 38.655 138.815 38.825 138.905 ;
        RECT 38.535 138.485 38.825 138.815 ;
        RECT 38.995 138.485 39.335 138.735 ;
        RECT 39.555 138.485 40.230 138.735 ;
        RECT 38.655 138.235 38.825 138.485 ;
        RECT 38.655 138.065 39.595 138.235 ;
        RECT 39.965 138.125 40.230 138.485 ;
        RECT 40.415 138.265 42.105 138.785 ;
        RECT 42.275 138.435 43.925 138.955 ;
        RECT 44.100 138.485 44.450 139.055 ;
        RECT 44.635 138.985 46.245 139.155 ;
        RECT 46.415 139.050 46.685 139.395 ;
        RECT 46.075 138.815 46.245 138.985 ;
        RECT 38.115 137.345 38.575 137.895 ;
        RECT 38.765 137.175 39.095 137.895 ;
        RECT 39.295 137.515 39.595 138.065 ;
        RECT 39.765 137.175 40.045 137.845 ;
        RECT 40.415 137.175 43.925 138.265 ;
        RECT 44.100 138.025 44.420 138.315 ;
        RECT 44.620 138.195 45.330 138.815 ;
        RECT 45.500 138.485 45.905 138.815 ;
        RECT 46.075 138.485 46.345 138.815 ;
        RECT 46.075 138.315 46.245 138.485 ;
        RECT 46.515 138.315 46.685 139.050 ;
        RECT 45.520 138.145 46.245 138.315 ;
        RECT 45.520 138.025 45.690 138.145 ;
        RECT 44.100 137.855 45.690 138.025 ;
        RECT 44.100 137.395 45.755 137.685 ;
        RECT 45.925 137.175 46.205 137.975 ;
        RECT 46.415 137.345 46.685 138.315 ;
        RECT 47.315 138.925 47.655 139.555 ;
        RECT 47.825 138.925 48.075 139.725 ;
        RECT 48.265 139.075 48.595 139.555 ;
        RECT 48.765 139.265 48.990 139.725 ;
        RECT 49.160 139.075 49.490 139.555 ;
        RECT 47.315 138.875 47.545 138.925 ;
        RECT 48.265 138.905 49.490 139.075 ;
        RECT 50.120 138.945 50.620 139.555 ;
        RECT 47.315 138.315 47.490 138.875 ;
        RECT 47.660 138.565 48.355 138.735 ;
        RECT 48.185 138.315 48.355 138.565 ;
        RECT 48.530 138.535 48.950 138.735 ;
        RECT 49.120 138.535 49.450 138.735 ;
        RECT 49.620 138.535 49.950 138.735 ;
        RECT 50.120 138.315 50.290 138.945 ;
        RECT 51.515 138.905 51.725 139.725 ;
        RECT 51.895 138.925 52.225 139.555 ;
        RECT 50.475 138.485 50.825 138.735 ;
        RECT 51.895 138.325 52.145 138.925 ;
        RECT 52.395 138.905 52.625 139.725 ;
        RECT 53.300 138.985 53.555 139.555 ;
        RECT 53.725 139.325 54.055 139.725 ;
        RECT 54.480 139.190 55.010 139.555 ;
        RECT 55.200 139.385 55.475 139.555 ;
        RECT 55.195 139.215 55.475 139.385 ;
        RECT 54.480 139.155 54.655 139.190 ;
        RECT 53.725 138.985 54.655 139.155 ;
        RECT 52.315 138.485 52.645 138.735 ;
        RECT 47.315 137.345 47.655 138.315 ;
        RECT 47.825 137.175 47.995 138.315 ;
        RECT 48.185 138.145 50.620 138.315 ;
        RECT 48.265 137.175 48.515 137.975 ;
        RECT 49.160 137.345 49.490 138.145 ;
        RECT 49.790 137.175 50.120 137.975 ;
        RECT 50.290 137.345 50.620 138.145 ;
        RECT 51.515 137.175 51.725 138.315 ;
        RECT 51.895 137.345 52.225 138.325 ;
        RECT 53.300 138.315 53.470 138.985 ;
        RECT 53.725 138.815 53.895 138.985 ;
        RECT 53.640 138.485 53.895 138.815 ;
        RECT 54.120 138.485 54.315 138.815 ;
        RECT 52.395 137.175 52.625 138.315 ;
        RECT 53.300 137.345 53.635 138.315 ;
        RECT 53.805 137.175 53.975 138.315 ;
        RECT 54.145 137.515 54.315 138.485 ;
        RECT 54.485 137.855 54.655 138.985 ;
        RECT 54.825 138.195 54.995 138.995 ;
        RECT 55.200 138.395 55.475 139.215 ;
        RECT 55.645 138.195 55.835 139.555 ;
        RECT 56.015 139.190 56.525 139.725 ;
        RECT 56.745 138.915 56.990 139.520 ;
        RECT 57.435 138.955 60.945 139.725 ;
        RECT 61.115 139.000 61.405 139.725 ;
        RECT 61.665 139.175 61.835 139.555 ;
        RECT 62.015 139.345 62.345 139.725 ;
        RECT 61.665 139.005 62.330 139.175 ;
        RECT 62.525 139.050 62.785 139.555 ;
        RECT 56.035 138.745 57.265 138.915 ;
        RECT 54.825 138.025 55.835 138.195 ;
        RECT 56.005 138.180 56.755 138.370 ;
        RECT 54.485 137.685 55.610 137.855 ;
        RECT 56.005 137.515 56.175 138.180 ;
        RECT 56.925 137.935 57.265 138.745 ;
        RECT 54.145 137.345 56.175 137.515 ;
        RECT 56.345 137.175 56.515 137.935 ;
        RECT 56.750 137.525 57.265 137.935 ;
        RECT 57.435 138.265 59.125 138.785 ;
        RECT 59.295 138.435 60.945 138.955 ;
        RECT 61.595 138.455 61.935 138.825 ;
        RECT 62.160 138.750 62.330 139.005 ;
        RECT 62.160 138.420 62.435 138.750 ;
        RECT 57.435 137.175 60.945 138.265 ;
        RECT 61.115 137.175 61.405 138.340 ;
        RECT 62.160 138.275 62.330 138.420 ;
        RECT 61.655 138.105 62.330 138.275 ;
        RECT 62.605 138.250 62.785 139.050 ;
        RECT 63.070 139.095 63.355 139.555 ;
        RECT 63.525 139.265 63.795 139.725 ;
        RECT 63.070 138.925 64.025 139.095 ;
        RECT 61.655 137.345 61.835 138.105 ;
        RECT 62.015 137.175 62.345 137.935 ;
        RECT 62.515 137.345 62.785 138.250 ;
        RECT 62.955 138.195 63.645 138.755 ;
        RECT 63.815 138.025 64.025 138.925 ;
        RECT 63.070 137.805 64.025 138.025 ;
        RECT 64.195 138.755 64.595 139.555 ;
        RECT 64.785 139.095 65.065 139.555 ;
        RECT 65.585 139.265 65.910 139.725 ;
        RECT 64.785 138.925 65.910 139.095 ;
        RECT 66.080 138.985 66.465 139.555 ;
        RECT 65.460 138.815 65.910 138.925 ;
        RECT 64.195 138.195 65.290 138.755 ;
        RECT 65.460 138.485 66.015 138.815 ;
        RECT 63.070 137.345 63.355 137.805 ;
        RECT 63.525 137.175 63.795 137.635 ;
        RECT 64.195 137.345 64.595 138.195 ;
        RECT 65.460 138.025 65.910 138.485 ;
        RECT 66.185 138.315 66.465 138.985 ;
        RECT 67.135 138.905 67.365 139.725 ;
        RECT 67.535 138.925 67.865 139.555 ;
        RECT 67.115 138.485 67.445 138.735 ;
        RECT 67.615 138.325 67.865 138.925 ;
        RECT 68.035 138.905 68.245 139.725 ;
        RECT 68.480 138.960 68.935 139.725 ;
        RECT 69.210 139.345 70.510 139.555 ;
        RECT 70.765 139.365 71.095 139.725 ;
        RECT 70.340 139.195 70.510 139.345 ;
        RECT 71.265 139.225 71.525 139.555 ;
        RECT 71.295 139.215 71.525 139.225 ;
        RECT 69.410 138.735 69.630 139.135 ;
        RECT 68.475 138.535 68.965 138.735 ;
        RECT 69.155 138.525 69.630 138.735 ;
        RECT 69.875 138.735 70.085 139.135 ;
        RECT 70.340 139.070 71.095 139.195 ;
        RECT 70.340 139.025 71.185 139.070 ;
        RECT 70.915 138.905 71.185 139.025 ;
        RECT 69.875 138.525 70.205 138.735 ;
        RECT 70.375 138.465 70.785 138.770 ;
        RECT 64.785 137.805 65.910 138.025 ;
        RECT 64.785 137.345 65.065 137.805 ;
        RECT 65.585 137.175 65.910 137.635 ;
        RECT 66.080 137.345 66.465 138.315 ;
        RECT 67.135 137.175 67.365 138.315 ;
        RECT 67.535 137.345 67.865 138.325 ;
        RECT 68.035 137.175 68.245 138.315 ;
        RECT 68.480 138.295 69.655 138.355 ;
        RECT 71.015 138.330 71.185 138.905 ;
        RECT 70.985 138.295 71.185 138.330 ;
        RECT 68.480 138.185 71.185 138.295 ;
        RECT 68.480 137.565 68.735 138.185 ;
        RECT 69.325 138.125 71.125 138.185 ;
        RECT 69.325 138.095 69.655 138.125 ;
        RECT 71.355 138.025 71.525 139.215 ;
        RECT 71.785 139.175 71.955 139.555 ;
        RECT 72.170 139.345 72.500 139.725 ;
        RECT 71.785 139.005 72.500 139.175 ;
        RECT 71.695 138.455 72.050 138.825 ;
        RECT 72.330 138.815 72.500 139.005 ;
        RECT 72.670 138.980 72.925 139.555 ;
        RECT 72.330 138.485 72.585 138.815 ;
        RECT 72.330 138.275 72.500 138.485 ;
        RECT 68.985 137.925 69.170 138.015 ;
        RECT 69.760 137.925 70.595 137.935 ;
        RECT 68.985 137.725 70.595 137.925 ;
        RECT 68.985 137.685 69.215 137.725 ;
        RECT 68.480 137.345 68.815 137.565 ;
        RECT 69.820 137.175 70.175 137.555 ;
        RECT 70.345 137.345 70.595 137.725 ;
        RECT 70.845 137.175 71.095 137.955 ;
        RECT 71.265 137.345 71.525 138.025 ;
        RECT 71.785 138.105 72.500 138.275 ;
        RECT 72.755 138.250 72.925 138.980 ;
        RECT 73.100 138.885 73.360 139.725 ;
        RECT 73.995 138.955 77.505 139.725 ;
        RECT 71.785 137.345 71.955 138.105 ;
        RECT 72.170 137.175 72.500 137.935 ;
        RECT 72.670 137.345 72.925 138.250 ;
        RECT 73.100 137.175 73.360 138.325 ;
        RECT 73.995 138.265 75.685 138.785 ;
        RECT 75.855 138.435 77.505 138.955 ;
        RECT 77.675 138.925 78.015 139.555 ;
        RECT 78.185 138.925 78.435 139.725 ;
        RECT 78.625 139.075 78.955 139.555 ;
        RECT 79.125 139.265 79.350 139.725 ;
        RECT 79.520 139.075 79.850 139.555 ;
        RECT 77.675 138.315 77.850 138.925 ;
        RECT 78.625 138.905 79.850 139.075 ;
        RECT 80.480 138.945 80.980 139.555 ;
        RECT 81.815 138.955 85.325 139.725 ;
        RECT 78.020 138.565 78.715 138.735 ;
        RECT 78.545 138.315 78.715 138.565 ;
        RECT 78.890 138.535 79.310 138.735 ;
        RECT 79.480 138.535 79.810 138.735 ;
        RECT 79.980 138.535 80.310 138.735 ;
        RECT 80.480 138.315 80.650 138.945 ;
        RECT 80.835 138.485 81.185 138.735 ;
        RECT 73.995 137.175 77.505 138.265 ;
        RECT 77.675 137.345 78.015 138.315 ;
        RECT 78.185 137.175 78.355 138.315 ;
        RECT 78.545 138.145 80.980 138.315 ;
        RECT 78.625 137.175 78.875 137.975 ;
        RECT 79.520 137.345 79.850 138.145 ;
        RECT 80.150 137.175 80.480 137.975 ;
        RECT 80.650 137.345 80.980 138.145 ;
        RECT 81.815 138.265 83.505 138.785 ;
        RECT 83.675 138.435 85.325 138.955 ;
        RECT 85.555 138.905 85.765 139.725 ;
        RECT 85.935 138.925 86.265 139.555 ;
        RECT 85.935 138.325 86.185 138.925 ;
        RECT 86.435 138.905 86.665 139.725 ;
        RECT 86.875 139.000 87.165 139.725 ;
        RECT 87.425 139.175 87.595 139.555 ;
        RECT 87.775 139.345 88.105 139.725 ;
        RECT 87.425 139.005 88.090 139.175 ;
        RECT 88.285 139.050 88.545 139.555 ;
        RECT 86.355 138.485 86.685 138.735 ;
        RECT 87.355 138.455 87.685 138.825 ;
        RECT 87.920 138.750 88.090 139.005 ;
        RECT 87.920 138.420 88.205 138.750 ;
        RECT 81.815 137.175 85.325 138.265 ;
        RECT 85.555 137.175 85.765 138.315 ;
        RECT 85.935 137.345 86.265 138.325 ;
        RECT 86.435 137.175 86.665 138.315 ;
        RECT 86.875 137.175 87.165 138.340 ;
        RECT 87.920 138.275 88.090 138.420 ;
        RECT 87.425 138.105 88.090 138.275 ;
        RECT 88.375 138.250 88.545 139.050 ;
        RECT 88.715 138.975 89.925 139.725 ;
        RECT 87.425 137.345 87.595 138.105 ;
        RECT 87.775 137.175 88.105 137.935 ;
        RECT 88.275 137.345 88.545 138.250 ;
        RECT 88.715 138.265 89.235 138.805 ;
        RECT 89.405 138.435 89.925 138.975 ;
        RECT 90.095 138.955 93.605 139.725 ;
        RECT 93.780 139.180 99.125 139.725 ;
        RECT 90.095 138.265 91.785 138.785 ;
        RECT 91.955 138.435 93.605 138.955 ;
        RECT 88.715 137.175 89.925 138.265 ;
        RECT 90.095 137.175 93.605 138.265 ;
        RECT 95.370 137.610 95.720 138.860 ;
        RECT 97.200 138.350 97.540 139.180 ;
        RECT 99.295 139.050 99.565 139.395 ;
        RECT 99.755 139.325 100.135 139.725 ;
        RECT 100.305 139.155 100.475 139.505 ;
        RECT 100.645 139.325 100.975 139.725 ;
        RECT 101.175 139.155 101.345 139.505 ;
        RECT 101.545 139.225 101.875 139.725 ;
        RECT 99.295 138.315 99.465 139.050 ;
        RECT 99.735 138.985 101.345 139.155 ;
        RECT 99.735 138.815 99.905 138.985 ;
        RECT 99.635 138.485 99.905 138.815 ;
        RECT 100.075 138.485 100.480 138.815 ;
        RECT 99.735 138.315 99.905 138.485 ;
        RECT 93.780 137.175 99.125 137.610 ;
        RECT 99.295 137.345 99.565 138.315 ;
        RECT 99.735 138.145 100.460 138.315 ;
        RECT 100.650 138.195 101.360 138.815 ;
        RECT 101.530 138.485 101.880 139.055 ;
        RECT 102.055 139.050 102.325 139.395 ;
        RECT 102.515 139.325 102.895 139.725 ;
        RECT 103.065 139.155 103.235 139.505 ;
        RECT 103.405 139.325 103.735 139.725 ;
        RECT 103.935 139.155 104.105 139.505 ;
        RECT 104.305 139.225 104.635 139.725 ;
        RECT 102.055 138.315 102.225 139.050 ;
        RECT 102.495 138.985 104.105 139.155 ;
        RECT 102.495 138.815 102.665 138.985 ;
        RECT 102.395 138.485 102.665 138.815 ;
        RECT 102.835 138.485 103.240 138.815 ;
        RECT 102.495 138.315 102.665 138.485 ;
        RECT 100.290 138.025 100.460 138.145 ;
        RECT 101.560 138.025 101.880 138.315 ;
        RECT 99.775 137.175 100.055 137.975 ;
        RECT 100.290 137.855 101.880 138.025 ;
        RECT 100.225 137.395 101.880 137.685 ;
        RECT 102.055 137.345 102.325 138.315 ;
        RECT 102.495 138.145 103.220 138.315 ;
        RECT 103.410 138.195 104.120 138.815 ;
        RECT 104.290 138.485 104.640 139.055 ;
        RECT 104.815 138.925 105.155 139.555 ;
        RECT 105.325 138.925 105.575 139.725 ;
        RECT 105.765 139.075 106.095 139.555 ;
        RECT 106.265 139.265 106.490 139.725 ;
        RECT 106.660 139.075 106.990 139.555 ;
        RECT 104.815 138.315 104.990 138.925 ;
        RECT 105.765 138.905 106.990 139.075 ;
        RECT 107.620 138.945 108.120 139.555 ;
        RECT 105.160 138.565 105.855 138.735 ;
        RECT 105.685 138.315 105.855 138.565 ;
        RECT 106.030 138.535 106.450 138.735 ;
        RECT 106.620 138.535 106.950 138.735 ;
        RECT 107.120 138.535 107.450 138.735 ;
        RECT 107.620 138.315 107.790 138.945 ;
        RECT 108.770 138.915 109.015 139.520 ;
        RECT 109.235 139.190 109.745 139.725 ;
        RECT 108.495 138.745 109.725 138.915 ;
        RECT 107.975 138.485 108.325 138.735 ;
        RECT 103.050 138.025 103.220 138.145 ;
        RECT 104.320 138.025 104.640 138.315 ;
        RECT 102.535 137.175 102.815 137.975 ;
        RECT 103.050 137.855 104.640 138.025 ;
        RECT 102.985 137.395 104.640 137.685 ;
        RECT 104.815 137.345 105.155 138.315 ;
        RECT 105.325 137.175 105.495 138.315 ;
        RECT 105.685 138.145 108.120 138.315 ;
        RECT 105.765 137.175 106.015 137.975 ;
        RECT 106.660 137.345 106.990 138.145 ;
        RECT 107.290 137.175 107.620 137.975 ;
        RECT 107.790 137.345 108.120 138.145 ;
        RECT 108.495 137.935 108.835 138.745 ;
        RECT 109.005 138.180 109.755 138.370 ;
        RECT 108.495 137.525 109.010 137.935 ;
        RECT 109.245 137.175 109.415 137.935 ;
        RECT 109.585 137.515 109.755 138.180 ;
        RECT 109.925 138.195 110.115 139.555 ;
        RECT 110.285 139.385 110.560 139.555 ;
        RECT 110.285 139.215 110.565 139.385 ;
        RECT 110.285 138.395 110.560 139.215 ;
        RECT 110.750 139.190 111.280 139.555 ;
        RECT 111.705 139.325 112.035 139.725 ;
        RECT 111.105 139.155 111.280 139.190 ;
        RECT 110.765 138.195 110.935 138.995 ;
        RECT 109.925 138.025 110.935 138.195 ;
        RECT 111.105 138.985 112.035 139.155 ;
        RECT 112.205 138.985 112.460 139.555 ;
        RECT 112.635 139.000 112.925 139.725 ;
        RECT 111.105 137.855 111.275 138.985 ;
        RECT 111.865 138.815 112.035 138.985 ;
        RECT 110.150 137.685 111.275 137.855 ;
        RECT 111.445 138.485 111.640 138.815 ;
        RECT 111.865 138.485 112.120 138.815 ;
        RECT 111.445 137.515 111.615 138.485 ;
        RECT 112.290 138.315 112.460 138.985 ;
        RECT 113.135 138.905 113.365 139.725 ;
        RECT 113.535 138.925 113.865 139.555 ;
        RECT 113.115 138.485 113.445 138.735 ;
        RECT 109.585 137.345 111.615 137.515 ;
        RECT 111.785 137.175 111.955 138.315 ;
        RECT 112.125 137.345 112.460 138.315 ;
        RECT 112.635 137.175 112.925 138.340 ;
        RECT 113.615 138.325 113.865 138.925 ;
        RECT 114.035 138.905 114.245 139.725 ;
        RECT 114.850 139.045 115.105 139.545 ;
        RECT 115.285 139.265 115.570 139.725 ;
        RECT 114.765 139.015 115.105 139.045 ;
        RECT 114.765 138.875 115.030 139.015 ;
        RECT 113.135 137.175 113.365 138.315 ;
        RECT 113.535 137.345 113.865 138.325 ;
        RECT 114.035 137.175 114.245 138.315 ;
        RECT 114.850 138.155 115.030 138.875 ;
        RECT 115.750 138.815 116.000 139.465 ;
        RECT 115.200 138.485 116.000 138.815 ;
        RECT 114.850 137.485 115.105 138.155 ;
        RECT 115.285 137.175 115.570 137.975 ;
        RECT 115.750 137.895 116.000 138.485 ;
        RECT 116.200 139.130 116.520 139.460 ;
        RECT 116.700 139.245 117.360 139.725 ;
        RECT 117.560 139.335 118.410 139.505 ;
        RECT 116.200 138.235 116.390 139.130 ;
        RECT 116.710 138.805 117.370 139.075 ;
        RECT 117.040 138.745 117.370 138.805 ;
        RECT 116.560 138.575 116.890 138.635 ;
        RECT 117.560 138.575 117.730 139.335 ;
        RECT 118.970 139.265 119.290 139.725 ;
        RECT 119.490 139.085 119.740 139.515 ;
        RECT 120.030 139.285 120.440 139.725 ;
        RECT 120.610 139.345 121.625 139.545 ;
        RECT 117.900 138.915 119.150 139.085 ;
        RECT 117.900 138.795 118.230 138.915 ;
        RECT 116.560 138.405 118.460 138.575 ;
        RECT 116.200 138.065 118.120 138.235 ;
        RECT 116.200 138.045 116.520 138.065 ;
        RECT 115.750 137.385 116.080 137.895 ;
        RECT 116.350 137.435 116.520 138.045 ;
        RECT 118.290 137.895 118.460 138.405 ;
        RECT 118.630 138.335 118.810 138.745 ;
        RECT 118.980 138.155 119.150 138.915 ;
        RECT 116.690 137.175 117.020 137.865 ;
        RECT 117.250 137.725 118.460 137.895 ;
        RECT 118.630 137.845 119.150 138.155 ;
        RECT 119.320 138.745 119.740 139.085 ;
        RECT 120.030 138.745 120.440 139.075 ;
        RECT 119.320 137.975 119.510 138.745 ;
        RECT 120.610 138.615 120.780 139.345 ;
        RECT 121.925 139.175 122.095 139.505 ;
        RECT 122.265 139.345 122.595 139.725 ;
        RECT 120.950 138.795 121.300 139.165 ;
        RECT 120.610 138.575 121.030 138.615 ;
        RECT 119.680 138.405 121.030 138.575 ;
        RECT 119.680 138.245 119.930 138.405 ;
        RECT 120.440 137.975 120.690 138.235 ;
        RECT 119.320 137.725 120.690 137.975 ;
        RECT 117.250 137.435 117.490 137.725 ;
        RECT 118.290 137.645 118.460 137.725 ;
        RECT 117.690 137.175 118.110 137.555 ;
        RECT 118.290 137.395 118.920 137.645 ;
        RECT 119.390 137.175 119.720 137.555 ;
        RECT 119.890 137.435 120.060 137.725 ;
        RECT 120.860 137.560 121.030 138.405 ;
        RECT 121.480 138.235 121.700 139.105 ;
        RECT 121.925 138.985 122.620 139.175 ;
        RECT 121.200 137.855 121.700 138.235 ;
        RECT 121.870 138.185 122.280 138.805 ;
        RECT 122.450 138.015 122.620 138.985 ;
        RECT 121.925 137.845 122.620 138.015 ;
        RECT 120.240 137.175 120.620 137.555 ;
        RECT 120.860 137.390 121.690 137.560 ;
        RECT 121.925 137.345 122.095 137.845 ;
        RECT 122.265 137.175 122.595 137.675 ;
        RECT 122.810 137.345 123.035 139.465 ;
        RECT 123.205 139.345 123.535 139.725 ;
        RECT 123.705 139.175 123.875 139.465 ;
        RECT 123.210 139.005 123.875 139.175 ;
        RECT 123.210 138.015 123.440 139.005 ;
        RECT 124.595 138.975 125.805 139.725 ;
        RECT 123.610 138.185 123.960 138.835 ;
        RECT 124.595 138.265 125.115 138.805 ;
        RECT 125.285 138.435 125.805 138.975 ;
        RECT 123.210 137.845 123.875 138.015 ;
        RECT 123.205 137.175 123.535 137.675 ;
        RECT 123.705 137.345 123.875 137.845 ;
        RECT 124.595 137.175 125.805 138.265 ;
        RECT 11.810 137.005 125.890 137.175 ;
        RECT 11.895 135.915 13.105 137.005 ;
        RECT 11.895 135.205 12.415 135.745 ;
        RECT 12.585 135.375 13.105 135.915 ;
        RECT 14.195 135.915 17.705 137.005 ;
        RECT 17.875 136.245 18.390 136.655 ;
        RECT 18.625 136.245 18.795 137.005 ;
        RECT 18.965 136.665 20.995 136.835 ;
        RECT 14.195 135.395 15.885 135.915 ;
        RECT 16.055 135.225 17.705 135.745 ;
        RECT 17.875 135.435 18.215 136.245 ;
        RECT 18.965 136.000 19.135 136.665 ;
        RECT 19.530 136.325 20.655 136.495 ;
        RECT 18.385 135.810 19.135 136.000 ;
        RECT 19.305 135.985 20.315 136.155 ;
        RECT 17.875 135.265 19.105 135.435 ;
        RECT 11.895 134.455 13.105 135.205 ;
        RECT 14.195 134.455 17.705 135.225 ;
        RECT 18.150 134.660 18.395 135.265 ;
        RECT 18.615 134.455 19.125 134.990 ;
        RECT 19.305 134.625 19.495 135.985 ;
        RECT 19.665 134.965 19.940 135.785 ;
        RECT 20.145 135.185 20.315 135.985 ;
        RECT 20.485 135.195 20.655 136.325 ;
        RECT 20.825 135.695 20.995 136.665 ;
        RECT 21.165 135.865 21.335 137.005 ;
        RECT 21.505 135.865 21.840 136.835 ;
        RECT 20.825 135.365 21.020 135.695 ;
        RECT 21.245 135.365 21.500 135.695 ;
        RECT 21.245 135.195 21.415 135.365 ;
        RECT 21.670 135.195 21.840 135.865 ;
        RECT 22.475 135.840 22.765 137.005 ;
        RECT 23.855 135.915 27.365 137.005 ;
        RECT 27.910 136.665 28.165 136.695 ;
        RECT 27.825 136.495 28.165 136.665 ;
        RECT 27.910 136.025 28.165 136.495 ;
        RECT 28.345 136.205 28.630 137.005 ;
        RECT 28.810 136.285 29.140 136.795 ;
        RECT 23.855 135.395 25.545 135.915 ;
        RECT 25.715 135.225 27.365 135.745 ;
        RECT 20.485 135.025 21.415 135.195 ;
        RECT 20.485 134.990 20.660 135.025 ;
        RECT 19.665 134.795 19.945 134.965 ;
        RECT 19.665 134.625 19.940 134.795 ;
        RECT 20.130 134.625 20.660 134.990 ;
        RECT 21.085 134.455 21.415 134.855 ;
        RECT 21.585 134.625 21.840 135.195 ;
        RECT 22.475 134.455 22.765 135.180 ;
        RECT 23.855 134.455 27.365 135.225 ;
        RECT 27.910 135.165 28.090 136.025 ;
        RECT 28.810 135.695 29.060 136.285 ;
        RECT 29.410 136.135 29.580 136.745 ;
        RECT 29.750 136.315 30.080 137.005 ;
        RECT 30.310 136.455 30.550 136.745 ;
        RECT 30.750 136.625 31.170 137.005 ;
        RECT 31.350 136.535 31.980 136.785 ;
        RECT 32.450 136.625 32.780 137.005 ;
        RECT 31.350 136.455 31.520 136.535 ;
        RECT 32.950 136.455 33.120 136.745 ;
        RECT 33.300 136.625 33.680 137.005 ;
        RECT 33.920 136.620 34.750 136.790 ;
        RECT 30.310 136.285 31.520 136.455 ;
        RECT 28.260 135.365 29.060 135.695 ;
        RECT 27.910 134.635 28.165 135.165 ;
        RECT 28.345 134.455 28.630 134.915 ;
        RECT 28.810 134.715 29.060 135.365 ;
        RECT 29.260 136.115 29.580 136.135 ;
        RECT 29.260 135.945 31.180 136.115 ;
        RECT 29.260 135.050 29.450 135.945 ;
        RECT 31.350 135.775 31.520 136.285 ;
        RECT 31.690 136.025 32.210 136.335 ;
        RECT 29.620 135.605 31.520 135.775 ;
        RECT 29.620 135.545 29.950 135.605 ;
        RECT 30.100 135.375 30.430 135.435 ;
        RECT 29.770 135.105 30.430 135.375 ;
        RECT 29.260 134.720 29.580 135.050 ;
        RECT 29.760 134.455 30.420 134.935 ;
        RECT 30.620 134.845 30.790 135.605 ;
        RECT 31.690 135.435 31.870 135.845 ;
        RECT 30.960 135.265 31.290 135.385 ;
        RECT 32.040 135.265 32.210 136.025 ;
        RECT 30.960 135.095 32.210 135.265 ;
        RECT 32.380 136.205 33.750 136.455 ;
        RECT 32.380 135.435 32.570 136.205 ;
        RECT 33.500 135.945 33.750 136.205 ;
        RECT 32.740 135.775 32.990 135.935 ;
        RECT 33.920 135.775 34.090 136.620 ;
        RECT 34.985 136.335 35.155 136.835 ;
        RECT 35.325 136.505 35.655 137.005 ;
        RECT 34.260 135.945 34.760 136.325 ;
        RECT 34.985 136.165 35.680 136.335 ;
        RECT 32.740 135.605 34.090 135.775 ;
        RECT 33.670 135.565 34.090 135.605 ;
        RECT 32.380 135.095 32.800 135.435 ;
        RECT 33.090 135.105 33.500 135.435 ;
        RECT 30.620 134.675 31.470 134.845 ;
        RECT 32.030 134.455 32.350 134.915 ;
        RECT 32.550 134.665 32.800 135.095 ;
        RECT 33.090 134.455 33.500 134.895 ;
        RECT 33.670 134.835 33.840 135.565 ;
        RECT 34.010 135.015 34.360 135.385 ;
        RECT 34.540 135.075 34.760 135.945 ;
        RECT 34.930 135.375 35.340 135.995 ;
        RECT 35.510 135.195 35.680 136.165 ;
        RECT 34.985 135.005 35.680 135.195 ;
        RECT 33.670 134.635 34.685 134.835 ;
        RECT 34.985 134.675 35.155 135.005 ;
        RECT 35.325 134.455 35.655 134.835 ;
        RECT 35.870 134.715 36.095 136.835 ;
        RECT 36.265 136.505 36.595 137.005 ;
        RECT 36.765 136.335 36.935 136.835 ;
        RECT 36.270 136.165 36.935 136.335 ;
        RECT 36.270 135.175 36.500 136.165 ;
        RECT 36.670 135.345 37.020 135.995 ;
        RECT 37.195 135.930 37.465 136.835 ;
        RECT 37.635 136.245 37.965 137.005 ;
        RECT 38.145 136.075 38.315 136.835 ;
        RECT 36.270 135.005 36.935 135.175 ;
        RECT 36.265 134.455 36.595 134.835 ;
        RECT 36.765 134.715 36.935 135.005 ;
        RECT 37.195 135.130 37.365 135.930 ;
        RECT 37.650 135.905 38.315 136.075 ;
        RECT 39.035 135.915 42.545 137.005 ;
        RECT 42.720 136.570 48.065 137.005 ;
        RECT 37.650 135.760 37.820 135.905 ;
        RECT 37.535 135.430 37.820 135.760 ;
        RECT 37.650 135.175 37.820 135.430 ;
        RECT 38.055 135.355 38.385 135.725 ;
        RECT 39.035 135.395 40.725 135.915 ;
        RECT 40.895 135.225 42.545 135.745 ;
        RECT 44.310 135.320 44.660 136.570 ;
        RECT 48.235 135.840 48.525 137.005 ;
        RECT 48.695 135.915 49.905 137.005 ;
        RECT 50.080 136.570 55.425 137.005 ;
        RECT 55.600 136.570 60.945 137.005 ;
        RECT 37.195 134.625 37.455 135.130 ;
        RECT 37.650 135.005 38.315 135.175 ;
        RECT 37.635 134.455 37.965 134.835 ;
        RECT 38.145 134.625 38.315 135.005 ;
        RECT 39.035 134.455 42.545 135.225 ;
        RECT 46.140 135.000 46.480 135.830 ;
        RECT 48.695 135.375 49.215 135.915 ;
        RECT 49.385 135.205 49.905 135.745 ;
        RECT 51.670 135.320 52.020 136.570 ;
        RECT 42.720 134.455 48.065 135.000 ;
        RECT 48.235 134.455 48.525 135.180 ;
        RECT 48.695 134.455 49.905 135.205 ;
        RECT 53.500 135.000 53.840 135.830 ;
        RECT 57.190 135.320 57.540 136.570 ;
        RECT 61.115 136.245 61.630 136.655 ;
        RECT 61.865 136.245 62.035 137.005 ;
        RECT 62.205 136.665 64.235 136.835 ;
        RECT 59.020 135.000 59.360 135.830 ;
        RECT 61.115 135.435 61.455 136.245 ;
        RECT 62.205 136.000 62.375 136.665 ;
        RECT 62.770 136.325 63.895 136.495 ;
        RECT 61.625 135.810 62.375 136.000 ;
        RECT 62.545 135.985 63.555 136.155 ;
        RECT 61.115 135.265 62.345 135.435 ;
        RECT 50.080 134.455 55.425 135.000 ;
        RECT 55.600 134.455 60.945 135.000 ;
        RECT 61.390 134.660 61.635 135.265 ;
        RECT 61.855 134.455 62.365 134.990 ;
        RECT 62.545 134.625 62.735 135.985 ;
        RECT 62.905 135.645 63.180 135.785 ;
        RECT 62.905 135.475 63.185 135.645 ;
        RECT 62.905 134.625 63.180 135.475 ;
        RECT 63.385 135.185 63.555 135.985 ;
        RECT 63.725 135.195 63.895 136.325 ;
        RECT 64.065 135.695 64.235 136.665 ;
        RECT 64.405 135.865 64.575 137.005 ;
        RECT 64.745 135.865 65.080 136.835 ;
        RECT 65.805 136.075 65.975 136.835 ;
        RECT 66.155 136.245 66.485 137.005 ;
        RECT 65.805 135.905 66.470 136.075 ;
        RECT 66.655 135.930 66.925 136.835 ;
        RECT 64.065 135.365 64.260 135.695 ;
        RECT 64.485 135.365 64.740 135.695 ;
        RECT 64.485 135.195 64.655 135.365 ;
        RECT 64.910 135.195 65.080 135.865 ;
        RECT 66.300 135.760 66.470 135.905 ;
        RECT 65.735 135.355 66.065 135.725 ;
        RECT 66.300 135.430 66.585 135.760 ;
        RECT 63.725 135.025 64.655 135.195 ;
        RECT 63.725 134.990 63.900 135.025 ;
        RECT 63.370 134.625 63.900 134.990 ;
        RECT 64.325 134.455 64.655 134.855 ;
        RECT 64.825 134.625 65.080 135.195 ;
        RECT 66.300 135.175 66.470 135.430 ;
        RECT 65.805 135.005 66.470 135.175 ;
        RECT 66.755 135.130 66.925 135.930 ;
        RECT 67.095 135.915 68.305 137.005 ;
        RECT 68.480 136.570 73.825 137.005 ;
        RECT 67.095 135.375 67.615 135.915 ;
        RECT 67.785 135.205 68.305 135.745 ;
        RECT 70.070 135.320 70.420 136.570 ;
        RECT 73.995 135.840 74.285 137.005 ;
        RECT 74.455 135.915 75.665 137.005 ;
        RECT 65.805 134.625 65.975 135.005 ;
        RECT 66.155 134.455 66.485 134.835 ;
        RECT 66.665 134.625 66.925 135.130 ;
        RECT 67.095 134.455 68.305 135.205 ;
        RECT 71.900 135.000 72.240 135.830 ;
        RECT 74.455 135.375 74.975 135.915 ;
        RECT 75.835 135.865 76.105 136.835 ;
        RECT 76.315 136.205 76.595 137.005 ;
        RECT 76.765 136.495 78.420 136.785 ;
        RECT 76.830 136.155 78.420 136.325 ;
        RECT 76.830 136.035 77.000 136.155 ;
        RECT 76.275 135.865 77.000 136.035 ;
        RECT 75.145 135.205 75.665 135.745 ;
        RECT 68.480 134.455 73.825 135.000 ;
        RECT 73.995 134.455 74.285 135.180 ;
        RECT 74.455 134.455 75.665 135.205 ;
        RECT 75.835 135.130 76.005 135.865 ;
        RECT 76.275 135.695 76.445 135.865 ;
        RECT 76.175 135.365 76.445 135.695 ;
        RECT 76.615 135.365 77.020 135.695 ;
        RECT 77.190 135.365 77.900 135.985 ;
        RECT 78.100 135.865 78.420 136.155 ;
        RECT 79.055 135.915 82.565 137.005 ;
        RECT 82.735 136.245 83.250 136.655 ;
        RECT 83.485 136.245 83.655 137.005 ;
        RECT 83.825 136.665 85.855 136.835 ;
        RECT 76.275 135.195 76.445 135.365 ;
        RECT 75.835 134.785 76.105 135.130 ;
        RECT 76.275 135.025 77.885 135.195 ;
        RECT 78.070 135.125 78.420 135.695 ;
        RECT 79.055 135.395 80.745 135.915 ;
        RECT 80.915 135.225 82.565 135.745 ;
        RECT 82.735 135.435 83.075 136.245 ;
        RECT 83.825 136.000 83.995 136.665 ;
        RECT 84.390 136.325 85.515 136.495 ;
        RECT 83.245 135.810 83.995 136.000 ;
        RECT 84.165 135.985 85.175 136.155 ;
        RECT 82.735 135.265 83.965 135.435 ;
        RECT 76.295 134.455 76.675 134.855 ;
        RECT 76.845 134.675 77.015 135.025 ;
        RECT 77.185 134.455 77.515 134.855 ;
        RECT 77.715 134.675 77.885 135.025 ;
        RECT 78.085 134.455 78.415 134.955 ;
        RECT 79.055 134.455 82.565 135.225 ;
        RECT 83.010 134.660 83.255 135.265 ;
        RECT 83.475 134.455 83.985 134.990 ;
        RECT 84.165 134.625 84.355 135.985 ;
        RECT 84.525 134.965 84.800 135.785 ;
        RECT 85.005 135.185 85.175 135.985 ;
        RECT 85.345 135.195 85.515 136.325 ;
        RECT 85.685 135.695 85.855 136.665 ;
        RECT 86.025 135.865 86.195 137.005 ;
        RECT 86.365 135.865 86.700 136.835 ;
        RECT 87.340 136.570 92.685 137.005 ;
        RECT 85.685 135.365 85.880 135.695 ;
        RECT 86.105 135.365 86.360 135.695 ;
        RECT 86.105 135.195 86.275 135.365 ;
        RECT 86.530 135.195 86.700 135.865 ;
        RECT 88.930 135.320 89.280 136.570 ;
        RECT 92.855 136.245 93.370 136.655 ;
        RECT 93.605 136.245 93.775 137.005 ;
        RECT 93.945 136.665 95.975 136.835 ;
        RECT 85.345 135.025 86.275 135.195 ;
        RECT 85.345 134.990 85.520 135.025 ;
        RECT 84.525 134.795 84.805 134.965 ;
        RECT 84.525 134.625 84.800 134.795 ;
        RECT 84.990 134.625 85.520 134.990 ;
        RECT 85.945 134.455 86.275 134.855 ;
        RECT 86.445 134.625 86.700 135.195 ;
        RECT 90.760 135.000 91.100 135.830 ;
        RECT 92.855 135.435 93.195 136.245 ;
        RECT 93.945 136.000 94.115 136.665 ;
        RECT 94.510 136.325 95.635 136.495 ;
        RECT 93.365 135.810 94.115 136.000 ;
        RECT 94.285 135.985 95.295 136.155 ;
        RECT 92.855 135.265 94.085 135.435 ;
        RECT 87.340 134.455 92.685 135.000 ;
        RECT 93.130 134.660 93.375 135.265 ;
        RECT 93.595 134.455 94.105 134.990 ;
        RECT 94.285 134.625 94.475 135.985 ;
        RECT 94.645 135.305 94.920 135.785 ;
        RECT 94.645 135.135 94.925 135.305 ;
        RECT 95.125 135.185 95.295 135.985 ;
        RECT 95.465 135.195 95.635 136.325 ;
        RECT 95.805 135.695 95.975 136.665 ;
        RECT 96.145 135.865 96.315 137.005 ;
        RECT 96.485 135.865 96.820 136.835 ;
        RECT 95.805 135.365 96.000 135.695 ;
        RECT 96.225 135.365 96.480 135.695 ;
        RECT 96.225 135.195 96.395 135.365 ;
        RECT 96.650 135.195 96.820 135.865 ;
        RECT 96.995 135.915 99.585 137.005 ;
        RECT 96.995 135.395 98.205 135.915 ;
        RECT 99.755 135.840 100.045 137.005 ;
        RECT 100.715 135.865 100.945 137.005 ;
        RECT 101.115 135.855 101.445 136.835 ;
        RECT 101.615 135.865 101.825 137.005 ;
        RECT 102.055 136.245 102.570 136.655 ;
        RECT 102.805 136.245 102.975 137.005 ;
        RECT 103.145 136.665 105.175 136.835 ;
        RECT 98.375 135.225 99.585 135.745 ;
        RECT 100.695 135.445 101.025 135.695 ;
        RECT 94.645 134.625 94.920 135.135 ;
        RECT 95.465 135.025 96.395 135.195 ;
        RECT 95.465 134.990 95.640 135.025 ;
        RECT 95.110 134.625 95.640 134.990 ;
        RECT 96.065 134.455 96.395 134.855 ;
        RECT 96.565 134.625 96.820 135.195 ;
        RECT 96.995 134.455 99.585 135.225 ;
        RECT 99.755 134.455 100.045 135.180 ;
        RECT 100.715 134.455 100.945 135.275 ;
        RECT 101.195 135.255 101.445 135.855 ;
        RECT 102.055 135.435 102.395 136.245 ;
        RECT 103.145 136.000 103.315 136.665 ;
        RECT 103.710 136.325 104.835 136.495 ;
        RECT 102.565 135.810 103.315 136.000 ;
        RECT 103.485 135.985 104.495 136.155 ;
        RECT 101.115 134.625 101.445 135.255 ;
        RECT 101.615 134.455 101.825 135.275 ;
        RECT 102.055 135.265 103.285 135.435 ;
        RECT 102.330 134.660 102.575 135.265 ;
        RECT 102.795 134.455 103.305 134.990 ;
        RECT 103.485 134.625 103.675 135.985 ;
        RECT 103.845 135.645 104.120 135.785 ;
        RECT 103.845 135.475 104.125 135.645 ;
        RECT 103.845 134.625 104.120 135.475 ;
        RECT 104.325 135.185 104.495 135.985 ;
        RECT 104.665 135.195 104.835 136.325 ;
        RECT 105.005 135.695 105.175 136.665 ;
        RECT 105.345 135.865 105.515 137.005 ;
        RECT 105.685 135.865 106.020 136.835 ;
        RECT 105.005 135.365 105.200 135.695 ;
        RECT 105.425 135.365 105.680 135.695 ;
        RECT 105.425 135.195 105.595 135.365 ;
        RECT 105.850 135.195 106.020 135.865 ;
        RECT 104.665 135.025 105.595 135.195 ;
        RECT 104.665 134.990 104.840 135.025 ;
        RECT 104.310 134.625 104.840 134.990 ;
        RECT 105.265 134.455 105.595 134.855 ;
        RECT 105.765 134.625 106.020 135.195 ;
        RECT 106.195 135.930 106.465 136.835 ;
        RECT 106.635 136.245 106.965 137.005 ;
        RECT 107.145 136.075 107.315 136.835 ;
        RECT 106.195 135.130 106.365 135.930 ;
        RECT 106.650 135.905 107.315 136.075 ;
        RECT 108.035 135.915 111.545 137.005 ;
        RECT 112.090 136.025 112.345 136.695 ;
        RECT 112.525 136.205 112.810 137.005 ;
        RECT 112.990 136.285 113.320 136.795 ;
        RECT 112.090 135.985 112.270 136.025 ;
        RECT 106.650 135.760 106.820 135.905 ;
        RECT 106.535 135.430 106.820 135.760 ;
        RECT 106.650 135.175 106.820 135.430 ;
        RECT 107.055 135.355 107.385 135.725 ;
        RECT 108.035 135.395 109.725 135.915 ;
        RECT 112.005 135.815 112.270 135.985 ;
        RECT 109.895 135.225 111.545 135.745 ;
        RECT 106.195 134.625 106.455 135.130 ;
        RECT 106.650 135.005 107.315 135.175 ;
        RECT 106.635 134.455 106.965 134.835 ;
        RECT 107.145 134.625 107.315 135.005 ;
        RECT 108.035 134.455 111.545 135.225 ;
        RECT 112.090 135.165 112.270 135.815 ;
        RECT 112.990 135.695 113.240 136.285 ;
        RECT 113.590 136.135 113.760 136.745 ;
        RECT 113.930 136.315 114.260 137.005 ;
        RECT 114.490 136.455 114.730 136.745 ;
        RECT 114.930 136.625 115.350 137.005 ;
        RECT 115.530 136.535 116.160 136.785 ;
        RECT 116.630 136.625 116.960 137.005 ;
        RECT 115.530 136.455 115.700 136.535 ;
        RECT 117.130 136.455 117.300 136.745 ;
        RECT 117.480 136.625 117.860 137.005 ;
        RECT 118.100 136.620 118.930 136.790 ;
        RECT 114.490 136.285 115.700 136.455 ;
        RECT 112.440 135.365 113.240 135.695 ;
        RECT 112.090 134.635 112.345 135.165 ;
        RECT 112.525 134.455 112.810 134.915 ;
        RECT 112.990 134.715 113.240 135.365 ;
        RECT 113.440 136.115 113.760 136.135 ;
        RECT 113.440 135.945 115.360 136.115 ;
        RECT 113.440 135.050 113.630 135.945 ;
        RECT 115.530 135.775 115.700 136.285 ;
        RECT 115.870 136.025 116.390 136.335 ;
        RECT 113.800 135.605 115.700 135.775 ;
        RECT 113.800 135.545 114.130 135.605 ;
        RECT 114.280 135.375 114.610 135.435 ;
        RECT 113.950 135.105 114.610 135.375 ;
        RECT 113.440 134.720 113.760 135.050 ;
        RECT 113.940 134.455 114.600 134.935 ;
        RECT 114.800 134.845 114.970 135.605 ;
        RECT 115.870 135.435 116.050 135.845 ;
        RECT 115.140 135.265 115.470 135.385 ;
        RECT 116.220 135.265 116.390 136.025 ;
        RECT 115.140 135.095 116.390 135.265 ;
        RECT 116.560 136.205 117.930 136.455 ;
        RECT 116.560 135.435 116.750 136.205 ;
        RECT 117.680 135.945 117.930 136.205 ;
        RECT 116.920 135.775 117.170 135.935 ;
        RECT 118.100 135.775 118.270 136.620 ;
        RECT 119.165 136.335 119.335 136.835 ;
        RECT 119.505 136.505 119.835 137.005 ;
        RECT 118.440 135.945 118.940 136.325 ;
        RECT 119.165 136.165 119.860 136.335 ;
        RECT 116.920 135.605 118.270 135.775 ;
        RECT 117.850 135.565 118.270 135.605 ;
        RECT 116.560 135.095 116.980 135.435 ;
        RECT 117.270 135.105 117.680 135.435 ;
        RECT 114.800 134.675 115.650 134.845 ;
        RECT 116.210 134.455 116.530 134.915 ;
        RECT 116.730 134.665 116.980 135.095 ;
        RECT 117.270 134.455 117.680 134.895 ;
        RECT 117.850 134.835 118.020 135.565 ;
        RECT 118.190 135.015 118.540 135.385 ;
        RECT 118.720 135.075 118.940 135.945 ;
        RECT 119.110 135.375 119.520 135.995 ;
        RECT 119.690 135.195 119.860 136.165 ;
        RECT 119.165 135.005 119.860 135.195 ;
        RECT 117.850 134.635 118.865 134.835 ;
        RECT 119.165 134.675 119.335 135.005 ;
        RECT 119.505 134.455 119.835 134.835 ;
        RECT 120.050 134.715 120.275 136.835 ;
        RECT 120.445 136.505 120.775 137.005 ;
        RECT 120.945 136.335 121.115 136.835 ;
        RECT 120.450 136.165 121.115 136.335 ;
        RECT 120.450 135.175 120.680 136.165 ;
        RECT 120.850 135.345 121.200 135.995 ;
        RECT 121.835 135.915 124.425 137.005 ;
        RECT 124.595 135.915 125.805 137.005 ;
        RECT 121.835 135.395 123.045 135.915 ;
        RECT 123.215 135.225 124.425 135.745 ;
        RECT 124.595 135.375 125.115 135.915 ;
        RECT 120.450 135.005 121.115 135.175 ;
        RECT 120.445 134.455 120.775 134.835 ;
        RECT 120.945 134.715 121.115 135.005 ;
        RECT 121.835 134.455 124.425 135.225 ;
        RECT 125.285 135.205 125.805 135.745 ;
        RECT 124.595 134.455 125.805 135.205 ;
        RECT 11.810 134.285 125.890 134.455 ;
        RECT 11.895 133.535 13.105 134.285 ;
        RECT 14.110 133.575 14.365 134.105 ;
        RECT 14.545 133.825 14.830 134.285 ;
        RECT 11.895 132.995 12.415 133.535 ;
        RECT 12.585 132.825 13.105 133.365 ;
        RECT 11.895 131.735 13.105 132.825 ;
        RECT 14.110 132.715 14.290 133.575 ;
        RECT 15.010 133.375 15.260 134.025 ;
        RECT 14.460 133.045 15.260 133.375 ;
        RECT 14.110 132.245 14.365 132.715 ;
        RECT 14.025 132.075 14.365 132.245 ;
        RECT 14.110 132.045 14.365 132.075 ;
        RECT 14.545 131.735 14.830 132.535 ;
        RECT 15.010 132.455 15.260 133.045 ;
        RECT 15.460 133.690 15.780 134.020 ;
        RECT 15.960 133.805 16.620 134.285 ;
        RECT 16.820 133.895 17.670 134.065 ;
        RECT 15.460 132.795 15.650 133.690 ;
        RECT 15.970 133.365 16.630 133.635 ;
        RECT 16.300 133.305 16.630 133.365 ;
        RECT 15.820 133.135 16.150 133.195 ;
        RECT 16.820 133.135 16.990 133.895 ;
        RECT 18.230 133.825 18.550 134.285 ;
        RECT 18.750 133.645 19.000 134.075 ;
        RECT 19.290 133.845 19.700 134.285 ;
        RECT 19.870 133.905 20.885 134.105 ;
        RECT 17.160 133.475 18.410 133.645 ;
        RECT 17.160 133.355 17.490 133.475 ;
        RECT 15.820 132.965 17.720 133.135 ;
        RECT 15.460 132.625 17.380 132.795 ;
        RECT 15.460 132.605 15.780 132.625 ;
        RECT 15.010 131.945 15.340 132.455 ;
        RECT 15.610 131.995 15.780 132.605 ;
        RECT 17.550 132.455 17.720 132.965 ;
        RECT 17.890 132.895 18.070 133.305 ;
        RECT 18.240 132.715 18.410 133.475 ;
        RECT 15.950 131.735 16.280 132.425 ;
        RECT 16.510 132.285 17.720 132.455 ;
        RECT 17.890 132.405 18.410 132.715 ;
        RECT 18.580 133.305 19.000 133.645 ;
        RECT 19.290 133.305 19.700 133.635 ;
        RECT 18.580 132.535 18.770 133.305 ;
        RECT 19.870 133.175 20.040 133.905 ;
        RECT 21.185 133.735 21.355 134.065 ;
        RECT 21.525 133.905 21.855 134.285 ;
        RECT 20.210 133.355 20.560 133.725 ;
        RECT 19.870 133.135 20.290 133.175 ;
        RECT 18.940 132.965 20.290 133.135 ;
        RECT 18.940 132.805 19.190 132.965 ;
        RECT 19.700 132.535 19.950 132.795 ;
        RECT 18.580 132.285 19.950 132.535 ;
        RECT 16.510 131.995 16.750 132.285 ;
        RECT 17.550 132.205 17.720 132.285 ;
        RECT 16.950 131.735 17.370 132.115 ;
        RECT 17.550 131.955 18.180 132.205 ;
        RECT 18.650 131.735 18.980 132.115 ;
        RECT 19.150 131.995 19.320 132.285 ;
        RECT 20.120 132.120 20.290 132.965 ;
        RECT 20.740 132.795 20.960 133.665 ;
        RECT 21.185 133.545 21.880 133.735 ;
        RECT 20.460 132.415 20.960 132.795 ;
        RECT 21.130 132.745 21.540 133.365 ;
        RECT 21.710 132.575 21.880 133.545 ;
        RECT 21.185 132.405 21.880 132.575 ;
        RECT 19.500 131.735 19.880 132.115 ;
        RECT 20.120 131.950 20.950 132.120 ;
        RECT 21.185 131.905 21.355 132.405 ;
        RECT 21.525 131.735 21.855 132.235 ;
        RECT 22.070 131.905 22.295 134.025 ;
        RECT 22.465 133.905 22.795 134.285 ;
        RECT 22.965 133.735 23.135 134.025 ;
        RECT 22.470 133.565 23.135 133.735 ;
        RECT 23.395 133.610 23.655 134.115 ;
        RECT 23.835 133.905 24.165 134.285 ;
        RECT 24.345 133.735 24.515 134.115 ;
        RECT 22.470 132.575 22.700 133.565 ;
        RECT 22.870 132.745 23.220 133.395 ;
        RECT 23.395 132.810 23.565 133.610 ;
        RECT 23.850 133.565 24.515 133.735 ;
        RECT 23.850 133.310 24.020 133.565 ;
        RECT 25.695 133.515 29.205 134.285 ;
        RECT 23.735 132.980 24.020 133.310 ;
        RECT 24.255 133.015 24.585 133.385 ;
        RECT 23.850 132.835 24.020 132.980 ;
        RECT 22.470 132.405 23.135 132.575 ;
        RECT 22.465 131.735 22.795 132.235 ;
        RECT 22.965 131.905 23.135 132.405 ;
        RECT 23.395 131.905 23.665 132.810 ;
        RECT 23.850 132.665 24.515 132.835 ;
        RECT 23.835 131.735 24.165 132.495 ;
        RECT 24.345 131.905 24.515 132.665 ;
        RECT 25.695 132.825 27.385 133.345 ;
        RECT 27.555 132.995 29.205 133.515 ;
        RECT 29.415 133.465 29.645 134.285 ;
        RECT 29.815 133.485 30.145 134.115 ;
        RECT 29.395 133.045 29.725 133.295 ;
        RECT 29.895 132.885 30.145 133.485 ;
        RECT 30.315 133.465 30.525 134.285 ;
        RECT 30.795 133.465 31.025 134.285 ;
        RECT 31.195 133.485 31.525 134.115 ;
        RECT 30.775 133.045 31.105 133.295 ;
        RECT 31.275 132.885 31.525 133.485 ;
        RECT 31.695 133.465 31.905 134.285 ;
        RECT 32.595 133.515 35.185 134.285 ;
        RECT 35.355 133.560 35.645 134.285 ;
        RECT 35.820 133.740 41.165 134.285 ;
        RECT 25.695 131.735 29.205 132.825 ;
        RECT 29.415 131.735 29.645 132.875 ;
        RECT 29.815 131.905 30.145 132.885 ;
        RECT 30.315 131.735 30.525 132.875 ;
        RECT 30.795 131.735 31.025 132.875 ;
        RECT 31.195 131.905 31.525 132.885 ;
        RECT 31.695 131.735 31.905 132.875 ;
        RECT 32.595 132.825 33.805 133.345 ;
        RECT 33.975 132.995 35.185 133.515 ;
        RECT 32.595 131.735 35.185 132.825 ;
        RECT 35.355 131.735 35.645 132.900 ;
        RECT 37.410 132.170 37.760 133.420 ;
        RECT 39.240 132.910 39.580 133.740 ;
        RECT 41.535 133.655 41.865 134.015 ;
        RECT 42.485 133.825 42.735 134.285 ;
        RECT 42.905 133.825 43.465 134.115 ;
        RECT 41.535 133.465 42.925 133.655 ;
        RECT 42.755 133.375 42.925 133.465 ;
        RECT 41.350 133.045 42.025 133.295 ;
        RECT 42.245 133.045 42.585 133.295 ;
        RECT 42.755 133.045 43.045 133.375 ;
        RECT 41.350 132.685 41.615 133.045 ;
        RECT 42.755 132.795 42.925 133.045 ;
        RECT 41.985 132.625 42.925 132.795 ;
        RECT 35.820 131.735 41.165 132.170 ;
        RECT 41.535 131.735 41.815 132.405 ;
        RECT 41.985 132.075 42.285 132.625 ;
        RECT 43.215 132.455 43.465 133.825 ;
        RECT 42.485 131.735 42.815 132.455 ;
        RECT 43.005 131.905 43.465 132.455 ;
        RECT 43.635 133.610 43.905 133.955 ;
        RECT 44.095 133.885 44.475 134.285 ;
        RECT 44.645 133.715 44.815 134.065 ;
        RECT 44.985 133.885 45.315 134.285 ;
        RECT 45.515 133.715 45.685 134.065 ;
        RECT 45.885 133.785 46.215 134.285 ;
        RECT 43.635 132.875 43.805 133.610 ;
        RECT 44.075 133.545 45.685 133.715 ;
        RECT 44.075 133.375 44.245 133.545 ;
        RECT 43.975 133.045 44.245 133.375 ;
        RECT 44.415 133.045 44.820 133.375 ;
        RECT 44.075 132.875 44.245 133.045 ;
        RECT 44.990 132.925 45.700 133.375 ;
        RECT 45.870 133.045 46.220 133.615 ;
        RECT 46.395 133.515 48.065 134.285 ;
        RECT 43.635 131.905 43.905 132.875 ;
        RECT 44.075 132.705 44.800 132.875 ;
        RECT 44.990 132.755 45.705 132.925 ;
        RECT 44.630 132.585 44.800 132.705 ;
        RECT 45.900 132.585 46.220 132.875 ;
        RECT 44.115 131.735 44.395 132.535 ;
        RECT 44.630 132.415 46.220 132.585 ;
        RECT 46.395 132.825 47.145 133.345 ;
        RECT 47.315 132.995 48.065 133.515 ;
        RECT 48.235 133.485 48.575 134.115 ;
        RECT 48.745 133.485 48.995 134.285 ;
        RECT 49.185 133.635 49.515 134.115 ;
        RECT 49.685 133.825 49.910 134.285 ;
        RECT 50.080 133.635 50.410 134.115 ;
        RECT 48.235 133.435 48.465 133.485 ;
        RECT 49.185 133.465 50.410 133.635 ;
        RECT 51.040 133.505 51.540 134.115 ;
        RECT 51.915 133.535 53.125 134.285 ;
        RECT 48.235 132.875 48.410 133.435 ;
        RECT 48.580 133.125 49.275 133.295 ;
        RECT 49.105 132.875 49.275 133.125 ;
        RECT 49.450 133.095 49.870 133.295 ;
        RECT 50.040 133.095 50.370 133.295 ;
        RECT 50.540 133.095 50.870 133.295 ;
        RECT 51.040 132.875 51.210 133.505 ;
        RECT 51.395 133.045 51.745 133.295 ;
        RECT 44.565 131.955 46.220 132.245 ;
        RECT 46.395 131.735 48.065 132.825 ;
        RECT 48.235 131.905 48.575 132.875 ;
        RECT 48.745 131.735 48.915 132.875 ;
        RECT 49.105 132.705 51.540 132.875 ;
        RECT 49.185 131.735 49.435 132.535 ;
        RECT 50.080 131.905 50.410 132.705 ;
        RECT 50.710 131.735 51.040 132.535 ;
        RECT 51.210 131.905 51.540 132.705 ;
        RECT 51.915 132.825 52.435 133.365 ;
        RECT 52.605 132.995 53.125 133.535 ;
        RECT 53.570 133.475 53.815 134.080 ;
        RECT 54.035 133.750 54.545 134.285 ;
        RECT 53.295 133.305 54.525 133.475 ;
        RECT 51.915 131.735 53.125 132.825 ;
        RECT 53.295 132.495 53.635 133.305 ;
        RECT 53.805 132.740 54.555 132.930 ;
        RECT 53.295 132.085 53.810 132.495 ;
        RECT 54.045 131.735 54.215 132.495 ;
        RECT 54.385 132.075 54.555 132.740 ;
        RECT 54.725 132.755 54.915 134.115 ;
        RECT 55.085 133.945 55.360 134.115 ;
        RECT 55.085 133.775 55.365 133.945 ;
        RECT 55.085 132.955 55.360 133.775 ;
        RECT 55.550 133.750 56.080 134.115 ;
        RECT 56.505 133.885 56.835 134.285 ;
        RECT 55.905 133.715 56.080 133.750 ;
        RECT 55.565 132.755 55.735 133.555 ;
        RECT 54.725 132.585 55.735 132.755 ;
        RECT 55.905 133.545 56.835 133.715 ;
        RECT 57.005 133.545 57.260 134.115 ;
        RECT 57.985 133.735 58.155 134.115 ;
        RECT 58.335 133.905 58.665 134.285 ;
        RECT 57.985 133.565 58.650 133.735 ;
        RECT 58.845 133.610 59.105 134.115 ;
        RECT 55.905 132.415 56.075 133.545 ;
        RECT 56.665 133.375 56.835 133.545 ;
        RECT 54.950 132.245 56.075 132.415 ;
        RECT 56.245 133.045 56.440 133.375 ;
        RECT 56.665 133.045 56.920 133.375 ;
        RECT 56.245 132.075 56.415 133.045 ;
        RECT 57.090 132.875 57.260 133.545 ;
        RECT 57.915 133.015 58.245 133.385 ;
        RECT 58.480 133.310 58.650 133.565 ;
        RECT 54.385 131.905 56.415 132.075 ;
        RECT 56.585 131.735 56.755 132.875 ;
        RECT 56.925 131.905 57.260 132.875 ;
        RECT 58.480 132.980 58.765 133.310 ;
        RECT 58.480 132.835 58.650 132.980 ;
        RECT 57.985 132.665 58.650 132.835 ;
        RECT 58.935 132.810 59.105 133.610 ;
        RECT 59.275 133.515 60.945 134.285 ;
        RECT 61.115 133.560 61.405 134.285 ;
        RECT 61.950 133.945 62.205 134.105 ;
        RECT 61.865 133.775 62.205 133.945 ;
        RECT 62.385 133.825 62.670 134.285 ;
        RECT 61.950 133.575 62.205 133.775 ;
        RECT 57.985 131.905 58.155 132.665 ;
        RECT 58.335 131.735 58.665 132.495 ;
        RECT 58.835 131.905 59.105 132.810 ;
        RECT 59.275 132.825 60.025 133.345 ;
        RECT 60.195 132.995 60.945 133.515 ;
        RECT 59.275 131.735 60.945 132.825 ;
        RECT 61.115 131.735 61.405 132.900 ;
        RECT 61.950 132.715 62.130 133.575 ;
        RECT 62.850 133.375 63.100 134.025 ;
        RECT 62.300 133.045 63.100 133.375 ;
        RECT 61.950 132.045 62.205 132.715 ;
        RECT 62.385 131.735 62.670 132.535 ;
        RECT 62.850 132.455 63.100 133.045 ;
        RECT 63.300 133.690 63.620 134.020 ;
        RECT 63.800 133.805 64.460 134.285 ;
        RECT 64.660 133.895 65.510 134.065 ;
        RECT 63.300 132.795 63.490 133.690 ;
        RECT 63.810 133.365 64.470 133.635 ;
        RECT 64.140 133.305 64.470 133.365 ;
        RECT 63.660 133.135 63.990 133.195 ;
        RECT 64.660 133.135 64.830 133.895 ;
        RECT 66.070 133.825 66.390 134.285 ;
        RECT 66.590 133.645 66.840 134.075 ;
        RECT 67.130 133.845 67.540 134.285 ;
        RECT 67.710 133.905 68.725 134.105 ;
        RECT 65.000 133.475 66.250 133.645 ;
        RECT 65.000 133.355 65.330 133.475 ;
        RECT 63.660 132.965 65.560 133.135 ;
        RECT 63.300 132.625 65.220 132.795 ;
        RECT 63.300 132.605 63.620 132.625 ;
        RECT 62.850 131.945 63.180 132.455 ;
        RECT 63.450 131.995 63.620 132.605 ;
        RECT 65.390 132.455 65.560 132.965 ;
        RECT 65.730 132.895 65.910 133.305 ;
        RECT 66.080 132.715 66.250 133.475 ;
        RECT 63.790 131.735 64.120 132.425 ;
        RECT 64.350 132.285 65.560 132.455 ;
        RECT 65.730 132.405 66.250 132.715 ;
        RECT 66.420 133.305 66.840 133.645 ;
        RECT 67.130 133.305 67.540 133.635 ;
        RECT 66.420 132.535 66.610 133.305 ;
        RECT 67.710 133.175 67.880 133.905 ;
        RECT 69.025 133.735 69.195 134.065 ;
        RECT 69.365 133.905 69.695 134.285 ;
        RECT 68.050 133.355 68.400 133.725 ;
        RECT 67.710 133.135 68.130 133.175 ;
        RECT 66.780 132.965 68.130 133.135 ;
        RECT 66.780 132.805 67.030 132.965 ;
        RECT 67.540 132.535 67.790 132.795 ;
        RECT 66.420 132.285 67.790 132.535 ;
        RECT 64.350 131.995 64.590 132.285 ;
        RECT 65.390 132.205 65.560 132.285 ;
        RECT 64.790 131.735 65.210 132.115 ;
        RECT 65.390 131.955 66.020 132.205 ;
        RECT 66.490 131.735 66.820 132.115 ;
        RECT 66.990 131.995 67.160 132.285 ;
        RECT 67.960 132.120 68.130 132.965 ;
        RECT 68.580 132.795 68.800 133.665 ;
        RECT 69.025 133.545 69.720 133.735 ;
        RECT 68.300 132.415 68.800 132.795 ;
        RECT 68.970 132.745 69.380 133.365 ;
        RECT 69.550 132.575 69.720 133.545 ;
        RECT 69.025 132.405 69.720 132.575 ;
        RECT 67.340 131.735 67.720 132.115 ;
        RECT 67.960 131.950 68.790 132.120 ;
        RECT 69.025 131.905 69.195 132.405 ;
        RECT 69.365 131.735 69.695 132.235 ;
        RECT 69.910 131.905 70.135 134.025 ;
        RECT 70.305 133.905 70.635 134.285 ;
        RECT 70.805 133.735 70.975 134.025 ;
        RECT 72.160 133.740 77.505 134.285 ;
        RECT 70.310 133.565 70.975 133.735 ;
        RECT 70.310 132.575 70.540 133.565 ;
        RECT 70.710 132.745 71.060 133.395 ;
        RECT 70.310 132.405 70.975 132.575 ;
        RECT 70.305 131.735 70.635 132.235 ;
        RECT 70.805 131.905 70.975 132.405 ;
        RECT 73.750 132.170 74.100 133.420 ;
        RECT 75.580 132.910 75.920 133.740 ;
        RECT 77.675 133.485 78.015 134.115 ;
        RECT 78.185 133.485 78.435 134.285 ;
        RECT 78.625 133.635 78.955 134.115 ;
        RECT 79.125 133.825 79.350 134.285 ;
        RECT 79.520 133.635 79.850 134.115 ;
        RECT 77.675 132.875 77.850 133.485 ;
        RECT 78.625 133.465 79.850 133.635 ;
        RECT 80.480 133.505 80.980 134.115 ;
        RECT 81.355 133.535 82.565 134.285 ;
        RECT 78.020 133.125 78.715 133.295 ;
        RECT 78.545 132.875 78.715 133.125 ;
        RECT 78.890 133.095 79.310 133.295 ;
        RECT 79.480 133.095 79.810 133.295 ;
        RECT 79.980 133.095 80.310 133.295 ;
        RECT 80.480 132.875 80.650 133.505 ;
        RECT 80.835 133.045 81.185 133.295 ;
        RECT 72.160 131.735 77.505 132.170 ;
        RECT 77.675 131.905 78.015 132.875 ;
        RECT 78.185 131.735 78.355 132.875 ;
        RECT 78.545 132.705 80.980 132.875 ;
        RECT 78.625 131.735 78.875 132.535 ;
        RECT 79.520 131.905 79.850 132.705 ;
        RECT 80.150 131.735 80.480 132.535 ;
        RECT 80.650 131.905 80.980 132.705 ;
        RECT 81.355 132.825 81.875 133.365 ;
        RECT 82.045 132.995 82.565 133.535 ;
        RECT 83.010 133.475 83.255 134.080 ;
        RECT 83.475 133.750 83.985 134.285 ;
        RECT 82.735 133.305 83.965 133.475 ;
        RECT 81.355 131.735 82.565 132.825 ;
        RECT 82.735 132.495 83.075 133.305 ;
        RECT 83.245 132.740 83.995 132.930 ;
        RECT 82.735 132.085 83.250 132.495 ;
        RECT 83.485 131.735 83.655 132.495 ;
        RECT 83.825 132.075 83.995 132.740 ;
        RECT 84.165 132.755 84.355 134.115 ;
        RECT 84.525 133.265 84.800 134.115 ;
        RECT 84.990 133.750 85.520 134.115 ;
        RECT 85.945 133.885 86.275 134.285 ;
        RECT 85.345 133.715 85.520 133.750 ;
        RECT 84.525 133.095 84.805 133.265 ;
        RECT 84.525 132.955 84.800 133.095 ;
        RECT 85.005 132.755 85.175 133.555 ;
        RECT 84.165 132.585 85.175 132.755 ;
        RECT 85.345 133.545 86.275 133.715 ;
        RECT 86.445 133.545 86.700 134.115 ;
        RECT 86.875 133.560 87.165 134.285 ;
        RECT 87.425 133.735 87.595 134.115 ;
        RECT 87.775 133.905 88.105 134.285 ;
        RECT 87.425 133.565 88.090 133.735 ;
        RECT 88.285 133.610 88.545 134.115 ;
        RECT 85.345 132.415 85.515 133.545 ;
        RECT 86.105 133.375 86.275 133.545 ;
        RECT 84.390 132.245 85.515 132.415 ;
        RECT 85.685 133.045 85.880 133.375 ;
        RECT 86.105 133.045 86.360 133.375 ;
        RECT 85.685 132.075 85.855 133.045 ;
        RECT 86.530 132.875 86.700 133.545 ;
        RECT 87.355 133.015 87.685 133.385 ;
        RECT 87.920 133.310 88.090 133.565 ;
        RECT 87.920 132.980 88.205 133.310 ;
        RECT 83.825 131.905 85.855 132.075 ;
        RECT 86.025 131.735 86.195 132.875 ;
        RECT 86.365 131.905 86.700 132.875 ;
        RECT 86.875 131.735 87.165 132.900 ;
        RECT 87.920 132.835 88.090 132.980 ;
        RECT 87.425 132.665 88.090 132.835 ;
        RECT 88.375 132.810 88.545 133.610 ;
        RECT 89.090 133.575 89.345 134.105 ;
        RECT 89.525 133.825 89.810 134.285 ;
        RECT 89.090 132.925 89.270 133.575 ;
        RECT 89.990 133.375 90.240 134.025 ;
        RECT 89.440 133.045 90.240 133.375 ;
        RECT 87.425 131.905 87.595 132.665 ;
        RECT 87.775 131.735 88.105 132.495 ;
        RECT 88.275 131.905 88.545 132.810 ;
        RECT 89.005 132.755 89.270 132.925 ;
        RECT 89.090 132.715 89.270 132.755 ;
        RECT 89.090 132.045 89.345 132.715 ;
        RECT 89.525 131.735 89.810 132.535 ;
        RECT 89.990 132.455 90.240 133.045 ;
        RECT 90.440 133.690 90.760 134.020 ;
        RECT 90.940 133.805 91.600 134.285 ;
        RECT 91.800 133.895 92.650 134.065 ;
        RECT 90.440 132.795 90.630 133.690 ;
        RECT 90.950 133.365 91.610 133.635 ;
        RECT 91.280 133.305 91.610 133.365 ;
        RECT 90.800 133.135 91.130 133.195 ;
        RECT 91.800 133.135 91.970 133.895 ;
        RECT 93.210 133.825 93.530 134.285 ;
        RECT 93.730 133.645 93.980 134.075 ;
        RECT 94.270 133.845 94.680 134.285 ;
        RECT 94.850 133.905 95.865 134.105 ;
        RECT 92.140 133.475 93.390 133.645 ;
        RECT 92.140 133.355 92.470 133.475 ;
        RECT 90.800 132.965 92.700 133.135 ;
        RECT 90.440 132.625 92.360 132.795 ;
        RECT 90.440 132.605 90.760 132.625 ;
        RECT 89.990 131.945 90.320 132.455 ;
        RECT 90.590 131.995 90.760 132.605 ;
        RECT 92.530 132.455 92.700 132.965 ;
        RECT 92.870 132.895 93.050 133.305 ;
        RECT 93.220 132.715 93.390 133.475 ;
        RECT 90.930 131.735 91.260 132.425 ;
        RECT 91.490 132.285 92.700 132.455 ;
        RECT 92.870 132.405 93.390 132.715 ;
        RECT 93.560 133.305 93.980 133.645 ;
        RECT 94.270 133.305 94.680 133.635 ;
        RECT 93.560 132.535 93.750 133.305 ;
        RECT 94.850 133.175 95.020 133.905 ;
        RECT 96.165 133.735 96.335 134.065 ;
        RECT 96.505 133.905 96.835 134.285 ;
        RECT 95.190 133.355 95.540 133.725 ;
        RECT 94.850 133.135 95.270 133.175 ;
        RECT 93.920 132.965 95.270 133.135 ;
        RECT 93.920 132.805 94.170 132.965 ;
        RECT 94.680 132.535 94.930 132.795 ;
        RECT 93.560 132.285 94.930 132.535 ;
        RECT 91.490 131.995 91.730 132.285 ;
        RECT 92.530 132.205 92.700 132.285 ;
        RECT 91.930 131.735 92.350 132.115 ;
        RECT 92.530 131.955 93.160 132.205 ;
        RECT 93.630 131.735 93.960 132.115 ;
        RECT 94.130 131.995 94.300 132.285 ;
        RECT 95.100 132.120 95.270 132.965 ;
        RECT 95.720 132.795 95.940 133.665 ;
        RECT 96.165 133.545 96.860 133.735 ;
        RECT 95.440 132.415 95.940 132.795 ;
        RECT 96.110 132.745 96.520 133.365 ;
        RECT 96.690 132.575 96.860 133.545 ;
        RECT 96.165 132.405 96.860 132.575 ;
        RECT 94.480 131.735 94.860 132.115 ;
        RECT 95.100 131.950 95.930 132.120 ;
        RECT 96.165 131.905 96.335 132.405 ;
        RECT 96.505 131.735 96.835 132.235 ;
        RECT 97.050 131.905 97.275 134.025 ;
        RECT 97.445 133.905 97.775 134.285 ;
        RECT 97.945 133.735 98.115 134.025 ;
        RECT 98.750 133.945 99.005 134.105 ;
        RECT 98.665 133.775 99.005 133.945 ;
        RECT 99.185 133.825 99.470 134.285 ;
        RECT 97.450 133.565 98.115 133.735 ;
        RECT 98.750 133.575 99.005 133.775 ;
        RECT 97.450 132.575 97.680 133.565 ;
        RECT 97.850 132.745 98.200 133.395 ;
        RECT 98.750 132.715 98.930 133.575 ;
        RECT 99.650 133.375 99.900 134.025 ;
        RECT 99.100 133.045 99.900 133.375 ;
        RECT 97.450 132.405 98.115 132.575 ;
        RECT 97.445 131.735 97.775 132.235 ;
        RECT 97.945 131.905 98.115 132.405 ;
        RECT 98.750 132.045 99.005 132.715 ;
        RECT 99.185 131.735 99.470 132.535 ;
        RECT 99.650 132.455 99.900 133.045 ;
        RECT 100.100 133.690 100.420 134.020 ;
        RECT 100.600 133.805 101.260 134.285 ;
        RECT 101.460 133.895 102.310 134.065 ;
        RECT 100.100 132.795 100.290 133.690 ;
        RECT 100.610 133.365 101.270 133.635 ;
        RECT 100.940 133.305 101.270 133.365 ;
        RECT 100.460 133.135 100.790 133.195 ;
        RECT 101.460 133.135 101.630 133.895 ;
        RECT 102.870 133.825 103.190 134.285 ;
        RECT 103.390 133.645 103.640 134.075 ;
        RECT 103.930 133.845 104.340 134.285 ;
        RECT 104.510 133.905 105.525 134.105 ;
        RECT 101.800 133.475 103.050 133.645 ;
        RECT 101.800 133.355 102.130 133.475 ;
        RECT 100.460 132.965 102.360 133.135 ;
        RECT 100.100 132.625 102.020 132.795 ;
        RECT 100.100 132.605 100.420 132.625 ;
        RECT 99.650 131.945 99.980 132.455 ;
        RECT 100.250 131.995 100.420 132.605 ;
        RECT 102.190 132.455 102.360 132.965 ;
        RECT 102.530 132.895 102.710 133.305 ;
        RECT 102.880 132.715 103.050 133.475 ;
        RECT 100.590 131.735 100.920 132.425 ;
        RECT 101.150 132.285 102.360 132.455 ;
        RECT 102.530 132.405 103.050 132.715 ;
        RECT 103.220 133.305 103.640 133.645 ;
        RECT 103.930 133.305 104.340 133.635 ;
        RECT 103.220 132.535 103.410 133.305 ;
        RECT 104.510 133.175 104.680 133.905 ;
        RECT 105.825 133.735 105.995 134.065 ;
        RECT 106.165 133.905 106.495 134.285 ;
        RECT 104.850 133.355 105.200 133.725 ;
        RECT 104.510 133.135 104.930 133.175 ;
        RECT 103.580 132.965 104.930 133.135 ;
        RECT 103.580 132.805 103.830 132.965 ;
        RECT 104.340 132.535 104.590 132.795 ;
        RECT 103.220 132.285 104.590 132.535 ;
        RECT 101.150 131.995 101.390 132.285 ;
        RECT 102.190 132.205 102.360 132.285 ;
        RECT 101.590 131.735 102.010 132.115 ;
        RECT 102.190 131.955 102.820 132.205 ;
        RECT 103.290 131.735 103.620 132.115 ;
        RECT 103.790 131.995 103.960 132.285 ;
        RECT 104.760 132.120 104.930 132.965 ;
        RECT 105.380 132.795 105.600 133.665 ;
        RECT 105.825 133.545 106.520 133.735 ;
        RECT 105.100 132.415 105.600 132.795 ;
        RECT 105.770 132.745 106.180 133.365 ;
        RECT 106.350 132.575 106.520 133.545 ;
        RECT 105.825 132.405 106.520 132.575 ;
        RECT 104.140 131.735 104.520 132.115 ;
        RECT 104.760 131.950 105.590 132.120 ;
        RECT 105.825 131.905 105.995 132.405 ;
        RECT 106.165 131.735 106.495 132.235 ;
        RECT 106.710 131.905 106.935 134.025 ;
        RECT 107.105 133.905 107.435 134.285 ;
        RECT 107.605 133.735 107.775 134.025 ;
        RECT 107.110 133.565 107.775 133.735 ;
        RECT 108.035 133.825 108.595 134.115 ;
        RECT 108.765 133.825 109.015 134.285 ;
        RECT 107.110 132.575 107.340 133.565 ;
        RECT 107.510 132.745 107.860 133.395 ;
        RECT 107.110 132.405 107.775 132.575 ;
        RECT 107.105 131.735 107.435 132.235 ;
        RECT 107.605 131.905 107.775 132.405 ;
        RECT 108.035 132.455 108.285 133.825 ;
        RECT 109.635 133.655 109.965 134.015 ;
        RECT 108.575 133.465 109.965 133.655 ;
        RECT 110.795 133.515 112.465 134.285 ;
        RECT 112.635 133.560 112.925 134.285 ;
        RECT 113.555 133.515 117.065 134.285 ;
        RECT 117.325 133.735 117.495 134.115 ;
        RECT 117.675 133.905 118.005 134.285 ;
        RECT 117.325 133.565 117.990 133.735 ;
        RECT 118.185 133.610 118.445 134.115 ;
        RECT 119.080 133.740 124.425 134.285 ;
        RECT 108.575 133.375 108.745 133.465 ;
        RECT 108.455 133.045 108.745 133.375 ;
        RECT 108.915 133.045 109.255 133.295 ;
        RECT 109.475 133.045 110.150 133.295 ;
        RECT 108.575 132.795 108.745 133.045 ;
        RECT 108.575 132.625 109.515 132.795 ;
        RECT 109.885 132.685 110.150 133.045 ;
        RECT 110.795 132.825 111.545 133.345 ;
        RECT 111.715 132.995 112.465 133.515 ;
        RECT 108.035 131.905 108.495 132.455 ;
        RECT 108.685 131.735 109.015 132.455 ;
        RECT 109.215 132.075 109.515 132.625 ;
        RECT 109.685 131.735 109.965 132.405 ;
        RECT 110.795 131.735 112.465 132.825 ;
        RECT 112.635 131.735 112.925 132.900 ;
        RECT 113.555 132.825 115.245 133.345 ;
        RECT 115.415 132.995 117.065 133.515 ;
        RECT 117.255 133.015 117.585 133.385 ;
        RECT 117.820 133.310 117.990 133.565 ;
        RECT 117.820 132.980 118.105 133.310 ;
        RECT 117.820 132.835 117.990 132.980 ;
        RECT 113.555 131.735 117.065 132.825 ;
        RECT 117.325 132.665 117.990 132.835 ;
        RECT 118.275 132.810 118.445 133.610 ;
        RECT 117.325 131.905 117.495 132.665 ;
        RECT 117.675 131.735 118.005 132.495 ;
        RECT 118.175 131.905 118.445 132.810 ;
        RECT 120.670 132.170 121.020 133.420 ;
        RECT 122.500 132.910 122.840 133.740 ;
        RECT 124.595 133.535 125.805 134.285 ;
        RECT 124.595 132.825 125.115 133.365 ;
        RECT 125.285 132.995 125.805 133.535 ;
        RECT 119.080 131.735 124.425 132.170 ;
        RECT 124.595 131.735 125.805 132.825 ;
        RECT 11.810 131.565 125.890 131.735 ;
        RECT 11.895 130.475 13.105 131.565 ;
        RECT 11.895 129.765 12.415 130.305 ;
        RECT 12.585 129.935 13.105 130.475 ;
        RECT 13.275 130.475 16.785 131.565 ;
        RECT 13.275 129.955 14.965 130.475 ;
        RECT 16.995 130.425 17.225 131.565 ;
        RECT 17.395 130.415 17.725 131.395 ;
        RECT 17.895 130.425 18.105 131.565 ;
        RECT 18.335 130.805 18.850 131.215 ;
        RECT 19.085 130.805 19.255 131.565 ;
        RECT 19.425 131.225 21.455 131.395 ;
        RECT 15.135 129.785 16.785 130.305 ;
        RECT 16.975 130.005 17.305 130.255 ;
        RECT 11.895 129.015 13.105 129.765 ;
        RECT 13.275 129.015 16.785 129.785 ;
        RECT 16.995 129.015 17.225 129.835 ;
        RECT 17.475 129.815 17.725 130.415 ;
        RECT 18.335 129.995 18.675 130.805 ;
        RECT 19.425 130.560 19.595 131.225 ;
        RECT 19.990 130.885 21.115 131.055 ;
        RECT 18.845 130.370 19.595 130.560 ;
        RECT 19.765 130.545 20.775 130.715 ;
        RECT 17.395 129.185 17.725 129.815 ;
        RECT 17.895 129.015 18.105 129.835 ;
        RECT 18.335 129.825 19.565 129.995 ;
        RECT 18.610 129.220 18.855 129.825 ;
        RECT 19.075 129.015 19.585 129.550 ;
        RECT 19.765 129.185 19.955 130.545 ;
        RECT 20.125 129.865 20.400 130.345 ;
        RECT 20.125 129.695 20.405 129.865 ;
        RECT 20.605 129.745 20.775 130.545 ;
        RECT 20.945 129.755 21.115 130.885 ;
        RECT 21.285 130.255 21.455 131.225 ;
        RECT 21.625 130.425 21.795 131.565 ;
        RECT 21.965 130.425 22.300 131.395 ;
        RECT 21.285 129.925 21.480 130.255 ;
        RECT 21.705 129.925 21.960 130.255 ;
        RECT 21.705 129.755 21.875 129.925 ;
        RECT 22.130 129.755 22.300 130.425 ;
        RECT 22.475 130.400 22.765 131.565 ;
        RECT 22.935 130.475 26.445 131.565 ;
        RECT 26.705 130.895 26.875 131.395 ;
        RECT 27.045 131.065 27.375 131.565 ;
        RECT 26.705 130.725 27.370 130.895 ;
        RECT 22.935 129.955 24.625 130.475 ;
        RECT 24.795 129.785 26.445 130.305 ;
        RECT 26.620 129.905 26.970 130.555 ;
        RECT 20.125 129.185 20.400 129.695 ;
        RECT 20.945 129.585 21.875 129.755 ;
        RECT 20.945 129.550 21.120 129.585 ;
        RECT 20.590 129.185 21.120 129.550 ;
        RECT 21.545 129.015 21.875 129.415 ;
        RECT 22.045 129.185 22.300 129.755 ;
        RECT 22.475 129.015 22.765 129.740 ;
        RECT 22.935 129.015 26.445 129.785 ;
        RECT 27.140 129.735 27.370 130.725 ;
        RECT 26.705 129.565 27.370 129.735 ;
        RECT 26.705 129.275 26.875 129.565 ;
        RECT 27.045 129.015 27.375 129.395 ;
        RECT 27.545 129.275 27.770 131.395 ;
        RECT 27.985 131.065 28.315 131.565 ;
        RECT 28.485 130.895 28.655 131.395 ;
        RECT 28.890 131.180 29.720 131.350 ;
        RECT 29.960 131.185 30.340 131.565 ;
        RECT 27.960 130.725 28.655 130.895 ;
        RECT 27.960 129.755 28.130 130.725 ;
        RECT 28.300 129.935 28.710 130.555 ;
        RECT 28.880 130.505 29.380 130.885 ;
        RECT 27.960 129.565 28.655 129.755 ;
        RECT 28.880 129.635 29.100 130.505 ;
        RECT 29.550 130.335 29.720 131.180 ;
        RECT 30.520 131.015 30.690 131.305 ;
        RECT 30.860 131.185 31.190 131.565 ;
        RECT 31.660 131.095 32.290 131.345 ;
        RECT 32.470 131.185 32.890 131.565 ;
        RECT 32.120 131.015 32.290 131.095 ;
        RECT 33.090 131.015 33.330 131.305 ;
        RECT 29.890 130.765 31.260 131.015 ;
        RECT 29.890 130.505 30.140 130.765 ;
        RECT 30.650 130.335 30.900 130.495 ;
        RECT 29.550 130.165 30.900 130.335 ;
        RECT 29.550 130.125 29.970 130.165 ;
        RECT 29.280 129.575 29.630 129.945 ;
        RECT 27.985 129.015 28.315 129.395 ;
        RECT 28.485 129.235 28.655 129.565 ;
        RECT 29.800 129.395 29.970 130.125 ;
        RECT 31.070 129.995 31.260 130.765 ;
        RECT 30.140 129.665 30.550 129.995 ;
        RECT 30.840 129.655 31.260 129.995 ;
        RECT 31.430 130.585 31.950 130.895 ;
        RECT 32.120 130.845 33.330 131.015 ;
        RECT 33.560 130.875 33.890 131.565 ;
        RECT 31.430 129.825 31.600 130.585 ;
        RECT 31.770 129.995 31.950 130.405 ;
        RECT 32.120 130.335 32.290 130.845 ;
        RECT 34.060 130.695 34.230 131.305 ;
        RECT 34.500 130.845 34.830 131.355 ;
        RECT 34.060 130.675 34.380 130.695 ;
        RECT 32.460 130.505 34.380 130.675 ;
        RECT 32.120 130.165 34.020 130.335 ;
        RECT 32.350 129.825 32.680 129.945 ;
        RECT 31.430 129.655 32.680 129.825 ;
        RECT 28.955 129.195 29.970 129.395 ;
        RECT 30.140 129.015 30.550 129.455 ;
        RECT 30.840 129.225 31.090 129.655 ;
        RECT 31.290 129.015 31.610 129.475 ;
        RECT 32.850 129.405 33.020 130.165 ;
        RECT 33.690 130.105 34.020 130.165 ;
        RECT 33.210 129.935 33.540 129.995 ;
        RECT 33.210 129.665 33.870 129.935 ;
        RECT 34.190 129.610 34.380 130.505 ;
        RECT 32.170 129.235 33.020 129.405 ;
        RECT 33.220 129.015 33.880 129.495 ;
        RECT 34.060 129.280 34.380 129.610 ;
        RECT 34.580 130.255 34.830 130.845 ;
        RECT 35.010 130.765 35.295 131.565 ;
        RECT 35.475 131.225 35.730 131.255 ;
        RECT 35.475 131.055 35.815 131.225 ;
        RECT 35.475 130.585 35.730 131.055 ;
        RECT 36.790 130.695 37.075 131.565 ;
        RECT 37.245 130.935 37.505 131.395 ;
        RECT 37.680 131.105 37.935 131.565 ;
        RECT 38.105 130.935 38.365 131.395 ;
        RECT 37.245 130.765 38.365 130.935 ;
        RECT 38.535 130.765 38.845 131.565 ;
        RECT 34.580 129.925 35.380 130.255 ;
        RECT 34.580 129.275 34.830 129.925 ;
        RECT 35.550 129.725 35.730 130.585 ;
        RECT 37.245 130.515 37.505 130.765 ;
        RECT 39.015 130.595 39.325 131.395 ;
        RECT 39.695 130.895 39.975 131.565 ;
        RECT 40.145 130.675 40.445 131.225 ;
        RECT 40.645 130.845 40.975 131.565 ;
        RECT 41.165 130.845 41.625 131.395 ;
        RECT 41.800 131.055 43.455 131.345 ;
        RECT 35.010 129.015 35.295 129.475 ;
        RECT 35.475 129.195 35.730 129.725 ;
        RECT 36.750 130.345 37.505 130.515 ;
        RECT 38.295 130.425 39.325 130.595 ;
        RECT 36.750 129.835 37.155 130.345 ;
        RECT 38.295 130.175 38.465 130.425 ;
        RECT 37.325 130.005 38.465 130.175 ;
        RECT 36.750 129.665 38.400 129.835 ;
        RECT 38.635 129.685 38.985 130.255 ;
        RECT 36.795 129.015 37.075 129.495 ;
        RECT 37.245 129.275 37.505 129.665 ;
        RECT 37.680 129.015 37.935 129.495 ;
        RECT 38.105 129.275 38.400 129.665 ;
        RECT 39.155 129.515 39.325 130.425 ;
        RECT 39.510 130.255 39.775 130.615 ;
        RECT 40.145 130.505 41.085 130.675 ;
        RECT 40.915 130.255 41.085 130.505 ;
        RECT 39.510 130.005 40.185 130.255 ;
        RECT 40.405 130.005 40.745 130.255 ;
        RECT 40.915 129.925 41.205 130.255 ;
        RECT 40.915 129.835 41.085 129.925 ;
        RECT 38.580 129.015 38.855 129.495 ;
        RECT 39.025 129.185 39.325 129.515 ;
        RECT 39.695 129.645 41.085 129.835 ;
        RECT 39.695 129.285 40.025 129.645 ;
        RECT 41.375 129.475 41.625 130.845 ;
        RECT 41.800 130.715 43.390 130.885 ;
        RECT 43.625 130.765 43.905 131.565 ;
        RECT 41.800 130.425 42.120 130.715 ;
        RECT 43.220 130.595 43.390 130.715 ;
        RECT 42.315 130.375 43.030 130.545 ;
        RECT 43.220 130.425 43.945 130.595 ;
        RECT 44.115 130.425 44.385 131.395 ;
        RECT 41.800 129.685 42.150 130.255 ;
        RECT 42.320 129.925 43.030 130.375 ;
        RECT 43.775 130.255 43.945 130.425 ;
        RECT 43.200 129.925 43.605 130.255 ;
        RECT 43.775 129.925 44.045 130.255 ;
        RECT 43.775 129.755 43.945 129.925 ;
        RECT 42.335 129.585 43.945 129.755 ;
        RECT 44.215 129.690 44.385 130.425 ;
        RECT 40.645 129.015 40.895 129.475 ;
        RECT 41.065 129.185 41.625 129.475 ;
        RECT 41.805 129.015 42.135 129.515 ;
        RECT 42.335 129.235 42.505 129.585 ;
        RECT 42.705 129.015 43.035 129.415 ;
        RECT 43.205 129.235 43.375 129.585 ;
        RECT 43.545 129.015 43.925 129.415 ;
        RECT 44.115 129.345 44.385 129.690 ;
        RECT 44.555 130.425 44.895 131.395 ;
        RECT 45.065 130.425 45.235 131.565 ;
        RECT 45.505 130.765 45.755 131.565 ;
        RECT 46.400 130.595 46.730 131.395 ;
        RECT 47.030 130.765 47.360 131.565 ;
        RECT 47.530 130.595 47.860 131.395 ;
        RECT 45.425 130.425 47.860 130.595 ;
        RECT 44.555 129.815 44.730 130.425 ;
        RECT 45.425 130.175 45.595 130.425 ;
        RECT 44.900 130.005 45.595 130.175 ;
        RECT 45.770 130.005 46.190 130.205 ;
        RECT 46.360 130.005 46.690 130.205 ;
        RECT 46.860 130.005 47.190 130.205 ;
        RECT 44.555 129.185 44.895 129.815 ;
        RECT 45.065 129.015 45.315 129.815 ;
        RECT 45.505 129.665 46.730 129.835 ;
        RECT 45.505 129.185 45.835 129.665 ;
        RECT 46.005 129.015 46.230 129.475 ;
        RECT 46.400 129.185 46.730 129.665 ;
        RECT 47.360 129.795 47.530 130.425 ;
        RECT 48.235 130.400 48.525 131.565 ;
        RECT 49.155 130.475 51.745 131.565 ;
        RECT 52.290 130.585 52.545 131.255 ;
        RECT 52.725 130.765 53.010 131.565 ;
        RECT 53.190 130.845 53.520 131.355 ;
        RECT 47.715 130.005 48.065 130.255 ;
        RECT 49.155 129.955 50.365 130.475 ;
        RECT 47.360 129.185 47.860 129.795 ;
        RECT 50.535 129.785 51.745 130.305 ;
        RECT 48.235 129.015 48.525 129.740 ;
        RECT 49.155 129.015 51.745 129.785 ;
        RECT 52.290 129.725 52.470 130.585 ;
        RECT 53.190 130.255 53.440 130.845 ;
        RECT 53.790 130.695 53.960 131.305 ;
        RECT 54.130 130.875 54.460 131.565 ;
        RECT 54.690 131.015 54.930 131.305 ;
        RECT 55.130 131.185 55.550 131.565 ;
        RECT 55.730 131.095 56.360 131.345 ;
        RECT 56.830 131.185 57.160 131.565 ;
        RECT 55.730 131.015 55.900 131.095 ;
        RECT 57.330 131.015 57.500 131.305 ;
        RECT 57.680 131.185 58.060 131.565 ;
        RECT 58.300 131.180 59.130 131.350 ;
        RECT 54.690 130.845 55.900 131.015 ;
        RECT 52.640 129.925 53.440 130.255 ;
        RECT 52.290 129.525 52.545 129.725 ;
        RECT 52.205 129.355 52.545 129.525 ;
        RECT 52.290 129.195 52.545 129.355 ;
        RECT 52.725 129.015 53.010 129.475 ;
        RECT 53.190 129.275 53.440 129.925 ;
        RECT 53.640 130.675 53.960 130.695 ;
        RECT 53.640 130.505 55.560 130.675 ;
        RECT 53.640 129.610 53.830 130.505 ;
        RECT 55.730 130.335 55.900 130.845 ;
        RECT 56.070 130.585 56.590 130.895 ;
        RECT 54.000 130.165 55.900 130.335 ;
        RECT 54.000 130.105 54.330 130.165 ;
        RECT 54.480 129.935 54.810 129.995 ;
        RECT 54.150 129.665 54.810 129.935 ;
        RECT 53.640 129.280 53.960 129.610 ;
        RECT 54.140 129.015 54.800 129.495 ;
        RECT 55.000 129.405 55.170 130.165 ;
        RECT 56.070 129.995 56.250 130.405 ;
        RECT 55.340 129.825 55.670 129.945 ;
        RECT 56.420 129.825 56.590 130.585 ;
        RECT 55.340 129.655 56.590 129.825 ;
        RECT 56.760 130.765 58.130 131.015 ;
        RECT 56.760 129.995 56.950 130.765 ;
        RECT 57.880 130.505 58.130 130.765 ;
        RECT 57.120 130.335 57.370 130.495 ;
        RECT 58.300 130.335 58.470 131.180 ;
        RECT 59.365 130.895 59.535 131.395 ;
        RECT 59.705 131.065 60.035 131.565 ;
        RECT 58.640 130.505 59.140 130.885 ;
        RECT 59.365 130.725 60.060 130.895 ;
        RECT 57.120 130.165 58.470 130.335 ;
        RECT 58.050 130.125 58.470 130.165 ;
        RECT 56.760 129.655 57.180 129.995 ;
        RECT 57.470 129.665 57.880 129.995 ;
        RECT 55.000 129.235 55.850 129.405 ;
        RECT 56.410 129.015 56.730 129.475 ;
        RECT 56.930 129.225 57.180 129.655 ;
        RECT 57.470 129.015 57.880 129.455 ;
        RECT 58.050 129.395 58.220 130.125 ;
        RECT 58.390 129.575 58.740 129.945 ;
        RECT 58.920 129.635 59.140 130.505 ;
        RECT 59.310 129.935 59.720 130.555 ;
        RECT 59.890 129.755 60.060 130.725 ;
        RECT 59.365 129.565 60.060 129.755 ;
        RECT 58.050 129.195 59.065 129.395 ;
        RECT 59.365 129.235 59.535 129.565 ;
        RECT 59.705 129.015 60.035 129.395 ;
        RECT 60.250 129.275 60.475 131.395 ;
        RECT 60.645 131.065 60.975 131.565 ;
        RECT 61.145 130.895 61.315 131.395 ;
        RECT 60.650 130.725 61.315 130.895 ;
        RECT 60.650 129.735 60.880 130.725 ;
        RECT 61.050 129.905 61.400 130.555 ;
        RECT 61.575 130.475 64.165 131.565 ;
        RECT 61.575 129.955 62.785 130.475 ;
        RECT 64.375 130.425 64.605 131.565 ;
        RECT 64.775 130.415 65.105 131.395 ;
        RECT 65.275 130.425 65.485 131.565 ;
        RECT 66.725 130.635 66.895 131.395 ;
        RECT 67.075 130.805 67.405 131.565 ;
        RECT 66.725 130.465 67.390 130.635 ;
        RECT 67.575 130.490 67.845 131.395 ;
        RECT 68.020 131.140 68.355 131.565 ;
        RECT 68.525 130.960 68.710 131.365 ;
        RECT 62.955 129.785 64.165 130.305 ;
        RECT 64.355 130.005 64.685 130.255 ;
        RECT 60.650 129.565 61.315 129.735 ;
        RECT 60.645 129.015 60.975 129.395 ;
        RECT 61.145 129.275 61.315 129.565 ;
        RECT 61.575 129.015 64.165 129.785 ;
        RECT 64.375 129.015 64.605 129.835 ;
        RECT 64.855 129.815 65.105 130.415 ;
        RECT 67.220 130.320 67.390 130.465 ;
        RECT 66.655 129.915 66.985 130.285 ;
        RECT 67.220 129.990 67.505 130.320 ;
        RECT 64.775 129.185 65.105 129.815 ;
        RECT 65.275 129.015 65.485 129.835 ;
        RECT 67.220 129.735 67.390 129.990 ;
        RECT 66.725 129.565 67.390 129.735 ;
        RECT 67.675 129.690 67.845 130.490 ;
        RECT 66.725 129.185 66.895 129.565 ;
        RECT 67.075 129.015 67.405 129.395 ;
        RECT 67.585 129.185 67.845 129.690 ;
        RECT 68.045 130.785 68.710 130.960 ;
        RECT 68.915 130.785 69.245 131.565 ;
        RECT 68.045 129.755 68.385 130.785 ;
        RECT 69.415 130.595 69.685 131.365 ;
        RECT 68.555 130.425 69.685 130.595 ;
        RECT 68.555 129.925 68.805 130.425 ;
        RECT 68.045 129.585 68.730 129.755 ;
        RECT 68.985 129.675 69.345 130.255 ;
        RECT 68.020 129.015 68.355 129.415 ;
        RECT 68.525 129.185 68.730 129.585 ;
        RECT 69.515 129.515 69.685 130.425 ;
        RECT 68.940 129.015 69.215 129.495 ;
        RECT 69.425 129.185 69.685 129.515 ;
        RECT 69.855 130.595 70.125 131.365 ;
        RECT 70.295 130.785 70.625 131.565 ;
        RECT 70.830 130.960 71.015 131.365 ;
        RECT 71.185 131.140 71.520 131.565 ;
        RECT 70.830 130.785 71.495 130.960 ;
        RECT 71.895 130.895 72.175 131.565 ;
        RECT 69.855 130.425 70.985 130.595 ;
        RECT 69.855 129.515 70.025 130.425 ;
        RECT 70.195 129.675 70.555 130.255 ;
        RECT 70.735 129.925 70.985 130.425 ;
        RECT 71.155 129.755 71.495 130.785 ;
        RECT 72.345 130.675 72.645 131.225 ;
        RECT 72.845 130.845 73.175 131.565 ;
        RECT 73.365 130.845 73.825 131.395 ;
        RECT 71.710 130.255 71.975 130.615 ;
        RECT 72.345 130.505 73.285 130.675 ;
        RECT 73.115 130.255 73.285 130.505 ;
        RECT 71.710 130.005 72.385 130.255 ;
        RECT 72.605 130.005 72.945 130.255 ;
        RECT 73.115 129.925 73.405 130.255 ;
        RECT 73.115 129.835 73.285 129.925 ;
        RECT 70.810 129.585 71.495 129.755 ;
        RECT 71.895 129.645 73.285 129.835 ;
        RECT 69.855 129.185 70.115 129.515 ;
        RECT 70.325 129.015 70.600 129.495 ;
        RECT 70.810 129.185 71.015 129.585 ;
        RECT 71.185 129.015 71.520 129.415 ;
        RECT 71.895 129.285 72.225 129.645 ;
        RECT 73.575 129.475 73.825 130.845 ;
        RECT 73.995 130.400 74.285 131.565 ;
        RECT 74.455 130.475 75.665 131.565 ;
        RECT 75.840 131.055 77.495 131.345 ;
        RECT 75.840 130.715 77.430 130.885 ;
        RECT 77.665 130.765 77.945 131.565 ;
        RECT 74.455 129.935 74.975 130.475 ;
        RECT 75.840 130.425 76.160 130.715 ;
        RECT 77.260 130.595 77.430 130.715 ;
        RECT 75.145 129.765 75.665 130.305 ;
        RECT 72.845 129.015 73.095 129.475 ;
        RECT 73.265 129.185 73.825 129.475 ;
        RECT 73.995 129.015 74.285 129.740 ;
        RECT 74.455 129.015 75.665 129.765 ;
        RECT 75.840 129.685 76.190 130.255 ;
        RECT 76.360 129.925 77.070 130.545 ;
        RECT 77.260 130.425 77.985 130.595 ;
        RECT 78.155 130.425 78.425 131.395 ;
        RECT 77.815 130.255 77.985 130.425 ;
        RECT 77.240 129.925 77.645 130.255 ;
        RECT 77.815 129.925 78.085 130.255 ;
        RECT 77.815 129.755 77.985 129.925 ;
        RECT 76.375 129.585 77.985 129.755 ;
        RECT 78.255 129.690 78.425 130.425 ;
        RECT 75.845 129.015 76.175 129.515 ;
        RECT 76.375 129.235 76.545 129.585 ;
        RECT 76.745 129.015 77.075 129.415 ;
        RECT 77.245 129.235 77.415 129.585 ;
        RECT 77.585 129.015 77.965 129.415 ;
        RECT 78.155 129.345 78.425 129.690 ;
        RECT 78.595 130.425 78.935 131.395 ;
        RECT 79.105 130.425 79.275 131.565 ;
        RECT 79.545 130.765 79.795 131.565 ;
        RECT 80.440 130.595 80.770 131.395 ;
        RECT 81.070 130.765 81.400 131.565 ;
        RECT 81.570 130.595 81.900 131.395 ;
        RECT 83.570 131.225 83.825 131.255 ;
        RECT 83.485 131.055 83.825 131.225 ;
        RECT 79.465 130.425 81.900 130.595 ;
        RECT 83.570 130.585 83.825 131.055 ;
        RECT 84.005 130.765 84.290 131.565 ;
        RECT 84.470 130.845 84.800 131.355 ;
        RECT 78.595 129.815 78.770 130.425 ;
        RECT 79.465 130.175 79.635 130.425 ;
        RECT 78.940 130.005 79.635 130.175 ;
        RECT 79.810 130.005 80.230 130.205 ;
        RECT 80.400 130.005 80.730 130.205 ;
        RECT 80.900 130.005 81.230 130.205 ;
        RECT 78.595 129.185 78.935 129.815 ;
        RECT 79.105 129.015 79.355 129.815 ;
        RECT 79.545 129.665 80.770 129.835 ;
        RECT 79.545 129.185 79.875 129.665 ;
        RECT 80.045 129.015 80.270 129.475 ;
        RECT 80.440 129.185 80.770 129.665 ;
        RECT 81.400 129.795 81.570 130.425 ;
        RECT 81.755 130.005 82.105 130.255 ;
        RECT 81.400 129.185 81.900 129.795 ;
        RECT 83.570 129.725 83.750 130.585 ;
        RECT 84.470 130.255 84.720 130.845 ;
        RECT 85.070 130.695 85.240 131.305 ;
        RECT 85.410 130.875 85.740 131.565 ;
        RECT 85.970 131.015 86.210 131.305 ;
        RECT 86.410 131.185 86.830 131.565 ;
        RECT 87.010 131.095 87.640 131.345 ;
        RECT 88.110 131.185 88.440 131.565 ;
        RECT 87.010 131.015 87.180 131.095 ;
        RECT 88.610 131.015 88.780 131.305 ;
        RECT 88.960 131.185 89.340 131.565 ;
        RECT 89.580 131.180 90.410 131.350 ;
        RECT 85.970 130.845 87.180 131.015 ;
        RECT 83.920 129.925 84.720 130.255 ;
        RECT 83.570 129.195 83.825 129.725 ;
        RECT 84.005 129.015 84.290 129.475 ;
        RECT 84.470 129.275 84.720 129.925 ;
        RECT 84.920 130.675 85.240 130.695 ;
        RECT 84.920 130.505 86.840 130.675 ;
        RECT 84.920 129.610 85.110 130.505 ;
        RECT 87.010 130.335 87.180 130.845 ;
        RECT 87.350 130.585 87.870 130.895 ;
        RECT 85.280 130.165 87.180 130.335 ;
        RECT 85.280 130.105 85.610 130.165 ;
        RECT 85.760 129.935 86.090 129.995 ;
        RECT 85.430 129.665 86.090 129.935 ;
        RECT 84.920 129.280 85.240 129.610 ;
        RECT 85.420 129.015 86.080 129.495 ;
        RECT 86.280 129.405 86.450 130.165 ;
        RECT 87.350 129.995 87.530 130.405 ;
        RECT 86.620 129.825 86.950 129.945 ;
        RECT 87.700 129.825 87.870 130.585 ;
        RECT 86.620 129.655 87.870 129.825 ;
        RECT 88.040 130.765 89.410 131.015 ;
        RECT 88.040 129.995 88.230 130.765 ;
        RECT 89.160 130.505 89.410 130.765 ;
        RECT 88.400 130.335 88.650 130.495 ;
        RECT 89.580 130.335 89.750 131.180 ;
        RECT 90.645 130.895 90.815 131.395 ;
        RECT 90.985 131.065 91.315 131.565 ;
        RECT 89.920 130.505 90.420 130.885 ;
        RECT 90.645 130.725 91.340 130.895 ;
        RECT 88.400 130.165 89.750 130.335 ;
        RECT 89.330 130.125 89.750 130.165 ;
        RECT 88.040 129.655 88.460 129.995 ;
        RECT 88.750 129.665 89.160 129.995 ;
        RECT 86.280 129.235 87.130 129.405 ;
        RECT 87.690 129.015 88.010 129.475 ;
        RECT 88.210 129.225 88.460 129.655 ;
        RECT 88.750 129.015 89.160 129.455 ;
        RECT 89.330 129.395 89.500 130.125 ;
        RECT 89.670 129.575 90.020 129.945 ;
        RECT 90.200 129.635 90.420 130.505 ;
        RECT 90.590 129.935 91.000 130.555 ;
        RECT 91.170 129.755 91.340 130.725 ;
        RECT 90.645 129.565 91.340 129.755 ;
        RECT 89.330 129.195 90.345 129.395 ;
        RECT 90.645 129.235 90.815 129.565 ;
        RECT 90.985 129.015 91.315 129.395 ;
        RECT 91.530 129.275 91.755 131.395 ;
        RECT 91.925 131.065 92.255 131.565 ;
        RECT 92.425 130.895 92.595 131.395 ;
        RECT 91.930 130.725 92.595 130.895 ;
        RECT 91.930 129.735 92.160 130.725 ;
        RECT 92.330 129.905 92.680 130.555 ;
        RECT 92.915 130.425 93.125 131.565 ;
        RECT 93.295 130.415 93.625 131.395 ;
        RECT 93.795 130.425 94.025 131.565 ;
        RECT 94.235 130.475 95.445 131.565 ;
        RECT 95.615 130.490 95.885 131.395 ;
        RECT 96.055 130.805 96.385 131.565 ;
        RECT 96.565 130.635 96.735 131.395 ;
        RECT 91.930 129.565 92.595 129.735 ;
        RECT 91.925 129.015 92.255 129.395 ;
        RECT 92.425 129.275 92.595 129.565 ;
        RECT 92.915 129.015 93.125 129.835 ;
        RECT 93.295 129.815 93.545 130.415 ;
        RECT 93.715 130.005 94.045 130.255 ;
        RECT 94.235 129.935 94.755 130.475 ;
        RECT 93.295 129.185 93.625 129.815 ;
        RECT 93.795 129.015 94.025 129.835 ;
        RECT 94.925 129.765 95.445 130.305 ;
        RECT 94.235 129.015 95.445 129.765 ;
        RECT 95.615 129.690 95.785 130.490 ;
        RECT 96.070 130.465 96.735 130.635 ;
        RECT 96.995 130.475 99.585 131.565 ;
        RECT 96.070 130.320 96.240 130.465 ;
        RECT 95.955 129.990 96.240 130.320 ;
        RECT 96.070 129.735 96.240 129.990 ;
        RECT 96.475 129.915 96.805 130.285 ;
        RECT 96.995 129.955 98.205 130.475 ;
        RECT 99.755 130.400 100.045 131.565 ;
        RECT 100.675 130.845 101.135 131.395 ;
        RECT 101.325 130.845 101.655 131.565 ;
        RECT 98.375 129.785 99.585 130.305 ;
        RECT 95.615 129.185 95.875 129.690 ;
        RECT 96.070 129.565 96.735 129.735 ;
        RECT 96.055 129.015 96.385 129.395 ;
        RECT 96.565 129.185 96.735 129.565 ;
        RECT 96.995 129.015 99.585 129.785 ;
        RECT 99.755 129.015 100.045 129.740 ;
        RECT 100.675 129.475 100.925 130.845 ;
        RECT 101.855 130.675 102.155 131.225 ;
        RECT 102.325 130.895 102.605 131.565 ;
        RECT 103.030 130.695 103.315 131.565 ;
        RECT 103.485 130.935 103.745 131.395 ;
        RECT 103.920 131.105 104.175 131.565 ;
        RECT 104.345 130.935 104.605 131.395 ;
        RECT 103.485 130.765 104.605 130.935 ;
        RECT 104.775 130.765 105.085 131.565 ;
        RECT 101.215 130.505 102.155 130.675 ;
        RECT 101.215 130.255 101.385 130.505 ;
        RECT 102.525 130.255 102.790 130.615 ;
        RECT 103.485 130.515 103.745 130.765 ;
        RECT 105.255 130.595 105.565 131.395 ;
        RECT 101.095 129.925 101.385 130.255 ;
        RECT 101.555 130.005 101.895 130.255 ;
        RECT 102.115 130.005 102.790 130.255 ;
        RECT 102.990 130.345 103.745 130.515 ;
        RECT 104.535 130.425 105.565 130.595 ;
        RECT 101.215 129.835 101.385 129.925 ;
        RECT 102.990 129.835 103.395 130.345 ;
        RECT 104.535 130.175 104.705 130.425 ;
        RECT 103.565 130.005 104.705 130.175 ;
        RECT 101.215 129.645 102.605 129.835 ;
        RECT 102.990 129.665 104.640 129.835 ;
        RECT 104.875 129.685 105.225 130.255 ;
        RECT 100.675 129.185 101.235 129.475 ;
        RECT 101.405 129.015 101.655 129.475 ;
        RECT 102.275 129.285 102.605 129.645 ;
        RECT 103.035 129.015 103.315 129.495 ;
        RECT 103.485 129.275 103.745 129.665 ;
        RECT 103.920 129.015 104.175 129.495 ;
        RECT 104.345 129.275 104.640 129.665 ;
        RECT 105.395 129.515 105.565 130.425 ;
        RECT 104.820 129.015 105.095 129.495 ;
        RECT 105.265 129.185 105.565 129.515 ;
        RECT 106.655 130.845 107.115 131.395 ;
        RECT 107.305 130.845 107.635 131.565 ;
        RECT 106.655 129.475 106.905 130.845 ;
        RECT 107.835 130.675 108.135 131.225 ;
        RECT 108.305 130.895 108.585 131.565 ;
        RECT 107.195 130.505 108.135 130.675 ;
        RECT 108.955 130.845 109.415 131.395 ;
        RECT 109.605 130.845 109.935 131.565 ;
        RECT 107.195 130.255 107.365 130.505 ;
        RECT 108.505 130.255 108.770 130.615 ;
        RECT 107.075 129.925 107.365 130.255 ;
        RECT 107.535 130.005 107.875 130.255 ;
        RECT 108.095 130.005 108.770 130.255 ;
        RECT 107.195 129.835 107.365 129.925 ;
        RECT 107.195 129.645 108.585 129.835 ;
        RECT 106.655 129.185 107.215 129.475 ;
        RECT 107.385 129.015 107.635 129.475 ;
        RECT 108.255 129.285 108.585 129.645 ;
        RECT 108.955 129.475 109.205 130.845 ;
        RECT 110.135 130.675 110.435 131.225 ;
        RECT 110.605 130.895 110.885 131.565 ;
        RECT 109.495 130.505 110.435 130.675 ;
        RECT 109.495 130.255 109.665 130.505 ;
        RECT 110.805 130.255 111.070 130.615 ;
        RECT 109.375 129.925 109.665 130.255 ;
        RECT 109.835 130.005 110.175 130.255 ;
        RECT 110.395 130.005 111.070 130.255 ;
        RECT 111.715 130.475 113.385 131.565 ;
        RECT 113.560 131.130 118.905 131.565 ;
        RECT 119.080 131.130 124.425 131.565 ;
        RECT 111.715 129.955 112.465 130.475 ;
        RECT 109.495 129.835 109.665 129.925 ;
        RECT 109.495 129.645 110.885 129.835 ;
        RECT 112.635 129.785 113.385 130.305 ;
        RECT 115.150 129.880 115.500 131.130 ;
        RECT 108.955 129.185 109.515 129.475 ;
        RECT 109.685 129.015 109.935 129.475 ;
        RECT 110.555 129.285 110.885 129.645 ;
        RECT 111.715 129.015 113.385 129.785 ;
        RECT 116.980 129.560 117.320 130.390 ;
        RECT 120.670 129.880 121.020 131.130 ;
        RECT 124.595 130.475 125.805 131.565 ;
        RECT 122.500 129.560 122.840 130.390 ;
        RECT 124.595 129.935 125.115 130.475 ;
        RECT 125.285 129.765 125.805 130.305 ;
        RECT 113.560 129.015 118.905 129.560 ;
        RECT 119.080 129.015 124.425 129.560 ;
        RECT 124.595 129.015 125.805 129.765 ;
        RECT 11.810 128.845 125.890 129.015 ;
        RECT 11.895 128.095 13.105 128.845 ;
        RECT 14.570 128.505 14.825 128.665 ;
        RECT 14.485 128.335 14.825 128.505 ;
        RECT 15.005 128.385 15.290 128.845 ;
        RECT 14.570 128.135 14.825 128.335 ;
        RECT 11.895 127.555 12.415 128.095 ;
        RECT 12.585 127.385 13.105 127.925 ;
        RECT 11.895 126.295 13.105 127.385 ;
        RECT 14.570 127.275 14.750 128.135 ;
        RECT 15.470 127.935 15.720 128.585 ;
        RECT 14.920 127.605 15.720 127.935 ;
        RECT 14.570 126.605 14.825 127.275 ;
        RECT 15.005 126.295 15.290 127.095 ;
        RECT 15.470 127.015 15.720 127.605 ;
        RECT 15.920 128.250 16.240 128.580 ;
        RECT 16.420 128.365 17.080 128.845 ;
        RECT 17.280 128.455 18.130 128.625 ;
        RECT 15.920 127.355 16.110 128.250 ;
        RECT 16.430 127.925 17.090 128.195 ;
        RECT 16.760 127.865 17.090 127.925 ;
        RECT 16.280 127.695 16.610 127.755 ;
        RECT 17.280 127.695 17.450 128.455 ;
        RECT 18.690 128.385 19.010 128.845 ;
        RECT 19.210 128.205 19.460 128.635 ;
        RECT 19.750 128.405 20.160 128.845 ;
        RECT 20.330 128.465 21.345 128.665 ;
        RECT 17.620 128.035 18.870 128.205 ;
        RECT 17.620 127.915 17.950 128.035 ;
        RECT 16.280 127.525 18.180 127.695 ;
        RECT 15.920 127.185 17.840 127.355 ;
        RECT 15.920 127.165 16.240 127.185 ;
        RECT 15.470 126.505 15.800 127.015 ;
        RECT 16.070 126.555 16.240 127.165 ;
        RECT 18.010 127.015 18.180 127.525 ;
        RECT 18.350 127.455 18.530 127.865 ;
        RECT 18.700 127.275 18.870 128.035 ;
        RECT 16.410 126.295 16.740 126.985 ;
        RECT 16.970 126.845 18.180 127.015 ;
        RECT 18.350 126.965 18.870 127.275 ;
        RECT 19.040 127.865 19.460 128.205 ;
        RECT 19.750 127.865 20.160 128.195 ;
        RECT 19.040 127.095 19.230 127.865 ;
        RECT 20.330 127.735 20.500 128.465 ;
        RECT 21.645 128.295 21.815 128.625 ;
        RECT 21.985 128.465 22.315 128.845 ;
        RECT 20.670 127.915 21.020 128.285 ;
        RECT 20.330 127.695 20.750 127.735 ;
        RECT 19.400 127.525 20.750 127.695 ;
        RECT 19.400 127.365 19.650 127.525 ;
        RECT 20.160 127.095 20.410 127.355 ;
        RECT 19.040 126.845 20.410 127.095 ;
        RECT 16.970 126.555 17.210 126.845 ;
        RECT 18.010 126.765 18.180 126.845 ;
        RECT 17.410 126.295 17.830 126.675 ;
        RECT 18.010 126.515 18.640 126.765 ;
        RECT 19.110 126.295 19.440 126.675 ;
        RECT 19.610 126.555 19.780 126.845 ;
        RECT 20.580 126.680 20.750 127.525 ;
        RECT 21.200 127.355 21.420 128.225 ;
        RECT 21.645 128.105 22.340 128.295 ;
        RECT 20.920 126.975 21.420 127.355 ;
        RECT 21.590 127.305 22.000 127.925 ;
        RECT 22.170 127.135 22.340 128.105 ;
        RECT 21.645 126.965 22.340 127.135 ;
        RECT 19.960 126.295 20.340 126.675 ;
        RECT 20.580 126.510 21.410 126.680 ;
        RECT 21.645 126.465 21.815 126.965 ;
        RECT 21.985 126.295 22.315 126.795 ;
        RECT 22.530 126.465 22.755 128.585 ;
        RECT 22.925 128.465 23.255 128.845 ;
        RECT 23.425 128.295 23.595 128.585 ;
        RECT 22.930 128.125 23.595 128.295 ;
        RECT 23.855 128.170 24.115 128.675 ;
        RECT 24.295 128.465 24.625 128.845 ;
        RECT 24.805 128.295 24.975 128.675 ;
        RECT 22.930 127.135 23.160 128.125 ;
        RECT 23.330 127.305 23.680 127.955 ;
        RECT 23.855 127.370 24.025 128.170 ;
        RECT 24.310 128.125 24.975 128.295 ;
        RECT 26.245 128.295 26.415 128.675 ;
        RECT 26.595 128.465 26.925 128.845 ;
        RECT 26.245 128.125 26.910 128.295 ;
        RECT 27.105 128.170 27.365 128.675 ;
        RECT 24.310 127.870 24.480 128.125 ;
        RECT 24.195 127.540 24.480 127.870 ;
        RECT 24.715 127.575 25.045 127.945 ;
        RECT 26.175 127.575 26.505 127.945 ;
        RECT 26.740 127.870 26.910 128.125 ;
        RECT 24.310 127.395 24.480 127.540 ;
        RECT 26.740 127.540 27.025 127.870 ;
        RECT 26.740 127.395 26.910 127.540 ;
        RECT 22.930 126.965 23.595 127.135 ;
        RECT 22.925 126.295 23.255 126.795 ;
        RECT 23.425 126.465 23.595 126.965 ;
        RECT 23.855 126.465 24.125 127.370 ;
        RECT 24.310 127.225 24.975 127.395 ;
        RECT 24.295 126.295 24.625 127.055 ;
        RECT 24.805 126.465 24.975 127.225 ;
        RECT 26.245 127.225 26.910 127.395 ;
        RECT 27.195 127.370 27.365 128.170 ;
        RECT 27.735 128.215 28.065 128.575 ;
        RECT 28.685 128.385 28.935 128.845 ;
        RECT 29.105 128.385 29.665 128.675 ;
        RECT 27.735 128.025 29.125 128.215 ;
        RECT 28.955 127.935 29.125 128.025 ;
        RECT 26.245 126.465 26.415 127.225 ;
        RECT 26.595 126.295 26.925 127.055 ;
        RECT 27.095 126.465 27.365 127.370 ;
        RECT 27.550 127.605 28.225 127.855 ;
        RECT 28.445 127.605 28.785 127.855 ;
        RECT 28.955 127.605 29.245 127.935 ;
        RECT 27.550 127.245 27.815 127.605 ;
        RECT 28.955 127.355 29.125 127.605 ;
        RECT 28.185 127.185 29.125 127.355 ;
        RECT 27.735 126.295 28.015 126.965 ;
        RECT 28.185 126.635 28.485 127.185 ;
        RECT 29.415 127.015 29.665 128.385 ;
        RECT 28.685 126.295 29.015 127.015 ;
        RECT 29.205 126.465 29.665 127.015 ;
        RECT 29.840 128.105 30.095 128.675 ;
        RECT 30.265 128.445 30.595 128.845 ;
        RECT 31.020 128.310 31.550 128.675 ;
        RECT 31.740 128.505 32.015 128.675 ;
        RECT 31.735 128.335 32.015 128.505 ;
        RECT 31.020 128.275 31.195 128.310 ;
        RECT 30.265 128.105 31.195 128.275 ;
        RECT 29.840 127.435 30.010 128.105 ;
        RECT 30.265 127.935 30.435 128.105 ;
        RECT 30.180 127.605 30.435 127.935 ;
        RECT 30.660 127.605 30.855 127.935 ;
        RECT 29.840 126.465 30.175 127.435 ;
        RECT 30.345 126.295 30.515 127.435 ;
        RECT 30.685 126.635 30.855 127.605 ;
        RECT 31.025 126.975 31.195 128.105 ;
        RECT 31.365 127.315 31.535 128.115 ;
        RECT 31.740 127.515 32.015 128.335 ;
        RECT 32.185 127.315 32.375 128.675 ;
        RECT 32.555 128.310 33.065 128.845 ;
        RECT 33.285 128.035 33.530 128.640 ;
        RECT 33.975 128.095 35.185 128.845 ;
        RECT 35.355 128.120 35.645 128.845 ;
        RECT 35.815 128.095 37.025 128.845 ;
        RECT 32.575 127.865 33.805 128.035 ;
        RECT 31.365 127.145 32.375 127.315 ;
        RECT 32.545 127.300 33.295 127.490 ;
        RECT 31.025 126.805 32.150 126.975 ;
        RECT 32.545 126.635 32.715 127.300 ;
        RECT 33.465 127.055 33.805 127.865 ;
        RECT 30.685 126.465 32.715 126.635 ;
        RECT 32.885 126.295 33.055 127.055 ;
        RECT 33.290 126.645 33.805 127.055 ;
        RECT 33.975 127.385 34.495 127.925 ;
        RECT 34.665 127.555 35.185 128.095 ;
        RECT 33.975 126.295 35.185 127.385 ;
        RECT 35.355 126.295 35.645 127.460 ;
        RECT 35.815 127.385 36.335 127.925 ;
        RECT 36.505 127.555 37.025 128.095 ;
        RECT 37.195 128.170 37.465 128.515 ;
        RECT 37.655 128.445 38.035 128.845 ;
        RECT 38.205 128.275 38.375 128.625 ;
        RECT 38.545 128.445 38.875 128.845 ;
        RECT 39.075 128.275 39.245 128.625 ;
        RECT 39.445 128.345 39.775 128.845 ;
        RECT 37.195 127.435 37.365 128.170 ;
        RECT 37.635 128.105 39.245 128.275 ;
        RECT 37.635 127.935 37.805 128.105 ;
        RECT 37.535 127.605 37.805 127.935 ;
        RECT 37.975 127.605 38.380 127.935 ;
        RECT 37.635 127.435 37.805 127.605 ;
        RECT 35.815 126.295 37.025 127.385 ;
        RECT 37.195 126.465 37.465 127.435 ;
        RECT 37.635 127.265 38.360 127.435 ;
        RECT 38.550 127.315 39.260 127.935 ;
        RECT 39.430 127.605 39.780 128.175 ;
        RECT 39.955 128.045 40.295 128.675 ;
        RECT 40.465 128.045 40.715 128.845 ;
        RECT 40.905 128.195 41.235 128.675 ;
        RECT 41.405 128.385 41.630 128.845 ;
        RECT 41.800 128.195 42.130 128.675 ;
        RECT 39.955 127.435 40.130 128.045 ;
        RECT 40.905 128.025 42.130 128.195 ;
        RECT 42.760 128.065 43.260 128.675 ;
        RECT 43.745 128.365 43.915 128.845 ;
        RECT 44.085 128.195 44.415 128.670 ;
        RECT 44.585 128.365 44.755 128.845 ;
        RECT 44.925 128.195 45.255 128.670 ;
        RECT 45.425 128.365 45.595 128.845 ;
        RECT 45.765 128.195 46.095 128.670 ;
        RECT 46.265 128.365 46.435 128.845 ;
        RECT 46.605 128.195 46.935 128.670 ;
        RECT 47.105 128.365 47.275 128.845 ;
        RECT 47.445 128.195 47.775 128.670 ;
        RECT 47.945 128.365 48.115 128.845 ;
        RECT 48.365 128.670 48.535 128.675 ;
        RECT 48.285 128.195 48.615 128.670 ;
        RECT 48.785 128.365 48.955 128.845 ;
        RECT 49.205 128.670 49.375 128.675 ;
        RECT 49.125 128.195 49.455 128.670 ;
        RECT 49.625 128.365 49.795 128.845 ;
        RECT 50.045 128.670 50.295 128.675 ;
        RECT 49.965 128.195 50.295 128.670 ;
        RECT 50.465 128.365 50.635 128.845 ;
        RECT 50.805 128.195 51.135 128.670 ;
        RECT 51.305 128.365 51.475 128.845 ;
        RECT 51.645 128.195 51.975 128.670 ;
        RECT 52.145 128.365 52.315 128.845 ;
        RECT 52.485 128.195 52.815 128.670 ;
        RECT 52.985 128.365 53.155 128.845 ;
        RECT 53.325 128.195 53.655 128.670 ;
        RECT 53.825 128.365 53.995 128.845 ;
        RECT 54.165 128.195 54.495 128.670 ;
        RECT 40.300 127.685 40.995 127.855 ;
        RECT 40.825 127.435 40.995 127.685 ;
        RECT 41.170 127.655 41.590 127.855 ;
        RECT 41.760 127.655 42.090 127.855 ;
        RECT 42.260 127.655 42.590 127.855 ;
        RECT 42.760 127.435 42.930 128.065 ;
        RECT 43.635 128.025 50.295 128.195 ;
        RECT 50.465 128.025 52.815 128.195 ;
        RECT 52.985 128.025 54.495 128.195 ;
        RECT 54.715 128.025 54.945 128.845 ;
        RECT 55.115 128.045 55.445 128.675 ;
        RECT 43.115 127.605 43.465 127.855 ;
        RECT 43.635 127.485 43.910 128.025 ;
        RECT 50.465 127.855 50.640 128.025 ;
        RECT 52.985 127.855 53.155 128.025 ;
        RECT 44.080 127.655 50.640 127.855 ;
        RECT 50.845 127.655 53.155 127.855 ;
        RECT 53.325 127.655 54.500 127.855 ;
        RECT 50.465 127.485 50.640 127.655 ;
        RECT 52.985 127.485 53.155 127.655 ;
        RECT 54.695 127.605 55.025 127.855 ;
        RECT 38.190 127.145 38.360 127.265 ;
        RECT 39.460 127.145 39.780 127.435 ;
        RECT 37.675 126.295 37.955 127.095 ;
        RECT 38.190 126.975 39.780 127.145 ;
        RECT 38.125 126.515 39.780 126.805 ;
        RECT 39.955 126.465 40.295 127.435 ;
        RECT 40.465 126.295 40.635 127.435 ;
        RECT 40.825 127.265 43.260 127.435 ;
        RECT 43.635 127.315 50.295 127.485 ;
        RECT 50.465 127.315 52.815 127.485 ;
        RECT 52.985 127.315 54.495 127.485 ;
        RECT 55.195 127.445 55.445 128.045 ;
        RECT 55.615 128.025 55.825 128.845 ;
        RECT 56.330 128.035 56.575 128.640 ;
        RECT 56.795 128.310 57.305 128.845 ;
        RECT 40.905 126.295 41.155 127.095 ;
        RECT 41.800 126.465 42.130 127.265 ;
        RECT 42.430 126.295 42.760 127.095 ;
        RECT 42.930 126.465 43.260 127.265 ;
        RECT 43.745 126.295 43.915 127.095 ;
        RECT 44.085 126.465 44.415 127.315 ;
        RECT 44.585 126.295 44.755 127.095 ;
        RECT 44.925 126.465 45.255 127.315 ;
        RECT 45.425 126.295 45.595 127.095 ;
        RECT 45.765 126.465 46.095 127.315 ;
        RECT 46.265 126.295 46.435 127.095 ;
        RECT 46.605 126.465 46.935 127.315 ;
        RECT 47.105 126.295 47.275 127.095 ;
        RECT 47.445 126.465 47.775 127.315 ;
        RECT 47.945 126.295 48.115 127.095 ;
        RECT 48.285 126.465 48.615 127.315 ;
        RECT 48.785 126.295 48.955 127.095 ;
        RECT 49.125 126.465 49.455 127.315 ;
        RECT 49.625 126.295 49.795 127.095 ;
        RECT 49.965 126.465 50.295 127.315 ;
        RECT 50.465 126.295 50.635 127.095 ;
        RECT 50.805 126.465 51.135 127.315 ;
        RECT 51.305 126.295 51.475 127.095 ;
        RECT 51.645 126.465 51.975 127.315 ;
        RECT 52.145 126.295 52.315 127.095 ;
        RECT 52.485 126.465 52.815 127.315 ;
        RECT 52.985 126.295 53.155 127.145 ;
        RECT 53.325 126.465 53.655 127.315 ;
        RECT 53.825 126.295 53.995 127.145 ;
        RECT 54.165 126.465 54.495 127.315 ;
        RECT 54.715 126.295 54.945 127.435 ;
        RECT 55.115 126.465 55.445 127.445 ;
        RECT 56.055 127.865 57.285 128.035 ;
        RECT 55.615 126.295 55.825 127.435 ;
        RECT 56.055 127.055 56.395 127.865 ;
        RECT 56.565 127.300 57.315 127.490 ;
        RECT 56.055 126.645 56.570 127.055 ;
        RECT 56.805 126.295 56.975 127.055 ;
        RECT 57.145 126.635 57.315 127.300 ;
        RECT 57.485 127.315 57.675 128.675 ;
        RECT 57.845 128.505 58.120 128.675 ;
        RECT 57.845 128.335 58.125 128.505 ;
        RECT 57.845 127.515 58.120 128.335 ;
        RECT 58.310 128.310 58.840 128.675 ;
        RECT 59.265 128.445 59.595 128.845 ;
        RECT 58.665 128.275 58.840 128.310 ;
        RECT 58.325 127.315 58.495 128.115 ;
        RECT 57.485 127.145 58.495 127.315 ;
        RECT 58.665 128.105 59.595 128.275 ;
        RECT 59.765 128.105 60.020 128.675 ;
        RECT 61.115 128.120 61.405 128.845 ;
        RECT 62.585 128.295 62.755 128.675 ;
        RECT 62.935 128.465 63.265 128.845 ;
        RECT 62.585 128.125 63.250 128.295 ;
        RECT 63.445 128.170 63.705 128.675 ;
        RECT 58.665 126.975 58.835 128.105 ;
        RECT 59.425 127.935 59.595 128.105 ;
        RECT 57.710 126.805 58.835 126.975 ;
        RECT 59.005 127.605 59.200 127.935 ;
        RECT 59.425 127.605 59.680 127.935 ;
        RECT 59.005 126.635 59.175 127.605 ;
        RECT 59.850 127.435 60.020 128.105 ;
        RECT 62.515 127.575 62.845 127.945 ;
        RECT 63.080 127.870 63.250 128.125 ;
        RECT 63.080 127.540 63.365 127.870 ;
        RECT 57.145 126.465 59.175 126.635 ;
        RECT 59.345 126.295 59.515 127.435 ;
        RECT 59.685 126.465 60.020 127.435 ;
        RECT 61.115 126.295 61.405 127.460 ;
        RECT 63.080 127.395 63.250 127.540 ;
        RECT 62.585 127.225 63.250 127.395 ;
        RECT 63.535 127.370 63.705 128.170 ;
        RECT 63.915 128.025 64.145 128.845 ;
        RECT 64.315 128.045 64.645 128.675 ;
        RECT 63.895 127.605 64.225 127.855 ;
        RECT 64.395 127.445 64.645 128.045 ;
        RECT 64.815 128.025 65.025 128.845 ;
        RECT 65.255 128.095 66.465 128.845 ;
        RECT 62.585 126.465 62.755 127.225 ;
        RECT 62.935 126.295 63.265 127.055 ;
        RECT 63.435 126.465 63.705 127.370 ;
        RECT 63.915 126.295 64.145 127.435 ;
        RECT 64.315 126.465 64.645 127.445 ;
        RECT 64.815 126.295 65.025 127.435 ;
        RECT 65.255 127.385 65.775 127.925 ;
        RECT 65.945 127.555 66.465 128.095 ;
        RECT 66.635 128.075 70.145 128.845 ;
        RECT 66.635 127.385 68.325 127.905 ;
        RECT 68.495 127.555 70.145 128.075 ;
        RECT 70.315 128.385 70.875 128.675 ;
        RECT 71.045 128.385 71.295 128.845 ;
        RECT 65.255 126.295 66.465 127.385 ;
        RECT 66.635 126.295 70.145 127.385 ;
        RECT 70.315 127.015 70.565 128.385 ;
        RECT 71.915 128.215 72.245 128.575 ;
        RECT 70.855 128.025 72.245 128.215 ;
        RECT 72.615 128.075 74.285 128.845 ;
        RECT 70.855 127.935 71.025 128.025 ;
        RECT 70.735 127.605 71.025 127.935 ;
        RECT 71.195 127.605 71.535 127.855 ;
        RECT 71.755 127.605 72.430 127.855 ;
        RECT 70.855 127.355 71.025 127.605 ;
        RECT 70.855 127.185 71.795 127.355 ;
        RECT 72.165 127.245 72.430 127.605 ;
        RECT 72.615 127.385 73.365 127.905 ;
        RECT 73.535 127.555 74.285 128.075 ;
        RECT 74.655 128.215 74.985 128.575 ;
        RECT 75.605 128.385 75.855 128.845 ;
        RECT 76.025 128.385 76.585 128.675 ;
        RECT 74.655 128.025 76.045 128.215 ;
        RECT 75.875 127.935 76.045 128.025 ;
        RECT 74.470 127.605 75.145 127.855 ;
        RECT 75.365 127.605 75.705 127.855 ;
        RECT 75.875 127.605 76.165 127.935 ;
        RECT 70.315 126.465 70.775 127.015 ;
        RECT 70.965 126.295 71.295 127.015 ;
        RECT 71.495 126.635 71.795 127.185 ;
        RECT 71.965 126.295 72.245 126.965 ;
        RECT 72.615 126.295 74.285 127.385 ;
        RECT 74.470 127.245 74.735 127.605 ;
        RECT 75.875 127.355 76.045 127.605 ;
        RECT 75.105 127.185 76.045 127.355 ;
        RECT 74.655 126.295 74.935 126.965 ;
        RECT 75.105 126.635 75.405 127.185 ;
        RECT 76.335 127.015 76.585 128.385 ;
        RECT 75.605 126.295 75.935 127.015 ;
        RECT 76.125 126.465 76.585 127.015 ;
        RECT 76.755 128.170 77.025 128.515 ;
        RECT 77.215 128.445 77.595 128.845 ;
        RECT 77.765 128.275 77.935 128.625 ;
        RECT 78.105 128.445 78.435 128.845 ;
        RECT 78.635 128.275 78.805 128.625 ;
        RECT 79.005 128.345 79.335 128.845 ;
        RECT 79.515 128.385 80.075 128.675 ;
        RECT 80.245 128.385 80.495 128.845 ;
        RECT 76.755 127.435 76.925 128.170 ;
        RECT 77.195 128.105 78.805 128.275 ;
        RECT 77.195 127.935 77.365 128.105 ;
        RECT 77.095 127.605 77.365 127.935 ;
        RECT 77.535 127.605 77.940 127.935 ;
        RECT 77.195 127.435 77.365 127.605 ;
        RECT 78.110 127.485 78.820 127.935 ;
        RECT 78.990 127.605 79.340 128.175 ;
        RECT 76.755 126.465 77.025 127.435 ;
        RECT 77.195 127.265 77.920 127.435 ;
        RECT 78.110 127.315 78.825 127.485 ;
        RECT 77.750 127.145 77.920 127.265 ;
        RECT 79.020 127.145 79.340 127.435 ;
        RECT 77.235 126.295 77.515 127.095 ;
        RECT 77.750 126.975 79.340 127.145 ;
        RECT 79.515 127.015 79.765 128.385 ;
        RECT 81.115 128.215 81.445 128.575 ;
        RECT 80.055 128.025 81.445 128.215 ;
        RECT 81.815 128.095 83.025 128.845 ;
        RECT 80.055 127.935 80.225 128.025 ;
        RECT 79.935 127.605 80.225 127.935 ;
        RECT 80.395 127.605 80.735 127.855 ;
        RECT 80.955 127.605 81.630 127.855 ;
        RECT 80.055 127.355 80.225 127.605 ;
        RECT 80.055 127.185 80.995 127.355 ;
        RECT 81.365 127.245 81.630 127.605 ;
        RECT 81.815 127.385 82.335 127.925 ;
        RECT 82.505 127.555 83.025 128.095 ;
        RECT 83.195 128.075 86.705 128.845 ;
        RECT 86.875 128.120 87.165 128.845 ;
        RECT 83.195 127.385 84.885 127.905 ;
        RECT 85.055 127.555 86.705 128.075 ;
        RECT 87.855 128.025 88.065 128.845 ;
        RECT 88.235 128.045 88.565 128.675 ;
        RECT 77.685 126.515 79.340 126.805 ;
        RECT 79.515 126.465 79.975 127.015 ;
        RECT 80.165 126.295 80.495 127.015 ;
        RECT 80.695 126.635 80.995 127.185 ;
        RECT 81.165 126.295 81.445 126.965 ;
        RECT 81.815 126.295 83.025 127.385 ;
        RECT 83.195 126.295 86.705 127.385 ;
        RECT 86.875 126.295 87.165 127.460 ;
        RECT 88.235 127.445 88.485 128.045 ;
        RECT 88.735 128.025 88.965 128.845 ;
        RECT 89.635 128.075 91.305 128.845 ;
        RECT 91.480 128.375 91.810 128.845 ;
        RECT 91.980 128.205 92.205 128.650 ;
        RECT 92.375 128.320 92.670 128.845 ;
        RECT 94.235 128.385 94.795 128.675 ;
        RECT 94.965 128.385 95.215 128.845 ;
        RECT 88.655 127.605 88.985 127.855 ;
        RECT 87.855 126.295 88.065 127.435 ;
        RECT 88.235 126.465 88.565 127.445 ;
        RECT 88.735 126.295 88.965 127.435 ;
        RECT 89.635 127.385 90.385 127.905 ;
        RECT 90.555 127.555 91.305 128.075 ;
        RECT 91.475 128.035 92.205 128.205 ;
        RECT 91.475 127.470 91.755 128.035 ;
        RECT 91.925 127.640 93.145 127.865 ;
        RECT 89.635 126.295 91.305 127.385 ;
        RECT 91.475 127.300 93.075 127.470 ;
        RECT 91.535 126.295 91.790 127.130 ;
        RECT 91.960 126.495 92.220 127.300 ;
        RECT 92.390 126.295 92.650 127.130 ;
        RECT 92.820 126.495 93.075 127.300 ;
        RECT 94.235 127.015 94.485 128.385 ;
        RECT 95.835 128.215 96.165 128.575 ;
        RECT 96.535 128.335 96.840 128.845 ;
        RECT 94.775 128.025 96.165 128.215 ;
        RECT 94.775 127.935 94.945 128.025 ;
        RECT 94.655 127.605 94.945 127.935 ;
        RECT 95.115 127.605 95.455 127.855 ;
        RECT 95.675 127.605 96.350 127.855 ;
        RECT 96.535 127.605 96.850 128.165 ;
        RECT 97.020 127.855 97.270 128.665 ;
        RECT 97.440 128.320 97.700 128.845 ;
        RECT 97.880 127.855 98.130 128.665 ;
        RECT 98.300 128.285 98.560 128.845 ;
        RECT 98.730 128.195 98.990 128.650 ;
        RECT 99.160 128.365 99.420 128.845 ;
        RECT 99.590 128.195 99.850 128.650 ;
        RECT 100.020 128.365 100.280 128.845 ;
        RECT 100.450 128.195 100.710 128.650 ;
        RECT 100.880 128.365 101.125 128.845 ;
        RECT 101.295 128.195 101.570 128.650 ;
        RECT 101.740 128.365 101.985 128.845 ;
        RECT 102.155 128.195 102.415 128.650 ;
        RECT 102.595 128.365 102.845 128.845 ;
        RECT 103.015 128.195 103.275 128.650 ;
        RECT 103.455 128.365 103.705 128.845 ;
        RECT 103.875 128.195 104.135 128.650 ;
        RECT 104.315 128.365 104.575 128.845 ;
        RECT 104.745 128.195 105.005 128.650 ;
        RECT 105.175 128.365 105.475 128.845 ;
        RECT 105.735 128.385 106.295 128.675 ;
        RECT 106.465 128.385 106.715 128.845 ;
        RECT 98.730 128.165 105.475 128.195 ;
        RECT 98.730 128.025 105.505 128.165 ;
        RECT 104.310 127.995 105.505 128.025 ;
        RECT 97.020 127.605 104.140 127.855 ;
        RECT 94.775 127.355 94.945 127.605 ;
        RECT 94.775 127.185 95.715 127.355 ;
        RECT 96.085 127.245 96.350 127.605 ;
        RECT 94.235 126.465 94.695 127.015 ;
        RECT 94.885 126.295 95.215 127.015 ;
        RECT 95.415 126.635 95.715 127.185 ;
        RECT 95.885 126.295 96.165 126.965 ;
        RECT 96.545 126.295 96.840 127.105 ;
        RECT 97.020 126.465 97.265 127.605 ;
        RECT 97.440 126.295 97.700 127.105 ;
        RECT 97.880 126.470 98.130 127.605 ;
        RECT 104.310 127.435 105.475 127.995 ;
        RECT 98.730 127.210 105.475 127.435 ;
        RECT 98.730 127.195 104.135 127.210 ;
        RECT 98.300 126.300 98.560 127.095 ;
        RECT 98.730 126.470 98.990 127.195 ;
        RECT 99.160 126.300 99.420 127.025 ;
        RECT 99.590 126.470 99.850 127.195 ;
        RECT 100.020 126.300 100.280 127.025 ;
        RECT 100.450 126.470 100.710 127.195 ;
        RECT 100.880 126.300 101.140 127.025 ;
        RECT 101.310 126.470 101.570 127.195 ;
        RECT 101.740 126.300 101.985 127.025 ;
        RECT 102.155 126.470 102.415 127.195 ;
        RECT 102.600 126.300 102.845 127.025 ;
        RECT 103.015 126.470 103.275 127.195 ;
        RECT 103.460 126.300 103.705 127.025 ;
        RECT 103.875 126.470 104.135 127.195 ;
        RECT 104.320 126.300 104.575 127.025 ;
        RECT 104.745 126.470 105.035 127.210 ;
        RECT 98.300 126.295 104.575 126.300 ;
        RECT 105.205 126.295 105.475 127.040 ;
        RECT 105.735 127.015 105.985 128.385 ;
        RECT 107.335 128.215 107.665 128.575 ;
        RECT 106.275 128.025 107.665 128.215 ;
        RECT 108.770 128.035 109.015 128.640 ;
        RECT 109.235 128.310 109.745 128.845 ;
        RECT 106.275 127.935 106.445 128.025 ;
        RECT 106.155 127.605 106.445 127.935 ;
        RECT 108.495 127.865 109.725 128.035 ;
        RECT 106.615 127.605 106.955 127.855 ;
        RECT 107.175 127.605 107.850 127.855 ;
        RECT 106.275 127.355 106.445 127.605 ;
        RECT 106.275 127.185 107.215 127.355 ;
        RECT 107.585 127.245 107.850 127.605 ;
        RECT 105.735 126.465 106.195 127.015 ;
        RECT 106.385 126.295 106.715 127.015 ;
        RECT 106.915 126.635 107.215 127.185 ;
        RECT 108.495 127.055 108.835 127.865 ;
        RECT 109.005 127.300 109.755 127.490 ;
        RECT 107.385 126.295 107.665 126.965 ;
        RECT 108.495 126.645 109.010 127.055 ;
        RECT 109.245 126.295 109.415 127.055 ;
        RECT 109.585 126.635 109.755 127.300 ;
        RECT 109.925 127.315 110.115 128.675 ;
        RECT 110.285 127.825 110.560 128.675 ;
        RECT 110.750 128.310 111.280 128.675 ;
        RECT 111.705 128.445 112.035 128.845 ;
        RECT 111.105 128.275 111.280 128.310 ;
        RECT 110.285 127.655 110.565 127.825 ;
        RECT 110.285 127.515 110.560 127.655 ;
        RECT 110.765 127.315 110.935 128.115 ;
        RECT 109.925 127.145 110.935 127.315 ;
        RECT 111.105 128.105 112.035 128.275 ;
        RECT 112.205 128.105 112.460 128.675 ;
        RECT 112.635 128.120 112.925 128.845 ;
        RECT 114.390 128.135 114.645 128.665 ;
        RECT 114.825 128.385 115.110 128.845 ;
        RECT 111.105 126.975 111.275 128.105 ;
        RECT 111.865 127.935 112.035 128.105 ;
        RECT 110.150 126.805 111.275 126.975 ;
        RECT 111.445 127.605 111.640 127.935 ;
        RECT 111.865 127.605 112.120 127.935 ;
        RECT 111.445 126.635 111.615 127.605 ;
        RECT 112.290 127.435 112.460 128.105 ;
        RECT 114.390 127.825 114.570 128.135 ;
        RECT 115.290 127.935 115.540 128.585 ;
        RECT 114.305 127.655 114.570 127.825 ;
        RECT 109.585 126.465 111.615 126.635 ;
        RECT 111.785 126.295 111.955 127.435 ;
        RECT 112.125 126.465 112.460 127.435 ;
        RECT 112.635 126.295 112.925 127.460 ;
        RECT 114.390 127.275 114.570 127.655 ;
        RECT 114.740 127.605 115.540 127.935 ;
        RECT 114.390 126.605 114.645 127.275 ;
        RECT 114.825 126.295 115.110 127.095 ;
        RECT 115.290 127.015 115.540 127.605 ;
        RECT 115.740 128.250 116.060 128.580 ;
        RECT 116.240 128.365 116.900 128.845 ;
        RECT 117.100 128.455 117.950 128.625 ;
        RECT 115.740 127.355 115.930 128.250 ;
        RECT 116.250 127.925 116.910 128.195 ;
        RECT 116.580 127.865 116.910 127.925 ;
        RECT 116.100 127.695 116.430 127.755 ;
        RECT 117.100 127.695 117.270 128.455 ;
        RECT 118.510 128.385 118.830 128.845 ;
        RECT 119.030 128.205 119.280 128.635 ;
        RECT 119.570 128.405 119.980 128.845 ;
        RECT 120.150 128.465 121.165 128.665 ;
        RECT 117.440 128.035 118.690 128.205 ;
        RECT 117.440 127.915 117.770 128.035 ;
        RECT 116.100 127.525 118.000 127.695 ;
        RECT 115.740 127.185 117.660 127.355 ;
        RECT 115.740 127.165 116.060 127.185 ;
        RECT 115.290 126.505 115.620 127.015 ;
        RECT 115.890 126.555 116.060 127.165 ;
        RECT 117.830 127.015 118.000 127.525 ;
        RECT 118.170 127.455 118.350 127.865 ;
        RECT 118.520 127.275 118.690 128.035 ;
        RECT 116.230 126.295 116.560 126.985 ;
        RECT 116.790 126.845 118.000 127.015 ;
        RECT 118.170 126.965 118.690 127.275 ;
        RECT 118.860 127.865 119.280 128.205 ;
        RECT 119.570 127.865 119.980 128.195 ;
        RECT 118.860 127.095 119.050 127.865 ;
        RECT 120.150 127.735 120.320 128.465 ;
        RECT 121.465 128.295 121.635 128.625 ;
        RECT 121.805 128.465 122.135 128.845 ;
        RECT 120.490 127.915 120.840 128.285 ;
        RECT 120.150 127.695 120.570 127.735 ;
        RECT 119.220 127.525 120.570 127.695 ;
        RECT 119.220 127.365 119.470 127.525 ;
        RECT 119.980 127.095 120.230 127.355 ;
        RECT 118.860 126.845 120.230 127.095 ;
        RECT 116.790 126.555 117.030 126.845 ;
        RECT 117.830 126.765 118.000 126.845 ;
        RECT 117.230 126.295 117.650 126.675 ;
        RECT 117.830 126.515 118.460 126.765 ;
        RECT 118.930 126.295 119.260 126.675 ;
        RECT 119.430 126.555 119.600 126.845 ;
        RECT 120.400 126.680 120.570 127.525 ;
        RECT 121.020 127.355 121.240 128.225 ;
        RECT 121.465 128.105 122.160 128.295 ;
        RECT 120.740 126.975 121.240 127.355 ;
        RECT 121.410 127.305 121.820 127.925 ;
        RECT 121.990 127.135 122.160 128.105 ;
        RECT 121.465 126.965 122.160 127.135 ;
        RECT 119.780 126.295 120.160 126.675 ;
        RECT 120.400 126.510 121.230 126.680 ;
        RECT 121.465 126.465 121.635 126.965 ;
        RECT 121.805 126.295 122.135 126.795 ;
        RECT 122.350 126.465 122.575 128.585 ;
        RECT 122.745 128.465 123.075 128.845 ;
        RECT 123.245 128.295 123.415 128.585 ;
        RECT 122.750 128.125 123.415 128.295 ;
        RECT 122.750 127.135 122.980 128.125 ;
        RECT 124.595 128.095 125.805 128.845 ;
        RECT 123.150 127.305 123.500 127.955 ;
        RECT 124.595 127.385 125.115 127.925 ;
        RECT 125.285 127.555 125.805 128.095 ;
        RECT 122.750 126.965 123.415 127.135 ;
        RECT 122.745 126.295 123.075 126.795 ;
        RECT 123.245 126.465 123.415 126.965 ;
        RECT 124.595 126.295 125.805 127.385 ;
        RECT 11.810 126.125 125.890 126.295 ;
        RECT 11.895 125.035 13.105 126.125 ;
        RECT 11.895 124.325 12.415 124.865 ;
        RECT 12.585 124.495 13.105 125.035 ;
        RECT 13.275 125.035 16.785 126.125 ;
        RECT 13.275 124.515 14.965 125.035 ;
        RECT 16.995 124.985 17.225 126.125 ;
        RECT 17.395 124.975 17.725 125.955 ;
        RECT 17.895 124.985 18.105 126.125 ;
        RECT 18.335 125.365 18.850 125.775 ;
        RECT 19.085 125.365 19.255 126.125 ;
        RECT 19.425 125.785 21.455 125.955 ;
        RECT 15.135 124.345 16.785 124.865 ;
        RECT 16.975 124.565 17.305 124.815 ;
        RECT 11.895 123.575 13.105 124.325 ;
        RECT 13.275 123.575 16.785 124.345 ;
        RECT 16.995 123.575 17.225 124.395 ;
        RECT 17.475 124.375 17.725 124.975 ;
        RECT 18.335 124.555 18.675 125.365 ;
        RECT 19.425 125.120 19.595 125.785 ;
        RECT 19.990 125.445 21.115 125.615 ;
        RECT 18.845 124.930 19.595 125.120 ;
        RECT 19.765 125.105 20.775 125.275 ;
        RECT 17.395 123.745 17.725 124.375 ;
        RECT 17.895 123.575 18.105 124.395 ;
        RECT 18.335 124.385 19.565 124.555 ;
        RECT 18.610 123.780 18.855 124.385 ;
        RECT 19.075 123.575 19.585 124.110 ;
        RECT 19.765 123.745 19.955 125.105 ;
        RECT 20.125 124.085 20.400 124.905 ;
        RECT 20.605 124.305 20.775 125.105 ;
        RECT 20.945 124.315 21.115 125.445 ;
        RECT 21.285 124.815 21.455 125.785 ;
        RECT 21.625 124.985 21.795 126.125 ;
        RECT 21.965 124.985 22.300 125.955 ;
        RECT 21.285 124.485 21.480 124.815 ;
        RECT 21.705 124.485 21.960 124.815 ;
        RECT 21.705 124.315 21.875 124.485 ;
        RECT 22.130 124.315 22.300 124.985 ;
        RECT 22.475 124.960 22.765 126.125 ;
        RECT 23.025 125.195 23.195 125.955 ;
        RECT 23.375 125.365 23.705 126.125 ;
        RECT 23.025 125.025 23.690 125.195 ;
        RECT 23.875 125.050 24.145 125.955 ;
        RECT 23.520 124.880 23.690 125.025 ;
        RECT 22.955 124.475 23.285 124.845 ;
        RECT 23.520 124.550 23.805 124.880 ;
        RECT 20.945 124.145 21.875 124.315 ;
        RECT 20.945 124.110 21.120 124.145 ;
        RECT 20.125 123.915 20.405 124.085 ;
        RECT 20.125 123.745 20.400 123.915 ;
        RECT 20.590 123.745 21.120 124.110 ;
        RECT 21.545 123.575 21.875 123.975 ;
        RECT 22.045 123.745 22.300 124.315 ;
        RECT 22.475 123.575 22.765 124.300 ;
        RECT 23.520 124.295 23.690 124.550 ;
        RECT 23.025 124.125 23.690 124.295 ;
        RECT 23.975 124.250 24.145 125.050 ;
        RECT 24.315 125.035 26.905 126.125 ;
        RECT 27.275 125.455 27.555 126.125 ;
        RECT 27.725 125.235 28.025 125.785 ;
        RECT 28.225 125.405 28.555 126.125 ;
        RECT 28.745 125.405 29.205 125.955 ;
        RECT 24.315 124.515 25.525 125.035 ;
        RECT 25.695 124.345 26.905 124.865 ;
        RECT 27.090 124.815 27.355 125.175 ;
        RECT 27.725 125.065 28.665 125.235 ;
        RECT 28.495 124.815 28.665 125.065 ;
        RECT 27.090 124.565 27.765 124.815 ;
        RECT 27.985 124.565 28.325 124.815 ;
        RECT 28.495 124.485 28.785 124.815 ;
        RECT 28.495 124.395 28.665 124.485 ;
        RECT 23.025 123.745 23.195 124.125 ;
        RECT 23.375 123.575 23.705 123.955 ;
        RECT 23.885 123.745 24.145 124.250 ;
        RECT 24.315 123.575 26.905 124.345 ;
        RECT 27.275 124.205 28.665 124.395 ;
        RECT 27.275 123.845 27.605 124.205 ;
        RECT 28.955 124.035 29.205 125.405 ;
        RECT 29.465 125.380 29.735 126.125 ;
        RECT 30.365 126.120 36.640 126.125 ;
        RECT 29.905 125.210 30.195 125.950 ;
        RECT 30.365 125.395 30.620 126.120 ;
        RECT 30.805 125.225 31.065 125.950 ;
        RECT 31.235 125.395 31.480 126.120 ;
        RECT 31.665 125.225 31.925 125.950 ;
        RECT 32.095 125.395 32.340 126.120 ;
        RECT 32.525 125.225 32.785 125.950 ;
        RECT 32.955 125.395 33.200 126.120 ;
        RECT 33.370 125.225 33.630 125.950 ;
        RECT 33.800 125.395 34.060 126.120 ;
        RECT 34.230 125.225 34.490 125.950 ;
        RECT 34.660 125.395 34.920 126.120 ;
        RECT 35.090 125.225 35.350 125.950 ;
        RECT 35.520 125.395 35.780 126.120 ;
        RECT 35.950 125.225 36.210 125.950 ;
        RECT 36.380 125.325 36.640 126.120 ;
        RECT 30.805 125.210 36.210 125.225 ;
        RECT 29.465 124.985 36.210 125.210 ;
        RECT 29.465 124.395 30.630 124.985 ;
        RECT 36.810 124.815 37.060 125.950 ;
        RECT 37.240 125.315 37.500 126.125 ;
        RECT 37.675 124.815 37.920 125.955 ;
        RECT 38.100 125.315 38.395 126.125 ;
        RECT 39.040 125.615 40.695 125.905 ;
        RECT 39.040 125.275 40.630 125.445 ;
        RECT 40.865 125.325 41.145 126.125 ;
        RECT 39.040 124.985 39.360 125.275 ;
        RECT 40.460 125.155 40.630 125.275 ;
        RECT 39.555 124.935 40.270 125.105 ;
        RECT 40.460 124.985 41.185 125.155 ;
        RECT 41.355 124.985 41.625 125.955 ;
        RECT 30.800 124.565 37.920 124.815 ;
        RECT 29.465 124.225 36.210 124.395 ;
        RECT 28.225 123.575 28.475 124.035 ;
        RECT 28.645 123.745 29.205 124.035 ;
        RECT 29.465 123.575 29.765 124.055 ;
        RECT 29.935 123.770 30.195 124.225 ;
        RECT 30.365 123.575 30.625 124.055 ;
        RECT 30.805 123.770 31.065 124.225 ;
        RECT 31.235 123.575 31.485 124.055 ;
        RECT 31.665 123.770 31.925 124.225 ;
        RECT 32.095 123.575 32.345 124.055 ;
        RECT 32.525 123.770 32.785 124.225 ;
        RECT 32.955 123.575 33.200 124.055 ;
        RECT 33.370 123.770 33.645 124.225 ;
        RECT 33.815 123.575 34.060 124.055 ;
        RECT 34.230 123.770 34.490 124.225 ;
        RECT 34.660 123.575 34.920 124.055 ;
        RECT 35.090 123.770 35.350 124.225 ;
        RECT 35.520 123.575 35.780 124.055 ;
        RECT 35.950 123.770 36.210 124.225 ;
        RECT 36.380 123.575 36.640 124.135 ;
        RECT 36.810 123.755 37.060 124.565 ;
        RECT 37.240 123.575 37.500 124.100 ;
        RECT 37.670 123.755 37.920 124.565 ;
        RECT 38.090 124.255 38.405 124.815 ;
        RECT 39.040 124.245 39.390 124.815 ;
        RECT 39.560 124.485 40.270 124.935 ;
        RECT 41.015 124.815 41.185 124.985 ;
        RECT 40.440 124.485 40.845 124.815 ;
        RECT 41.015 124.485 41.285 124.815 ;
        RECT 41.015 124.315 41.185 124.485 ;
        RECT 39.575 124.145 41.185 124.315 ;
        RECT 41.455 124.250 41.625 124.985 ;
        RECT 38.100 123.575 38.405 124.085 ;
        RECT 39.045 123.575 39.375 124.075 ;
        RECT 39.575 123.795 39.745 124.145 ;
        RECT 39.945 123.575 40.275 123.975 ;
        RECT 40.445 123.795 40.615 124.145 ;
        RECT 40.785 123.575 41.165 123.975 ;
        RECT 41.355 123.905 41.625 124.250 ;
        RECT 41.795 124.985 42.065 125.955 ;
        RECT 42.275 125.325 42.555 126.125 ;
        RECT 42.725 125.615 44.380 125.905 ;
        RECT 42.790 125.275 44.380 125.445 ;
        RECT 42.790 125.155 42.960 125.275 ;
        RECT 42.235 124.985 42.960 125.155 ;
        RECT 41.795 124.250 41.965 124.985 ;
        RECT 42.235 124.815 42.405 124.985 ;
        RECT 43.150 124.935 43.865 125.105 ;
        RECT 44.060 124.985 44.380 125.275 ;
        RECT 44.555 124.985 44.895 125.955 ;
        RECT 45.065 124.985 45.235 126.125 ;
        RECT 45.505 125.325 45.755 126.125 ;
        RECT 46.400 125.155 46.730 125.955 ;
        RECT 47.030 125.325 47.360 126.125 ;
        RECT 47.530 125.155 47.860 125.955 ;
        RECT 45.425 124.985 47.860 125.155 ;
        RECT 42.135 124.485 42.405 124.815 ;
        RECT 42.575 124.485 42.980 124.815 ;
        RECT 43.150 124.485 43.860 124.935 ;
        RECT 42.235 124.315 42.405 124.485 ;
        RECT 41.795 123.905 42.065 124.250 ;
        RECT 42.235 124.145 43.845 124.315 ;
        RECT 44.030 124.245 44.380 124.815 ;
        RECT 44.555 124.425 44.730 124.985 ;
        RECT 45.425 124.735 45.595 124.985 ;
        RECT 44.900 124.565 45.595 124.735 ;
        RECT 45.770 124.565 46.190 124.765 ;
        RECT 46.360 124.565 46.690 124.765 ;
        RECT 46.860 124.565 47.190 124.765 ;
        RECT 44.555 124.375 44.785 124.425 ;
        RECT 42.255 123.575 42.635 123.975 ;
        RECT 42.805 123.795 42.975 124.145 ;
        RECT 43.145 123.575 43.475 123.975 ;
        RECT 43.675 123.795 43.845 124.145 ;
        RECT 44.045 123.575 44.375 124.075 ;
        RECT 44.555 123.745 44.895 124.375 ;
        RECT 45.065 123.575 45.315 124.375 ;
        RECT 45.505 124.225 46.730 124.395 ;
        RECT 45.505 123.745 45.835 124.225 ;
        RECT 46.005 123.575 46.230 124.035 ;
        RECT 46.400 123.745 46.730 124.225 ;
        RECT 47.360 124.355 47.530 124.985 ;
        RECT 48.235 124.960 48.525 126.125 ;
        RECT 49.615 124.985 49.955 125.955 ;
        RECT 50.125 124.985 50.295 126.125 ;
        RECT 50.565 125.325 50.815 126.125 ;
        RECT 51.460 125.155 51.790 125.955 ;
        RECT 52.090 125.325 52.420 126.125 ;
        RECT 52.590 125.155 52.920 125.955 ;
        RECT 50.485 124.985 52.920 125.155 ;
        RECT 54.215 125.035 57.725 126.125 ;
        RECT 58.270 125.145 58.525 125.815 ;
        RECT 58.705 125.325 58.990 126.125 ;
        RECT 59.170 125.405 59.500 125.915 ;
        RECT 58.270 125.105 58.450 125.145 ;
        RECT 47.715 124.565 48.065 124.815 ;
        RECT 49.615 124.375 49.790 124.985 ;
        RECT 50.485 124.735 50.655 124.985 ;
        RECT 49.960 124.565 50.655 124.735 ;
        RECT 50.830 124.565 51.250 124.765 ;
        RECT 51.420 124.565 51.750 124.765 ;
        RECT 51.920 124.565 52.250 124.765 ;
        RECT 47.360 123.745 47.860 124.355 ;
        RECT 48.235 123.575 48.525 124.300 ;
        RECT 49.615 123.745 49.955 124.375 ;
        RECT 50.125 123.575 50.375 124.375 ;
        RECT 50.565 124.225 51.790 124.395 ;
        RECT 50.565 123.745 50.895 124.225 ;
        RECT 51.065 123.575 51.290 124.035 ;
        RECT 51.460 123.745 51.790 124.225 ;
        RECT 52.420 124.355 52.590 124.985 ;
        RECT 52.775 124.565 53.125 124.815 ;
        RECT 54.215 124.515 55.905 125.035 ;
        RECT 58.185 124.935 58.450 125.105 ;
        RECT 52.420 123.745 52.920 124.355 ;
        RECT 56.075 124.345 57.725 124.865 ;
        RECT 54.215 123.575 57.725 124.345 ;
        RECT 58.270 124.285 58.450 124.935 ;
        RECT 59.170 124.815 59.420 125.405 ;
        RECT 59.770 125.255 59.940 125.865 ;
        RECT 60.110 125.435 60.440 126.125 ;
        RECT 60.670 125.575 60.910 125.865 ;
        RECT 61.110 125.745 61.530 126.125 ;
        RECT 61.710 125.655 62.340 125.905 ;
        RECT 62.810 125.745 63.140 126.125 ;
        RECT 61.710 125.575 61.880 125.655 ;
        RECT 63.310 125.575 63.480 125.865 ;
        RECT 63.660 125.745 64.040 126.125 ;
        RECT 64.280 125.740 65.110 125.910 ;
        RECT 60.670 125.405 61.880 125.575 ;
        RECT 58.620 124.485 59.420 124.815 ;
        RECT 58.270 123.755 58.525 124.285 ;
        RECT 58.705 123.575 58.990 124.035 ;
        RECT 59.170 123.835 59.420 124.485 ;
        RECT 59.620 125.235 59.940 125.255 ;
        RECT 59.620 125.065 61.540 125.235 ;
        RECT 59.620 124.170 59.810 125.065 ;
        RECT 61.710 124.895 61.880 125.405 ;
        RECT 62.050 125.145 62.570 125.455 ;
        RECT 59.980 124.725 61.880 124.895 ;
        RECT 59.980 124.665 60.310 124.725 ;
        RECT 60.460 124.495 60.790 124.555 ;
        RECT 60.130 124.225 60.790 124.495 ;
        RECT 59.620 123.840 59.940 124.170 ;
        RECT 60.120 123.575 60.780 124.055 ;
        RECT 60.980 123.965 61.150 124.725 ;
        RECT 62.050 124.555 62.230 124.965 ;
        RECT 61.320 124.385 61.650 124.505 ;
        RECT 62.400 124.385 62.570 125.145 ;
        RECT 61.320 124.215 62.570 124.385 ;
        RECT 62.740 125.325 64.110 125.575 ;
        RECT 62.740 124.555 62.930 125.325 ;
        RECT 63.860 125.065 64.110 125.325 ;
        RECT 63.100 124.895 63.350 125.055 ;
        RECT 64.280 124.895 64.450 125.740 ;
        RECT 65.345 125.455 65.515 125.955 ;
        RECT 65.685 125.625 66.015 126.125 ;
        RECT 64.620 125.065 65.120 125.445 ;
        RECT 65.345 125.285 66.040 125.455 ;
        RECT 63.100 124.725 64.450 124.895 ;
        RECT 64.030 124.685 64.450 124.725 ;
        RECT 62.740 124.215 63.160 124.555 ;
        RECT 63.450 124.225 63.860 124.555 ;
        RECT 60.980 123.795 61.830 123.965 ;
        RECT 62.390 123.575 62.710 124.035 ;
        RECT 62.910 123.785 63.160 124.215 ;
        RECT 63.450 123.575 63.860 124.015 ;
        RECT 64.030 123.955 64.200 124.685 ;
        RECT 64.370 124.135 64.720 124.505 ;
        RECT 64.900 124.195 65.120 125.065 ;
        RECT 65.290 124.495 65.700 125.115 ;
        RECT 65.870 124.315 66.040 125.285 ;
        RECT 65.345 124.125 66.040 124.315 ;
        RECT 64.030 123.755 65.045 123.955 ;
        RECT 65.345 123.795 65.515 124.125 ;
        RECT 65.685 123.575 66.015 123.955 ;
        RECT 66.230 123.835 66.455 125.955 ;
        RECT 66.625 125.625 66.955 126.125 ;
        RECT 67.125 125.455 67.295 125.955 ;
        RECT 66.630 125.285 67.295 125.455 ;
        RECT 66.630 124.295 66.860 125.285 ;
        RECT 67.030 124.465 67.380 125.115 ;
        RECT 68.015 125.035 70.605 126.125 ;
        RECT 70.775 125.155 71.085 125.955 ;
        RECT 71.255 125.325 71.565 126.125 ;
        RECT 71.735 125.495 71.995 125.955 ;
        RECT 72.165 125.665 72.420 126.125 ;
        RECT 72.595 125.495 72.855 125.955 ;
        RECT 71.735 125.325 72.855 125.495 ;
        RECT 68.015 124.515 69.225 125.035 ;
        RECT 70.775 124.985 71.805 125.155 ;
        RECT 69.395 124.345 70.605 124.865 ;
        RECT 66.630 124.125 67.295 124.295 ;
        RECT 66.625 123.575 66.955 123.955 ;
        RECT 67.125 123.835 67.295 124.125 ;
        RECT 68.015 123.575 70.605 124.345 ;
        RECT 70.775 124.075 70.945 124.985 ;
        RECT 71.115 124.245 71.465 124.815 ;
        RECT 71.635 124.735 71.805 124.985 ;
        RECT 72.595 125.075 72.855 125.325 ;
        RECT 73.025 125.255 73.310 126.125 ;
        RECT 72.595 124.905 73.350 125.075 ;
        RECT 73.995 124.960 74.285 126.125 ;
        RECT 74.915 125.035 77.505 126.125 ;
        RECT 77.675 125.405 78.135 125.955 ;
        RECT 78.325 125.405 78.655 126.125 ;
        RECT 71.635 124.565 72.775 124.735 ;
        RECT 72.945 124.395 73.350 124.905 ;
        RECT 74.915 124.515 76.125 125.035 ;
        RECT 71.700 124.225 73.350 124.395 ;
        RECT 76.295 124.345 77.505 124.865 ;
        RECT 70.775 123.745 71.075 124.075 ;
        RECT 71.245 123.575 71.520 124.055 ;
        RECT 71.700 123.835 71.995 124.225 ;
        RECT 72.165 123.575 72.420 124.055 ;
        RECT 72.595 123.835 72.855 124.225 ;
        RECT 73.025 123.575 73.305 124.055 ;
        RECT 73.995 123.575 74.285 124.300 ;
        RECT 74.915 123.575 77.505 124.345 ;
        RECT 77.675 124.035 77.925 125.405 ;
        RECT 78.855 125.235 79.155 125.785 ;
        RECT 79.325 125.455 79.605 126.125 ;
        RECT 78.215 125.065 79.155 125.235 ;
        RECT 78.215 124.815 78.385 125.065 ;
        RECT 79.525 124.815 79.790 125.175 ;
        RECT 78.095 124.485 78.385 124.815 ;
        RECT 78.555 124.565 78.895 124.815 ;
        RECT 79.115 124.565 79.790 124.815 ;
        RECT 80.435 125.035 83.945 126.125 ;
        RECT 84.205 125.380 84.475 126.125 ;
        RECT 85.105 126.120 91.380 126.125 ;
        RECT 84.645 125.210 84.935 125.950 ;
        RECT 85.105 125.395 85.360 126.120 ;
        RECT 85.545 125.225 85.805 125.950 ;
        RECT 85.975 125.395 86.220 126.120 ;
        RECT 86.405 125.225 86.665 125.950 ;
        RECT 86.835 125.395 87.080 126.120 ;
        RECT 87.265 125.225 87.525 125.950 ;
        RECT 87.695 125.395 87.940 126.120 ;
        RECT 88.110 125.225 88.370 125.950 ;
        RECT 88.540 125.395 88.800 126.120 ;
        RECT 88.970 125.225 89.230 125.950 ;
        RECT 89.400 125.395 89.660 126.120 ;
        RECT 89.830 125.225 90.090 125.950 ;
        RECT 90.260 125.395 90.520 126.120 ;
        RECT 90.690 125.225 90.950 125.950 ;
        RECT 91.120 125.325 91.380 126.120 ;
        RECT 85.545 125.210 90.950 125.225 ;
        RECT 80.435 124.515 82.125 125.035 ;
        RECT 84.205 124.985 90.950 125.210 ;
        RECT 78.215 124.395 78.385 124.485 ;
        RECT 78.215 124.205 79.605 124.395 ;
        RECT 82.295 124.345 83.945 124.865 ;
        RECT 77.675 123.745 78.235 124.035 ;
        RECT 78.405 123.575 78.655 124.035 ;
        RECT 79.275 123.845 79.605 124.205 ;
        RECT 80.435 123.575 83.945 124.345 ;
        RECT 84.205 124.395 85.370 124.985 ;
        RECT 91.550 124.815 91.800 125.950 ;
        RECT 91.980 125.315 92.240 126.125 ;
        RECT 92.415 124.815 92.660 125.955 ;
        RECT 92.840 125.315 93.135 126.125 ;
        RECT 94.240 125.690 99.585 126.125 ;
        RECT 85.540 124.565 92.660 124.815 ;
        RECT 84.205 124.225 90.950 124.395 ;
        RECT 84.205 123.575 84.505 124.055 ;
        RECT 84.675 123.770 84.935 124.225 ;
        RECT 85.105 123.575 85.365 124.055 ;
        RECT 85.545 123.770 85.805 124.225 ;
        RECT 85.975 123.575 86.225 124.055 ;
        RECT 86.405 123.770 86.665 124.225 ;
        RECT 86.835 123.575 87.085 124.055 ;
        RECT 87.265 123.770 87.525 124.225 ;
        RECT 87.695 123.575 87.940 124.055 ;
        RECT 88.110 123.770 88.385 124.225 ;
        RECT 88.555 123.575 88.800 124.055 ;
        RECT 88.970 123.770 89.230 124.225 ;
        RECT 89.400 123.575 89.660 124.055 ;
        RECT 89.830 123.770 90.090 124.225 ;
        RECT 90.260 123.575 90.520 124.055 ;
        RECT 90.690 123.770 90.950 124.225 ;
        RECT 91.120 123.575 91.380 124.135 ;
        RECT 91.550 123.755 91.800 124.565 ;
        RECT 91.980 123.575 92.240 124.100 ;
        RECT 92.410 123.755 92.660 124.565 ;
        RECT 92.830 124.255 93.145 124.815 ;
        RECT 95.830 124.440 96.180 125.690 ;
        RECT 99.755 124.960 100.045 126.125 ;
        RECT 100.215 125.365 100.730 125.775 ;
        RECT 100.965 125.365 101.135 126.125 ;
        RECT 101.305 125.785 103.335 125.955 ;
        RECT 97.660 124.120 98.000 124.950 ;
        RECT 100.215 124.555 100.555 125.365 ;
        RECT 101.305 125.120 101.475 125.785 ;
        RECT 101.870 125.445 102.995 125.615 ;
        RECT 100.725 124.930 101.475 125.120 ;
        RECT 101.645 125.105 102.655 125.275 ;
        RECT 100.215 124.385 101.445 124.555 ;
        RECT 92.840 123.575 93.145 124.085 ;
        RECT 94.240 123.575 99.585 124.120 ;
        RECT 99.755 123.575 100.045 124.300 ;
        RECT 100.490 123.780 100.735 124.385 ;
        RECT 100.955 123.575 101.465 124.110 ;
        RECT 101.645 123.745 101.835 125.105 ;
        RECT 102.005 124.085 102.280 124.905 ;
        RECT 102.485 124.305 102.655 125.105 ;
        RECT 102.825 124.315 102.995 125.445 ;
        RECT 103.165 124.815 103.335 125.785 ;
        RECT 103.505 124.985 103.675 126.125 ;
        RECT 103.845 124.985 104.180 125.955 ;
        RECT 104.905 125.195 105.075 125.955 ;
        RECT 105.255 125.365 105.585 126.125 ;
        RECT 104.905 125.025 105.570 125.195 ;
        RECT 105.755 125.050 106.025 125.955 ;
        RECT 103.165 124.485 103.360 124.815 ;
        RECT 103.585 124.485 103.840 124.815 ;
        RECT 103.585 124.315 103.755 124.485 ;
        RECT 104.010 124.315 104.180 124.985 ;
        RECT 105.400 124.880 105.570 125.025 ;
        RECT 104.835 124.475 105.165 124.845 ;
        RECT 105.400 124.550 105.685 124.880 ;
        RECT 102.825 124.145 103.755 124.315 ;
        RECT 102.825 124.110 103.000 124.145 ;
        RECT 102.005 123.915 102.285 124.085 ;
        RECT 102.005 123.745 102.280 123.915 ;
        RECT 102.470 123.745 103.000 124.110 ;
        RECT 103.425 123.575 103.755 123.975 ;
        RECT 103.925 123.745 104.180 124.315 ;
        RECT 105.400 124.295 105.570 124.550 ;
        RECT 104.905 124.125 105.570 124.295 ;
        RECT 105.855 124.250 106.025 125.050 ;
        RECT 106.195 125.035 107.865 126.125 ;
        RECT 108.035 125.365 108.550 125.775 ;
        RECT 108.785 125.365 108.955 126.125 ;
        RECT 109.125 125.785 111.155 125.955 ;
        RECT 106.195 124.515 106.945 125.035 ;
        RECT 107.115 124.345 107.865 124.865 ;
        RECT 108.035 124.555 108.375 125.365 ;
        RECT 109.125 125.120 109.295 125.785 ;
        RECT 109.690 125.445 110.815 125.615 ;
        RECT 108.545 124.930 109.295 125.120 ;
        RECT 109.465 125.105 110.475 125.275 ;
        RECT 108.035 124.385 109.265 124.555 ;
        RECT 104.905 123.745 105.075 124.125 ;
        RECT 105.255 123.575 105.585 123.955 ;
        RECT 105.765 123.745 106.025 124.250 ;
        RECT 106.195 123.575 107.865 124.345 ;
        RECT 108.310 123.780 108.555 124.385 ;
        RECT 108.775 123.575 109.285 124.110 ;
        RECT 109.465 123.745 109.655 125.105 ;
        RECT 109.825 124.765 110.100 124.905 ;
        RECT 109.825 124.595 110.105 124.765 ;
        RECT 109.825 123.745 110.100 124.595 ;
        RECT 110.305 124.305 110.475 125.105 ;
        RECT 110.645 124.315 110.815 125.445 ;
        RECT 110.985 124.815 111.155 125.785 ;
        RECT 111.325 124.985 111.495 126.125 ;
        RECT 111.665 124.985 112.000 125.955 ;
        RECT 110.985 124.485 111.180 124.815 ;
        RECT 111.405 124.485 111.660 124.815 ;
        RECT 111.405 124.315 111.575 124.485 ;
        RECT 111.830 124.315 112.000 124.985 ;
        RECT 112.550 125.145 112.805 125.815 ;
        RECT 112.985 125.325 113.270 126.125 ;
        RECT 113.450 125.405 113.780 125.915 ;
        RECT 112.550 124.765 112.730 125.145 ;
        RECT 113.450 124.815 113.700 125.405 ;
        RECT 114.050 125.255 114.220 125.865 ;
        RECT 114.390 125.435 114.720 126.125 ;
        RECT 114.950 125.575 115.190 125.865 ;
        RECT 115.390 125.745 115.810 126.125 ;
        RECT 115.990 125.655 116.620 125.905 ;
        RECT 117.090 125.745 117.420 126.125 ;
        RECT 115.990 125.575 116.160 125.655 ;
        RECT 117.590 125.575 117.760 125.865 ;
        RECT 117.940 125.745 118.320 126.125 ;
        RECT 118.560 125.740 119.390 125.910 ;
        RECT 114.950 125.405 116.160 125.575 ;
        RECT 112.465 124.595 112.730 124.765 ;
        RECT 110.645 124.145 111.575 124.315 ;
        RECT 110.645 124.110 110.820 124.145 ;
        RECT 110.290 123.745 110.820 124.110 ;
        RECT 111.245 123.575 111.575 123.975 ;
        RECT 111.745 123.745 112.000 124.315 ;
        RECT 112.550 124.285 112.730 124.595 ;
        RECT 112.900 124.485 113.700 124.815 ;
        RECT 112.550 123.755 112.805 124.285 ;
        RECT 112.985 123.575 113.270 124.035 ;
        RECT 113.450 123.835 113.700 124.485 ;
        RECT 113.900 125.235 114.220 125.255 ;
        RECT 113.900 125.065 115.820 125.235 ;
        RECT 113.900 124.170 114.090 125.065 ;
        RECT 115.990 124.895 116.160 125.405 ;
        RECT 116.330 125.145 116.850 125.455 ;
        RECT 114.260 124.725 116.160 124.895 ;
        RECT 114.260 124.665 114.590 124.725 ;
        RECT 114.740 124.495 115.070 124.555 ;
        RECT 114.410 124.225 115.070 124.495 ;
        RECT 113.900 123.840 114.220 124.170 ;
        RECT 114.400 123.575 115.060 124.055 ;
        RECT 115.260 123.965 115.430 124.725 ;
        RECT 116.330 124.555 116.510 124.965 ;
        RECT 115.600 124.385 115.930 124.505 ;
        RECT 116.680 124.385 116.850 125.145 ;
        RECT 115.600 124.215 116.850 124.385 ;
        RECT 117.020 125.325 118.390 125.575 ;
        RECT 117.020 124.555 117.210 125.325 ;
        RECT 118.140 125.065 118.390 125.325 ;
        RECT 117.380 124.895 117.630 125.055 ;
        RECT 118.560 124.895 118.730 125.740 ;
        RECT 119.625 125.455 119.795 125.955 ;
        RECT 119.965 125.625 120.295 126.125 ;
        RECT 118.900 125.065 119.400 125.445 ;
        RECT 119.625 125.285 120.320 125.455 ;
        RECT 117.380 124.725 118.730 124.895 ;
        RECT 118.310 124.685 118.730 124.725 ;
        RECT 117.020 124.215 117.440 124.555 ;
        RECT 117.730 124.225 118.140 124.555 ;
        RECT 115.260 123.795 116.110 123.965 ;
        RECT 116.670 123.575 116.990 124.035 ;
        RECT 117.190 123.785 117.440 124.215 ;
        RECT 117.730 123.575 118.140 124.015 ;
        RECT 118.310 123.955 118.480 124.685 ;
        RECT 118.650 124.135 119.000 124.505 ;
        RECT 119.180 124.195 119.400 125.065 ;
        RECT 119.570 124.495 119.980 125.115 ;
        RECT 120.150 124.315 120.320 125.285 ;
        RECT 119.625 124.125 120.320 124.315 ;
        RECT 118.310 123.755 119.325 123.955 ;
        RECT 119.625 123.795 119.795 124.125 ;
        RECT 119.965 123.575 120.295 123.955 ;
        RECT 120.510 123.835 120.735 125.955 ;
        RECT 120.905 125.625 121.235 126.125 ;
        RECT 121.405 125.455 121.575 125.955 ;
        RECT 120.910 125.285 121.575 125.455 ;
        RECT 120.910 124.295 121.140 125.285 ;
        RECT 121.310 124.465 121.660 125.115 ;
        RECT 121.835 125.050 122.105 125.955 ;
        RECT 122.275 125.365 122.605 126.125 ;
        RECT 122.785 125.195 122.955 125.955 ;
        RECT 120.910 124.125 121.575 124.295 ;
        RECT 120.905 123.575 121.235 123.955 ;
        RECT 121.405 123.835 121.575 124.125 ;
        RECT 121.835 124.250 122.005 125.050 ;
        RECT 122.290 125.025 122.955 125.195 ;
        RECT 123.215 125.050 123.485 125.955 ;
        RECT 123.655 125.365 123.985 126.125 ;
        RECT 124.165 125.195 124.335 125.955 ;
        RECT 122.290 124.880 122.460 125.025 ;
        RECT 122.175 124.550 122.460 124.880 ;
        RECT 122.290 124.295 122.460 124.550 ;
        RECT 122.695 124.475 123.025 124.845 ;
        RECT 121.835 123.745 122.095 124.250 ;
        RECT 122.290 124.125 122.955 124.295 ;
        RECT 122.275 123.575 122.605 123.955 ;
        RECT 122.785 123.745 122.955 124.125 ;
        RECT 123.215 124.250 123.385 125.050 ;
        RECT 123.670 125.025 124.335 125.195 ;
        RECT 124.595 125.035 125.805 126.125 ;
        RECT 123.670 124.880 123.840 125.025 ;
        RECT 123.555 124.550 123.840 124.880 ;
        RECT 123.670 124.295 123.840 124.550 ;
        RECT 124.075 124.475 124.405 124.845 ;
        RECT 124.595 124.495 125.115 125.035 ;
        RECT 125.285 124.325 125.805 124.865 ;
        RECT 123.215 123.745 123.475 124.250 ;
        RECT 123.670 124.125 124.335 124.295 ;
        RECT 123.655 123.575 123.985 123.955 ;
        RECT 124.165 123.745 124.335 124.125 ;
        RECT 124.595 123.575 125.805 124.325 ;
        RECT 11.810 123.405 125.890 123.575 ;
        RECT 11.895 122.655 13.105 123.405 ;
        RECT 13.275 122.655 14.485 123.405 ;
        RECT 11.895 122.115 12.415 122.655 ;
        RECT 12.585 121.945 13.105 122.485 ;
        RECT 11.895 120.855 13.105 121.945 ;
        RECT 13.275 121.945 13.795 122.485 ;
        RECT 13.965 122.115 14.485 122.655 ;
        RECT 15.030 122.695 15.285 123.225 ;
        RECT 15.465 122.945 15.750 123.405 ;
        RECT 15.030 122.385 15.210 122.695 ;
        RECT 15.930 122.495 16.180 123.145 ;
        RECT 14.945 122.215 15.210 122.385 ;
        RECT 13.275 120.855 14.485 121.945 ;
        RECT 15.030 121.835 15.210 122.215 ;
        RECT 15.380 122.165 16.180 122.495 ;
        RECT 15.030 121.165 15.285 121.835 ;
        RECT 15.465 120.855 15.750 121.655 ;
        RECT 15.930 121.575 16.180 122.165 ;
        RECT 16.380 122.810 16.700 123.140 ;
        RECT 16.880 122.925 17.540 123.405 ;
        RECT 17.740 123.015 18.590 123.185 ;
        RECT 16.380 121.915 16.570 122.810 ;
        RECT 16.890 122.485 17.550 122.755 ;
        RECT 17.220 122.425 17.550 122.485 ;
        RECT 16.740 122.255 17.070 122.315 ;
        RECT 17.740 122.255 17.910 123.015 ;
        RECT 19.150 122.945 19.470 123.405 ;
        RECT 19.670 122.765 19.920 123.195 ;
        RECT 20.210 122.965 20.620 123.405 ;
        RECT 20.790 123.025 21.805 123.225 ;
        RECT 18.080 122.595 19.330 122.765 ;
        RECT 18.080 122.475 18.410 122.595 ;
        RECT 16.740 122.085 18.640 122.255 ;
        RECT 16.380 121.745 18.300 121.915 ;
        RECT 16.380 121.725 16.700 121.745 ;
        RECT 15.930 121.065 16.260 121.575 ;
        RECT 16.530 121.115 16.700 121.725 ;
        RECT 18.470 121.575 18.640 122.085 ;
        RECT 18.810 122.015 18.990 122.425 ;
        RECT 19.160 121.835 19.330 122.595 ;
        RECT 16.870 120.855 17.200 121.545 ;
        RECT 17.430 121.405 18.640 121.575 ;
        RECT 18.810 121.525 19.330 121.835 ;
        RECT 19.500 122.425 19.920 122.765 ;
        RECT 20.210 122.425 20.620 122.755 ;
        RECT 19.500 121.655 19.690 122.425 ;
        RECT 20.790 122.295 20.960 123.025 ;
        RECT 22.105 122.855 22.275 123.185 ;
        RECT 22.445 123.025 22.775 123.405 ;
        RECT 21.130 122.475 21.480 122.845 ;
        RECT 20.790 122.255 21.210 122.295 ;
        RECT 19.860 122.085 21.210 122.255 ;
        RECT 19.860 121.925 20.110 122.085 ;
        RECT 20.620 121.655 20.870 121.915 ;
        RECT 19.500 121.405 20.870 121.655 ;
        RECT 17.430 121.115 17.670 121.405 ;
        RECT 18.470 121.325 18.640 121.405 ;
        RECT 17.870 120.855 18.290 121.235 ;
        RECT 18.470 121.075 19.100 121.325 ;
        RECT 19.570 120.855 19.900 121.235 ;
        RECT 20.070 121.115 20.240 121.405 ;
        RECT 21.040 121.240 21.210 122.085 ;
        RECT 21.660 121.915 21.880 122.785 ;
        RECT 22.105 122.665 22.800 122.855 ;
        RECT 21.380 121.535 21.880 121.915 ;
        RECT 22.050 121.865 22.460 122.485 ;
        RECT 22.630 121.695 22.800 122.665 ;
        RECT 22.105 121.525 22.800 121.695 ;
        RECT 20.420 120.855 20.800 121.235 ;
        RECT 21.040 121.070 21.870 121.240 ;
        RECT 22.105 121.025 22.275 121.525 ;
        RECT 22.445 120.855 22.775 121.355 ;
        RECT 22.990 121.025 23.215 123.145 ;
        RECT 23.385 123.025 23.715 123.405 ;
        RECT 23.885 122.855 24.055 123.145 ;
        RECT 23.390 122.685 24.055 122.855 ;
        RECT 25.610 122.695 25.865 123.225 ;
        RECT 26.045 122.945 26.330 123.405 ;
        RECT 23.390 121.695 23.620 122.685 ;
        RECT 23.790 121.865 24.140 122.515 ;
        RECT 25.610 122.045 25.790 122.695 ;
        RECT 26.510 122.495 26.760 123.145 ;
        RECT 25.960 122.165 26.760 122.495 ;
        RECT 25.525 121.875 25.790 122.045 ;
        RECT 25.610 121.835 25.790 121.875 ;
        RECT 23.390 121.525 24.055 121.695 ;
        RECT 23.385 120.855 23.715 121.355 ;
        RECT 23.885 121.025 24.055 121.525 ;
        RECT 25.610 121.165 25.865 121.835 ;
        RECT 26.045 120.855 26.330 121.655 ;
        RECT 26.510 121.575 26.760 122.165 ;
        RECT 26.960 122.810 27.280 123.140 ;
        RECT 27.460 122.925 28.120 123.405 ;
        RECT 28.320 123.015 29.170 123.185 ;
        RECT 26.960 121.915 27.150 122.810 ;
        RECT 27.470 122.485 28.130 122.755 ;
        RECT 27.800 122.425 28.130 122.485 ;
        RECT 27.320 122.255 27.650 122.315 ;
        RECT 28.320 122.255 28.490 123.015 ;
        RECT 29.730 122.945 30.050 123.405 ;
        RECT 30.250 122.765 30.500 123.195 ;
        RECT 30.790 122.965 31.200 123.405 ;
        RECT 31.370 123.025 32.385 123.225 ;
        RECT 28.660 122.595 29.910 122.765 ;
        RECT 28.660 122.475 28.990 122.595 ;
        RECT 27.320 122.085 29.220 122.255 ;
        RECT 26.960 121.745 28.880 121.915 ;
        RECT 26.960 121.725 27.280 121.745 ;
        RECT 26.510 121.065 26.840 121.575 ;
        RECT 27.110 121.115 27.280 121.725 ;
        RECT 29.050 121.575 29.220 122.085 ;
        RECT 29.390 122.015 29.570 122.425 ;
        RECT 29.740 121.835 29.910 122.595 ;
        RECT 27.450 120.855 27.780 121.545 ;
        RECT 28.010 121.405 29.220 121.575 ;
        RECT 29.390 121.525 29.910 121.835 ;
        RECT 30.080 122.425 30.500 122.765 ;
        RECT 30.790 122.425 31.200 122.755 ;
        RECT 30.080 121.655 30.270 122.425 ;
        RECT 31.370 122.295 31.540 123.025 ;
        RECT 32.685 122.855 32.855 123.185 ;
        RECT 33.025 123.025 33.355 123.405 ;
        RECT 31.710 122.475 32.060 122.845 ;
        RECT 31.370 122.255 31.790 122.295 ;
        RECT 30.440 122.085 31.790 122.255 ;
        RECT 30.440 121.925 30.690 122.085 ;
        RECT 31.200 121.655 31.450 121.915 ;
        RECT 30.080 121.405 31.450 121.655 ;
        RECT 28.010 121.115 28.250 121.405 ;
        RECT 29.050 121.325 29.220 121.405 ;
        RECT 28.450 120.855 28.870 121.235 ;
        RECT 29.050 121.075 29.680 121.325 ;
        RECT 30.150 120.855 30.480 121.235 ;
        RECT 30.650 121.115 30.820 121.405 ;
        RECT 31.620 121.240 31.790 122.085 ;
        RECT 32.240 121.915 32.460 122.785 ;
        RECT 32.685 122.665 33.380 122.855 ;
        RECT 31.960 121.535 32.460 121.915 ;
        RECT 32.630 121.865 33.040 122.485 ;
        RECT 33.210 121.695 33.380 122.665 ;
        RECT 32.685 121.525 33.380 121.695 ;
        RECT 31.000 120.855 31.380 121.235 ;
        RECT 31.620 121.070 32.450 121.240 ;
        RECT 32.685 121.025 32.855 121.525 ;
        RECT 33.025 120.855 33.355 121.355 ;
        RECT 33.570 121.025 33.795 123.145 ;
        RECT 33.965 123.025 34.295 123.405 ;
        RECT 34.465 122.855 34.635 123.145 ;
        RECT 33.970 122.685 34.635 122.855 ;
        RECT 33.970 121.695 34.200 122.685 ;
        RECT 35.355 122.680 35.645 123.405 ;
        RECT 35.965 122.605 36.295 123.405 ;
        RECT 36.465 122.755 36.635 123.235 ;
        RECT 36.805 122.925 37.135 123.405 ;
        RECT 37.305 122.755 37.475 123.235 ;
        RECT 37.725 122.925 37.965 123.405 ;
        RECT 38.145 122.755 38.315 123.235 ;
        RECT 36.465 122.585 37.475 122.755 ;
        RECT 37.680 122.585 38.315 122.755 ;
        RECT 38.665 122.855 38.835 123.235 ;
        RECT 39.015 123.025 39.345 123.405 ;
        RECT 38.665 122.685 39.330 122.855 ;
        RECT 39.525 122.730 39.785 123.235 ;
        RECT 36.465 122.555 36.965 122.585 ;
        RECT 34.370 121.865 34.720 122.515 ;
        RECT 36.465 122.045 36.960 122.555 ;
        RECT 37.680 122.415 37.850 122.585 ;
        RECT 37.350 122.245 37.850 122.415 ;
        RECT 33.970 121.525 34.635 121.695 ;
        RECT 33.965 120.855 34.295 121.355 ;
        RECT 34.465 121.025 34.635 121.525 ;
        RECT 35.355 120.855 35.645 122.020 ;
        RECT 35.965 120.855 36.295 122.005 ;
        RECT 36.465 121.875 37.475 122.045 ;
        RECT 36.465 121.025 36.635 121.875 ;
        RECT 36.805 120.855 37.135 121.655 ;
        RECT 37.305 121.025 37.475 121.875 ;
        RECT 37.680 122.005 37.850 122.245 ;
        RECT 38.020 122.175 38.400 122.415 ;
        RECT 38.595 122.135 38.925 122.505 ;
        RECT 39.160 122.430 39.330 122.685 ;
        RECT 39.160 122.100 39.445 122.430 ;
        RECT 37.680 121.835 38.395 122.005 ;
        RECT 39.160 121.955 39.330 122.100 ;
        RECT 37.655 120.855 37.895 121.655 ;
        RECT 38.065 121.025 38.395 121.835 ;
        RECT 38.665 121.785 39.330 121.955 ;
        RECT 39.615 121.930 39.785 122.730 ;
        RECT 38.665 121.025 38.835 121.785 ;
        RECT 39.015 120.855 39.345 121.615 ;
        RECT 39.515 121.025 39.785 121.930 ;
        RECT 40.415 122.945 40.975 123.235 ;
        RECT 41.145 122.945 41.395 123.405 ;
        RECT 40.415 121.575 40.665 122.945 ;
        RECT 42.015 122.775 42.345 123.135 ;
        RECT 40.955 122.585 42.345 122.775 ;
        RECT 42.915 122.775 43.245 123.135 ;
        RECT 43.865 122.945 44.115 123.405 ;
        RECT 44.285 122.945 44.845 123.235 ;
        RECT 42.915 122.585 44.305 122.775 ;
        RECT 40.955 122.495 41.125 122.585 ;
        RECT 40.835 122.165 41.125 122.495 ;
        RECT 44.135 122.495 44.305 122.585 ;
        RECT 41.295 122.165 41.635 122.415 ;
        RECT 41.855 122.165 42.530 122.415 ;
        RECT 40.955 121.915 41.125 122.165 ;
        RECT 40.955 121.745 41.895 121.915 ;
        RECT 42.265 121.805 42.530 122.165 ;
        RECT 42.730 122.165 43.405 122.415 ;
        RECT 43.625 122.165 43.965 122.415 ;
        RECT 44.135 122.165 44.425 122.495 ;
        RECT 42.730 121.805 42.995 122.165 ;
        RECT 44.135 121.915 44.305 122.165 ;
        RECT 40.415 121.025 40.875 121.575 ;
        RECT 41.065 120.855 41.395 121.575 ;
        RECT 41.595 121.195 41.895 121.745 ;
        RECT 43.365 121.745 44.305 121.915 ;
        RECT 42.065 120.855 42.345 121.525 ;
        RECT 42.915 120.855 43.195 121.525 ;
        RECT 43.365 121.195 43.665 121.745 ;
        RECT 44.595 121.575 44.845 122.945 ;
        RECT 45.475 122.895 45.780 123.405 ;
        RECT 45.475 122.165 45.790 122.725 ;
        RECT 45.960 122.415 46.210 123.225 ;
        RECT 46.380 122.880 46.640 123.405 ;
        RECT 46.820 122.415 47.070 123.225 ;
        RECT 47.240 122.845 47.500 123.405 ;
        RECT 47.670 122.755 47.930 123.210 ;
        RECT 48.100 122.925 48.360 123.405 ;
        RECT 48.530 122.755 48.790 123.210 ;
        RECT 48.960 122.925 49.220 123.405 ;
        RECT 49.390 122.755 49.650 123.210 ;
        RECT 49.820 122.925 50.065 123.405 ;
        RECT 50.235 122.755 50.510 123.210 ;
        RECT 50.680 122.925 50.925 123.405 ;
        RECT 51.095 122.755 51.355 123.210 ;
        RECT 51.535 122.925 51.785 123.405 ;
        RECT 51.955 122.755 52.215 123.210 ;
        RECT 52.395 122.925 52.645 123.405 ;
        RECT 52.815 122.755 53.075 123.210 ;
        RECT 53.255 122.925 53.515 123.405 ;
        RECT 53.685 122.755 53.945 123.210 ;
        RECT 54.115 122.925 54.415 123.405 ;
        RECT 47.670 122.585 54.415 122.755 ;
        RECT 54.675 122.635 56.345 123.405 ;
        RECT 45.960 122.165 53.080 122.415 ;
        RECT 43.865 120.855 44.195 121.575 ;
        RECT 44.385 121.025 44.845 121.575 ;
        RECT 45.485 120.855 45.780 121.665 ;
        RECT 45.960 121.025 46.205 122.165 ;
        RECT 46.380 120.855 46.640 121.665 ;
        RECT 46.820 121.030 47.070 122.165 ;
        RECT 53.250 121.995 54.415 122.585 ;
        RECT 47.670 121.770 54.415 121.995 ;
        RECT 54.675 121.945 55.425 122.465 ;
        RECT 55.595 122.115 56.345 122.635 ;
        RECT 56.790 122.595 57.035 123.200 ;
        RECT 57.255 122.870 57.765 123.405 ;
        RECT 56.515 122.425 57.745 122.595 ;
        RECT 47.670 121.755 53.075 121.770 ;
        RECT 47.240 120.860 47.500 121.655 ;
        RECT 47.670 121.030 47.930 121.755 ;
        RECT 48.100 120.860 48.360 121.585 ;
        RECT 48.530 121.030 48.790 121.755 ;
        RECT 48.960 120.860 49.220 121.585 ;
        RECT 49.390 121.030 49.650 121.755 ;
        RECT 49.820 120.860 50.080 121.585 ;
        RECT 50.250 121.030 50.510 121.755 ;
        RECT 50.680 120.860 50.925 121.585 ;
        RECT 51.095 121.030 51.355 121.755 ;
        RECT 51.540 120.860 51.785 121.585 ;
        RECT 51.955 121.030 52.215 121.755 ;
        RECT 52.400 120.860 52.645 121.585 ;
        RECT 52.815 121.030 53.075 121.755 ;
        RECT 53.260 120.860 53.515 121.585 ;
        RECT 53.685 121.030 53.975 121.770 ;
        RECT 47.240 120.855 53.515 120.860 ;
        RECT 54.145 120.855 54.415 121.600 ;
        RECT 54.675 120.855 56.345 121.945 ;
        RECT 56.515 121.615 56.855 122.425 ;
        RECT 57.025 121.860 57.775 122.050 ;
        RECT 56.515 121.205 57.030 121.615 ;
        RECT 57.265 120.855 57.435 121.615 ;
        RECT 57.605 121.195 57.775 121.860 ;
        RECT 57.945 121.875 58.135 123.235 ;
        RECT 58.305 123.065 58.580 123.235 ;
        RECT 58.305 122.895 58.585 123.065 ;
        RECT 58.305 122.075 58.580 122.895 ;
        RECT 58.770 122.870 59.300 123.235 ;
        RECT 59.725 123.005 60.055 123.405 ;
        RECT 59.125 122.835 59.300 122.870 ;
        RECT 58.785 121.875 58.955 122.675 ;
        RECT 57.945 121.705 58.955 121.875 ;
        RECT 59.125 122.665 60.055 122.835 ;
        RECT 60.225 122.665 60.480 123.235 ;
        RECT 61.115 122.680 61.405 123.405 ;
        RECT 61.665 122.855 61.835 123.235 ;
        RECT 62.015 123.025 62.345 123.405 ;
        RECT 61.665 122.685 62.330 122.855 ;
        RECT 62.525 122.730 62.785 123.235 ;
        RECT 59.125 121.535 59.295 122.665 ;
        RECT 59.885 122.495 60.055 122.665 ;
        RECT 58.170 121.365 59.295 121.535 ;
        RECT 59.465 122.165 59.660 122.495 ;
        RECT 59.885 122.165 60.140 122.495 ;
        RECT 59.465 121.195 59.635 122.165 ;
        RECT 60.310 121.995 60.480 122.665 ;
        RECT 61.595 122.135 61.925 122.505 ;
        RECT 62.160 122.430 62.330 122.685 ;
        RECT 62.160 122.100 62.445 122.430 ;
        RECT 57.605 121.025 59.635 121.195 ;
        RECT 59.805 120.855 59.975 121.995 ;
        RECT 60.145 121.025 60.480 121.995 ;
        RECT 61.115 120.855 61.405 122.020 ;
        RECT 62.160 121.955 62.330 122.100 ;
        RECT 61.665 121.785 62.330 121.955 ;
        RECT 62.615 121.930 62.785 122.730 ;
        RECT 63.415 122.635 66.005 123.405 ;
        RECT 66.180 122.860 71.525 123.405 ;
        RECT 72.070 123.065 72.325 123.225 ;
        RECT 71.985 122.895 72.325 123.065 ;
        RECT 72.505 122.945 72.790 123.405 ;
        RECT 61.665 121.025 61.835 121.785 ;
        RECT 62.015 120.855 62.345 121.615 ;
        RECT 62.515 121.025 62.785 121.930 ;
        RECT 63.415 121.945 64.625 122.465 ;
        RECT 64.795 122.115 66.005 122.635 ;
        RECT 63.415 120.855 66.005 121.945 ;
        RECT 67.770 121.290 68.120 122.540 ;
        RECT 69.600 122.030 69.940 122.860 ;
        RECT 72.070 122.695 72.325 122.895 ;
        RECT 72.070 121.835 72.250 122.695 ;
        RECT 72.970 122.495 73.220 123.145 ;
        RECT 72.420 122.165 73.220 122.495 ;
        RECT 66.180 120.855 71.525 121.290 ;
        RECT 72.070 121.165 72.325 121.835 ;
        RECT 72.505 120.855 72.790 121.655 ;
        RECT 72.970 121.575 73.220 122.165 ;
        RECT 73.420 122.810 73.740 123.140 ;
        RECT 73.920 122.925 74.580 123.405 ;
        RECT 74.780 123.015 75.630 123.185 ;
        RECT 73.420 121.915 73.610 122.810 ;
        RECT 73.930 122.485 74.590 122.755 ;
        RECT 74.260 122.425 74.590 122.485 ;
        RECT 73.780 122.255 74.110 122.315 ;
        RECT 74.780 122.255 74.950 123.015 ;
        RECT 76.190 122.945 76.510 123.405 ;
        RECT 76.710 122.765 76.960 123.195 ;
        RECT 77.250 122.965 77.660 123.405 ;
        RECT 77.830 123.025 78.845 123.225 ;
        RECT 75.120 122.595 76.370 122.765 ;
        RECT 75.120 122.475 75.450 122.595 ;
        RECT 73.780 122.085 75.680 122.255 ;
        RECT 73.420 121.745 75.340 121.915 ;
        RECT 73.420 121.725 73.740 121.745 ;
        RECT 72.970 121.065 73.300 121.575 ;
        RECT 73.570 121.115 73.740 121.725 ;
        RECT 75.510 121.575 75.680 122.085 ;
        RECT 75.850 122.015 76.030 122.425 ;
        RECT 76.200 121.835 76.370 122.595 ;
        RECT 73.910 120.855 74.240 121.545 ;
        RECT 74.470 121.405 75.680 121.575 ;
        RECT 75.850 121.525 76.370 121.835 ;
        RECT 76.540 122.425 76.960 122.765 ;
        RECT 77.250 122.425 77.660 122.755 ;
        RECT 76.540 121.655 76.730 122.425 ;
        RECT 77.830 122.295 78.000 123.025 ;
        RECT 79.145 122.855 79.315 123.185 ;
        RECT 79.485 123.025 79.815 123.405 ;
        RECT 78.170 122.475 78.520 122.845 ;
        RECT 77.830 122.255 78.250 122.295 ;
        RECT 76.900 122.085 78.250 122.255 ;
        RECT 76.900 121.925 77.150 122.085 ;
        RECT 77.660 121.655 77.910 121.915 ;
        RECT 76.540 121.405 77.910 121.655 ;
        RECT 74.470 121.115 74.710 121.405 ;
        RECT 75.510 121.325 75.680 121.405 ;
        RECT 74.910 120.855 75.330 121.235 ;
        RECT 75.510 121.075 76.140 121.325 ;
        RECT 76.610 120.855 76.940 121.235 ;
        RECT 77.110 121.115 77.280 121.405 ;
        RECT 78.080 121.240 78.250 122.085 ;
        RECT 78.700 121.915 78.920 122.785 ;
        RECT 79.145 122.665 79.840 122.855 ;
        RECT 78.420 121.535 78.920 121.915 ;
        RECT 79.090 121.865 79.500 122.485 ;
        RECT 79.670 121.695 79.840 122.665 ;
        RECT 79.145 121.525 79.840 121.695 ;
        RECT 77.460 120.855 77.840 121.235 ;
        RECT 78.080 121.070 78.910 121.240 ;
        RECT 79.145 121.025 79.315 121.525 ;
        RECT 79.485 120.855 79.815 121.355 ;
        RECT 80.030 121.025 80.255 123.145 ;
        RECT 80.425 123.025 80.755 123.405 ;
        RECT 80.925 122.855 81.095 123.145 ;
        RECT 80.430 122.685 81.095 122.855 ;
        RECT 80.430 121.695 80.660 122.685 ;
        RECT 81.630 122.595 81.875 123.200 ;
        RECT 82.095 122.870 82.605 123.405 ;
        RECT 80.830 121.865 81.180 122.515 ;
        RECT 81.355 122.425 82.585 122.595 ;
        RECT 80.430 121.525 81.095 121.695 ;
        RECT 80.425 120.855 80.755 121.355 ;
        RECT 80.925 121.025 81.095 121.525 ;
        RECT 81.355 121.615 81.695 122.425 ;
        RECT 81.865 121.860 82.615 122.050 ;
        RECT 81.355 121.205 81.870 121.615 ;
        RECT 82.105 120.855 82.275 121.615 ;
        RECT 82.445 121.195 82.615 121.860 ;
        RECT 82.785 121.875 82.975 123.235 ;
        RECT 83.145 123.065 83.420 123.235 ;
        RECT 83.145 122.895 83.425 123.065 ;
        RECT 83.145 122.075 83.420 122.895 ;
        RECT 83.610 122.870 84.140 123.235 ;
        RECT 84.565 123.005 84.895 123.405 ;
        RECT 83.965 122.835 84.140 122.870 ;
        RECT 83.625 121.875 83.795 122.675 ;
        RECT 82.785 121.705 83.795 121.875 ;
        RECT 83.965 122.665 84.895 122.835 ;
        RECT 85.065 122.665 85.320 123.235 ;
        RECT 83.965 121.535 84.135 122.665 ;
        RECT 84.725 122.495 84.895 122.665 ;
        RECT 83.010 121.365 84.135 121.535 ;
        RECT 84.305 122.165 84.500 122.495 ;
        RECT 84.725 122.165 84.980 122.495 ;
        RECT 84.305 121.195 84.475 122.165 ;
        RECT 85.150 121.995 85.320 122.665 ;
        RECT 85.535 122.585 85.765 123.405 ;
        RECT 85.935 122.605 86.265 123.235 ;
        RECT 85.515 122.165 85.845 122.415 ;
        RECT 86.015 122.005 86.265 122.605 ;
        RECT 86.435 122.585 86.645 123.405 ;
        RECT 86.875 122.680 87.165 123.405 ;
        RECT 87.710 123.065 87.965 123.225 ;
        RECT 87.625 122.895 87.965 123.065 ;
        RECT 88.145 122.945 88.430 123.405 ;
        RECT 87.710 122.695 87.965 122.895 ;
        RECT 82.445 121.025 84.475 121.195 ;
        RECT 84.645 120.855 84.815 121.995 ;
        RECT 84.985 121.025 85.320 121.995 ;
        RECT 85.535 120.855 85.765 121.995 ;
        RECT 85.935 121.025 86.265 122.005 ;
        RECT 86.435 120.855 86.645 121.995 ;
        RECT 86.875 120.855 87.165 122.020 ;
        RECT 87.710 121.835 87.890 122.695 ;
        RECT 88.610 122.495 88.860 123.145 ;
        RECT 88.060 122.165 88.860 122.495 ;
        RECT 87.710 121.165 87.965 121.835 ;
        RECT 88.145 120.855 88.430 121.655 ;
        RECT 88.610 121.575 88.860 122.165 ;
        RECT 89.060 122.810 89.380 123.140 ;
        RECT 89.560 122.925 90.220 123.405 ;
        RECT 90.420 123.015 91.270 123.185 ;
        RECT 89.060 121.915 89.250 122.810 ;
        RECT 89.570 122.485 90.230 122.755 ;
        RECT 89.900 122.425 90.230 122.485 ;
        RECT 89.420 122.255 89.750 122.315 ;
        RECT 90.420 122.255 90.590 123.015 ;
        RECT 91.830 122.945 92.150 123.405 ;
        RECT 92.350 122.765 92.600 123.195 ;
        RECT 92.890 122.965 93.300 123.405 ;
        RECT 93.470 123.025 94.485 123.225 ;
        RECT 90.760 122.595 92.010 122.765 ;
        RECT 90.760 122.475 91.090 122.595 ;
        RECT 89.420 122.085 91.320 122.255 ;
        RECT 89.060 121.745 90.980 121.915 ;
        RECT 89.060 121.725 89.380 121.745 ;
        RECT 88.610 121.065 88.940 121.575 ;
        RECT 89.210 121.115 89.380 121.725 ;
        RECT 91.150 121.575 91.320 122.085 ;
        RECT 91.490 122.015 91.670 122.425 ;
        RECT 91.840 121.835 92.010 122.595 ;
        RECT 89.550 120.855 89.880 121.545 ;
        RECT 90.110 121.405 91.320 121.575 ;
        RECT 91.490 121.525 92.010 121.835 ;
        RECT 92.180 122.425 92.600 122.765 ;
        RECT 92.890 122.425 93.300 122.755 ;
        RECT 92.180 121.655 92.370 122.425 ;
        RECT 93.470 122.295 93.640 123.025 ;
        RECT 94.785 122.855 94.955 123.185 ;
        RECT 95.125 123.025 95.455 123.405 ;
        RECT 93.810 122.475 94.160 122.845 ;
        RECT 93.470 122.255 93.890 122.295 ;
        RECT 92.540 122.085 93.890 122.255 ;
        RECT 92.540 121.925 92.790 122.085 ;
        RECT 93.300 121.655 93.550 121.915 ;
        RECT 92.180 121.405 93.550 121.655 ;
        RECT 90.110 121.115 90.350 121.405 ;
        RECT 91.150 121.325 91.320 121.405 ;
        RECT 90.550 120.855 90.970 121.235 ;
        RECT 91.150 121.075 91.780 121.325 ;
        RECT 92.250 120.855 92.580 121.235 ;
        RECT 92.750 121.115 92.920 121.405 ;
        RECT 93.720 121.240 93.890 122.085 ;
        RECT 94.340 121.915 94.560 122.785 ;
        RECT 94.785 122.665 95.480 122.855 ;
        RECT 94.060 121.535 94.560 121.915 ;
        RECT 94.730 121.865 95.140 122.485 ;
        RECT 95.310 121.695 95.480 122.665 ;
        RECT 94.785 121.525 95.480 121.695 ;
        RECT 93.100 120.855 93.480 121.235 ;
        RECT 93.720 121.070 94.550 121.240 ;
        RECT 94.785 121.025 94.955 121.525 ;
        RECT 95.125 120.855 95.455 121.355 ;
        RECT 95.670 121.025 95.895 123.145 ;
        RECT 96.065 123.025 96.395 123.405 ;
        RECT 96.565 122.855 96.735 123.145 ;
        RECT 96.070 122.685 96.735 122.855 ;
        RECT 96.070 121.695 96.300 122.685 ;
        RECT 97.955 122.585 98.185 123.405 ;
        RECT 98.355 122.605 98.685 123.235 ;
        RECT 96.470 121.865 96.820 122.515 ;
        RECT 97.935 122.165 98.265 122.415 ;
        RECT 98.435 122.005 98.685 122.605 ;
        RECT 98.855 122.585 99.065 123.405 ;
        RECT 99.670 123.065 99.925 123.225 ;
        RECT 99.585 122.895 99.925 123.065 ;
        RECT 100.105 122.945 100.390 123.405 ;
        RECT 99.670 122.695 99.925 122.895 ;
        RECT 96.070 121.525 96.735 121.695 ;
        RECT 96.065 120.855 96.395 121.355 ;
        RECT 96.565 121.025 96.735 121.525 ;
        RECT 97.955 120.855 98.185 121.995 ;
        RECT 98.355 121.025 98.685 122.005 ;
        RECT 98.855 120.855 99.065 121.995 ;
        RECT 99.670 121.835 99.850 122.695 ;
        RECT 100.570 122.495 100.820 123.145 ;
        RECT 100.020 122.165 100.820 122.495 ;
        RECT 99.670 121.165 99.925 121.835 ;
        RECT 100.105 120.855 100.390 121.655 ;
        RECT 100.570 121.575 100.820 122.165 ;
        RECT 101.020 122.810 101.340 123.140 ;
        RECT 101.520 122.925 102.180 123.405 ;
        RECT 102.380 123.015 103.230 123.185 ;
        RECT 101.020 121.915 101.210 122.810 ;
        RECT 101.530 122.485 102.190 122.755 ;
        RECT 101.860 122.425 102.190 122.485 ;
        RECT 101.380 122.255 101.710 122.315 ;
        RECT 102.380 122.255 102.550 123.015 ;
        RECT 103.790 122.945 104.110 123.405 ;
        RECT 104.310 122.765 104.560 123.195 ;
        RECT 104.850 122.965 105.260 123.405 ;
        RECT 105.430 123.025 106.445 123.225 ;
        RECT 102.720 122.595 103.970 122.765 ;
        RECT 102.720 122.475 103.050 122.595 ;
        RECT 101.380 122.085 103.280 122.255 ;
        RECT 101.020 121.745 102.940 121.915 ;
        RECT 101.020 121.725 101.340 121.745 ;
        RECT 100.570 121.065 100.900 121.575 ;
        RECT 101.170 121.115 101.340 121.725 ;
        RECT 103.110 121.575 103.280 122.085 ;
        RECT 103.450 122.015 103.630 122.425 ;
        RECT 103.800 121.835 103.970 122.595 ;
        RECT 101.510 120.855 101.840 121.545 ;
        RECT 102.070 121.405 103.280 121.575 ;
        RECT 103.450 121.525 103.970 121.835 ;
        RECT 104.140 122.425 104.560 122.765 ;
        RECT 104.850 122.425 105.260 122.755 ;
        RECT 104.140 121.655 104.330 122.425 ;
        RECT 105.430 122.295 105.600 123.025 ;
        RECT 106.745 122.855 106.915 123.185 ;
        RECT 107.085 123.025 107.415 123.405 ;
        RECT 105.770 122.475 106.120 122.845 ;
        RECT 105.430 122.255 105.850 122.295 ;
        RECT 104.500 122.085 105.850 122.255 ;
        RECT 104.500 121.925 104.750 122.085 ;
        RECT 105.260 121.655 105.510 121.915 ;
        RECT 104.140 121.405 105.510 121.655 ;
        RECT 102.070 121.115 102.310 121.405 ;
        RECT 103.110 121.325 103.280 121.405 ;
        RECT 102.510 120.855 102.930 121.235 ;
        RECT 103.110 121.075 103.740 121.325 ;
        RECT 104.210 120.855 104.540 121.235 ;
        RECT 104.710 121.115 104.880 121.405 ;
        RECT 105.680 121.240 105.850 122.085 ;
        RECT 106.300 121.915 106.520 122.785 ;
        RECT 106.745 122.665 107.440 122.855 ;
        RECT 106.020 121.535 106.520 121.915 ;
        RECT 106.690 121.865 107.100 122.485 ;
        RECT 107.270 121.695 107.440 122.665 ;
        RECT 106.745 121.525 107.440 121.695 ;
        RECT 105.060 120.855 105.440 121.235 ;
        RECT 105.680 121.070 106.510 121.240 ;
        RECT 106.745 121.025 106.915 121.525 ;
        RECT 107.085 120.855 107.415 121.355 ;
        RECT 107.630 121.025 107.855 123.145 ;
        RECT 108.025 123.025 108.355 123.405 ;
        RECT 108.525 122.855 108.695 123.145 ;
        RECT 108.030 122.685 108.695 122.855 ;
        RECT 108.030 121.695 108.260 122.685 ;
        RECT 108.955 122.635 112.465 123.405 ;
        RECT 112.635 122.680 112.925 123.405 ;
        RECT 108.430 121.865 108.780 122.515 ;
        RECT 108.955 121.945 110.645 122.465 ;
        RECT 110.815 122.115 112.465 122.635 ;
        RECT 113.370 122.595 113.615 123.200 ;
        RECT 113.835 122.870 114.345 123.405 ;
        RECT 113.095 122.425 114.325 122.595 ;
        RECT 108.030 121.525 108.695 121.695 ;
        RECT 108.025 120.855 108.355 121.355 ;
        RECT 108.525 121.025 108.695 121.525 ;
        RECT 108.955 120.855 112.465 121.945 ;
        RECT 112.635 120.855 112.925 122.020 ;
        RECT 113.095 121.615 113.435 122.425 ;
        RECT 113.605 121.860 114.355 122.050 ;
        RECT 113.095 121.205 113.610 121.615 ;
        RECT 113.845 120.855 114.015 121.615 ;
        RECT 114.185 121.195 114.355 121.860 ;
        RECT 114.525 121.875 114.715 123.235 ;
        RECT 114.885 122.385 115.160 123.235 ;
        RECT 115.350 122.870 115.880 123.235 ;
        RECT 116.305 123.005 116.635 123.405 ;
        RECT 115.705 122.835 115.880 122.870 ;
        RECT 114.885 122.215 115.165 122.385 ;
        RECT 114.885 122.075 115.160 122.215 ;
        RECT 115.365 121.875 115.535 122.675 ;
        RECT 114.525 121.705 115.535 121.875 ;
        RECT 115.705 122.665 116.635 122.835 ;
        RECT 116.805 122.665 117.060 123.235 ;
        RECT 115.705 121.535 115.875 122.665 ;
        RECT 116.465 122.495 116.635 122.665 ;
        RECT 114.750 121.365 115.875 121.535 ;
        RECT 116.045 122.165 116.240 122.495 ;
        RECT 116.465 122.165 116.720 122.495 ;
        RECT 116.045 121.195 116.215 122.165 ;
        RECT 116.890 121.995 117.060 122.665 ;
        RECT 117.295 122.585 117.505 123.405 ;
        RECT 117.675 122.605 118.005 123.235 ;
        RECT 117.675 122.005 117.925 122.605 ;
        RECT 118.175 122.585 118.405 123.405 ;
        RECT 118.655 122.585 118.885 123.405 ;
        RECT 119.055 122.605 119.385 123.235 ;
        RECT 118.095 122.165 118.425 122.415 ;
        RECT 118.635 122.165 118.965 122.415 ;
        RECT 119.135 122.005 119.385 122.605 ;
        RECT 119.555 122.585 119.765 123.405 ;
        RECT 120.915 122.635 124.425 123.405 ;
        RECT 124.595 122.655 125.805 123.405 ;
        RECT 114.185 121.025 116.215 121.195 ;
        RECT 116.385 120.855 116.555 121.995 ;
        RECT 116.725 121.025 117.060 121.995 ;
        RECT 117.295 120.855 117.505 121.995 ;
        RECT 117.675 121.025 118.005 122.005 ;
        RECT 118.175 120.855 118.405 121.995 ;
        RECT 118.655 120.855 118.885 121.995 ;
        RECT 119.055 121.025 119.385 122.005 ;
        RECT 119.555 120.855 119.765 121.995 ;
        RECT 120.915 121.945 122.605 122.465 ;
        RECT 122.775 122.115 124.425 122.635 ;
        RECT 124.595 121.945 125.115 122.485 ;
        RECT 125.285 122.115 125.805 122.655 ;
        RECT 120.915 120.855 124.425 121.945 ;
        RECT 124.595 120.855 125.805 121.945 ;
        RECT 11.810 120.685 125.890 120.855 ;
        RECT 11.895 119.595 13.105 120.685 ;
        RECT 11.895 118.885 12.415 119.425 ;
        RECT 12.585 119.055 13.105 119.595 ;
        RECT 13.735 119.595 15.405 120.685 ;
        RECT 13.735 119.075 14.485 119.595 ;
        RECT 15.615 119.545 15.845 120.685 ;
        RECT 16.015 119.535 16.345 120.515 ;
        RECT 16.515 119.545 16.725 120.685 ;
        RECT 16.995 119.545 17.225 120.685 ;
        RECT 17.395 119.535 17.725 120.515 ;
        RECT 17.895 119.545 18.105 120.685 ;
        RECT 18.335 119.925 18.850 120.335 ;
        RECT 19.085 119.925 19.255 120.685 ;
        RECT 19.425 120.345 21.455 120.515 ;
        RECT 14.655 118.905 15.405 119.425 ;
        RECT 15.595 119.125 15.925 119.375 ;
        RECT 11.895 118.135 13.105 118.885 ;
        RECT 13.735 118.135 15.405 118.905 ;
        RECT 15.615 118.135 15.845 118.955 ;
        RECT 16.095 118.935 16.345 119.535 ;
        RECT 16.975 119.125 17.305 119.375 ;
        RECT 16.015 118.305 16.345 118.935 ;
        RECT 16.515 118.135 16.725 118.955 ;
        RECT 16.995 118.135 17.225 118.955 ;
        RECT 17.475 118.935 17.725 119.535 ;
        RECT 18.335 119.115 18.675 119.925 ;
        RECT 19.425 119.680 19.595 120.345 ;
        RECT 19.990 120.005 21.115 120.175 ;
        RECT 18.845 119.490 19.595 119.680 ;
        RECT 19.765 119.665 20.775 119.835 ;
        RECT 17.395 118.305 17.725 118.935 ;
        RECT 17.895 118.135 18.105 118.955 ;
        RECT 18.335 118.945 19.565 119.115 ;
        RECT 18.610 118.340 18.855 118.945 ;
        RECT 19.075 118.135 19.585 118.670 ;
        RECT 19.765 118.305 19.955 119.665 ;
        RECT 20.125 118.645 20.400 119.465 ;
        RECT 20.605 118.865 20.775 119.665 ;
        RECT 20.945 118.875 21.115 120.005 ;
        RECT 21.285 119.375 21.455 120.345 ;
        RECT 21.625 119.545 21.795 120.685 ;
        RECT 21.965 119.545 22.300 120.515 ;
        RECT 21.285 119.045 21.480 119.375 ;
        RECT 21.705 119.045 21.960 119.375 ;
        RECT 21.705 118.875 21.875 119.045 ;
        RECT 22.130 118.875 22.300 119.545 ;
        RECT 22.475 119.520 22.765 120.685 ;
        RECT 22.935 119.610 23.205 120.515 ;
        RECT 23.375 119.925 23.705 120.685 ;
        RECT 23.885 119.755 24.055 120.515 ;
        RECT 20.945 118.705 21.875 118.875 ;
        RECT 20.945 118.670 21.120 118.705 ;
        RECT 20.125 118.475 20.405 118.645 ;
        RECT 20.125 118.305 20.400 118.475 ;
        RECT 20.590 118.305 21.120 118.670 ;
        RECT 21.545 118.135 21.875 118.535 ;
        RECT 22.045 118.305 22.300 118.875 ;
        RECT 22.475 118.135 22.765 118.860 ;
        RECT 22.935 118.810 23.105 119.610 ;
        RECT 23.390 119.585 24.055 119.755 ;
        RECT 23.390 119.440 23.560 119.585 ;
        RECT 24.815 119.545 25.045 120.685 ;
        RECT 25.215 119.535 25.545 120.515 ;
        RECT 25.715 119.545 25.925 120.685 ;
        RECT 26.195 119.545 26.425 120.685 ;
        RECT 26.595 119.535 26.925 120.515 ;
        RECT 27.095 119.545 27.305 120.685 ;
        RECT 27.535 119.925 28.050 120.335 ;
        RECT 28.285 119.925 28.455 120.685 ;
        RECT 28.625 120.345 30.655 120.515 ;
        RECT 23.275 119.110 23.560 119.440 ;
        RECT 23.390 118.855 23.560 119.110 ;
        RECT 23.795 119.035 24.125 119.405 ;
        RECT 24.795 119.125 25.125 119.375 ;
        RECT 22.935 118.305 23.195 118.810 ;
        RECT 23.390 118.685 24.055 118.855 ;
        RECT 23.375 118.135 23.705 118.515 ;
        RECT 23.885 118.305 24.055 118.685 ;
        RECT 24.815 118.135 25.045 118.955 ;
        RECT 25.295 118.935 25.545 119.535 ;
        RECT 26.175 119.125 26.505 119.375 ;
        RECT 25.215 118.305 25.545 118.935 ;
        RECT 25.715 118.135 25.925 118.955 ;
        RECT 26.195 118.135 26.425 118.955 ;
        RECT 26.675 118.935 26.925 119.535 ;
        RECT 27.535 119.115 27.875 119.925 ;
        RECT 28.625 119.680 28.795 120.345 ;
        RECT 29.190 120.005 30.315 120.175 ;
        RECT 28.045 119.490 28.795 119.680 ;
        RECT 28.965 119.665 29.975 119.835 ;
        RECT 26.595 118.305 26.925 118.935 ;
        RECT 27.095 118.135 27.305 118.955 ;
        RECT 27.535 118.945 28.765 119.115 ;
        RECT 27.810 118.340 28.055 118.945 ;
        RECT 28.275 118.135 28.785 118.670 ;
        RECT 28.965 118.305 29.155 119.665 ;
        RECT 29.325 118.645 29.600 119.465 ;
        RECT 29.805 118.865 29.975 119.665 ;
        RECT 30.145 118.875 30.315 120.005 ;
        RECT 30.485 119.375 30.655 120.345 ;
        RECT 30.825 119.545 30.995 120.685 ;
        RECT 31.165 119.545 31.500 120.515 ;
        RECT 32.050 119.705 32.305 120.375 ;
        RECT 32.485 119.885 32.770 120.685 ;
        RECT 32.950 119.965 33.280 120.475 ;
        RECT 32.050 119.665 32.230 119.705 ;
        RECT 30.485 119.045 30.680 119.375 ;
        RECT 30.905 119.045 31.160 119.375 ;
        RECT 30.905 118.875 31.075 119.045 ;
        RECT 31.330 118.875 31.500 119.545 ;
        RECT 31.965 119.495 32.230 119.665 ;
        RECT 30.145 118.705 31.075 118.875 ;
        RECT 30.145 118.670 30.320 118.705 ;
        RECT 29.325 118.475 29.605 118.645 ;
        RECT 29.325 118.305 29.600 118.475 ;
        RECT 29.790 118.305 30.320 118.670 ;
        RECT 30.745 118.135 31.075 118.535 ;
        RECT 31.245 118.305 31.500 118.875 ;
        RECT 32.050 118.845 32.230 119.495 ;
        RECT 32.950 119.375 33.200 119.965 ;
        RECT 33.550 119.815 33.720 120.425 ;
        RECT 33.890 119.995 34.220 120.685 ;
        RECT 34.450 120.135 34.690 120.425 ;
        RECT 34.890 120.305 35.310 120.685 ;
        RECT 35.490 120.215 36.120 120.465 ;
        RECT 36.590 120.305 36.920 120.685 ;
        RECT 35.490 120.135 35.660 120.215 ;
        RECT 37.090 120.135 37.260 120.425 ;
        RECT 37.440 120.305 37.820 120.685 ;
        RECT 38.060 120.300 38.890 120.470 ;
        RECT 34.450 119.965 35.660 120.135 ;
        RECT 32.400 119.045 33.200 119.375 ;
        RECT 32.050 118.315 32.305 118.845 ;
        RECT 32.485 118.135 32.770 118.595 ;
        RECT 32.950 118.395 33.200 119.045 ;
        RECT 33.400 119.795 33.720 119.815 ;
        RECT 33.400 119.625 35.320 119.795 ;
        RECT 33.400 118.730 33.590 119.625 ;
        RECT 35.490 119.455 35.660 119.965 ;
        RECT 35.830 119.705 36.350 120.015 ;
        RECT 33.760 119.285 35.660 119.455 ;
        RECT 33.760 119.225 34.090 119.285 ;
        RECT 34.240 119.055 34.570 119.115 ;
        RECT 33.910 118.785 34.570 119.055 ;
        RECT 33.400 118.400 33.720 118.730 ;
        RECT 33.900 118.135 34.560 118.615 ;
        RECT 34.760 118.525 34.930 119.285 ;
        RECT 35.830 119.115 36.010 119.525 ;
        RECT 35.100 118.945 35.430 119.065 ;
        RECT 36.180 118.945 36.350 119.705 ;
        RECT 35.100 118.775 36.350 118.945 ;
        RECT 36.520 119.885 37.890 120.135 ;
        RECT 36.520 119.115 36.710 119.885 ;
        RECT 37.640 119.625 37.890 119.885 ;
        RECT 36.880 119.455 37.130 119.615 ;
        RECT 38.060 119.455 38.230 120.300 ;
        RECT 39.125 120.015 39.295 120.515 ;
        RECT 39.465 120.185 39.795 120.685 ;
        RECT 38.400 119.625 38.900 120.005 ;
        RECT 39.125 119.845 39.820 120.015 ;
        RECT 36.880 119.285 38.230 119.455 ;
        RECT 37.810 119.245 38.230 119.285 ;
        RECT 36.520 118.775 36.940 119.115 ;
        RECT 37.230 118.785 37.640 119.115 ;
        RECT 34.760 118.355 35.610 118.525 ;
        RECT 36.170 118.135 36.490 118.595 ;
        RECT 36.690 118.345 36.940 118.775 ;
        RECT 37.230 118.135 37.640 118.575 ;
        RECT 37.810 118.515 37.980 119.245 ;
        RECT 38.150 118.695 38.500 119.065 ;
        RECT 38.680 118.755 38.900 119.625 ;
        RECT 39.070 119.055 39.480 119.675 ;
        RECT 39.650 118.875 39.820 119.845 ;
        RECT 39.125 118.685 39.820 118.875 ;
        RECT 37.810 118.315 38.825 118.515 ;
        RECT 39.125 118.355 39.295 118.685 ;
        RECT 39.465 118.135 39.795 118.515 ;
        RECT 40.010 118.395 40.235 120.515 ;
        RECT 40.405 120.185 40.735 120.685 ;
        RECT 40.905 120.015 41.075 120.515 ;
        RECT 40.410 119.845 41.075 120.015 ;
        RECT 40.410 118.855 40.640 119.845 ;
        RECT 40.810 119.025 41.160 119.675 ;
        RECT 41.335 119.595 42.545 120.685 ;
        RECT 42.720 120.250 48.065 120.685 ;
        RECT 41.335 119.055 41.855 119.595 ;
        RECT 42.025 118.885 42.545 119.425 ;
        RECT 44.310 119.000 44.660 120.250 ;
        RECT 48.235 119.520 48.525 120.685 ;
        RECT 49.675 119.545 49.885 120.685 ;
        RECT 50.055 119.535 50.385 120.515 ;
        RECT 50.555 119.545 50.785 120.685 ;
        RECT 50.995 119.925 51.510 120.335 ;
        RECT 51.745 119.925 51.915 120.685 ;
        RECT 52.085 120.345 54.115 120.515 ;
        RECT 40.410 118.685 41.075 118.855 ;
        RECT 40.405 118.135 40.735 118.515 ;
        RECT 40.905 118.395 41.075 118.685 ;
        RECT 41.335 118.135 42.545 118.885 ;
        RECT 46.140 118.680 46.480 119.510 ;
        RECT 42.720 118.135 48.065 118.680 ;
        RECT 48.235 118.135 48.525 118.860 ;
        RECT 49.675 118.135 49.885 118.955 ;
        RECT 50.055 118.935 50.305 119.535 ;
        RECT 50.475 119.125 50.805 119.375 ;
        RECT 50.995 119.115 51.335 119.925 ;
        RECT 52.085 119.680 52.255 120.345 ;
        RECT 52.650 120.005 53.775 120.175 ;
        RECT 51.505 119.490 52.255 119.680 ;
        RECT 52.425 119.665 53.435 119.835 ;
        RECT 50.055 118.305 50.385 118.935 ;
        RECT 50.555 118.135 50.785 118.955 ;
        RECT 50.995 118.945 52.225 119.115 ;
        RECT 51.270 118.340 51.515 118.945 ;
        RECT 51.735 118.135 52.245 118.670 ;
        RECT 52.425 118.305 52.615 119.665 ;
        RECT 52.785 119.325 53.060 119.465 ;
        RECT 52.785 119.155 53.065 119.325 ;
        RECT 52.785 118.305 53.060 119.155 ;
        RECT 53.265 118.865 53.435 119.665 ;
        RECT 53.605 118.875 53.775 120.005 ;
        RECT 53.945 119.375 54.115 120.345 ;
        RECT 54.285 119.545 54.455 120.685 ;
        RECT 54.625 119.545 54.960 120.515 ;
        RECT 53.945 119.045 54.140 119.375 ;
        RECT 54.365 119.045 54.620 119.375 ;
        RECT 54.365 118.875 54.535 119.045 ;
        RECT 54.790 118.875 54.960 119.545 ;
        RECT 55.135 119.595 56.345 120.685 ;
        RECT 56.890 119.705 57.145 120.375 ;
        RECT 57.325 119.885 57.610 120.685 ;
        RECT 57.790 119.965 58.120 120.475 ;
        RECT 55.135 119.055 55.655 119.595 ;
        RECT 55.825 118.885 56.345 119.425 ;
        RECT 56.890 119.325 57.070 119.705 ;
        RECT 57.790 119.375 58.040 119.965 ;
        RECT 58.390 119.815 58.560 120.425 ;
        RECT 58.730 119.995 59.060 120.685 ;
        RECT 59.290 120.135 59.530 120.425 ;
        RECT 59.730 120.305 60.150 120.685 ;
        RECT 60.330 120.215 60.960 120.465 ;
        RECT 61.430 120.305 61.760 120.685 ;
        RECT 60.330 120.135 60.500 120.215 ;
        RECT 61.930 120.135 62.100 120.425 ;
        RECT 62.280 120.305 62.660 120.685 ;
        RECT 62.900 120.300 63.730 120.470 ;
        RECT 59.290 119.965 60.500 120.135 ;
        RECT 56.805 119.155 57.070 119.325 ;
        RECT 53.605 118.705 54.535 118.875 ;
        RECT 53.605 118.670 53.780 118.705 ;
        RECT 53.250 118.305 53.780 118.670 ;
        RECT 54.205 118.135 54.535 118.535 ;
        RECT 54.705 118.305 54.960 118.875 ;
        RECT 55.135 118.135 56.345 118.885 ;
        RECT 56.890 118.845 57.070 119.155 ;
        RECT 57.240 119.045 58.040 119.375 ;
        RECT 56.890 118.315 57.145 118.845 ;
        RECT 57.325 118.135 57.610 118.595 ;
        RECT 57.790 118.395 58.040 119.045 ;
        RECT 58.240 119.795 58.560 119.815 ;
        RECT 58.240 119.625 60.160 119.795 ;
        RECT 58.240 118.730 58.430 119.625 ;
        RECT 60.330 119.455 60.500 119.965 ;
        RECT 60.670 119.705 61.190 120.015 ;
        RECT 58.600 119.285 60.500 119.455 ;
        RECT 58.600 119.225 58.930 119.285 ;
        RECT 59.080 119.055 59.410 119.115 ;
        RECT 58.750 118.785 59.410 119.055 ;
        RECT 58.240 118.400 58.560 118.730 ;
        RECT 58.740 118.135 59.400 118.615 ;
        RECT 59.600 118.525 59.770 119.285 ;
        RECT 60.670 119.115 60.850 119.525 ;
        RECT 59.940 118.945 60.270 119.065 ;
        RECT 61.020 118.945 61.190 119.705 ;
        RECT 59.940 118.775 61.190 118.945 ;
        RECT 61.360 119.885 62.730 120.135 ;
        RECT 61.360 119.115 61.550 119.885 ;
        RECT 62.480 119.625 62.730 119.885 ;
        RECT 61.720 119.455 61.970 119.615 ;
        RECT 62.900 119.455 63.070 120.300 ;
        RECT 63.965 120.015 64.135 120.515 ;
        RECT 64.305 120.185 64.635 120.685 ;
        RECT 63.240 119.625 63.740 120.005 ;
        RECT 63.965 119.845 64.660 120.015 ;
        RECT 61.720 119.285 63.070 119.455 ;
        RECT 62.650 119.245 63.070 119.285 ;
        RECT 61.360 118.775 61.780 119.115 ;
        RECT 62.070 118.785 62.480 119.115 ;
        RECT 59.600 118.355 60.450 118.525 ;
        RECT 61.010 118.135 61.330 118.595 ;
        RECT 61.530 118.345 61.780 118.775 ;
        RECT 62.070 118.135 62.480 118.575 ;
        RECT 62.650 118.515 62.820 119.245 ;
        RECT 62.990 118.695 63.340 119.065 ;
        RECT 63.520 118.755 63.740 119.625 ;
        RECT 63.910 119.055 64.320 119.675 ;
        RECT 64.490 118.875 64.660 119.845 ;
        RECT 63.965 118.685 64.660 118.875 ;
        RECT 62.650 118.315 63.665 118.515 ;
        RECT 63.965 118.355 64.135 118.685 ;
        RECT 64.305 118.135 64.635 118.515 ;
        RECT 64.850 118.395 65.075 120.515 ;
        RECT 65.245 120.185 65.575 120.685 ;
        RECT 65.745 120.015 65.915 120.515 ;
        RECT 65.250 119.845 65.915 120.015 ;
        RECT 65.250 118.855 65.480 119.845 ;
        RECT 65.650 119.025 66.000 119.675 ;
        RECT 66.635 119.595 68.305 120.685 ;
        RECT 66.635 119.075 67.385 119.595 ;
        RECT 68.515 119.545 68.745 120.685 ;
        RECT 68.915 119.535 69.245 120.515 ;
        RECT 69.415 119.545 69.625 120.685 ;
        RECT 69.855 119.925 70.370 120.335 ;
        RECT 70.605 119.925 70.775 120.685 ;
        RECT 70.945 120.345 72.975 120.515 ;
        RECT 67.555 118.905 68.305 119.425 ;
        RECT 68.495 119.125 68.825 119.375 ;
        RECT 65.250 118.685 65.915 118.855 ;
        RECT 65.245 118.135 65.575 118.515 ;
        RECT 65.745 118.395 65.915 118.685 ;
        RECT 66.635 118.135 68.305 118.905 ;
        RECT 68.515 118.135 68.745 118.955 ;
        RECT 68.995 118.935 69.245 119.535 ;
        RECT 69.855 119.115 70.195 119.925 ;
        RECT 70.945 119.680 71.115 120.345 ;
        RECT 71.510 120.005 72.635 120.175 ;
        RECT 70.365 119.490 71.115 119.680 ;
        RECT 71.285 119.665 72.295 119.835 ;
        RECT 68.915 118.305 69.245 118.935 ;
        RECT 69.415 118.135 69.625 118.955 ;
        RECT 69.855 118.945 71.085 119.115 ;
        RECT 70.130 118.340 70.375 118.945 ;
        RECT 70.595 118.135 71.105 118.670 ;
        RECT 71.285 118.305 71.475 119.665 ;
        RECT 71.645 119.325 71.920 119.465 ;
        RECT 71.645 119.155 71.925 119.325 ;
        RECT 71.645 118.305 71.920 119.155 ;
        RECT 72.125 118.865 72.295 119.665 ;
        RECT 72.465 118.875 72.635 120.005 ;
        RECT 72.805 119.375 72.975 120.345 ;
        RECT 73.145 119.545 73.315 120.685 ;
        RECT 73.485 119.545 73.820 120.515 ;
        RECT 72.805 119.045 73.000 119.375 ;
        RECT 73.225 119.045 73.480 119.375 ;
        RECT 73.225 118.875 73.395 119.045 ;
        RECT 73.650 118.875 73.820 119.545 ;
        RECT 73.995 119.520 74.285 120.685 ;
        RECT 74.915 119.925 75.430 120.335 ;
        RECT 75.665 119.925 75.835 120.685 ;
        RECT 76.005 120.345 78.035 120.515 ;
        RECT 74.915 119.115 75.255 119.925 ;
        RECT 76.005 119.680 76.175 120.345 ;
        RECT 76.570 120.005 77.695 120.175 ;
        RECT 75.425 119.490 76.175 119.680 ;
        RECT 76.345 119.665 77.355 119.835 ;
        RECT 74.915 118.945 76.145 119.115 ;
        RECT 72.465 118.705 73.395 118.875 ;
        RECT 72.465 118.670 72.640 118.705 ;
        RECT 72.110 118.305 72.640 118.670 ;
        RECT 73.065 118.135 73.395 118.535 ;
        RECT 73.565 118.305 73.820 118.875 ;
        RECT 73.995 118.135 74.285 118.860 ;
        RECT 75.190 118.340 75.435 118.945 ;
        RECT 75.655 118.135 76.165 118.670 ;
        RECT 76.345 118.305 76.535 119.665 ;
        RECT 76.705 118.985 76.980 119.465 ;
        RECT 76.705 118.815 76.985 118.985 ;
        RECT 77.185 118.865 77.355 119.665 ;
        RECT 77.525 118.875 77.695 120.005 ;
        RECT 77.865 119.375 78.035 120.345 ;
        RECT 78.205 119.545 78.375 120.685 ;
        RECT 78.545 119.545 78.880 120.515 ;
        RECT 79.115 119.545 79.325 120.685 ;
        RECT 77.865 119.045 78.060 119.375 ;
        RECT 78.285 119.045 78.540 119.375 ;
        RECT 78.285 118.875 78.455 119.045 ;
        RECT 78.710 118.875 78.880 119.545 ;
        RECT 79.495 119.535 79.825 120.515 ;
        RECT 79.995 119.545 80.225 120.685 ;
        RECT 80.495 119.545 80.705 120.685 ;
        RECT 80.875 119.535 81.205 120.515 ;
        RECT 81.375 119.545 81.605 120.685 ;
        RECT 82.650 120.345 82.905 120.375 ;
        RECT 82.565 120.175 82.905 120.345 ;
        RECT 82.650 119.705 82.905 120.175 ;
        RECT 83.085 119.885 83.370 120.685 ;
        RECT 83.550 119.965 83.880 120.475 ;
        RECT 76.705 118.305 76.980 118.815 ;
        RECT 77.525 118.705 78.455 118.875 ;
        RECT 77.525 118.670 77.700 118.705 ;
        RECT 77.170 118.305 77.700 118.670 ;
        RECT 78.125 118.135 78.455 118.535 ;
        RECT 78.625 118.305 78.880 118.875 ;
        RECT 79.115 118.135 79.325 118.955 ;
        RECT 79.495 118.935 79.745 119.535 ;
        RECT 79.915 119.125 80.245 119.375 ;
        RECT 79.495 118.305 79.825 118.935 ;
        RECT 79.995 118.135 80.225 118.955 ;
        RECT 80.495 118.135 80.705 118.955 ;
        RECT 80.875 118.935 81.125 119.535 ;
        RECT 81.295 119.125 81.625 119.375 ;
        RECT 80.875 118.305 81.205 118.935 ;
        RECT 81.375 118.135 81.605 118.955 ;
        RECT 82.650 118.845 82.830 119.705 ;
        RECT 83.550 119.375 83.800 119.965 ;
        RECT 84.150 119.815 84.320 120.425 ;
        RECT 84.490 119.995 84.820 120.685 ;
        RECT 85.050 120.135 85.290 120.425 ;
        RECT 85.490 120.305 85.910 120.685 ;
        RECT 86.090 120.215 86.720 120.465 ;
        RECT 87.190 120.305 87.520 120.685 ;
        RECT 86.090 120.135 86.260 120.215 ;
        RECT 87.690 120.135 87.860 120.425 ;
        RECT 88.040 120.305 88.420 120.685 ;
        RECT 88.660 120.300 89.490 120.470 ;
        RECT 85.050 119.965 86.260 120.135 ;
        RECT 83.000 119.045 83.800 119.375 ;
        RECT 82.650 118.315 82.905 118.845 ;
        RECT 83.085 118.135 83.370 118.595 ;
        RECT 83.550 118.395 83.800 119.045 ;
        RECT 84.000 119.795 84.320 119.815 ;
        RECT 84.000 119.625 85.920 119.795 ;
        RECT 84.000 118.730 84.190 119.625 ;
        RECT 86.090 119.455 86.260 119.965 ;
        RECT 86.430 119.705 86.950 120.015 ;
        RECT 84.360 119.285 86.260 119.455 ;
        RECT 84.360 119.225 84.690 119.285 ;
        RECT 84.840 119.055 85.170 119.115 ;
        RECT 84.510 118.785 85.170 119.055 ;
        RECT 84.000 118.400 84.320 118.730 ;
        RECT 84.500 118.135 85.160 118.615 ;
        RECT 85.360 118.525 85.530 119.285 ;
        RECT 86.430 119.115 86.610 119.525 ;
        RECT 85.700 118.945 86.030 119.065 ;
        RECT 86.780 118.945 86.950 119.705 ;
        RECT 85.700 118.775 86.950 118.945 ;
        RECT 87.120 119.885 88.490 120.135 ;
        RECT 87.120 119.115 87.310 119.885 ;
        RECT 88.240 119.625 88.490 119.885 ;
        RECT 87.480 119.455 87.730 119.615 ;
        RECT 88.660 119.455 88.830 120.300 ;
        RECT 89.725 120.015 89.895 120.515 ;
        RECT 90.065 120.185 90.395 120.685 ;
        RECT 89.000 119.625 89.500 120.005 ;
        RECT 89.725 119.845 90.420 120.015 ;
        RECT 87.480 119.285 88.830 119.455 ;
        RECT 88.410 119.245 88.830 119.285 ;
        RECT 87.120 118.775 87.540 119.115 ;
        RECT 87.830 118.785 88.240 119.115 ;
        RECT 85.360 118.355 86.210 118.525 ;
        RECT 86.770 118.135 87.090 118.595 ;
        RECT 87.290 118.345 87.540 118.775 ;
        RECT 87.830 118.135 88.240 118.575 ;
        RECT 88.410 118.515 88.580 119.245 ;
        RECT 88.750 118.695 89.100 119.065 ;
        RECT 89.280 118.755 89.500 119.625 ;
        RECT 89.670 119.055 90.080 119.675 ;
        RECT 90.250 118.875 90.420 119.845 ;
        RECT 89.725 118.685 90.420 118.875 ;
        RECT 88.410 118.315 89.425 118.515 ;
        RECT 89.725 118.355 89.895 118.685 ;
        RECT 90.065 118.135 90.395 118.515 ;
        RECT 90.610 118.395 90.835 120.515 ;
        RECT 91.005 120.185 91.335 120.685 ;
        RECT 91.505 120.015 91.675 120.515 ;
        RECT 91.010 119.845 91.675 120.015 ;
        RECT 91.935 119.925 92.450 120.335 ;
        RECT 92.685 119.925 92.855 120.685 ;
        RECT 93.025 120.345 95.055 120.515 ;
        RECT 91.010 118.855 91.240 119.845 ;
        RECT 91.410 119.025 91.760 119.675 ;
        RECT 91.935 119.115 92.275 119.925 ;
        RECT 93.025 119.680 93.195 120.345 ;
        RECT 93.590 120.005 94.715 120.175 ;
        RECT 92.445 119.490 93.195 119.680 ;
        RECT 93.365 119.665 94.375 119.835 ;
        RECT 91.935 118.945 93.165 119.115 ;
        RECT 91.010 118.685 91.675 118.855 ;
        RECT 91.005 118.135 91.335 118.515 ;
        RECT 91.505 118.395 91.675 118.685 ;
        RECT 92.210 118.340 92.455 118.945 ;
        RECT 92.675 118.135 93.185 118.670 ;
        RECT 93.365 118.305 93.555 119.665 ;
        RECT 93.725 119.325 94.000 119.465 ;
        RECT 93.725 119.155 94.005 119.325 ;
        RECT 93.725 118.305 94.000 119.155 ;
        RECT 94.205 118.865 94.375 119.665 ;
        RECT 94.545 118.875 94.715 120.005 ;
        RECT 94.885 119.375 95.055 120.345 ;
        RECT 95.225 119.545 95.395 120.685 ;
        RECT 95.565 119.545 95.900 120.515 ;
        RECT 94.885 119.045 95.080 119.375 ;
        RECT 95.305 119.045 95.560 119.375 ;
        RECT 95.305 118.875 95.475 119.045 ;
        RECT 95.730 118.875 95.900 119.545 ;
        RECT 94.545 118.705 95.475 118.875 ;
        RECT 94.545 118.670 94.720 118.705 ;
        RECT 94.190 118.305 94.720 118.670 ;
        RECT 95.145 118.135 95.475 118.535 ;
        RECT 95.645 118.305 95.900 118.875 ;
        RECT 96.075 119.610 96.345 120.515 ;
        RECT 96.515 119.925 96.845 120.685 ;
        RECT 97.025 119.755 97.195 120.515 ;
        RECT 96.075 118.810 96.245 119.610 ;
        RECT 96.530 119.585 97.195 119.755 ;
        RECT 98.375 119.610 98.645 120.515 ;
        RECT 98.815 119.925 99.145 120.685 ;
        RECT 99.325 119.755 99.495 120.515 ;
        RECT 96.530 119.440 96.700 119.585 ;
        RECT 96.415 119.110 96.700 119.440 ;
        RECT 96.530 118.855 96.700 119.110 ;
        RECT 96.935 119.035 97.265 119.405 ;
        RECT 96.075 118.305 96.335 118.810 ;
        RECT 96.530 118.685 97.195 118.855 ;
        RECT 96.515 118.135 96.845 118.515 ;
        RECT 97.025 118.305 97.195 118.685 ;
        RECT 98.375 118.810 98.545 119.610 ;
        RECT 98.830 119.585 99.495 119.755 ;
        RECT 98.830 119.440 99.000 119.585 ;
        RECT 99.755 119.520 100.045 120.685 ;
        RECT 100.220 119.545 100.555 120.515 ;
        RECT 100.725 119.545 100.895 120.685 ;
        RECT 101.065 120.345 103.095 120.515 ;
        RECT 98.715 119.110 99.000 119.440 ;
        RECT 98.830 118.855 99.000 119.110 ;
        RECT 99.235 119.035 99.565 119.405 ;
        RECT 100.220 118.875 100.390 119.545 ;
        RECT 101.065 119.375 101.235 120.345 ;
        RECT 100.560 119.045 100.815 119.375 ;
        RECT 101.040 119.045 101.235 119.375 ;
        RECT 101.405 120.005 102.530 120.175 ;
        RECT 100.645 118.875 100.815 119.045 ;
        RECT 101.405 118.875 101.575 120.005 ;
        RECT 98.375 118.305 98.635 118.810 ;
        RECT 98.830 118.685 99.495 118.855 ;
        RECT 98.815 118.135 99.145 118.515 ;
        RECT 99.325 118.305 99.495 118.685 ;
        RECT 99.755 118.135 100.045 118.860 ;
        RECT 100.220 118.305 100.475 118.875 ;
        RECT 100.645 118.705 101.575 118.875 ;
        RECT 101.745 119.665 102.755 119.835 ;
        RECT 101.745 118.865 101.915 119.665 ;
        RECT 102.120 118.985 102.395 119.465 ;
        RECT 102.115 118.815 102.395 118.985 ;
        RECT 101.400 118.670 101.575 118.705 ;
        RECT 100.645 118.135 100.975 118.535 ;
        RECT 101.400 118.305 101.930 118.670 ;
        RECT 102.120 118.305 102.395 118.815 ;
        RECT 102.565 118.305 102.755 119.665 ;
        RECT 102.925 119.680 103.095 120.345 ;
        RECT 103.265 119.925 103.435 120.685 ;
        RECT 103.670 119.925 104.185 120.335 ;
        RECT 102.925 119.490 103.675 119.680 ;
        RECT 103.845 119.115 104.185 119.925 ;
        RECT 104.395 119.545 104.625 120.685 ;
        RECT 104.795 119.535 105.125 120.515 ;
        RECT 105.295 119.545 105.505 120.685 ;
        RECT 105.735 119.925 106.250 120.335 ;
        RECT 106.485 119.925 106.655 120.685 ;
        RECT 106.825 120.345 108.855 120.515 ;
        RECT 104.375 119.125 104.705 119.375 ;
        RECT 102.955 118.945 104.185 119.115 ;
        RECT 102.935 118.135 103.445 118.670 ;
        RECT 103.665 118.340 103.910 118.945 ;
        RECT 104.395 118.135 104.625 118.955 ;
        RECT 104.875 118.935 105.125 119.535 ;
        RECT 105.735 119.115 106.075 119.925 ;
        RECT 106.825 119.680 106.995 120.345 ;
        RECT 107.390 120.005 108.515 120.175 ;
        RECT 106.245 119.490 106.995 119.680 ;
        RECT 107.165 119.665 108.175 119.835 ;
        RECT 104.795 118.305 105.125 118.935 ;
        RECT 105.295 118.135 105.505 118.955 ;
        RECT 105.735 118.945 106.965 119.115 ;
        RECT 106.010 118.340 106.255 118.945 ;
        RECT 106.475 118.135 106.985 118.670 ;
        RECT 107.165 118.305 107.355 119.665 ;
        RECT 107.525 119.325 107.800 119.465 ;
        RECT 107.525 119.155 107.805 119.325 ;
        RECT 107.525 118.305 107.800 119.155 ;
        RECT 108.005 118.865 108.175 119.665 ;
        RECT 108.345 118.875 108.515 120.005 ;
        RECT 108.685 119.375 108.855 120.345 ;
        RECT 109.025 119.545 109.195 120.685 ;
        RECT 109.365 119.545 109.700 120.515 ;
        RECT 108.685 119.045 108.880 119.375 ;
        RECT 109.105 119.045 109.360 119.375 ;
        RECT 109.105 118.875 109.275 119.045 ;
        RECT 109.530 118.875 109.700 119.545 ;
        RECT 110.335 119.595 112.925 120.685 ;
        RECT 113.470 119.705 113.725 120.375 ;
        RECT 113.905 119.885 114.190 120.685 ;
        RECT 114.370 119.965 114.700 120.475 ;
        RECT 113.470 119.665 113.650 119.705 ;
        RECT 110.335 119.075 111.545 119.595 ;
        RECT 113.385 119.495 113.650 119.665 ;
        RECT 111.715 118.905 112.925 119.425 ;
        RECT 108.345 118.705 109.275 118.875 ;
        RECT 108.345 118.670 108.520 118.705 ;
        RECT 107.990 118.305 108.520 118.670 ;
        RECT 108.945 118.135 109.275 118.535 ;
        RECT 109.445 118.305 109.700 118.875 ;
        RECT 110.335 118.135 112.925 118.905 ;
        RECT 113.470 118.845 113.650 119.495 ;
        RECT 114.370 119.375 114.620 119.965 ;
        RECT 114.970 119.815 115.140 120.425 ;
        RECT 115.310 119.995 115.640 120.685 ;
        RECT 115.870 120.135 116.110 120.425 ;
        RECT 116.310 120.305 116.730 120.685 ;
        RECT 116.910 120.215 117.540 120.465 ;
        RECT 118.010 120.305 118.340 120.685 ;
        RECT 116.910 120.135 117.080 120.215 ;
        RECT 118.510 120.135 118.680 120.425 ;
        RECT 118.860 120.305 119.240 120.685 ;
        RECT 119.480 120.300 120.310 120.470 ;
        RECT 115.870 119.965 117.080 120.135 ;
        RECT 113.820 119.045 114.620 119.375 ;
        RECT 113.470 118.315 113.725 118.845 ;
        RECT 113.905 118.135 114.190 118.595 ;
        RECT 114.370 118.395 114.620 119.045 ;
        RECT 114.820 119.795 115.140 119.815 ;
        RECT 114.820 119.625 116.740 119.795 ;
        RECT 114.820 118.730 115.010 119.625 ;
        RECT 116.910 119.455 117.080 119.965 ;
        RECT 117.250 119.705 117.770 120.015 ;
        RECT 115.180 119.285 117.080 119.455 ;
        RECT 115.180 119.225 115.510 119.285 ;
        RECT 115.660 119.055 115.990 119.115 ;
        RECT 115.330 118.785 115.990 119.055 ;
        RECT 114.820 118.400 115.140 118.730 ;
        RECT 115.320 118.135 115.980 118.615 ;
        RECT 116.180 118.525 116.350 119.285 ;
        RECT 117.250 119.115 117.430 119.525 ;
        RECT 116.520 118.945 116.850 119.065 ;
        RECT 117.600 118.945 117.770 119.705 ;
        RECT 116.520 118.775 117.770 118.945 ;
        RECT 117.940 119.885 119.310 120.135 ;
        RECT 117.940 119.115 118.130 119.885 ;
        RECT 119.060 119.625 119.310 119.885 ;
        RECT 118.300 119.455 118.550 119.615 ;
        RECT 119.480 119.455 119.650 120.300 ;
        RECT 120.545 120.015 120.715 120.515 ;
        RECT 120.885 120.185 121.215 120.685 ;
        RECT 119.820 119.625 120.320 120.005 ;
        RECT 120.545 119.845 121.240 120.015 ;
        RECT 118.300 119.285 119.650 119.455 ;
        RECT 119.230 119.245 119.650 119.285 ;
        RECT 117.940 118.775 118.360 119.115 ;
        RECT 118.650 118.785 119.060 119.115 ;
        RECT 116.180 118.355 117.030 118.525 ;
        RECT 117.590 118.135 117.910 118.595 ;
        RECT 118.110 118.345 118.360 118.775 ;
        RECT 118.650 118.135 119.060 118.575 ;
        RECT 119.230 118.515 119.400 119.245 ;
        RECT 119.570 118.695 119.920 119.065 ;
        RECT 120.100 118.755 120.320 119.625 ;
        RECT 120.490 119.055 120.900 119.675 ;
        RECT 121.070 118.875 121.240 119.845 ;
        RECT 120.545 118.685 121.240 118.875 ;
        RECT 119.230 118.315 120.245 118.515 ;
        RECT 120.545 118.355 120.715 118.685 ;
        RECT 120.885 118.135 121.215 118.515 ;
        RECT 121.430 118.395 121.655 120.515 ;
        RECT 121.825 120.185 122.155 120.685 ;
        RECT 122.325 120.015 122.495 120.515 ;
        RECT 121.830 119.845 122.495 120.015 ;
        RECT 121.830 118.855 122.060 119.845 ;
        RECT 122.230 119.025 122.580 119.675 ;
        RECT 122.755 119.595 124.425 120.685 ;
        RECT 124.595 119.595 125.805 120.685 ;
        RECT 122.755 119.075 123.505 119.595 ;
        RECT 123.675 118.905 124.425 119.425 ;
        RECT 124.595 119.055 125.115 119.595 ;
        RECT 121.830 118.685 122.495 118.855 ;
        RECT 121.825 118.135 122.155 118.515 ;
        RECT 122.325 118.395 122.495 118.685 ;
        RECT 122.755 118.135 124.425 118.905 ;
        RECT 125.285 118.885 125.805 119.425 ;
        RECT 124.595 118.135 125.805 118.885 ;
        RECT 11.810 117.965 125.890 118.135 ;
        RECT 11.895 117.215 13.105 117.965 ;
        RECT 11.895 116.675 12.415 117.215 ;
        RECT 13.275 117.195 15.865 117.965 ;
        RECT 16.410 117.625 16.665 117.785 ;
        RECT 16.325 117.455 16.665 117.625 ;
        RECT 16.845 117.505 17.130 117.965 ;
        RECT 12.585 116.505 13.105 117.045 ;
        RECT 11.895 115.415 13.105 116.505 ;
        RECT 13.275 116.505 14.485 117.025 ;
        RECT 14.655 116.675 15.865 117.195 ;
        RECT 16.410 117.255 16.665 117.455 ;
        RECT 13.275 115.415 15.865 116.505 ;
        RECT 16.410 116.395 16.590 117.255 ;
        RECT 17.310 117.055 17.560 117.705 ;
        RECT 16.760 116.725 17.560 117.055 ;
        RECT 16.410 115.725 16.665 116.395 ;
        RECT 16.845 115.415 17.130 116.215 ;
        RECT 17.310 116.135 17.560 116.725 ;
        RECT 17.760 117.370 18.080 117.700 ;
        RECT 18.260 117.485 18.920 117.965 ;
        RECT 19.120 117.575 19.970 117.745 ;
        RECT 17.760 116.475 17.950 117.370 ;
        RECT 18.270 117.045 18.930 117.315 ;
        RECT 18.600 116.985 18.930 117.045 ;
        RECT 18.120 116.815 18.450 116.875 ;
        RECT 19.120 116.815 19.290 117.575 ;
        RECT 20.530 117.505 20.850 117.965 ;
        RECT 21.050 117.325 21.300 117.755 ;
        RECT 21.590 117.525 22.000 117.965 ;
        RECT 22.170 117.585 23.185 117.785 ;
        RECT 19.460 117.155 20.710 117.325 ;
        RECT 19.460 117.035 19.790 117.155 ;
        RECT 18.120 116.645 20.020 116.815 ;
        RECT 17.760 116.305 19.680 116.475 ;
        RECT 17.760 116.285 18.080 116.305 ;
        RECT 17.310 115.625 17.640 116.135 ;
        RECT 17.910 115.675 18.080 116.285 ;
        RECT 19.850 116.135 20.020 116.645 ;
        RECT 20.190 116.575 20.370 116.985 ;
        RECT 20.540 116.395 20.710 117.155 ;
        RECT 18.250 115.415 18.580 116.105 ;
        RECT 18.810 115.965 20.020 116.135 ;
        RECT 20.190 116.085 20.710 116.395 ;
        RECT 20.880 116.985 21.300 117.325 ;
        RECT 21.590 116.985 22.000 117.315 ;
        RECT 20.880 116.215 21.070 116.985 ;
        RECT 22.170 116.855 22.340 117.585 ;
        RECT 23.485 117.415 23.655 117.745 ;
        RECT 23.825 117.585 24.155 117.965 ;
        RECT 22.510 117.035 22.860 117.405 ;
        RECT 22.170 116.815 22.590 116.855 ;
        RECT 21.240 116.645 22.590 116.815 ;
        RECT 21.240 116.485 21.490 116.645 ;
        RECT 22.000 116.215 22.250 116.475 ;
        RECT 20.880 115.965 22.250 116.215 ;
        RECT 18.810 115.675 19.050 115.965 ;
        RECT 19.850 115.885 20.020 115.965 ;
        RECT 19.250 115.415 19.670 115.795 ;
        RECT 19.850 115.635 20.480 115.885 ;
        RECT 20.950 115.415 21.280 115.795 ;
        RECT 21.450 115.675 21.620 115.965 ;
        RECT 22.420 115.800 22.590 116.645 ;
        RECT 23.040 116.475 23.260 117.345 ;
        RECT 23.485 117.225 24.180 117.415 ;
        RECT 22.760 116.095 23.260 116.475 ;
        RECT 23.430 116.425 23.840 117.045 ;
        RECT 24.010 116.255 24.180 117.225 ;
        RECT 23.485 116.085 24.180 116.255 ;
        RECT 21.800 115.415 22.180 115.795 ;
        RECT 22.420 115.630 23.250 115.800 ;
        RECT 23.485 115.585 23.655 116.085 ;
        RECT 23.825 115.415 24.155 115.915 ;
        RECT 24.370 115.585 24.595 117.705 ;
        RECT 24.765 117.585 25.095 117.965 ;
        RECT 25.265 117.415 25.435 117.705 ;
        RECT 24.770 117.245 25.435 117.415 ;
        RECT 24.770 116.255 25.000 117.245 ;
        RECT 26.155 117.195 29.665 117.965 ;
        RECT 29.925 117.415 30.095 117.795 ;
        RECT 30.275 117.585 30.605 117.965 ;
        RECT 29.925 117.245 30.590 117.415 ;
        RECT 30.785 117.290 31.045 117.795 ;
        RECT 25.170 116.425 25.520 117.075 ;
        RECT 26.155 116.505 27.845 117.025 ;
        RECT 28.015 116.675 29.665 117.195 ;
        RECT 29.855 116.695 30.185 117.065 ;
        RECT 30.420 116.990 30.590 117.245 ;
        RECT 30.420 116.660 30.705 116.990 ;
        RECT 30.420 116.515 30.590 116.660 ;
        RECT 24.770 116.085 25.435 116.255 ;
        RECT 24.765 115.415 25.095 115.915 ;
        RECT 25.265 115.585 25.435 116.085 ;
        RECT 26.155 115.415 29.665 116.505 ;
        RECT 29.925 116.345 30.590 116.515 ;
        RECT 30.875 116.490 31.045 117.290 ;
        RECT 31.490 117.155 31.735 117.760 ;
        RECT 31.955 117.430 32.465 117.965 ;
        RECT 29.925 115.585 30.095 116.345 ;
        RECT 30.275 115.415 30.605 116.175 ;
        RECT 30.775 115.585 31.045 116.490 ;
        RECT 31.215 116.985 32.445 117.155 ;
        RECT 31.215 116.175 31.555 116.985 ;
        RECT 31.725 116.420 32.475 116.610 ;
        RECT 31.215 115.765 31.730 116.175 ;
        RECT 31.965 115.415 32.135 116.175 ;
        RECT 32.305 115.755 32.475 116.420 ;
        RECT 32.645 116.435 32.835 117.795 ;
        RECT 33.005 117.285 33.280 117.795 ;
        RECT 33.470 117.430 34.000 117.795 ;
        RECT 34.425 117.565 34.755 117.965 ;
        RECT 33.825 117.395 34.000 117.430 ;
        RECT 33.005 117.115 33.285 117.285 ;
        RECT 33.005 116.635 33.280 117.115 ;
        RECT 33.485 116.435 33.655 117.235 ;
        RECT 32.645 116.265 33.655 116.435 ;
        RECT 33.825 117.225 34.755 117.395 ;
        RECT 34.925 117.225 35.180 117.795 ;
        RECT 35.355 117.240 35.645 117.965 ;
        RECT 33.825 116.095 33.995 117.225 ;
        RECT 34.585 117.055 34.755 117.225 ;
        RECT 32.870 115.925 33.995 116.095 ;
        RECT 34.165 116.725 34.360 117.055 ;
        RECT 34.585 116.725 34.840 117.055 ;
        RECT 34.165 115.755 34.335 116.725 ;
        RECT 35.010 116.555 35.180 117.225 ;
        RECT 35.815 117.215 37.025 117.965 ;
        RECT 32.305 115.585 34.335 115.755 ;
        RECT 34.505 115.415 34.675 116.555 ;
        RECT 34.845 115.585 35.180 116.555 ;
        RECT 35.355 115.415 35.645 116.580 ;
        RECT 35.815 116.505 36.335 117.045 ;
        RECT 36.505 116.675 37.025 117.215 ;
        RECT 37.195 117.195 40.705 117.965 ;
        RECT 40.880 117.420 46.225 117.965 ;
        RECT 37.195 116.505 38.885 117.025 ;
        RECT 39.055 116.675 40.705 117.195 ;
        RECT 35.815 115.415 37.025 116.505 ;
        RECT 37.195 115.415 40.705 116.505 ;
        RECT 42.470 115.850 42.820 117.100 ;
        RECT 44.300 116.590 44.640 117.420 ;
        RECT 46.395 117.290 46.655 117.795 ;
        RECT 46.835 117.585 47.165 117.965 ;
        RECT 47.345 117.415 47.515 117.795 ;
        RECT 48.150 117.625 48.405 117.785 ;
        RECT 48.065 117.455 48.405 117.625 ;
        RECT 48.585 117.505 48.870 117.965 ;
        RECT 46.395 116.490 46.565 117.290 ;
        RECT 46.850 117.245 47.515 117.415 ;
        RECT 48.150 117.255 48.405 117.455 ;
        RECT 46.850 116.990 47.020 117.245 ;
        RECT 46.735 116.660 47.020 116.990 ;
        RECT 47.255 116.695 47.585 117.065 ;
        RECT 46.850 116.515 47.020 116.660 ;
        RECT 40.880 115.415 46.225 115.850 ;
        RECT 46.395 115.585 46.665 116.490 ;
        RECT 46.850 116.345 47.515 116.515 ;
        RECT 46.835 115.415 47.165 116.175 ;
        RECT 47.345 115.585 47.515 116.345 ;
        RECT 48.150 116.395 48.330 117.255 ;
        RECT 49.050 117.055 49.300 117.705 ;
        RECT 48.500 116.725 49.300 117.055 ;
        RECT 48.150 115.725 48.405 116.395 ;
        RECT 48.585 115.415 48.870 116.215 ;
        RECT 49.050 116.135 49.300 116.725 ;
        RECT 49.500 117.370 49.820 117.700 ;
        RECT 50.000 117.485 50.660 117.965 ;
        RECT 50.860 117.575 51.710 117.745 ;
        RECT 49.500 116.475 49.690 117.370 ;
        RECT 50.010 117.045 50.670 117.315 ;
        RECT 50.340 116.985 50.670 117.045 ;
        RECT 49.860 116.815 50.190 116.875 ;
        RECT 50.860 116.815 51.030 117.575 ;
        RECT 52.270 117.505 52.590 117.965 ;
        RECT 52.790 117.325 53.040 117.755 ;
        RECT 53.330 117.525 53.740 117.965 ;
        RECT 53.910 117.585 54.925 117.785 ;
        RECT 51.200 117.155 52.450 117.325 ;
        RECT 51.200 117.035 51.530 117.155 ;
        RECT 49.860 116.645 51.760 116.815 ;
        RECT 49.500 116.305 51.420 116.475 ;
        RECT 49.500 116.285 49.820 116.305 ;
        RECT 49.050 115.625 49.380 116.135 ;
        RECT 49.650 115.675 49.820 116.285 ;
        RECT 51.590 116.135 51.760 116.645 ;
        RECT 51.930 116.575 52.110 116.985 ;
        RECT 52.280 116.395 52.450 117.155 ;
        RECT 49.990 115.415 50.320 116.105 ;
        RECT 50.550 115.965 51.760 116.135 ;
        RECT 51.930 116.085 52.450 116.395 ;
        RECT 52.620 116.985 53.040 117.325 ;
        RECT 53.330 116.985 53.740 117.315 ;
        RECT 52.620 116.215 52.810 116.985 ;
        RECT 53.910 116.855 54.080 117.585 ;
        RECT 55.225 117.415 55.395 117.745 ;
        RECT 55.565 117.585 55.895 117.965 ;
        RECT 54.250 117.035 54.600 117.405 ;
        RECT 53.910 116.815 54.330 116.855 ;
        RECT 52.980 116.645 54.330 116.815 ;
        RECT 52.980 116.485 53.230 116.645 ;
        RECT 53.740 116.215 53.990 116.475 ;
        RECT 52.620 115.965 53.990 116.215 ;
        RECT 50.550 115.675 50.790 115.965 ;
        RECT 51.590 115.885 51.760 115.965 ;
        RECT 50.990 115.415 51.410 115.795 ;
        RECT 51.590 115.635 52.220 115.885 ;
        RECT 52.690 115.415 53.020 115.795 ;
        RECT 53.190 115.675 53.360 115.965 ;
        RECT 54.160 115.800 54.330 116.645 ;
        RECT 54.780 116.475 55.000 117.345 ;
        RECT 55.225 117.225 55.920 117.415 ;
        RECT 54.500 116.095 55.000 116.475 ;
        RECT 55.170 116.425 55.580 117.045 ;
        RECT 55.750 116.255 55.920 117.225 ;
        RECT 55.225 116.085 55.920 116.255 ;
        RECT 53.540 115.415 53.920 115.795 ;
        RECT 54.160 115.630 54.990 115.800 ;
        RECT 55.225 115.585 55.395 116.085 ;
        RECT 55.565 115.415 55.895 115.915 ;
        RECT 56.110 115.585 56.335 117.705 ;
        RECT 56.505 117.585 56.835 117.965 ;
        RECT 57.005 117.415 57.175 117.705 ;
        RECT 56.510 117.245 57.175 117.415 ;
        RECT 56.510 116.255 56.740 117.245 ;
        RECT 57.895 117.195 59.565 117.965 ;
        RECT 56.910 116.425 57.260 117.075 ;
        RECT 57.895 116.505 58.645 117.025 ;
        RECT 58.815 116.675 59.565 117.195 ;
        RECT 59.775 117.145 60.005 117.965 ;
        RECT 60.175 117.165 60.505 117.795 ;
        RECT 59.755 116.725 60.085 116.975 ;
        RECT 60.255 116.565 60.505 117.165 ;
        RECT 60.675 117.145 60.885 117.965 ;
        RECT 61.115 117.240 61.405 117.965 ;
        RECT 61.850 117.155 62.095 117.760 ;
        RECT 62.315 117.430 62.825 117.965 ;
        RECT 61.575 116.985 62.805 117.155 ;
        RECT 56.510 116.085 57.175 116.255 ;
        RECT 56.505 115.415 56.835 115.915 ;
        RECT 57.005 115.585 57.175 116.085 ;
        RECT 57.895 115.415 59.565 116.505 ;
        RECT 59.775 115.415 60.005 116.555 ;
        RECT 60.175 115.585 60.505 116.565 ;
        RECT 60.675 115.415 60.885 116.555 ;
        RECT 61.115 115.415 61.405 116.580 ;
        RECT 61.575 116.175 61.915 116.985 ;
        RECT 62.085 116.420 62.835 116.610 ;
        RECT 61.575 115.765 62.090 116.175 ;
        RECT 62.325 115.415 62.495 116.175 ;
        RECT 62.665 115.755 62.835 116.420 ;
        RECT 63.005 116.435 63.195 117.795 ;
        RECT 63.365 117.285 63.640 117.795 ;
        RECT 63.830 117.430 64.360 117.795 ;
        RECT 64.785 117.565 65.115 117.965 ;
        RECT 64.185 117.395 64.360 117.430 ;
        RECT 63.365 117.115 63.645 117.285 ;
        RECT 63.365 116.635 63.640 117.115 ;
        RECT 63.845 116.435 64.015 117.235 ;
        RECT 63.005 116.265 64.015 116.435 ;
        RECT 64.185 117.225 65.115 117.395 ;
        RECT 65.285 117.225 65.540 117.795 ;
        RECT 65.805 117.415 65.975 117.795 ;
        RECT 66.155 117.585 66.485 117.965 ;
        RECT 65.805 117.245 66.470 117.415 ;
        RECT 66.665 117.290 66.925 117.795 ;
        RECT 64.185 116.095 64.355 117.225 ;
        RECT 64.945 117.055 65.115 117.225 ;
        RECT 63.230 115.925 64.355 116.095 ;
        RECT 64.525 116.725 64.720 117.055 ;
        RECT 64.945 116.725 65.200 117.055 ;
        RECT 64.525 115.755 64.695 116.725 ;
        RECT 65.370 116.555 65.540 117.225 ;
        RECT 65.735 116.695 66.065 117.065 ;
        RECT 66.300 116.990 66.470 117.245 ;
        RECT 62.665 115.585 64.695 115.755 ;
        RECT 64.865 115.415 65.035 116.555 ;
        RECT 65.205 115.585 65.540 116.555 ;
        RECT 66.300 116.660 66.585 116.990 ;
        RECT 66.300 116.515 66.470 116.660 ;
        RECT 65.805 116.345 66.470 116.515 ;
        RECT 66.755 116.490 66.925 117.290 ;
        RECT 68.015 117.195 71.525 117.965 ;
        RECT 65.805 115.585 65.975 116.345 ;
        RECT 66.155 115.415 66.485 116.175 ;
        RECT 66.655 115.585 66.925 116.490 ;
        RECT 68.015 116.505 69.705 117.025 ;
        RECT 69.875 116.675 71.525 117.195 ;
        RECT 72.070 117.255 72.325 117.785 ;
        RECT 72.505 117.505 72.790 117.965 ;
        RECT 72.070 116.605 72.250 117.255 ;
        RECT 72.970 117.055 73.220 117.705 ;
        RECT 72.420 116.725 73.220 117.055 ;
        RECT 68.015 115.415 71.525 116.505 ;
        RECT 71.985 116.435 72.250 116.605 ;
        RECT 72.070 116.395 72.250 116.435 ;
        RECT 72.070 115.725 72.325 116.395 ;
        RECT 72.505 115.415 72.790 116.215 ;
        RECT 72.970 116.135 73.220 116.725 ;
        RECT 73.420 117.370 73.740 117.700 ;
        RECT 73.920 117.485 74.580 117.965 ;
        RECT 74.780 117.575 75.630 117.745 ;
        RECT 73.420 116.475 73.610 117.370 ;
        RECT 73.930 117.045 74.590 117.315 ;
        RECT 74.260 116.985 74.590 117.045 ;
        RECT 73.780 116.815 74.110 116.875 ;
        RECT 74.780 116.815 74.950 117.575 ;
        RECT 76.190 117.505 76.510 117.965 ;
        RECT 76.710 117.325 76.960 117.755 ;
        RECT 77.250 117.525 77.660 117.965 ;
        RECT 77.830 117.585 78.845 117.785 ;
        RECT 75.120 117.155 76.370 117.325 ;
        RECT 75.120 117.035 75.450 117.155 ;
        RECT 73.780 116.645 75.680 116.815 ;
        RECT 73.420 116.305 75.340 116.475 ;
        RECT 73.420 116.285 73.740 116.305 ;
        RECT 72.970 115.625 73.300 116.135 ;
        RECT 73.570 115.675 73.740 116.285 ;
        RECT 75.510 116.135 75.680 116.645 ;
        RECT 75.850 116.575 76.030 116.985 ;
        RECT 76.200 116.395 76.370 117.155 ;
        RECT 73.910 115.415 74.240 116.105 ;
        RECT 74.470 115.965 75.680 116.135 ;
        RECT 75.850 116.085 76.370 116.395 ;
        RECT 76.540 116.985 76.960 117.325 ;
        RECT 77.250 116.985 77.660 117.315 ;
        RECT 76.540 116.215 76.730 116.985 ;
        RECT 77.830 116.855 78.000 117.585 ;
        RECT 79.145 117.415 79.315 117.745 ;
        RECT 79.485 117.585 79.815 117.965 ;
        RECT 78.170 117.035 78.520 117.405 ;
        RECT 77.830 116.815 78.250 116.855 ;
        RECT 76.900 116.645 78.250 116.815 ;
        RECT 76.900 116.485 77.150 116.645 ;
        RECT 77.660 116.215 77.910 116.475 ;
        RECT 76.540 115.965 77.910 116.215 ;
        RECT 74.470 115.675 74.710 115.965 ;
        RECT 75.510 115.885 75.680 115.965 ;
        RECT 74.910 115.415 75.330 115.795 ;
        RECT 75.510 115.635 76.140 115.885 ;
        RECT 76.610 115.415 76.940 115.795 ;
        RECT 77.110 115.675 77.280 115.965 ;
        RECT 78.080 115.800 78.250 116.645 ;
        RECT 78.700 116.475 78.920 117.345 ;
        RECT 79.145 117.225 79.840 117.415 ;
        RECT 78.420 116.095 78.920 116.475 ;
        RECT 79.090 116.425 79.500 117.045 ;
        RECT 79.670 116.255 79.840 117.225 ;
        RECT 79.145 116.085 79.840 116.255 ;
        RECT 77.460 115.415 77.840 115.795 ;
        RECT 78.080 115.630 78.910 115.800 ;
        RECT 79.145 115.585 79.315 116.085 ;
        RECT 79.485 115.415 79.815 115.915 ;
        RECT 80.030 115.585 80.255 117.705 ;
        RECT 80.425 117.585 80.755 117.965 ;
        RECT 80.925 117.415 81.095 117.705 ;
        RECT 80.430 117.245 81.095 117.415 ;
        RECT 81.355 117.290 81.615 117.795 ;
        RECT 81.795 117.585 82.125 117.965 ;
        RECT 82.305 117.415 82.475 117.795 ;
        RECT 80.430 116.255 80.660 117.245 ;
        RECT 80.830 116.425 81.180 117.075 ;
        RECT 81.355 116.490 81.525 117.290 ;
        RECT 81.810 117.245 82.475 117.415 ;
        RECT 81.810 116.990 81.980 117.245 ;
        RECT 82.735 117.195 85.325 117.965 ;
        RECT 85.585 117.415 85.755 117.795 ;
        RECT 85.935 117.585 86.265 117.965 ;
        RECT 85.585 117.245 86.250 117.415 ;
        RECT 86.445 117.290 86.705 117.795 ;
        RECT 81.695 116.660 81.980 116.990 ;
        RECT 82.215 116.695 82.545 117.065 ;
        RECT 81.810 116.515 81.980 116.660 ;
        RECT 80.430 116.085 81.095 116.255 ;
        RECT 80.425 115.415 80.755 115.915 ;
        RECT 80.925 115.585 81.095 116.085 ;
        RECT 81.355 115.585 81.625 116.490 ;
        RECT 81.810 116.345 82.475 116.515 ;
        RECT 81.795 115.415 82.125 116.175 ;
        RECT 82.305 115.585 82.475 116.345 ;
        RECT 82.735 116.505 83.945 117.025 ;
        RECT 84.115 116.675 85.325 117.195 ;
        RECT 85.515 116.695 85.845 117.065 ;
        RECT 86.080 116.990 86.250 117.245 ;
        RECT 86.080 116.660 86.365 116.990 ;
        RECT 86.080 116.515 86.250 116.660 ;
        RECT 82.735 115.415 85.325 116.505 ;
        RECT 85.585 116.345 86.250 116.515 ;
        RECT 86.535 116.490 86.705 117.290 ;
        RECT 86.875 117.240 87.165 117.965 ;
        RECT 87.375 117.145 87.605 117.965 ;
        RECT 87.775 117.165 88.105 117.795 ;
        RECT 87.355 116.725 87.685 116.975 ;
        RECT 85.585 115.585 85.755 116.345 ;
        RECT 85.935 115.415 86.265 116.175 ;
        RECT 86.435 115.585 86.705 116.490 ;
        RECT 86.875 115.415 87.165 116.580 ;
        RECT 87.855 116.565 88.105 117.165 ;
        RECT 88.275 117.145 88.485 117.965 ;
        RECT 88.755 117.145 88.985 117.965 ;
        RECT 89.155 117.165 89.485 117.795 ;
        RECT 88.735 116.725 89.065 116.975 ;
        RECT 89.235 116.565 89.485 117.165 ;
        RECT 89.655 117.145 89.865 117.965 ;
        RECT 90.930 117.625 91.185 117.785 ;
        RECT 90.845 117.455 91.185 117.625 ;
        RECT 91.365 117.505 91.650 117.965 ;
        RECT 90.930 117.255 91.185 117.455 ;
        RECT 87.375 115.415 87.605 116.555 ;
        RECT 87.775 115.585 88.105 116.565 ;
        RECT 88.275 115.415 88.485 116.555 ;
        RECT 88.755 115.415 88.985 116.555 ;
        RECT 89.155 115.585 89.485 116.565 ;
        RECT 89.655 115.415 89.865 116.555 ;
        RECT 90.930 116.395 91.110 117.255 ;
        RECT 91.830 117.055 92.080 117.705 ;
        RECT 91.280 116.725 92.080 117.055 ;
        RECT 90.930 115.725 91.185 116.395 ;
        RECT 91.365 115.415 91.650 116.215 ;
        RECT 91.830 116.135 92.080 116.725 ;
        RECT 92.280 117.370 92.600 117.700 ;
        RECT 92.780 117.485 93.440 117.965 ;
        RECT 93.640 117.575 94.490 117.745 ;
        RECT 92.280 116.475 92.470 117.370 ;
        RECT 92.790 117.045 93.450 117.315 ;
        RECT 93.120 116.985 93.450 117.045 ;
        RECT 92.640 116.815 92.970 116.875 ;
        RECT 93.640 116.815 93.810 117.575 ;
        RECT 95.050 117.505 95.370 117.965 ;
        RECT 95.570 117.325 95.820 117.755 ;
        RECT 96.110 117.525 96.520 117.965 ;
        RECT 96.690 117.585 97.705 117.785 ;
        RECT 93.980 117.155 95.230 117.325 ;
        RECT 93.980 117.035 94.310 117.155 ;
        RECT 92.640 116.645 94.540 116.815 ;
        RECT 92.280 116.305 94.200 116.475 ;
        RECT 92.280 116.285 92.600 116.305 ;
        RECT 91.830 115.625 92.160 116.135 ;
        RECT 92.430 115.675 92.600 116.285 ;
        RECT 94.370 116.135 94.540 116.645 ;
        RECT 94.710 116.575 94.890 116.985 ;
        RECT 95.060 116.395 95.230 117.155 ;
        RECT 92.770 115.415 93.100 116.105 ;
        RECT 93.330 115.965 94.540 116.135 ;
        RECT 94.710 116.085 95.230 116.395 ;
        RECT 95.400 116.985 95.820 117.325 ;
        RECT 96.110 116.985 96.520 117.315 ;
        RECT 95.400 116.215 95.590 116.985 ;
        RECT 96.690 116.855 96.860 117.585 ;
        RECT 98.005 117.415 98.175 117.745 ;
        RECT 98.345 117.585 98.675 117.965 ;
        RECT 97.030 117.035 97.380 117.405 ;
        RECT 96.690 116.815 97.110 116.855 ;
        RECT 95.760 116.645 97.110 116.815 ;
        RECT 95.760 116.485 96.010 116.645 ;
        RECT 96.520 116.215 96.770 116.475 ;
        RECT 95.400 115.965 96.770 116.215 ;
        RECT 93.330 115.675 93.570 115.965 ;
        RECT 94.370 115.885 94.540 115.965 ;
        RECT 93.770 115.415 94.190 115.795 ;
        RECT 94.370 115.635 95.000 115.885 ;
        RECT 95.470 115.415 95.800 115.795 ;
        RECT 95.970 115.675 96.140 115.965 ;
        RECT 96.940 115.800 97.110 116.645 ;
        RECT 97.560 116.475 97.780 117.345 ;
        RECT 98.005 117.225 98.700 117.415 ;
        RECT 97.280 116.095 97.780 116.475 ;
        RECT 97.950 116.425 98.360 117.045 ;
        RECT 98.530 116.255 98.700 117.225 ;
        RECT 98.005 116.085 98.700 116.255 ;
        RECT 96.320 115.415 96.700 115.795 ;
        RECT 96.940 115.630 97.770 115.800 ;
        RECT 98.005 115.585 98.175 116.085 ;
        RECT 98.345 115.415 98.675 115.915 ;
        RECT 98.890 115.585 99.115 117.705 ;
        RECT 99.285 117.585 99.615 117.965 ;
        RECT 99.785 117.415 99.955 117.705 ;
        RECT 101.510 117.625 101.765 117.785 ;
        RECT 101.425 117.455 101.765 117.625 ;
        RECT 101.945 117.505 102.230 117.965 ;
        RECT 99.290 117.245 99.955 117.415 ;
        RECT 101.510 117.255 101.765 117.455 ;
        RECT 99.290 116.255 99.520 117.245 ;
        RECT 99.690 116.425 100.040 117.075 ;
        RECT 101.510 116.395 101.690 117.255 ;
        RECT 102.410 117.055 102.660 117.705 ;
        RECT 101.860 116.725 102.660 117.055 ;
        RECT 99.290 116.085 99.955 116.255 ;
        RECT 99.285 115.415 99.615 115.915 ;
        RECT 99.785 115.585 99.955 116.085 ;
        RECT 101.510 115.725 101.765 116.395 ;
        RECT 101.945 115.415 102.230 116.215 ;
        RECT 102.410 116.135 102.660 116.725 ;
        RECT 102.860 117.370 103.180 117.700 ;
        RECT 103.360 117.485 104.020 117.965 ;
        RECT 104.220 117.575 105.070 117.745 ;
        RECT 102.860 116.475 103.050 117.370 ;
        RECT 103.370 117.045 104.030 117.315 ;
        RECT 103.700 116.985 104.030 117.045 ;
        RECT 103.220 116.815 103.550 116.875 ;
        RECT 104.220 116.815 104.390 117.575 ;
        RECT 105.630 117.505 105.950 117.965 ;
        RECT 106.150 117.325 106.400 117.755 ;
        RECT 106.690 117.525 107.100 117.965 ;
        RECT 107.270 117.585 108.285 117.785 ;
        RECT 104.560 117.155 105.810 117.325 ;
        RECT 104.560 117.035 104.890 117.155 ;
        RECT 103.220 116.645 105.120 116.815 ;
        RECT 102.860 116.305 104.780 116.475 ;
        RECT 102.860 116.285 103.180 116.305 ;
        RECT 102.410 115.625 102.740 116.135 ;
        RECT 103.010 115.675 103.180 116.285 ;
        RECT 104.950 116.135 105.120 116.645 ;
        RECT 105.290 116.575 105.470 116.985 ;
        RECT 105.640 116.395 105.810 117.155 ;
        RECT 103.350 115.415 103.680 116.105 ;
        RECT 103.910 115.965 105.120 116.135 ;
        RECT 105.290 116.085 105.810 116.395 ;
        RECT 105.980 116.985 106.400 117.325 ;
        RECT 106.690 116.985 107.100 117.315 ;
        RECT 105.980 116.215 106.170 116.985 ;
        RECT 107.270 116.855 107.440 117.585 ;
        RECT 108.585 117.415 108.755 117.745 ;
        RECT 108.925 117.585 109.255 117.965 ;
        RECT 107.610 117.035 107.960 117.405 ;
        RECT 107.270 116.815 107.690 116.855 ;
        RECT 106.340 116.645 107.690 116.815 ;
        RECT 106.340 116.485 106.590 116.645 ;
        RECT 107.100 116.215 107.350 116.475 ;
        RECT 105.980 115.965 107.350 116.215 ;
        RECT 103.910 115.675 104.150 115.965 ;
        RECT 104.950 115.885 105.120 115.965 ;
        RECT 104.350 115.415 104.770 115.795 ;
        RECT 104.950 115.635 105.580 115.885 ;
        RECT 106.050 115.415 106.380 115.795 ;
        RECT 106.550 115.675 106.720 115.965 ;
        RECT 107.520 115.800 107.690 116.645 ;
        RECT 108.140 116.475 108.360 117.345 ;
        RECT 108.585 117.225 109.280 117.415 ;
        RECT 107.860 116.095 108.360 116.475 ;
        RECT 108.530 116.425 108.940 117.045 ;
        RECT 109.110 116.255 109.280 117.225 ;
        RECT 108.585 116.085 109.280 116.255 ;
        RECT 106.900 115.415 107.280 115.795 ;
        RECT 107.520 115.630 108.350 115.800 ;
        RECT 108.585 115.585 108.755 116.085 ;
        RECT 108.925 115.415 109.255 115.915 ;
        RECT 109.470 115.585 109.695 117.705 ;
        RECT 109.865 117.585 110.195 117.965 ;
        RECT 110.365 117.415 110.535 117.705 ;
        RECT 109.870 117.245 110.535 117.415 ;
        RECT 110.795 117.290 111.055 117.795 ;
        RECT 111.235 117.585 111.565 117.965 ;
        RECT 111.745 117.415 111.915 117.795 ;
        RECT 109.870 116.255 110.100 117.245 ;
        RECT 110.270 116.425 110.620 117.075 ;
        RECT 110.795 116.490 110.965 117.290 ;
        RECT 111.250 117.245 111.915 117.415 ;
        RECT 111.250 116.990 111.420 117.245 ;
        RECT 112.635 117.240 112.925 117.965 ;
        RECT 113.555 117.195 116.145 117.965 ;
        RECT 111.135 116.660 111.420 116.990 ;
        RECT 111.655 116.695 111.985 117.065 ;
        RECT 111.250 116.515 111.420 116.660 ;
        RECT 109.870 116.085 110.535 116.255 ;
        RECT 109.865 115.415 110.195 115.915 ;
        RECT 110.365 115.585 110.535 116.085 ;
        RECT 110.795 115.585 111.065 116.490 ;
        RECT 111.250 116.345 111.915 116.515 ;
        RECT 111.235 115.415 111.565 116.175 ;
        RECT 111.745 115.585 111.915 116.345 ;
        RECT 112.635 115.415 112.925 116.580 ;
        RECT 113.555 116.505 114.765 117.025 ;
        RECT 114.935 116.675 116.145 117.195 ;
        RECT 116.355 117.145 116.585 117.965 ;
        RECT 116.755 117.165 117.085 117.795 ;
        RECT 116.335 116.725 116.665 116.975 ;
        RECT 116.835 116.565 117.085 117.165 ;
        RECT 117.255 117.145 117.465 117.965 ;
        RECT 118.245 117.415 118.415 117.795 ;
        RECT 118.595 117.585 118.925 117.965 ;
        RECT 118.245 117.245 118.910 117.415 ;
        RECT 119.105 117.290 119.365 117.795 ;
        RECT 118.175 116.695 118.505 117.065 ;
        RECT 118.740 116.990 118.910 117.245 ;
        RECT 113.555 115.415 116.145 116.505 ;
        RECT 116.355 115.415 116.585 116.555 ;
        RECT 116.755 115.585 117.085 116.565 ;
        RECT 118.740 116.660 119.025 116.990 ;
        RECT 117.255 115.415 117.465 116.555 ;
        RECT 118.740 116.515 118.910 116.660 ;
        RECT 118.245 116.345 118.910 116.515 ;
        RECT 119.195 116.490 119.365 117.290 ;
        RECT 119.535 117.215 120.745 117.965 ;
        RECT 118.245 115.585 118.415 116.345 ;
        RECT 118.595 115.415 118.925 116.175 ;
        RECT 119.095 115.585 119.365 116.490 ;
        RECT 119.535 116.505 120.055 117.045 ;
        RECT 120.225 116.675 120.745 117.215 ;
        RECT 120.915 117.195 124.425 117.965 ;
        RECT 124.595 117.215 125.805 117.965 ;
        RECT 120.915 116.505 122.605 117.025 ;
        RECT 122.775 116.675 124.425 117.195 ;
        RECT 124.595 116.505 125.115 117.045 ;
        RECT 125.285 116.675 125.805 117.215 ;
        RECT 119.535 115.415 120.745 116.505 ;
        RECT 120.915 115.415 124.425 116.505 ;
        RECT 124.595 115.415 125.805 116.505 ;
        RECT 11.810 115.245 125.890 115.415 ;
        RECT 11.895 114.155 13.105 115.245 ;
        RECT 11.895 113.445 12.415 113.985 ;
        RECT 12.585 113.615 13.105 114.155 ;
        RECT 13.275 114.155 16.785 115.245 ;
        RECT 16.960 114.810 22.305 115.245 ;
        RECT 13.275 113.635 14.965 114.155 ;
        RECT 15.135 113.465 16.785 113.985 ;
        RECT 18.550 113.560 18.900 114.810 ;
        RECT 22.475 114.080 22.765 115.245 ;
        RECT 22.935 114.155 24.605 115.245 ;
        RECT 24.865 114.315 25.035 115.075 ;
        RECT 25.215 114.485 25.545 115.245 ;
        RECT 11.895 112.695 13.105 113.445 ;
        RECT 13.275 112.695 16.785 113.465 ;
        RECT 20.380 113.240 20.720 114.070 ;
        RECT 22.935 113.635 23.685 114.155 ;
        RECT 24.865 114.145 25.530 114.315 ;
        RECT 25.715 114.170 25.985 115.075 ;
        RECT 25.360 114.000 25.530 114.145 ;
        RECT 23.855 113.465 24.605 113.985 ;
        RECT 24.795 113.595 25.125 113.965 ;
        RECT 25.360 113.670 25.645 114.000 ;
        RECT 16.960 112.695 22.305 113.240 ;
        RECT 22.475 112.695 22.765 113.420 ;
        RECT 22.935 112.695 24.605 113.465 ;
        RECT 25.360 113.415 25.530 113.670 ;
        RECT 24.865 113.245 25.530 113.415 ;
        RECT 25.815 113.370 25.985 114.170 ;
        RECT 26.615 114.155 30.125 115.245 ;
        RECT 30.300 114.810 35.645 115.245 ;
        RECT 35.820 114.810 41.165 115.245 ;
        RECT 41.340 114.810 46.685 115.245 ;
        RECT 26.615 113.635 28.305 114.155 ;
        RECT 28.475 113.465 30.125 113.985 ;
        RECT 31.890 113.560 32.240 114.810 ;
        RECT 24.865 112.865 25.035 113.245 ;
        RECT 25.215 112.695 25.545 113.075 ;
        RECT 25.725 112.865 25.985 113.370 ;
        RECT 26.615 112.695 30.125 113.465 ;
        RECT 33.720 113.240 34.060 114.070 ;
        RECT 37.410 113.560 37.760 114.810 ;
        RECT 39.240 113.240 39.580 114.070 ;
        RECT 42.930 113.560 43.280 114.810 ;
        RECT 46.895 114.105 47.125 115.245 ;
        RECT 47.295 114.095 47.625 115.075 ;
        RECT 47.795 114.105 48.005 115.245 ;
        RECT 44.760 113.240 45.100 114.070 ;
        RECT 46.875 113.685 47.205 113.935 ;
        RECT 30.300 112.695 35.645 113.240 ;
        RECT 35.820 112.695 41.165 113.240 ;
        RECT 41.340 112.695 46.685 113.240 ;
        RECT 46.895 112.695 47.125 113.515 ;
        RECT 47.375 113.495 47.625 114.095 ;
        RECT 48.235 114.080 48.525 115.245 ;
        RECT 49.620 114.105 49.955 115.075 ;
        RECT 50.125 114.105 50.295 115.245 ;
        RECT 50.465 114.905 52.495 115.075 ;
        RECT 47.295 112.865 47.625 113.495 ;
        RECT 47.795 112.695 48.005 113.515 ;
        RECT 49.620 113.435 49.790 114.105 ;
        RECT 50.465 113.935 50.635 114.905 ;
        RECT 49.960 113.605 50.215 113.935 ;
        RECT 50.440 113.605 50.635 113.935 ;
        RECT 50.805 114.565 51.930 114.735 ;
        RECT 50.045 113.435 50.215 113.605 ;
        RECT 50.805 113.435 50.975 114.565 ;
        RECT 48.235 112.695 48.525 113.420 ;
        RECT 49.620 112.865 49.875 113.435 ;
        RECT 50.045 113.265 50.975 113.435 ;
        RECT 51.145 114.225 52.155 114.395 ;
        RECT 51.145 113.425 51.315 114.225 ;
        RECT 51.520 113.885 51.795 114.025 ;
        RECT 51.515 113.715 51.795 113.885 ;
        RECT 50.800 113.230 50.975 113.265 ;
        RECT 50.045 112.695 50.375 113.095 ;
        RECT 50.800 112.865 51.330 113.230 ;
        RECT 51.520 112.865 51.795 113.715 ;
        RECT 51.965 112.865 52.155 114.225 ;
        RECT 52.325 114.240 52.495 114.905 ;
        RECT 52.665 114.485 52.835 115.245 ;
        RECT 53.070 114.485 53.585 114.895 ;
        RECT 52.325 114.050 53.075 114.240 ;
        RECT 53.245 113.675 53.585 114.485 ;
        RECT 54.305 114.315 54.475 115.075 ;
        RECT 54.655 114.485 54.985 115.245 ;
        RECT 54.305 114.145 54.970 114.315 ;
        RECT 55.155 114.170 55.425 115.075 ;
        RECT 54.800 114.000 54.970 114.145 ;
        RECT 52.355 113.505 53.585 113.675 ;
        RECT 54.235 113.595 54.565 113.965 ;
        RECT 54.800 113.670 55.085 114.000 ;
        RECT 52.335 112.695 52.845 113.230 ;
        RECT 53.065 112.900 53.310 113.505 ;
        RECT 54.800 113.415 54.970 113.670 ;
        RECT 54.305 113.245 54.970 113.415 ;
        RECT 55.255 113.370 55.425 114.170 ;
        RECT 55.595 114.155 56.805 115.245 ;
        RECT 56.975 114.155 60.485 115.245 ;
        RECT 61.030 114.905 61.285 114.935 ;
        RECT 60.945 114.735 61.285 114.905 ;
        RECT 61.030 114.265 61.285 114.735 ;
        RECT 61.465 114.445 61.750 115.245 ;
        RECT 61.930 114.525 62.260 115.035 ;
        RECT 55.595 113.615 56.115 114.155 ;
        RECT 56.285 113.445 56.805 113.985 ;
        RECT 56.975 113.635 58.665 114.155 ;
        RECT 58.835 113.465 60.485 113.985 ;
        RECT 54.305 112.865 54.475 113.245 ;
        RECT 54.655 112.695 54.985 113.075 ;
        RECT 55.165 112.865 55.425 113.370 ;
        RECT 55.595 112.695 56.805 113.445 ;
        RECT 56.975 112.695 60.485 113.465 ;
        RECT 61.030 113.405 61.210 114.265 ;
        RECT 61.930 113.935 62.180 114.525 ;
        RECT 62.530 114.375 62.700 114.985 ;
        RECT 62.870 114.555 63.200 115.245 ;
        RECT 63.430 114.695 63.670 114.985 ;
        RECT 63.870 114.865 64.290 115.245 ;
        RECT 64.470 114.775 65.100 115.025 ;
        RECT 65.570 114.865 65.900 115.245 ;
        RECT 64.470 114.695 64.640 114.775 ;
        RECT 66.070 114.695 66.240 114.985 ;
        RECT 66.420 114.865 66.800 115.245 ;
        RECT 67.040 114.860 67.870 115.030 ;
        RECT 63.430 114.525 64.640 114.695 ;
        RECT 61.380 113.605 62.180 113.935 ;
        RECT 61.030 112.875 61.285 113.405 ;
        RECT 61.465 112.695 61.750 113.155 ;
        RECT 61.930 112.955 62.180 113.605 ;
        RECT 62.380 114.355 62.700 114.375 ;
        RECT 62.380 114.185 64.300 114.355 ;
        RECT 62.380 113.290 62.570 114.185 ;
        RECT 64.470 114.015 64.640 114.525 ;
        RECT 64.810 114.265 65.330 114.575 ;
        RECT 62.740 113.845 64.640 114.015 ;
        RECT 62.740 113.785 63.070 113.845 ;
        RECT 63.220 113.615 63.550 113.675 ;
        RECT 62.890 113.345 63.550 113.615 ;
        RECT 62.380 112.960 62.700 113.290 ;
        RECT 62.880 112.695 63.540 113.175 ;
        RECT 63.740 113.085 63.910 113.845 ;
        RECT 64.810 113.675 64.990 114.085 ;
        RECT 64.080 113.505 64.410 113.625 ;
        RECT 65.160 113.505 65.330 114.265 ;
        RECT 64.080 113.335 65.330 113.505 ;
        RECT 65.500 114.445 66.870 114.695 ;
        RECT 65.500 113.675 65.690 114.445 ;
        RECT 66.620 114.185 66.870 114.445 ;
        RECT 65.860 114.015 66.110 114.175 ;
        RECT 67.040 114.015 67.210 114.860 ;
        RECT 68.105 114.575 68.275 115.075 ;
        RECT 68.445 114.745 68.775 115.245 ;
        RECT 67.380 114.185 67.880 114.565 ;
        RECT 68.105 114.405 68.800 114.575 ;
        RECT 65.860 113.845 67.210 114.015 ;
        RECT 66.790 113.805 67.210 113.845 ;
        RECT 65.500 113.335 65.920 113.675 ;
        RECT 66.210 113.345 66.620 113.675 ;
        RECT 63.740 112.915 64.590 113.085 ;
        RECT 65.150 112.695 65.470 113.155 ;
        RECT 65.670 112.905 65.920 113.335 ;
        RECT 66.210 112.695 66.620 113.135 ;
        RECT 66.790 113.075 66.960 113.805 ;
        RECT 67.130 113.255 67.480 113.625 ;
        RECT 67.660 113.315 67.880 114.185 ;
        RECT 68.050 113.615 68.460 114.235 ;
        RECT 68.630 113.435 68.800 114.405 ;
        RECT 68.105 113.245 68.800 113.435 ;
        RECT 66.790 112.875 67.805 113.075 ;
        RECT 68.105 112.915 68.275 113.245 ;
        RECT 68.445 112.695 68.775 113.075 ;
        RECT 68.990 112.955 69.215 115.075 ;
        RECT 69.385 114.745 69.715 115.245 ;
        RECT 69.885 114.575 70.055 115.075 ;
        RECT 69.390 114.405 70.055 114.575 ;
        RECT 69.390 113.415 69.620 114.405 ;
        RECT 69.790 113.585 70.140 114.235 ;
        RECT 70.315 114.155 73.825 115.245 ;
        RECT 70.315 113.635 72.005 114.155 ;
        RECT 73.995 114.080 74.285 115.245 ;
        RECT 74.455 114.155 77.965 115.245 ;
        RECT 78.225 114.315 78.395 115.075 ;
        RECT 78.575 114.485 78.905 115.245 ;
        RECT 72.175 113.465 73.825 113.985 ;
        RECT 74.455 113.635 76.145 114.155 ;
        RECT 78.225 114.145 78.890 114.315 ;
        RECT 79.075 114.170 79.345 115.075 ;
        RECT 78.720 114.000 78.890 114.145 ;
        RECT 76.315 113.465 77.965 113.985 ;
        RECT 78.155 113.595 78.485 113.965 ;
        RECT 78.720 113.670 79.005 114.000 ;
        RECT 69.390 113.245 70.055 113.415 ;
        RECT 69.385 112.695 69.715 113.075 ;
        RECT 69.885 112.955 70.055 113.245 ;
        RECT 70.315 112.695 73.825 113.465 ;
        RECT 73.995 112.695 74.285 113.420 ;
        RECT 74.455 112.695 77.965 113.465 ;
        RECT 78.720 113.415 78.890 113.670 ;
        RECT 78.225 113.245 78.890 113.415 ;
        RECT 79.175 113.370 79.345 114.170 ;
        RECT 79.515 114.155 83.025 115.245 ;
        RECT 83.200 114.810 88.545 115.245 ;
        RECT 88.720 114.810 94.065 115.245 ;
        RECT 94.240 114.810 99.585 115.245 ;
        RECT 79.515 113.635 81.205 114.155 ;
        RECT 81.375 113.465 83.025 113.985 ;
        RECT 84.790 113.560 85.140 114.810 ;
        RECT 78.225 112.865 78.395 113.245 ;
        RECT 78.575 112.695 78.905 113.075 ;
        RECT 79.085 112.865 79.345 113.370 ;
        RECT 79.515 112.695 83.025 113.465 ;
        RECT 86.620 113.240 86.960 114.070 ;
        RECT 90.310 113.560 90.660 114.810 ;
        RECT 92.140 113.240 92.480 114.070 ;
        RECT 95.830 113.560 96.180 114.810 ;
        RECT 99.755 114.080 100.045 115.245 ;
        RECT 100.215 114.155 101.425 115.245 ;
        RECT 101.595 114.155 105.105 115.245 ;
        RECT 105.280 114.810 110.625 115.245 ;
        RECT 110.800 114.810 116.145 115.245 ;
        RECT 97.660 113.240 98.000 114.070 ;
        RECT 100.215 113.615 100.735 114.155 ;
        RECT 100.905 113.445 101.425 113.985 ;
        RECT 101.595 113.635 103.285 114.155 ;
        RECT 103.455 113.465 105.105 113.985 ;
        RECT 106.870 113.560 107.220 114.810 ;
        RECT 83.200 112.695 88.545 113.240 ;
        RECT 88.720 112.695 94.065 113.240 ;
        RECT 94.240 112.695 99.585 113.240 ;
        RECT 99.755 112.695 100.045 113.420 ;
        RECT 100.215 112.695 101.425 113.445 ;
        RECT 101.595 112.695 105.105 113.465 ;
        RECT 108.700 113.240 109.040 114.070 ;
        RECT 112.390 113.560 112.740 114.810 ;
        RECT 116.355 114.105 116.585 115.245 ;
        RECT 116.755 114.095 117.085 115.075 ;
        RECT 117.255 114.105 117.465 115.245 ;
        RECT 117.695 114.170 117.965 115.075 ;
        RECT 118.135 114.485 118.465 115.245 ;
        RECT 118.645 114.315 118.815 115.075 ;
        RECT 114.220 113.240 114.560 114.070 ;
        RECT 116.335 113.685 116.665 113.935 ;
        RECT 105.280 112.695 110.625 113.240 ;
        RECT 110.800 112.695 116.145 113.240 ;
        RECT 116.355 112.695 116.585 113.515 ;
        RECT 116.835 113.495 117.085 114.095 ;
        RECT 116.755 112.865 117.085 113.495 ;
        RECT 117.255 112.695 117.465 113.515 ;
        RECT 117.695 113.370 117.865 114.170 ;
        RECT 118.150 114.145 118.815 114.315 ;
        RECT 119.165 114.315 119.335 115.075 ;
        RECT 119.515 114.485 119.845 115.245 ;
        RECT 119.165 114.145 119.830 114.315 ;
        RECT 120.015 114.170 120.285 115.075 ;
        RECT 118.150 114.000 118.320 114.145 ;
        RECT 118.035 113.670 118.320 114.000 ;
        RECT 119.660 114.000 119.830 114.145 ;
        RECT 118.150 113.415 118.320 113.670 ;
        RECT 118.555 113.595 118.885 113.965 ;
        RECT 119.095 113.595 119.425 113.965 ;
        RECT 119.660 113.670 119.945 114.000 ;
        RECT 119.660 113.415 119.830 113.670 ;
        RECT 117.695 112.865 117.955 113.370 ;
        RECT 118.150 113.245 118.815 113.415 ;
        RECT 118.135 112.695 118.465 113.075 ;
        RECT 118.645 112.865 118.815 113.245 ;
        RECT 119.165 113.245 119.830 113.415 ;
        RECT 120.115 113.370 120.285 114.170 ;
        RECT 120.455 114.155 123.045 115.245 ;
        RECT 123.215 114.170 123.485 115.075 ;
        RECT 123.655 114.485 123.985 115.245 ;
        RECT 124.165 114.315 124.345 115.075 ;
        RECT 120.455 113.635 121.665 114.155 ;
        RECT 121.835 113.465 123.045 113.985 ;
        RECT 119.165 112.865 119.335 113.245 ;
        RECT 119.515 112.695 119.845 113.075 ;
        RECT 120.025 112.865 120.285 113.370 ;
        RECT 120.455 112.695 123.045 113.465 ;
        RECT 123.215 113.370 123.395 114.170 ;
        RECT 123.670 114.145 124.345 114.315 ;
        RECT 124.595 114.155 125.805 115.245 ;
        RECT 123.670 114.000 123.840 114.145 ;
        RECT 123.565 113.670 123.840 114.000 ;
        RECT 123.670 113.415 123.840 113.670 ;
        RECT 124.065 113.595 124.405 113.965 ;
        RECT 124.595 113.615 125.115 114.155 ;
        RECT 125.285 113.445 125.805 113.985 ;
        RECT 123.215 112.865 123.475 113.370 ;
        RECT 123.670 113.245 124.335 113.415 ;
        RECT 123.655 112.695 123.985 113.075 ;
        RECT 124.165 112.865 124.335 113.245 ;
        RECT 124.595 112.695 125.805 113.445 ;
        RECT 11.810 112.525 125.890 112.695 ;
        RECT 11.895 111.775 13.105 112.525 ;
        RECT 11.895 111.235 12.415 111.775 ;
        RECT 13.275 111.755 16.785 112.525 ;
        RECT 17.265 112.055 17.435 112.525 ;
        RECT 17.605 111.875 17.935 112.355 ;
        RECT 18.105 112.055 18.275 112.525 ;
        RECT 18.445 111.875 18.775 112.355 ;
        RECT 12.585 111.065 13.105 111.605 ;
        RECT 11.895 109.975 13.105 111.065 ;
        RECT 13.275 111.065 14.965 111.585 ;
        RECT 15.135 111.235 16.785 111.755 ;
        RECT 17.010 111.705 18.775 111.875 ;
        RECT 18.945 111.715 19.115 112.525 ;
        RECT 19.315 112.145 20.385 112.315 ;
        RECT 19.315 111.790 19.635 112.145 ;
        RECT 17.010 111.155 17.420 111.705 ;
        RECT 19.310 111.535 19.635 111.790 ;
        RECT 17.605 111.325 19.635 111.535 ;
        RECT 19.290 111.315 19.635 111.325 ;
        RECT 19.805 111.575 20.045 111.975 ;
        RECT 20.215 111.915 20.385 112.145 ;
        RECT 20.555 112.085 20.745 112.525 ;
        RECT 20.915 112.075 21.865 112.355 ;
        RECT 22.085 112.165 22.435 112.335 ;
        RECT 20.215 111.745 20.745 111.915 ;
        RECT 13.275 109.975 16.785 111.065 ;
        RECT 17.010 110.985 18.735 111.155 ;
        RECT 17.265 109.975 17.435 110.815 ;
        RECT 17.645 110.145 17.895 110.985 ;
        RECT 18.105 109.975 18.275 110.815 ;
        RECT 18.445 110.145 18.735 110.985 ;
        RECT 18.945 109.975 19.115 111.035 ;
        RECT 19.290 110.695 19.460 111.315 ;
        RECT 19.805 111.205 20.345 111.575 ;
        RECT 20.525 111.465 20.745 111.745 ;
        RECT 20.915 111.295 21.085 112.075 ;
        RECT 20.680 111.125 21.085 111.295 ;
        RECT 21.255 111.285 21.605 111.905 ;
        RECT 20.680 111.035 20.850 111.125 ;
        RECT 21.775 111.115 21.985 111.905 ;
        RECT 19.630 110.865 20.850 111.035 ;
        RECT 21.310 110.955 21.985 111.115 ;
        RECT 19.290 110.525 20.090 110.695 ;
        RECT 19.410 109.975 19.740 110.355 ;
        RECT 19.920 110.235 20.090 110.525 ;
        RECT 20.680 110.485 20.850 110.865 ;
        RECT 21.020 110.945 21.985 110.955 ;
        RECT 22.175 111.775 22.435 112.165 ;
        RECT 22.645 112.065 22.975 112.525 ;
        RECT 23.850 112.135 24.705 112.305 ;
        RECT 24.910 112.135 25.405 112.305 ;
        RECT 25.575 112.165 25.905 112.525 ;
        RECT 22.175 111.085 22.345 111.775 ;
        RECT 22.515 111.425 22.685 111.605 ;
        RECT 22.855 111.595 23.645 111.845 ;
        RECT 23.850 111.425 24.020 112.135 ;
        RECT 24.190 111.625 24.545 111.845 ;
        RECT 22.515 111.255 24.205 111.425 ;
        RECT 21.020 110.655 21.480 110.945 ;
        RECT 22.175 110.915 23.675 111.085 ;
        RECT 22.175 110.775 22.345 110.915 ;
        RECT 21.785 110.605 22.345 110.775 ;
        RECT 20.260 109.975 20.510 110.435 ;
        RECT 20.680 110.145 21.550 110.485 ;
        RECT 21.785 110.145 21.955 110.605 ;
        RECT 22.790 110.575 23.865 110.745 ;
        RECT 22.125 109.975 22.495 110.435 ;
        RECT 22.790 110.235 22.960 110.575 ;
        RECT 23.130 109.975 23.460 110.405 ;
        RECT 23.695 110.235 23.865 110.575 ;
        RECT 24.035 110.475 24.205 111.255 ;
        RECT 24.375 111.035 24.545 111.625 ;
        RECT 24.715 111.225 25.065 111.845 ;
        RECT 24.375 110.645 24.840 111.035 ;
        RECT 25.235 110.775 25.405 112.135 ;
        RECT 25.575 110.945 26.035 111.995 ;
        RECT 25.010 110.605 25.405 110.775 ;
        RECT 25.010 110.475 25.180 110.605 ;
        RECT 24.035 110.145 24.715 110.475 ;
        RECT 24.930 110.145 25.180 110.475 ;
        RECT 25.350 109.975 25.600 110.435 ;
        RECT 25.770 110.160 26.095 110.945 ;
        RECT 26.265 110.145 26.435 112.265 ;
        RECT 26.605 112.145 26.935 112.525 ;
        RECT 27.105 111.975 27.360 112.265 ;
        RECT 26.610 111.805 27.360 111.975 ;
        RECT 26.610 110.815 26.840 111.805 ;
        RECT 27.535 111.775 28.745 112.525 ;
        RECT 27.010 110.985 27.360 111.635 ;
        RECT 27.535 111.065 28.055 111.605 ;
        RECT 28.225 111.235 28.745 111.775 ;
        RECT 28.915 111.850 29.175 112.355 ;
        RECT 29.355 112.145 29.685 112.525 ;
        RECT 29.865 111.975 30.035 112.355 ;
        RECT 26.610 110.645 27.360 110.815 ;
        RECT 26.605 109.975 26.935 110.475 ;
        RECT 27.105 110.145 27.360 110.645 ;
        RECT 27.535 109.975 28.745 111.065 ;
        RECT 28.915 111.050 29.085 111.850 ;
        RECT 29.370 111.805 30.035 111.975 ;
        RECT 29.370 111.550 29.540 111.805 ;
        RECT 30.355 111.705 30.565 112.525 ;
        RECT 30.735 111.725 31.065 112.355 ;
        RECT 29.255 111.220 29.540 111.550 ;
        RECT 29.775 111.255 30.105 111.625 ;
        RECT 29.370 111.075 29.540 111.220 ;
        RECT 30.735 111.125 30.985 111.725 ;
        RECT 31.235 111.705 31.465 112.525 ;
        RECT 32.595 111.850 32.855 112.355 ;
        RECT 33.035 112.145 33.365 112.525 ;
        RECT 33.545 111.975 33.715 112.355 ;
        RECT 31.155 111.285 31.485 111.535 ;
        RECT 28.915 110.145 29.185 111.050 ;
        RECT 29.370 110.905 30.035 111.075 ;
        RECT 29.355 109.975 29.685 110.735 ;
        RECT 29.865 110.145 30.035 110.905 ;
        RECT 30.355 109.975 30.565 111.115 ;
        RECT 30.735 110.145 31.065 111.125 ;
        RECT 31.235 109.975 31.465 111.115 ;
        RECT 32.595 111.050 32.765 111.850 ;
        RECT 33.050 111.805 33.715 111.975 ;
        RECT 34.065 111.975 34.235 112.355 ;
        RECT 34.415 112.145 34.745 112.525 ;
        RECT 34.065 111.805 34.730 111.975 ;
        RECT 34.925 111.850 35.185 112.355 ;
        RECT 33.050 111.550 33.220 111.805 ;
        RECT 32.935 111.220 33.220 111.550 ;
        RECT 33.455 111.255 33.785 111.625 ;
        RECT 33.995 111.255 34.325 111.625 ;
        RECT 34.560 111.550 34.730 111.805 ;
        RECT 33.050 111.075 33.220 111.220 ;
        RECT 34.560 111.220 34.845 111.550 ;
        RECT 34.560 111.075 34.730 111.220 ;
        RECT 32.595 110.145 32.865 111.050 ;
        RECT 33.050 110.905 33.715 111.075 ;
        RECT 33.035 109.975 33.365 110.735 ;
        RECT 33.545 110.145 33.715 110.905 ;
        RECT 34.065 110.905 34.730 111.075 ;
        RECT 35.015 111.050 35.185 111.850 ;
        RECT 35.355 111.800 35.645 112.525 ;
        RECT 36.425 111.725 36.755 112.525 ;
        RECT 36.925 111.875 37.095 112.355 ;
        RECT 37.265 112.045 37.595 112.525 ;
        RECT 37.765 111.875 37.935 112.355 ;
        RECT 38.185 112.045 38.425 112.525 ;
        RECT 38.605 111.875 38.775 112.355 ;
        RECT 36.925 111.705 37.935 111.875 ;
        RECT 38.140 111.705 38.775 111.875 ;
        RECT 39.535 111.705 39.765 112.525 ;
        RECT 39.935 111.725 40.265 112.355 ;
        RECT 36.925 111.675 37.425 111.705 ;
        RECT 36.925 111.165 37.420 111.675 ;
        RECT 38.140 111.535 38.310 111.705 ;
        RECT 37.810 111.365 38.310 111.535 ;
        RECT 34.065 110.145 34.235 110.905 ;
        RECT 34.415 109.975 34.745 110.735 ;
        RECT 34.915 110.145 35.185 111.050 ;
        RECT 35.355 109.975 35.645 111.140 ;
        RECT 36.425 109.975 36.755 111.125 ;
        RECT 36.925 110.995 37.935 111.165 ;
        RECT 36.925 110.145 37.095 110.995 ;
        RECT 37.265 109.975 37.595 110.775 ;
        RECT 37.765 110.145 37.935 110.995 ;
        RECT 38.140 111.125 38.310 111.365 ;
        RECT 38.480 111.295 38.860 111.535 ;
        RECT 39.515 111.285 39.845 111.535 ;
        RECT 40.015 111.125 40.265 111.725 ;
        RECT 40.435 111.705 40.645 112.525 ;
        RECT 40.875 111.850 41.135 112.355 ;
        RECT 41.315 112.145 41.645 112.525 ;
        RECT 41.825 111.975 41.995 112.355 ;
        RECT 38.140 110.955 38.855 111.125 ;
        RECT 38.115 109.975 38.355 110.775 ;
        RECT 38.525 110.145 38.855 110.955 ;
        RECT 39.535 109.975 39.765 111.115 ;
        RECT 39.935 110.145 40.265 111.125 ;
        RECT 40.435 109.975 40.645 111.115 ;
        RECT 40.875 111.050 41.045 111.850 ;
        RECT 41.330 111.805 41.995 111.975 ;
        RECT 42.805 111.975 42.975 112.355 ;
        RECT 43.155 112.145 43.485 112.525 ;
        RECT 42.805 111.805 43.470 111.975 ;
        RECT 43.665 111.850 43.925 112.355 ;
        RECT 41.330 111.550 41.500 111.805 ;
        RECT 41.215 111.220 41.500 111.550 ;
        RECT 41.735 111.255 42.065 111.625 ;
        RECT 42.735 111.255 43.065 111.625 ;
        RECT 43.300 111.550 43.470 111.805 ;
        RECT 41.330 111.075 41.500 111.220 ;
        RECT 43.300 111.220 43.585 111.550 ;
        RECT 43.300 111.075 43.470 111.220 ;
        RECT 40.875 110.145 41.145 111.050 ;
        RECT 41.330 110.905 41.995 111.075 ;
        RECT 41.315 109.975 41.645 110.735 ;
        RECT 41.825 110.145 41.995 110.905 ;
        RECT 42.805 110.905 43.470 111.075 ;
        RECT 43.755 111.050 43.925 111.850 ;
        RECT 44.645 111.975 44.815 112.265 ;
        RECT 44.985 112.145 45.315 112.525 ;
        RECT 44.645 111.805 45.310 111.975 ;
        RECT 42.805 110.145 42.975 110.905 ;
        RECT 43.155 109.975 43.485 110.735 ;
        RECT 43.655 110.145 43.925 111.050 ;
        RECT 44.560 110.985 44.910 111.635 ;
        RECT 45.080 110.815 45.310 111.805 ;
        RECT 44.645 110.645 45.310 110.815 ;
        RECT 44.645 110.145 44.815 110.645 ;
        RECT 44.985 109.975 45.315 110.475 ;
        RECT 45.485 110.145 45.710 112.265 ;
        RECT 45.925 112.145 46.255 112.525 ;
        RECT 46.425 111.975 46.595 112.305 ;
        RECT 46.895 112.145 47.910 112.345 ;
        RECT 45.900 111.785 46.595 111.975 ;
        RECT 45.900 110.815 46.070 111.785 ;
        RECT 46.240 110.985 46.650 111.605 ;
        RECT 46.820 111.035 47.040 111.905 ;
        RECT 47.220 111.595 47.570 111.965 ;
        RECT 47.740 111.415 47.910 112.145 ;
        RECT 48.080 112.085 48.490 112.525 ;
        RECT 48.780 111.885 49.030 112.315 ;
        RECT 49.230 112.065 49.550 112.525 ;
        RECT 50.110 112.135 50.960 112.305 ;
        RECT 48.080 111.545 48.490 111.875 ;
        RECT 48.780 111.545 49.200 111.885 ;
        RECT 47.490 111.375 47.910 111.415 ;
        RECT 47.490 111.205 48.840 111.375 ;
        RECT 45.900 110.645 46.595 110.815 ;
        RECT 46.820 110.655 47.320 111.035 ;
        RECT 45.925 109.975 46.255 110.475 ;
        RECT 46.425 110.145 46.595 110.645 ;
        RECT 47.490 110.360 47.660 111.205 ;
        RECT 48.590 111.045 48.840 111.205 ;
        RECT 47.830 110.775 48.080 111.035 ;
        RECT 49.010 110.775 49.200 111.545 ;
        RECT 47.830 110.525 49.200 110.775 ;
        RECT 49.370 111.715 50.620 111.885 ;
        RECT 49.370 110.955 49.540 111.715 ;
        RECT 50.290 111.595 50.620 111.715 ;
        RECT 49.710 111.135 49.890 111.545 ;
        RECT 50.790 111.375 50.960 112.135 ;
        RECT 51.160 112.045 51.820 112.525 ;
        RECT 52.000 111.930 52.320 112.260 ;
        RECT 51.150 111.605 51.810 111.875 ;
        RECT 51.150 111.545 51.480 111.605 ;
        RECT 51.630 111.375 51.960 111.435 ;
        RECT 50.060 111.205 51.960 111.375 ;
        RECT 49.370 110.645 49.890 110.955 ;
        RECT 50.060 110.695 50.230 111.205 ;
        RECT 52.130 111.035 52.320 111.930 ;
        RECT 50.400 110.865 52.320 111.035 ;
        RECT 52.000 110.845 52.320 110.865 ;
        RECT 52.520 111.615 52.770 112.265 ;
        RECT 52.950 112.065 53.235 112.525 ;
        RECT 53.415 112.185 53.670 112.345 ;
        RECT 53.415 112.015 53.755 112.185 ;
        RECT 53.415 111.815 53.670 112.015 ;
        RECT 52.520 111.285 53.320 111.615 ;
        RECT 50.060 110.525 51.270 110.695 ;
        RECT 46.830 110.190 47.660 110.360 ;
        RECT 47.900 109.975 48.280 110.355 ;
        RECT 48.460 110.235 48.630 110.525 ;
        RECT 50.060 110.445 50.230 110.525 ;
        RECT 48.800 109.975 49.130 110.355 ;
        RECT 49.600 110.195 50.230 110.445 ;
        RECT 50.410 109.975 50.830 110.355 ;
        RECT 51.030 110.235 51.270 110.525 ;
        RECT 51.500 109.975 51.830 110.665 ;
        RECT 52.000 110.235 52.170 110.845 ;
        RECT 52.520 110.695 52.770 111.285 ;
        RECT 53.490 110.955 53.670 111.815 ;
        RECT 54.215 111.775 55.425 112.525 ;
        RECT 55.600 111.980 60.945 112.525 ;
        RECT 52.440 110.185 52.770 110.695 ;
        RECT 52.950 109.975 53.235 110.775 ;
        RECT 53.415 110.285 53.670 110.955 ;
        RECT 54.215 111.065 54.735 111.605 ;
        RECT 54.905 111.235 55.425 111.775 ;
        RECT 54.215 109.975 55.425 111.065 ;
        RECT 57.190 110.410 57.540 111.660 ;
        RECT 59.020 111.150 59.360 111.980 ;
        RECT 61.115 111.800 61.405 112.525 ;
        RECT 61.665 111.975 61.835 112.355 ;
        RECT 62.015 112.145 62.345 112.525 ;
        RECT 61.665 111.805 62.330 111.975 ;
        RECT 62.525 111.850 62.785 112.355 ;
        RECT 61.595 111.255 61.925 111.625 ;
        RECT 62.160 111.550 62.330 111.805 ;
        RECT 62.160 111.220 62.445 111.550 ;
        RECT 55.600 109.975 60.945 110.410 ;
        RECT 61.115 109.975 61.405 111.140 ;
        RECT 62.160 111.075 62.330 111.220 ;
        RECT 61.665 110.905 62.330 111.075 ;
        RECT 62.615 111.050 62.785 111.850 ;
        RECT 62.955 111.775 64.165 112.525 ;
        RECT 61.665 110.145 61.835 110.905 ;
        RECT 62.015 109.975 62.345 110.735 ;
        RECT 62.515 110.145 62.785 111.050 ;
        RECT 62.955 111.065 63.475 111.605 ;
        RECT 63.645 111.235 64.165 111.775 ;
        RECT 64.395 111.705 64.605 112.525 ;
        RECT 64.775 111.725 65.105 112.355 ;
        RECT 64.775 111.125 65.025 111.725 ;
        RECT 65.275 111.705 65.505 112.525 ;
        RECT 66.175 111.755 68.765 112.525 ;
        RECT 68.940 111.980 74.285 112.525 ;
        RECT 65.195 111.285 65.525 111.535 ;
        RECT 62.955 109.975 64.165 111.065 ;
        RECT 64.395 109.975 64.605 111.115 ;
        RECT 64.775 110.145 65.105 111.125 ;
        RECT 65.275 109.975 65.505 111.115 ;
        RECT 66.175 111.065 67.385 111.585 ;
        RECT 67.555 111.235 68.765 111.755 ;
        RECT 66.175 109.975 68.765 111.065 ;
        RECT 70.530 110.410 70.880 111.660 ;
        RECT 72.360 111.150 72.700 111.980 ;
        RECT 74.545 111.975 74.715 112.355 ;
        RECT 74.895 112.145 75.225 112.525 ;
        RECT 74.545 111.805 75.210 111.975 ;
        RECT 75.405 111.850 75.665 112.355 ;
        RECT 74.475 111.255 74.805 111.625 ;
        RECT 75.040 111.550 75.210 111.805 ;
        RECT 75.040 111.220 75.325 111.550 ;
        RECT 75.040 111.075 75.210 111.220 ;
        RECT 74.545 110.905 75.210 111.075 ;
        RECT 75.495 111.050 75.665 111.850 ;
        RECT 75.925 111.875 76.095 112.355 ;
        RECT 76.275 112.045 76.515 112.525 ;
        RECT 76.765 111.875 76.935 112.355 ;
        RECT 77.105 112.045 77.435 112.525 ;
        RECT 77.605 111.875 77.775 112.355 ;
        RECT 75.925 111.705 76.560 111.875 ;
        RECT 76.765 111.705 77.775 111.875 ;
        RECT 77.945 111.725 78.275 112.525 ;
        RECT 78.595 111.755 81.185 112.525 ;
        RECT 81.360 111.980 86.705 112.525 ;
        RECT 76.390 111.535 76.560 111.705 ;
        RECT 75.840 111.295 76.220 111.535 ;
        RECT 76.390 111.365 76.890 111.535 ;
        RECT 76.390 111.125 76.560 111.365 ;
        RECT 77.280 111.165 77.775 111.705 ;
        RECT 68.940 109.975 74.285 110.410 ;
        RECT 74.545 110.145 74.715 110.905 ;
        RECT 74.895 109.975 75.225 110.735 ;
        RECT 75.395 110.145 75.665 111.050 ;
        RECT 75.845 110.955 76.560 111.125 ;
        RECT 76.765 110.995 77.775 111.165 ;
        RECT 75.845 110.145 76.175 110.955 ;
        RECT 76.345 109.975 76.585 110.775 ;
        RECT 76.765 110.145 76.935 110.995 ;
        RECT 77.105 109.975 77.435 110.775 ;
        RECT 77.605 110.145 77.775 110.995 ;
        RECT 77.945 109.975 78.275 111.125 ;
        RECT 78.595 111.065 79.805 111.585 ;
        RECT 79.975 111.235 81.185 111.755 ;
        RECT 78.595 109.975 81.185 111.065 ;
        RECT 82.950 110.410 83.300 111.660 ;
        RECT 84.780 111.150 85.120 111.980 ;
        RECT 86.875 111.800 87.165 112.525 ;
        RECT 88.255 111.755 91.765 112.525 ;
        RECT 91.940 111.980 97.285 112.525 ;
        RECT 81.360 109.975 86.705 110.410 ;
        RECT 86.875 109.975 87.165 111.140 ;
        RECT 88.255 111.065 89.945 111.585 ;
        RECT 90.115 111.235 91.765 111.755 ;
        RECT 88.255 109.975 91.765 111.065 ;
        RECT 93.530 110.410 93.880 111.660 ;
        RECT 95.360 111.150 95.700 111.980 ;
        RECT 97.545 111.975 97.715 112.355 ;
        RECT 97.895 112.145 98.225 112.525 ;
        RECT 97.545 111.805 98.210 111.975 ;
        RECT 98.405 111.850 98.665 112.355 ;
        RECT 97.475 111.255 97.805 111.625 ;
        RECT 98.040 111.550 98.210 111.805 ;
        RECT 98.040 111.220 98.325 111.550 ;
        RECT 98.040 111.075 98.210 111.220 ;
        RECT 97.545 110.905 98.210 111.075 ;
        RECT 98.495 111.050 98.665 111.850 ;
        RECT 98.835 111.755 101.425 112.525 ;
        RECT 91.940 109.975 97.285 110.410 ;
        RECT 97.545 110.145 97.715 110.905 ;
        RECT 97.895 109.975 98.225 110.735 ;
        RECT 98.395 110.145 98.665 111.050 ;
        RECT 98.835 111.065 100.045 111.585 ;
        RECT 100.215 111.235 101.425 111.755 ;
        RECT 101.635 111.705 101.865 112.525 ;
        RECT 102.035 111.725 102.365 112.355 ;
        RECT 101.615 111.285 101.945 111.535 ;
        RECT 102.115 111.125 102.365 111.725 ;
        RECT 102.535 111.705 102.745 112.525 ;
        RECT 103.985 111.975 104.155 112.355 ;
        RECT 104.335 112.145 104.665 112.525 ;
        RECT 103.985 111.805 104.650 111.975 ;
        RECT 104.845 111.850 105.105 112.355 ;
        RECT 103.915 111.255 104.245 111.625 ;
        RECT 104.480 111.550 104.650 111.805 ;
        RECT 98.835 109.975 101.425 111.065 ;
        RECT 101.635 109.975 101.865 111.115 ;
        RECT 102.035 110.145 102.365 111.125 ;
        RECT 104.480 111.220 104.765 111.550 ;
        RECT 102.535 109.975 102.745 111.115 ;
        RECT 104.480 111.075 104.650 111.220 ;
        RECT 103.985 110.905 104.650 111.075 ;
        RECT 104.935 111.050 105.105 111.850 ;
        RECT 105.335 111.705 105.545 112.525 ;
        RECT 105.715 111.725 106.045 112.355 ;
        RECT 105.715 111.125 105.965 111.725 ;
        RECT 106.215 111.705 106.445 112.525 ;
        RECT 106.745 111.975 106.915 112.355 ;
        RECT 107.095 112.145 107.425 112.525 ;
        RECT 106.745 111.805 107.410 111.975 ;
        RECT 107.605 111.850 107.865 112.355 ;
        RECT 106.135 111.285 106.465 111.535 ;
        RECT 106.675 111.255 107.005 111.625 ;
        RECT 107.240 111.550 107.410 111.805 ;
        RECT 107.240 111.220 107.525 111.550 ;
        RECT 103.985 110.145 104.155 110.905 ;
        RECT 104.335 109.975 104.665 110.735 ;
        RECT 104.835 110.145 105.105 111.050 ;
        RECT 105.335 109.975 105.545 111.115 ;
        RECT 105.715 110.145 106.045 111.125 ;
        RECT 106.215 109.975 106.445 111.115 ;
        RECT 107.240 111.075 107.410 111.220 ;
        RECT 106.745 110.905 107.410 111.075 ;
        RECT 107.695 111.050 107.865 111.850 ;
        RECT 108.495 111.755 111.085 112.525 ;
        RECT 106.745 110.145 106.915 110.905 ;
        RECT 107.095 109.975 107.425 110.735 ;
        RECT 107.595 110.145 107.865 111.050 ;
        RECT 108.495 111.065 109.705 111.585 ;
        RECT 109.875 111.235 111.085 111.755 ;
        RECT 111.295 111.705 111.525 112.525 ;
        RECT 111.695 111.725 112.025 112.355 ;
        RECT 111.275 111.285 111.605 111.535 ;
        RECT 111.775 111.125 112.025 111.725 ;
        RECT 112.195 111.705 112.405 112.525 ;
        RECT 112.635 111.800 112.925 112.525 ;
        RECT 114.020 111.975 114.275 112.265 ;
        RECT 114.445 112.145 114.775 112.525 ;
        RECT 114.020 111.805 114.770 111.975 ;
        RECT 108.495 109.975 111.085 111.065 ;
        RECT 111.295 109.975 111.525 111.115 ;
        RECT 111.695 110.145 112.025 111.125 ;
        RECT 112.195 109.975 112.405 111.115 ;
        RECT 112.635 109.975 112.925 111.140 ;
        RECT 114.020 110.985 114.370 111.635 ;
        RECT 114.540 110.815 114.770 111.805 ;
        RECT 114.020 110.645 114.770 110.815 ;
        RECT 114.020 110.145 114.275 110.645 ;
        RECT 114.445 109.975 114.775 110.475 ;
        RECT 114.945 110.145 115.115 112.265 ;
        RECT 115.475 112.165 115.805 112.525 ;
        RECT 115.975 112.135 116.470 112.305 ;
        RECT 116.675 112.135 117.530 112.305 ;
        RECT 115.345 110.945 115.805 111.995 ;
        RECT 115.285 110.160 115.610 110.945 ;
        RECT 115.975 110.775 116.145 112.135 ;
        RECT 116.315 111.225 116.665 111.845 ;
        RECT 116.835 111.625 117.190 111.845 ;
        RECT 116.835 111.035 117.005 111.625 ;
        RECT 117.360 111.425 117.530 112.135 ;
        RECT 118.405 112.065 118.735 112.525 ;
        RECT 118.945 112.165 119.295 112.335 ;
        RECT 117.735 111.595 118.525 111.845 ;
        RECT 118.945 111.775 119.205 112.165 ;
        RECT 119.515 112.075 120.465 112.355 ;
        RECT 120.635 112.085 120.825 112.525 ;
        RECT 120.995 112.145 122.065 112.315 ;
        RECT 118.695 111.425 118.865 111.605 ;
        RECT 115.975 110.605 116.370 110.775 ;
        RECT 116.540 110.645 117.005 111.035 ;
        RECT 117.175 111.255 118.865 111.425 ;
        RECT 116.200 110.475 116.370 110.605 ;
        RECT 117.175 110.475 117.345 111.255 ;
        RECT 119.035 111.085 119.205 111.775 ;
        RECT 117.705 110.915 119.205 111.085 ;
        RECT 119.395 111.115 119.605 111.905 ;
        RECT 119.775 111.285 120.125 111.905 ;
        RECT 120.295 111.295 120.465 112.075 ;
        RECT 120.995 111.915 121.165 112.145 ;
        RECT 120.635 111.745 121.165 111.915 ;
        RECT 120.635 111.465 120.855 111.745 ;
        RECT 121.335 111.575 121.575 111.975 ;
        RECT 120.295 111.125 120.700 111.295 ;
        RECT 121.035 111.205 121.575 111.575 ;
        RECT 121.745 111.790 122.065 112.145 ;
        RECT 121.745 111.535 122.070 111.790 ;
        RECT 122.265 111.715 122.435 112.525 ;
        RECT 122.605 111.875 122.935 112.355 ;
        RECT 123.105 112.055 123.275 112.525 ;
        RECT 123.445 111.875 123.775 112.355 ;
        RECT 123.945 112.055 124.115 112.525 ;
        RECT 122.605 111.705 124.370 111.875 ;
        RECT 124.595 111.775 125.805 112.525 ;
        RECT 121.745 111.325 123.775 111.535 ;
        RECT 121.745 111.315 122.090 111.325 ;
        RECT 119.395 110.955 120.070 111.115 ;
        RECT 120.530 111.035 120.700 111.125 ;
        RECT 119.395 110.945 120.360 110.955 ;
        RECT 119.035 110.775 119.205 110.915 ;
        RECT 115.780 109.975 116.030 110.435 ;
        RECT 116.200 110.145 116.450 110.475 ;
        RECT 116.665 110.145 117.345 110.475 ;
        RECT 117.515 110.575 118.590 110.745 ;
        RECT 119.035 110.605 119.595 110.775 ;
        RECT 119.900 110.655 120.360 110.945 ;
        RECT 120.530 110.865 121.750 111.035 ;
        RECT 117.515 110.235 117.685 110.575 ;
        RECT 117.920 109.975 118.250 110.405 ;
        RECT 118.420 110.235 118.590 110.575 ;
        RECT 118.885 109.975 119.255 110.435 ;
        RECT 119.425 110.145 119.595 110.605 ;
        RECT 120.530 110.485 120.700 110.865 ;
        RECT 121.920 110.695 122.090 111.315 ;
        RECT 123.960 111.155 124.370 111.705 ;
        RECT 119.830 110.145 120.700 110.485 ;
        RECT 121.290 110.525 122.090 110.695 ;
        RECT 120.870 109.975 121.120 110.435 ;
        RECT 121.290 110.235 121.460 110.525 ;
        RECT 121.640 109.975 121.970 110.355 ;
        RECT 122.265 109.975 122.435 111.035 ;
        RECT 122.645 110.985 124.370 111.155 ;
        RECT 124.595 111.065 125.115 111.605 ;
        RECT 125.285 111.235 125.805 111.775 ;
        RECT 122.645 110.145 122.935 110.985 ;
        RECT 123.105 109.975 123.275 110.815 ;
        RECT 123.485 110.145 123.735 110.985 ;
        RECT 123.945 109.975 124.115 110.815 ;
        RECT 124.595 109.975 125.805 111.065 ;
        RECT 11.810 109.805 125.890 109.975 ;
        RECT 11.895 108.715 13.105 109.805 ;
        RECT 13.280 109.370 18.625 109.805 ;
        RECT 11.895 108.005 12.415 108.545 ;
        RECT 12.585 108.175 13.105 108.715 ;
        RECT 14.870 108.120 15.220 109.370 ;
        RECT 18.855 108.665 19.065 109.805 ;
        RECT 19.235 108.655 19.565 109.635 ;
        RECT 19.735 108.665 19.965 109.805 ;
        RECT 21.155 108.665 21.365 109.805 ;
        RECT 21.535 108.655 21.865 109.635 ;
        RECT 22.035 108.665 22.265 109.805 ;
        RECT 11.895 107.255 13.105 108.005 ;
        RECT 16.700 107.800 17.040 108.630 ;
        RECT 13.280 107.255 18.625 107.800 ;
        RECT 18.855 107.255 19.065 108.075 ;
        RECT 19.235 108.055 19.485 108.655 ;
        RECT 19.655 108.245 19.985 108.495 ;
        RECT 19.235 107.425 19.565 108.055 ;
        RECT 19.735 107.255 19.965 108.075 ;
        RECT 21.155 107.255 21.365 108.075 ;
        RECT 21.535 108.055 21.785 108.655 ;
        RECT 22.475 108.640 22.765 109.805 ;
        RECT 22.935 108.715 24.145 109.805 ;
        RECT 21.955 108.245 22.285 108.495 ;
        RECT 22.935 108.175 23.455 108.715 ;
        RECT 24.375 108.665 24.585 109.805 ;
        RECT 24.755 108.655 25.085 109.635 ;
        RECT 25.255 108.665 25.485 109.805 ;
        RECT 26.005 108.965 26.175 109.805 ;
        RECT 26.385 108.795 26.635 109.635 ;
        RECT 26.845 108.965 27.015 109.805 ;
        RECT 27.185 108.795 27.475 109.635 ;
        RECT 21.535 107.425 21.865 108.055 ;
        RECT 22.035 107.255 22.265 108.075 ;
        RECT 23.625 108.005 24.145 108.545 ;
        RECT 22.475 107.255 22.765 107.980 ;
        RECT 22.935 107.255 24.145 108.005 ;
        RECT 24.375 107.255 24.585 108.075 ;
        RECT 24.755 108.055 25.005 108.655 ;
        RECT 25.750 108.625 27.475 108.795 ;
        RECT 27.685 108.745 27.855 109.805 ;
        RECT 28.150 109.425 28.480 109.805 ;
        RECT 28.660 109.255 28.830 109.545 ;
        RECT 29.000 109.345 29.250 109.805 ;
        RECT 28.030 109.085 28.830 109.255 ;
        RECT 29.420 109.295 30.290 109.635 ;
        RECT 25.175 108.245 25.505 108.495 ;
        RECT 25.750 108.075 26.160 108.625 ;
        RECT 28.030 108.465 28.200 109.085 ;
        RECT 29.420 108.915 29.590 109.295 ;
        RECT 30.525 109.175 30.695 109.635 ;
        RECT 30.865 109.345 31.235 109.805 ;
        RECT 31.530 109.205 31.700 109.545 ;
        RECT 31.870 109.375 32.200 109.805 ;
        RECT 32.435 109.205 32.605 109.545 ;
        RECT 28.370 108.745 29.590 108.915 ;
        RECT 29.760 108.835 30.220 109.125 ;
        RECT 30.525 109.005 31.085 109.175 ;
        RECT 31.530 109.035 32.605 109.205 ;
        RECT 32.775 109.305 33.455 109.635 ;
        RECT 33.670 109.305 33.920 109.635 ;
        RECT 34.090 109.345 34.340 109.805 ;
        RECT 30.915 108.865 31.085 109.005 ;
        RECT 29.760 108.825 30.725 108.835 ;
        RECT 29.420 108.655 29.590 108.745 ;
        RECT 30.050 108.665 30.725 108.825 ;
        RECT 28.030 108.455 28.375 108.465 ;
        RECT 26.345 108.245 28.375 108.455 ;
        RECT 24.755 107.425 25.085 108.055 ;
        RECT 25.255 107.255 25.485 108.075 ;
        RECT 25.750 107.905 27.515 108.075 ;
        RECT 26.005 107.255 26.175 107.725 ;
        RECT 26.345 107.425 26.675 107.905 ;
        RECT 26.845 107.255 27.015 107.725 ;
        RECT 27.185 107.425 27.515 107.905 ;
        RECT 27.685 107.255 27.855 108.065 ;
        RECT 28.050 107.990 28.375 108.245 ;
        RECT 28.055 107.635 28.375 107.990 ;
        RECT 28.545 108.205 29.085 108.575 ;
        RECT 29.420 108.485 29.825 108.655 ;
        RECT 28.545 107.805 28.785 108.205 ;
        RECT 29.265 108.035 29.485 108.315 ;
        RECT 28.955 107.865 29.485 108.035 ;
        RECT 28.955 107.635 29.125 107.865 ;
        RECT 29.655 107.705 29.825 108.485 ;
        RECT 29.995 107.875 30.345 108.495 ;
        RECT 30.515 107.875 30.725 108.665 ;
        RECT 30.915 108.695 32.415 108.865 ;
        RECT 30.915 108.005 31.085 108.695 ;
        RECT 32.775 108.525 32.945 109.305 ;
        RECT 33.750 109.175 33.920 109.305 ;
        RECT 31.255 108.355 32.945 108.525 ;
        RECT 33.115 108.745 33.580 109.135 ;
        RECT 33.750 109.005 34.145 109.175 ;
        RECT 31.255 108.175 31.425 108.355 ;
        RECT 28.055 107.465 29.125 107.635 ;
        RECT 29.295 107.255 29.485 107.695 ;
        RECT 29.655 107.425 30.605 107.705 ;
        RECT 30.915 107.615 31.175 108.005 ;
        RECT 31.595 107.935 32.385 108.185 ;
        RECT 30.825 107.445 31.175 107.615 ;
        RECT 31.385 107.255 31.715 107.715 ;
        RECT 32.590 107.645 32.760 108.355 ;
        RECT 33.115 108.155 33.285 108.745 ;
        RECT 32.930 107.935 33.285 108.155 ;
        RECT 33.455 107.935 33.805 108.555 ;
        RECT 33.975 107.645 34.145 109.005 ;
        RECT 34.510 108.835 34.835 109.620 ;
        RECT 34.315 107.785 34.775 108.835 ;
        RECT 32.590 107.475 33.445 107.645 ;
        RECT 33.650 107.475 34.145 107.645 ;
        RECT 34.315 107.255 34.645 107.615 ;
        RECT 35.005 107.515 35.175 109.635 ;
        RECT 35.345 109.305 35.675 109.805 ;
        RECT 35.845 109.135 36.100 109.635 ;
        RECT 35.350 108.965 36.100 109.135 ;
        RECT 36.585 108.965 36.755 109.805 ;
        RECT 35.350 107.975 35.580 108.965 ;
        RECT 36.965 108.795 37.215 109.635 ;
        RECT 37.425 108.965 37.595 109.805 ;
        RECT 37.765 108.795 38.055 109.635 ;
        RECT 35.750 108.145 36.100 108.795 ;
        RECT 36.330 108.625 38.055 108.795 ;
        RECT 38.265 108.745 38.435 109.805 ;
        RECT 38.730 109.425 39.060 109.805 ;
        RECT 39.240 109.255 39.410 109.545 ;
        RECT 39.580 109.345 39.830 109.805 ;
        RECT 38.610 109.085 39.410 109.255 ;
        RECT 40.000 109.295 40.870 109.635 ;
        RECT 36.330 108.075 36.740 108.625 ;
        RECT 38.610 108.465 38.780 109.085 ;
        RECT 40.000 108.915 40.170 109.295 ;
        RECT 41.105 109.175 41.275 109.635 ;
        RECT 41.445 109.345 41.815 109.805 ;
        RECT 42.110 109.205 42.280 109.545 ;
        RECT 42.450 109.375 42.780 109.805 ;
        RECT 43.015 109.205 43.185 109.545 ;
        RECT 38.950 108.745 40.170 108.915 ;
        RECT 40.340 108.835 40.800 109.125 ;
        RECT 41.105 109.005 41.665 109.175 ;
        RECT 42.110 109.035 43.185 109.205 ;
        RECT 43.355 109.305 44.035 109.635 ;
        RECT 44.250 109.305 44.500 109.635 ;
        RECT 44.670 109.345 44.920 109.805 ;
        RECT 41.495 108.865 41.665 109.005 ;
        RECT 40.340 108.825 41.305 108.835 ;
        RECT 40.000 108.655 40.170 108.745 ;
        RECT 40.630 108.665 41.305 108.825 ;
        RECT 38.610 108.455 38.955 108.465 ;
        RECT 36.925 108.245 38.955 108.455 ;
        RECT 35.350 107.805 36.100 107.975 ;
        RECT 36.330 107.905 38.095 108.075 ;
        RECT 35.345 107.255 35.675 107.635 ;
        RECT 35.845 107.515 36.100 107.805 ;
        RECT 36.585 107.255 36.755 107.725 ;
        RECT 36.925 107.425 37.255 107.905 ;
        RECT 37.425 107.255 37.595 107.725 ;
        RECT 37.765 107.425 38.095 107.905 ;
        RECT 38.265 107.255 38.435 108.065 ;
        RECT 38.630 107.990 38.955 108.245 ;
        RECT 38.635 107.635 38.955 107.990 ;
        RECT 39.125 108.205 39.665 108.575 ;
        RECT 40.000 108.485 40.405 108.655 ;
        RECT 39.125 107.805 39.365 108.205 ;
        RECT 39.845 108.035 40.065 108.315 ;
        RECT 39.535 107.865 40.065 108.035 ;
        RECT 39.535 107.635 39.705 107.865 ;
        RECT 40.235 107.705 40.405 108.485 ;
        RECT 40.575 107.875 40.925 108.495 ;
        RECT 41.095 107.875 41.305 108.665 ;
        RECT 41.495 108.695 42.995 108.865 ;
        RECT 41.495 108.005 41.665 108.695 ;
        RECT 43.355 108.525 43.525 109.305 ;
        RECT 44.330 109.175 44.500 109.305 ;
        RECT 41.835 108.355 43.525 108.525 ;
        RECT 43.695 108.745 44.160 109.135 ;
        RECT 44.330 109.005 44.725 109.175 ;
        RECT 41.835 108.175 42.005 108.355 ;
        RECT 38.635 107.465 39.705 107.635 ;
        RECT 39.875 107.255 40.065 107.695 ;
        RECT 40.235 107.425 41.185 107.705 ;
        RECT 41.495 107.615 41.755 108.005 ;
        RECT 42.175 107.935 42.965 108.185 ;
        RECT 41.405 107.445 41.755 107.615 ;
        RECT 41.965 107.255 42.295 107.715 ;
        RECT 43.170 107.645 43.340 108.355 ;
        RECT 43.695 108.155 43.865 108.745 ;
        RECT 43.510 107.935 43.865 108.155 ;
        RECT 44.035 107.935 44.385 108.555 ;
        RECT 44.555 107.645 44.725 109.005 ;
        RECT 45.090 108.835 45.415 109.620 ;
        RECT 44.895 107.785 45.355 108.835 ;
        RECT 43.170 107.475 44.025 107.645 ;
        RECT 44.230 107.475 44.725 107.645 ;
        RECT 44.895 107.255 45.225 107.615 ;
        RECT 45.585 107.515 45.755 109.635 ;
        RECT 45.925 109.305 46.255 109.805 ;
        RECT 46.425 109.135 46.680 109.635 ;
        RECT 45.930 108.965 46.680 109.135 ;
        RECT 45.930 107.975 46.160 108.965 ;
        RECT 46.945 108.875 47.115 109.635 ;
        RECT 47.295 109.045 47.625 109.805 ;
        RECT 46.330 108.145 46.680 108.795 ;
        RECT 46.945 108.705 47.610 108.875 ;
        RECT 47.795 108.730 48.065 109.635 ;
        RECT 47.440 108.560 47.610 108.705 ;
        RECT 46.875 108.155 47.205 108.525 ;
        RECT 47.440 108.230 47.725 108.560 ;
        RECT 47.440 107.975 47.610 108.230 ;
        RECT 45.930 107.805 46.680 107.975 ;
        RECT 45.925 107.255 46.255 107.635 ;
        RECT 46.425 107.515 46.680 107.805 ;
        RECT 46.945 107.805 47.610 107.975 ;
        RECT 47.895 107.930 48.065 108.730 ;
        RECT 48.235 108.640 48.525 109.805 ;
        RECT 48.695 108.715 50.365 109.805 ;
        RECT 50.625 108.875 50.795 109.635 ;
        RECT 50.975 109.045 51.305 109.805 ;
        RECT 48.695 108.195 49.445 108.715 ;
        RECT 50.625 108.705 51.290 108.875 ;
        RECT 51.475 108.730 51.745 109.635 ;
        RECT 51.120 108.560 51.290 108.705 ;
        RECT 49.615 108.025 50.365 108.545 ;
        RECT 50.555 108.155 50.885 108.525 ;
        RECT 51.120 108.230 51.405 108.560 ;
        RECT 46.945 107.425 47.115 107.805 ;
        RECT 47.295 107.255 47.625 107.635 ;
        RECT 47.805 107.425 48.065 107.930 ;
        RECT 48.235 107.255 48.525 107.980 ;
        RECT 48.695 107.255 50.365 108.025 ;
        RECT 51.120 107.975 51.290 108.230 ;
        RECT 50.625 107.805 51.290 107.975 ;
        RECT 51.575 107.930 51.745 108.730 ;
        RECT 52.375 108.715 54.965 109.805 ;
        RECT 52.375 108.195 53.585 108.715 ;
        RECT 55.175 108.665 55.405 109.805 ;
        RECT 55.575 108.655 55.905 109.635 ;
        RECT 56.075 108.665 56.285 109.805 ;
        RECT 56.825 108.965 56.995 109.805 ;
        RECT 57.205 108.795 57.455 109.635 ;
        RECT 57.665 108.965 57.835 109.805 ;
        RECT 58.005 108.795 58.295 109.635 ;
        RECT 53.755 108.025 54.965 108.545 ;
        RECT 55.155 108.245 55.485 108.495 ;
        RECT 50.625 107.425 50.795 107.805 ;
        RECT 50.975 107.255 51.305 107.635 ;
        RECT 51.485 107.425 51.745 107.930 ;
        RECT 52.375 107.255 54.965 108.025 ;
        RECT 55.175 107.255 55.405 108.075 ;
        RECT 55.655 108.055 55.905 108.655 ;
        RECT 56.570 108.625 58.295 108.795 ;
        RECT 58.505 108.745 58.675 109.805 ;
        RECT 58.970 109.425 59.300 109.805 ;
        RECT 59.480 109.255 59.650 109.545 ;
        RECT 59.820 109.345 60.070 109.805 ;
        RECT 58.850 109.085 59.650 109.255 ;
        RECT 60.240 109.295 61.110 109.635 ;
        RECT 56.570 108.075 56.980 108.625 ;
        RECT 58.850 108.465 59.020 109.085 ;
        RECT 60.240 108.915 60.410 109.295 ;
        RECT 61.345 109.175 61.515 109.635 ;
        RECT 61.685 109.345 62.055 109.805 ;
        RECT 62.350 109.205 62.520 109.545 ;
        RECT 62.690 109.375 63.020 109.805 ;
        RECT 63.255 109.205 63.425 109.545 ;
        RECT 59.190 108.745 60.410 108.915 ;
        RECT 60.580 108.835 61.040 109.125 ;
        RECT 61.345 109.005 61.905 109.175 ;
        RECT 62.350 109.035 63.425 109.205 ;
        RECT 63.595 109.305 64.275 109.635 ;
        RECT 64.490 109.305 64.740 109.635 ;
        RECT 64.910 109.345 65.160 109.805 ;
        RECT 61.735 108.865 61.905 109.005 ;
        RECT 60.580 108.825 61.545 108.835 ;
        RECT 60.240 108.655 60.410 108.745 ;
        RECT 60.870 108.665 61.545 108.825 ;
        RECT 58.850 108.455 59.195 108.465 ;
        RECT 57.165 108.245 59.195 108.455 ;
        RECT 55.575 107.425 55.905 108.055 ;
        RECT 56.075 107.255 56.285 108.075 ;
        RECT 56.570 107.905 58.335 108.075 ;
        RECT 56.825 107.255 56.995 107.725 ;
        RECT 57.165 107.425 57.495 107.905 ;
        RECT 57.665 107.255 57.835 107.725 ;
        RECT 58.005 107.425 58.335 107.905 ;
        RECT 58.505 107.255 58.675 108.065 ;
        RECT 58.870 107.990 59.195 108.245 ;
        RECT 58.875 107.635 59.195 107.990 ;
        RECT 59.365 108.205 59.905 108.575 ;
        RECT 60.240 108.485 60.645 108.655 ;
        RECT 59.365 107.805 59.605 108.205 ;
        RECT 60.085 108.035 60.305 108.315 ;
        RECT 59.775 107.865 60.305 108.035 ;
        RECT 59.775 107.635 59.945 107.865 ;
        RECT 60.475 107.705 60.645 108.485 ;
        RECT 60.815 107.875 61.165 108.495 ;
        RECT 61.335 107.875 61.545 108.665 ;
        RECT 61.735 108.695 63.235 108.865 ;
        RECT 61.735 108.005 61.905 108.695 ;
        RECT 63.595 108.525 63.765 109.305 ;
        RECT 64.570 109.175 64.740 109.305 ;
        RECT 62.075 108.355 63.765 108.525 ;
        RECT 63.935 108.745 64.400 109.135 ;
        RECT 64.570 109.005 64.965 109.175 ;
        RECT 62.075 108.175 62.245 108.355 ;
        RECT 58.875 107.465 59.945 107.635 ;
        RECT 60.115 107.255 60.305 107.695 ;
        RECT 60.475 107.425 61.425 107.705 ;
        RECT 61.735 107.615 61.995 108.005 ;
        RECT 62.415 107.935 63.205 108.185 ;
        RECT 61.645 107.445 61.995 107.615 ;
        RECT 62.205 107.255 62.535 107.715 ;
        RECT 63.410 107.645 63.580 108.355 ;
        RECT 63.935 108.155 64.105 108.745 ;
        RECT 63.750 107.935 64.105 108.155 ;
        RECT 64.275 107.935 64.625 108.555 ;
        RECT 64.795 107.645 64.965 109.005 ;
        RECT 65.330 108.835 65.655 109.620 ;
        RECT 65.135 107.785 65.595 108.835 ;
        RECT 63.410 107.475 64.265 107.645 ;
        RECT 64.470 107.475 64.965 107.645 ;
        RECT 65.135 107.255 65.465 107.615 ;
        RECT 65.825 107.515 65.995 109.635 ;
        RECT 66.165 109.305 66.495 109.805 ;
        RECT 66.665 109.135 66.920 109.635 ;
        RECT 66.170 108.965 66.920 109.135 ;
        RECT 66.170 107.975 66.400 108.965 ;
        RECT 67.185 108.875 67.355 109.635 ;
        RECT 67.535 109.045 67.865 109.805 ;
        RECT 66.570 108.145 66.920 108.795 ;
        RECT 67.185 108.705 67.850 108.875 ;
        RECT 68.035 108.730 68.305 109.635 ;
        RECT 67.680 108.560 67.850 108.705 ;
        RECT 67.115 108.155 67.445 108.525 ;
        RECT 67.680 108.230 67.965 108.560 ;
        RECT 67.680 107.975 67.850 108.230 ;
        RECT 66.170 107.805 66.920 107.975 ;
        RECT 66.165 107.255 66.495 107.635 ;
        RECT 66.665 107.515 66.920 107.805 ;
        RECT 67.185 107.805 67.850 107.975 ;
        RECT 68.135 107.930 68.305 108.730 ;
        RECT 68.935 108.715 72.445 109.805 ;
        RECT 72.705 108.875 72.875 109.635 ;
        RECT 73.055 109.045 73.385 109.805 ;
        RECT 68.935 108.195 70.625 108.715 ;
        RECT 72.705 108.705 73.370 108.875 ;
        RECT 73.555 108.730 73.825 109.635 ;
        RECT 73.200 108.560 73.370 108.705 ;
        RECT 70.795 108.025 72.445 108.545 ;
        RECT 72.635 108.155 72.965 108.525 ;
        RECT 73.200 108.230 73.485 108.560 ;
        RECT 67.185 107.425 67.355 107.805 ;
        RECT 67.535 107.255 67.865 107.635 ;
        RECT 68.045 107.425 68.305 107.930 ;
        RECT 68.935 107.255 72.445 108.025 ;
        RECT 73.200 107.975 73.370 108.230 ;
        RECT 72.705 107.805 73.370 107.975 ;
        RECT 73.655 107.930 73.825 108.730 ;
        RECT 73.995 108.640 74.285 109.805 ;
        RECT 74.765 108.965 74.935 109.805 ;
        RECT 75.145 108.795 75.395 109.635 ;
        RECT 75.605 108.965 75.775 109.805 ;
        RECT 75.945 108.795 76.235 109.635 ;
        RECT 74.510 108.625 76.235 108.795 ;
        RECT 76.445 108.745 76.615 109.805 ;
        RECT 76.910 109.425 77.240 109.805 ;
        RECT 77.420 109.255 77.590 109.545 ;
        RECT 77.760 109.345 78.010 109.805 ;
        RECT 76.790 109.085 77.590 109.255 ;
        RECT 78.180 109.295 79.050 109.635 ;
        RECT 74.510 108.075 74.920 108.625 ;
        RECT 76.790 108.465 76.960 109.085 ;
        RECT 78.180 108.915 78.350 109.295 ;
        RECT 79.285 109.175 79.455 109.635 ;
        RECT 79.625 109.345 79.995 109.805 ;
        RECT 80.290 109.205 80.460 109.545 ;
        RECT 80.630 109.375 80.960 109.805 ;
        RECT 81.195 109.205 81.365 109.545 ;
        RECT 77.130 108.745 78.350 108.915 ;
        RECT 78.520 108.835 78.980 109.125 ;
        RECT 79.285 109.005 79.845 109.175 ;
        RECT 80.290 109.035 81.365 109.205 ;
        RECT 81.535 109.305 82.215 109.635 ;
        RECT 82.430 109.305 82.680 109.635 ;
        RECT 82.850 109.345 83.100 109.805 ;
        RECT 79.675 108.865 79.845 109.005 ;
        RECT 78.520 108.825 79.485 108.835 ;
        RECT 78.180 108.655 78.350 108.745 ;
        RECT 78.810 108.665 79.485 108.825 ;
        RECT 76.790 108.455 77.135 108.465 ;
        RECT 75.105 108.245 77.135 108.455 ;
        RECT 72.705 107.425 72.875 107.805 ;
        RECT 73.055 107.255 73.385 107.635 ;
        RECT 73.565 107.425 73.825 107.930 ;
        RECT 73.995 107.255 74.285 107.980 ;
        RECT 74.510 107.905 76.275 108.075 ;
        RECT 74.765 107.255 74.935 107.725 ;
        RECT 75.105 107.425 75.435 107.905 ;
        RECT 75.605 107.255 75.775 107.725 ;
        RECT 75.945 107.425 76.275 107.905 ;
        RECT 76.445 107.255 76.615 108.065 ;
        RECT 76.810 107.990 77.135 108.245 ;
        RECT 76.815 107.635 77.135 107.990 ;
        RECT 77.305 108.205 77.845 108.575 ;
        RECT 78.180 108.485 78.585 108.655 ;
        RECT 77.305 107.805 77.545 108.205 ;
        RECT 78.025 108.035 78.245 108.315 ;
        RECT 77.715 107.865 78.245 108.035 ;
        RECT 77.715 107.635 77.885 107.865 ;
        RECT 78.415 107.705 78.585 108.485 ;
        RECT 78.755 107.875 79.105 108.495 ;
        RECT 79.275 107.875 79.485 108.665 ;
        RECT 79.675 108.695 81.175 108.865 ;
        RECT 79.675 108.005 79.845 108.695 ;
        RECT 81.535 108.525 81.705 109.305 ;
        RECT 82.510 109.175 82.680 109.305 ;
        RECT 80.015 108.355 81.705 108.525 ;
        RECT 81.875 108.745 82.340 109.135 ;
        RECT 82.510 109.005 82.905 109.175 ;
        RECT 80.015 108.175 80.185 108.355 ;
        RECT 76.815 107.465 77.885 107.635 ;
        RECT 78.055 107.255 78.245 107.695 ;
        RECT 78.415 107.425 79.365 107.705 ;
        RECT 79.675 107.615 79.935 108.005 ;
        RECT 80.355 107.935 81.145 108.185 ;
        RECT 79.585 107.445 79.935 107.615 ;
        RECT 80.145 107.255 80.475 107.715 ;
        RECT 81.350 107.645 81.520 108.355 ;
        RECT 81.875 108.155 82.045 108.745 ;
        RECT 81.690 107.935 82.045 108.155 ;
        RECT 82.215 107.935 82.565 108.555 ;
        RECT 82.735 107.645 82.905 109.005 ;
        RECT 83.270 108.835 83.595 109.620 ;
        RECT 83.075 107.785 83.535 108.835 ;
        RECT 81.350 107.475 82.205 107.645 ;
        RECT 82.410 107.475 82.905 107.645 ;
        RECT 83.075 107.255 83.405 107.615 ;
        RECT 83.765 107.515 83.935 109.635 ;
        RECT 84.105 109.305 84.435 109.805 ;
        RECT 84.605 109.135 84.860 109.635 ;
        RECT 84.110 108.965 84.860 109.135 ;
        RECT 84.110 107.975 84.340 108.965 ;
        RECT 84.510 108.145 84.860 108.795 ;
        RECT 85.035 108.730 85.305 109.635 ;
        RECT 85.475 109.045 85.805 109.805 ;
        RECT 85.985 108.875 86.155 109.635 ;
        RECT 84.110 107.805 84.860 107.975 ;
        RECT 84.105 107.255 84.435 107.635 ;
        RECT 84.605 107.515 84.860 107.805 ;
        RECT 85.035 107.930 85.205 108.730 ;
        RECT 85.490 108.705 86.155 108.875 ;
        RECT 86.415 108.715 87.625 109.805 ;
        RECT 87.885 108.875 88.055 109.635 ;
        RECT 88.235 109.045 88.565 109.805 ;
        RECT 85.490 108.560 85.660 108.705 ;
        RECT 85.375 108.230 85.660 108.560 ;
        RECT 85.490 107.975 85.660 108.230 ;
        RECT 85.895 108.155 86.225 108.525 ;
        RECT 86.415 108.175 86.935 108.715 ;
        RECT 87.885 108.705 88.550 108.875 ;
        RECT 88.735 108.730 89.005 109.635 ;
        RECT 89.485 108.965 89.655 109.805 ;
        RECT 89.865 108.795 90.115 109.635 ;
        RECT 90.325 108.965 90.495 109.805 ;
        RECT 90.665 108.795 90.955 109.635 ;
        RECT 88.380 108.560 88.550 108.705 ;
        RECT 87.105 108.005 87.625 108.545 ;
        RECT 87.815 108.155 88.145 108.525 ;
        RECT 88.380 108.230 88.665 108.560 ;
        RECT 85.035 107.425 85.295 107.930 ;
        RECT 85.490 107.805 86.155 107.975 ;
        RECT 85.475 107.255 85.805 107.635 ;
        RECT 85.985 107.425 86.155 107.805 ;
        RECT 86.415 107.255 87.625 108.005 ;
        RECT 88.380 107.975 88.550 108.230 ;
        RECT 87.885 107.805 88.550 107.975 ;
        RECT 88.835 107.930 89.005 108.730 ;
        RECT 87.885 107.425 88.055 107.805 ;
        RECT 88.235 107.255 88.565 107.635 ;
        RECT 88.745 107.425 89.005 107.930 ;
        RECT 89.230 108.625 90.955 108.795 ;
        RECT 91.165 108.745 91.335 109.805 ;
        RECT 91.630 109.425 91.960 109.805 ;
        RECT 92.140 109.255 92.310 109.545 ;
        RECT 92.480 109.345 92.730 109.805 ;
        RECT 91.510 109.085 92.310 109.255 ;
        RECT 92.900 109.295 93.770 109.635 ;
        RECT 89.230 108.075 89.640 108.625 ;
        RECT 91.510 108.465 91.680 109.085 ;
        RECT 92.900 108.915 93.070 109.295 ;
        RECT 94.005 109.175 94.175 109.635 ;
        RECT 94.345 109.345 94.715 109.805 ;
        RECT 95.010 109.205 95.180 109.545 ;
        RECT 95.350 109.375 95.680 109.805 ;
        RECT 95.915 109.205 96.085 109.545 ;
        RECT 91.850 108.745 93.070 108.915 ;
        RECT 93.240 108.835 93.700 109.125 ;
        RECT 94.005 109.005 94.565 109.175 ;
        RECT 95.010 109.035 96.085 109.205 ;
        RECT 96.255 109.305 96.935 109.635 ;
        RECT 97.150 109.305 97.400 109.635 ;
        RECT 97.570 109.345 97.820 109.805 ;
        RECT 94.395 108.865 94.565 109.005 ;
        RECT 93.240 108.825 94.205 108.835 ;
        RECT 92.900 108.655 93.070 108.745 ;
        RECT 93.530 108.665 94.205 108.825 ;
        RECT 91.510 108.455 91.855 108.465 ;
        RECT 89.825 108.245 91.855 108.455 ;
        RECT 89.230 107.905 90.995 108.075 ;
        RECT 89.485 107.255 89.655 107.725 ;
        RECT 89.825 107.425 90.155 107.905 ;
        RECT 90.325 107.255 90.495 107.725 ;
        RECT 90.665 107.425 90.995 107.905 ;
        RECT 91.165 107.255 91.335 108.065 ;
        RECT 91.530 107.990 91.855 108.245 ;
        RECT 91.535 107.635 91.855 107.990 ;
        RECT 92.025 108.205 92.565 108.575 ;
        RECT 92.900 108.485 93.305 108.655 ;
        RECT 92.025 107.805 92.265 108.205 ;
        RECT 92.745 108.035 92.965 108.315 ;
        RECT 92.435 107.865 92.965 108.035 ;
        RECT 92.435 107.635 92.605 107.865 ;
        RECT 93.135 107.705 93.305 108.485 ;
        RECT 93.475 107.875 93.825 108.495 ;
        RECT 93.995 107.875 94.205 108.665 ;
        RECT 94.395 108.695 95.895 108.865 ;
        RECT 94.395 108.005 94.565 108.695 ;
        RECT 96.255 108.525 96.425 109.305 ;
        RECT 97.230 109.175 97.400 109.305 ;
        RECT 94.735 108.355 96.425 108.525 ;
        RECT 96.595 108.745 97.060 109.135 ;
        RECT 97.230 109.005 97.625 109.175 ;
        RECT 94.735 108.175 94.905 108.355 ;
        RECT 91.535 107.465 92.605 107.635 ;
        RECT 92.775 107.255 92.965 107.695 ;
        RECT 93.135 107.425 94.085 107.705 ;
        RECT 94.395 107.615 94.655 108.005 ;
        RECT 95.075 107.935 95.865 108.185 ;
        RECT 94.305 107.445 94.655 107.615 ;
        RECT 94.865 107.255 95.195 107.715 ;
        RECT 96.070 107.645 96.240 108.355 ;
        RECT 96.595 108.155 96.765 108.745 ;
        RECT 96.410 107.935 96.765 108.155 ;
        RECT 96.935 107.935 97.285 108.555 ;
        RECT 97.455 107.645 97.625 109.005 ;
        RECT 97.990 108.835 98.315 109.620 ;
        RECT 97.795 107.785 98.255 108.835 ;
        RECT 96.070 107.475 96.925 107.645 ;
        RECT 97.130 107.475 97.625 107.645 ;
        RECT 97.795 107.255 98.125 107.615 ;
        RECT 98.485 107.515 98.655 109.635 ;
        RECT 98.825 109.305 99.155 109.805 ;
        RECT 99.325 109.135 99.580 109.635 ;
        RECT 98.830 108.965 99.580 109.135 ;
        RECT 98.830 107.975 99.060 108.965 ;
        RECT 99.230 108.145 99.580 108.795 ;
        RECT 99.755 108.640 100.045 109.805 ;
        RECT 100.985 108.965 101.155 109.805 ;
        RECT 101.365 108.795 101.615 109.635 ;
        RECT 101.825 108.965 101.995 109.805 ;
        RECT 102.165 108.795 102.455 109.635 ;
        RECT 100.730 108.625 102.455 108.795 ;
        RECT 102.665 108.745 102.835 109.805 ;
        RECT 103.130 109.425 103.460 109.805 ;
        RECT 103.640 109.255 103.810 109.545 ;
        RECT 103.980 109.345 104.230 109.805 ;
        RECT 103.010 109.085 103.810 109.255 ;
        RECT 104.400 109.295 105.270 109.635 ;
        RECT 100.730 108.075 101.140 108.625 ;
        RECT 103.010 108.465 103.180 109.085 ;
        RECT 104.400 108.915 104.570 109.295 ;
        RECT 105.505 109.175 105.675 109.635 ;
        RECT 105.845 109.345 106.215 109.805 ;
        RECT 106.510 109.205 106.680 109.545 ;
        RECT 106.850 109.375 107.180 109.805 ;
        RECT 107.415 109.205 107.585 109.545 ;
        RECT 103.350 108.745 104.570 108.915 ;
        RECT 104.740 108.835 105.200 109.125 ;
        RECT 105.505 109.005 106.065 109.175 ;
        RECT 106.510 109.035 107.585 109.205 ;
        RECT 107.755 109.305 108.435 109.635 ;
        RECT 108.650 109.305 108.900 109.635 ;
        RECT 109.070 109.345 109.320 109.805 ;
        RECT 105.895 108.865 106.065 109.005 ;
        RECT 104.740 108.825 105.705 108.835 ;
        RECT 104.400 108.655 104.570 108.745 ;
        RECT 105.030 108.665 105.705 108.825 ;
        RECT 103.010 108.455 103.355 108.465 ;
        RECT 101.325 108.245 103.355 108.455 ;
        RECT 98.830 107.805 99.580 107.975 ;
        RECT 98.825 107.255 99.155 107.635 ;
        RECT 99.325 107.515 99.580 107.805 ;
        RECT 99.755 107.255 100.045 107.980 ;
        RECT 100.730 107.905 102.495 108.075 ;
        RECT 100.985 107.255 101.155 107.725 ;
        RECT 101.325 107.425 101.655 107.905 ;
        RECT 101.825 107.255 101.995 107.725 ;
        RECT 102.165 107.425 102.495 107.905 ;
        RECT 102.665 107.255 102.835 108.065 ;
        RECT 103.030 107.990 103.355 108.245 ;
        RECT 103.035 107.635 103.355 107.990 ;
        RECT 103.525 108.205 104.065 108.575 ;
        RECT 104.400 108.485 104.805 108.655 ;
        RECT 103.525 107.805 103.765 108.205 ;
        RECT 104.245 108.035 104.465 108.315 ;
        RECT 103.935 107.865 104.465 108.035 ;
        RECT 103.935 107.635 104.105 107.865 ;
        RECT 104.635 107.705 104.805 108.485 ;
        RECT 104.975 107.875 105.325 108.495 ;
        RECT 105.495 107.875 105.705 108.665 ;
        RECT 105.895 108.695 107.395 108.865 ;
        RECT 105.895 108.005 106.065 108.695 ;
        RECT 107.755 108.525 107.925 109.305 ;
        RECT 108.730 109.175 108.900 109.305 ;
        RECT 106.235 108.355 107.925 108.525 ;
        RECT 108.095 108.745 108.560 109.135 ;
        RECT 108.730 109.005 109.125 109.175 ;
        RECT 106.235 108.175 106.405 108.355 ;
        RECT 103.035 107.465 104.105 107.635 ;
        RECT 104.275 107.255 104.465 107.695 ;
        RECT 104.635 107.425 105.585 107.705 ;
        RECT 105.895 107.615 106.155 108.005 ;
        RECT 106.575 107.935 107.365 108.185 ;
        RECT 105.805 107.445 106.155 107.615 ;
        RECT 106.365 107.255 106.695 107.715 ;
        RECT 107.570 107.645 107.740 108.355 ;
        RECT 108.095 108.155 108.265 108.745 ;
        RECT 107.910 107.935 108.265 108.155 ;
        RECT 108.435 107.935 108.785 108.555 ;
        RECT 108.955 107.645 109.125 109.005 ;
        RECT 109.490 108.835 109.815 109.620 ;
        RECT 109.295 107.785 109.755 108.835 ;
        RECT 107.570 107.475 108.425 107.645 ;
        RECT 108.630 107.475 109.125 107.645 ;
        RECT 109.295 107.255 109.625 107.615 ;
        RECT 109.985 107.515 110.155 109.635 ;
        RECT 110.325 109.305 110.655 109.805 ;
        RECT 110.825 109.135 111.080 109.635 ;
        RECT 110.330 108.965 111.080 109.135 ;
        RECT 110.330 107.975 110.560 108.965 ;
        RECT 111.345 108.875 111.515 109.635 ;
        RECT 111.695 109.045 112.025 109.805 ;
        RECT 110.730 108.145 111.080 108.795 ;
        RECT 111.345 108.705 112.010 108.875 ;
        RECT 112.195 108.730 112.465 109.635 ;
        RECT 113.865 108.965 114.035 109.805 ;
        RECT 114.245 108.795 114.495 109.635 ;
        RECT 114.705 108.965 114.875 109.805 ;
        RECT 115.045 108.795 115.335 109.635 ;
        RECT 111.840 108.560 112.010 108.705 ;
        RECT 111.275 108.155 111.605 108.525 ;
        RECT 111.840 108.230 112.125 108.560 ;
        RECT 111.840 107.975 112.010 108.230 ;
        RECT 110.330 107.805 111.080 107.975 ;
        RECT 110.325 107.255 110.655 107.635 ;
        RECT 110.825 107.515 111.080 107.805 ;
        RECT 111.345 107.805 112.010 107.975 ;
        RECT 112.295 107.930 112.465 108.730 ;
        RECT 111.345 107.425 111.515 107.805 ;
        RECT 111.695 107.255 112.025 107.635 ;
        RECT 112.205 107.425 112.465 107.930 ;
        RECT 113.610 108.625 115.335 108.795 ;
        RECT 115.545 108.745 115.715 109.805 ;
        RECT 116.010 109.425 116.340 109.805 ;
        RECT 116.520 109.255 116.690 109.545 ;
        RECT 116.860 109.345 117.110 109.805 ;
        RECT 115.890 109.085 116.690 109.255 ;
        RECT 117.280 109.295 118.150 109.635 ;
        RECT 113.610 108.075 114.020 108.625 ;
        RECT 115.890 108.465 116.060 109.085 ;
        RECT 117.280 108.915 117.450 109.295 ;
        RECT 118.385 109.175 118.555 109.635 ;
        RECT 118.725 109.345 119.095 109.805 ;
        RECT 119.390 109.205 119.560 109.545 ;
        RECT 119.730 109.375 120.060 109.805 ;
        RECT 120.295 109.205 120.465 109.545 ;
        RECT 116.230 108.745 117.450 108.915 ;
        RECT 117.620 108.835 118.080 109.125 ;
        RECT 118.385 109.005 118.945 109.175 ;
        RECT 119.390 109.035 120.465 109.205 ;
        RECT 120.635 109.305 121.315 109.635 ;
        RECT 121.530 109.305 121.780 109.635 ;
        RECT 121.950 109.345 122.200 109.805 ;
        RECT 118.775 108.865 118.945 109.005 ;
        RECT 117.620 108.825 118.585 108.835 ;
        RECT 117.280 108.655 117.450 108.745 ;
        RECT 117.910 108.665 118.585 108.825 ;
        RECT 115.890 108.455 116.235 108.465 ;
        RECT 114.205 108.245 116.235 108.455 ;
        RECT 113.610 107.905 115.375 108.075 ;
        RECT 113.865 107.255 114.035 107.725 ;
        RECT 114.205 107.425 114.535 107.905 ;
        RECT 114.705 107.255 114.875 107.725 ;
        RECT 115.045 107.425 115.375 107.905 ;
        RECT 115.545 107.255 115.715 108.065 ;
        RECT 115.910 107.990 116.235 108.245 ;
        RECT 115.915 107.635 116.235 107.990 ;
        RECT 116.405 108.205 116.945 108.575 ;
        RECT 117.280 108.485 117.685 108.655 ;
        RECT 116.405 107.805 116.645 108.205 ;
        RECT 117.125 108.035 117.345 108.315 ;
        RECT 116.815 107.865 117.345 108.035 ;
        RECT 116.815 107.635 116.985 107.865 ;
        RECT 117.515 107.705 117.685 108.485 ;
        RECT 117.855 107.875 118.205 108.495 ;
        RECT 118.375 107.875 118.585 108.665 ;
        RECT 118.775 108.695 120.275 108.865 ;
        RECT 118.775 108.005 118.945 108.695 ;
        RECT 120.635 108.525 120.805 109.305 ;
        RECT 121.610 109.175 121.780 109.305 ;
        RECT 119.115 108.355 120.805 108.525 ;
        RECT 120.975 108.745 121.440 109.135 ;
        RECT 121.610 109.005 122.005 109.175 ;
        RECT 119.115 108.175 119.285 108.355 ;
        RECT 115.915 107.465 116.985 107.635 ;
        RECT 117.155 107.255 117.345 107.695 ;
        RECT 117.515 107.425 118.465 107.705 ;
        RECT 118.775 107.615 119.035 108.005 ;
        RECT 119.455 107.935 120.245 108.185 ;
        RECT 118.685 107.445 119.035 107.615 ;
        RECT 119.245 107.255 119.575 107.715 ;
        RECT 120.450 107.645 120.620 108.355 ;
        RECT 120.975 108.155 121.145 108.745 ;
        RECT 120.790 107.935 121.145 108.155 ;
        RECT 121.315 107.935 121.665 108.555 ;
        RECT 121.835 107.645 122.005 109.005 ;
        RECT 122.370 108.835 122.695 109.620 ;
        RECT 122.175 107.785 122.635 108.835 ;
        RECT 120.450 107.475 121.305 107.645 ;
        RECT 121.510 107.475 122.005 107.645 ;
        RECT 122.175 107.255 122.505 107.615 ;
        RECT 122.865 107.515 123.035 109.635 ;
        RECT 123.205 109.305 123.535 109.805 ;
        RECT 123.705 109.135 123.960 109.635 ;
        RECT 123.210 108.965 123.960 109.135 ;
        RECT 123.210 107.975 123.440 108.965 ;
        RECT 123.610 108.145 123.960 108.795 ;
        RECT 124.595 108.715 125.805 109.805 ;
        RECT 124.595 108.175 125.115 108.715 ;
        RECT 125.285 108.005 125.805 108.545 ;
        RECT 123.210 107.805 123.960 107.975 ;
        RECT 123.205 107.255 123.535 107.635 ;
        RECT 123.705 107.515 123.960 107.805 ;
        RECT 124.595 107.255 125.805 108.005 ;
        RECT 11.810 107.085 125.890 107.255 ;
        RECT 11.895 106.335 13.105 107.085 ;
        RECT 14.505 106.615 14.675 107.085 ;
        RECT 14.845 106.435 15.175 106.915 ;
        RECT 15.345 106.615 15.515 107.085 ;
        RECT 15.685 106.435 16.015 106.915 ;
        RECT 11.895 105.795 12.415 106.335 ;
        RECT 14.250 106.265 16.015 106.435 ;
        RECT 16.185 106.275 16.355 107.085 ;
        RECT 16.555 106.705 17.625 106.875 ;
        RECT 16.555 106.350 16.875 106.705 ;
        RECT 12.585 105.625 13.105 106.165 ;
        RECT 11.895 104.535 13.105 105.625 ;
        RECT 14.250 105.715 14.660 106.265 ;
        RECT 16.550 106.095 16.875 106.350 ;
        RECT 14.845 105.885 16.875 106.095 ;
        RECT 16.530 105.875 16.875 105.885 ;
        RECT 17.045 106.135 17.285 106.535 ;
        RECT 17.455 106.475 17.625 106.705 ;
        RECT 17.795 106.645 17.985 107.085 ;
        RECT 18.155 106.635 19.105 106.915 ;
        RECT 19.325 106.725 19.675 106.895 ;
        RECT 17.455 106.305 17.985 106.475 ;
        RECT 14.250 105.545 15.975 105.715 ;
        RECT 14.505 104.535 14.675 105.375 ;
        RECT 14.885 104.705 15.135 105.545 ;
        RECT 15.345 104.535 15.515 105.375 ;
        RECT 15.685 104.705 15.975 105.545 ;
        RECT 16.185 104.535 16.355 105.595 ;
        RECT 16.530 105.255 16.700 105.875 ;
        RECT 17.045 105.765 17.585 106.135 ;
        RECT 17.765 106.025 17.985 106.305 ;
        RECT 18.155 105.855 18.325 106.635 ;
        RECT 17.920 105.685 18.325 105.855 ;
        RECT 18.495 105.845 18.845 106.465 ;
        RECT 17.920 105.595 18.090 105.685 ;
        RECT 19.015 105.675 19.225 106.465 ;
        RECT 16.870 105.425 18.090 105.595 ;
        RECT 18.550 105.515 19.225 105.675 ;
        RECT 16.530 105.085 17.330 105.255 ;
        RECT 16.650 104.535 16.980 104.915 ;
        RECT 17.160 104.795 17.330 105.085 ;
        RECT 17.920 105.045 18.090 105.425 ;
        RECT 18.260 105.505 19.225 105.515 ;
        RECT 19.415 106.335 19.675 106.725 ;
        RECT 19.885 106.625 20.215 107.085 ;
        RECT 21.090 106.695 21.945 106.865 ;
        RECT 22.150 106.695 22.645 106.865 ;
        RECT 22.815 106.725 23.145 107.085 ;
        RECT 19.415 105.645 19.585 106.335 ;
        RECT 19.755 105.985 19.925 106.165 ;
        RECT 20.095 106.155 20.885 106.405 ;
        RECT 21.090 105.985 21.260 106.695 ;
        RECT 21.430 106.185 21.785 106.405 ;
        RECT 19.755 105.815 21.445 105.985 ;
        RECT 18.260 105.215 18.720 105.505 ;
        RECT 19.415 105.475 20.915 105.645 ;
        RECT 19.415 105.335 19.585 105.475 ;
        RECT 19.025 105.165 19.585 105.335 ;
        RECT 17.500 104.535 17.750 104.995 ;
        RECT 17.920 104.705 18.790 105.045 ;
        RECT 19.025 104.705 19.195 105.165 ;
        RECT 20.030 105.135 21.105 105.305 ;
        RECT 19.365 104.535 19.735 104.995 ;
        RECT 20.030 104.795 20.200 105.135 ;
        RECT 20.370 104.535 20.700 104.965 ;
        RECT 20.935 104.795 21.105 105.135 ;
        RECT 21.275 105.035 21.445 105.815 ;
        RECT 21.615 105.595 21.785 106.185 ;
        RECT 21.955 105.785 22.305 106.405 ;
        RECT 21.615 105.205 22.080 105.595 ;
        RECT 22.475 105.335 22.645 106.695 ;
        RECT 22.815 105.505 23.275 106.555 ;
        RECT 22.250 105.165 22.645 105.335 ;
        RECT 22.250 105.035 22.420 105.165 ;
        RECT 21.275 104.705 21.955 105.035 ;
        RECT 22.170 104.705 22.420 105.035 ;
        RECT 22.590 104.535 22.840 104.995 ;
        RECT 23.010 104.720 23.335 105.505 ;
        RECT 23.505 104.705 23.675 106.825 ;
        RECT 23.845 106.705 24.175 107.085 ;
        RECT 24.345 106.535 24.600 106.825 ;
        RECT 23.850 106.365 24.600 106.535 ;
        RECT 24.780 106.535 25.035 106.825 ;
        RECT 25.205 106.705 25.535 107.085 ;
        RECT 24.780 106.365 25.530 106.535 ;
        RECT 23.850 105.375 24.080 106.365 ;
        RECT 24.250 105.545 24.600 106.195 ;
        RECT 24.780 105.545 25.130 106.195 ;
        RECT 25.300 105.375 25.530 106.365 ;
        RECT 23.850 105.205 24.600 105.375 ;
        RECT 23.845 104.535 24.175 105.035 ;
        RECT 24.345 104.705 24.600 105.205 ;
        RECT 24.780 105.205 25.530 105.375 ;
        RECT 24.780 104.705 25.035 105.205 ;
        RECT 25.205 104.535 25.535 105.035 ;
        RECT 25.705 104.705 25.875 106.825 ;
        RECT 26.235 106.725 26.565 107.085 ;
        RECT 26.735 106.695 27.230 106.865 ;
        RECT 27.435 106.695 28.290 106.865 ;
        RECT 26.105 105.505 26.565 106.555 ;
        RECT 26.045 104.720 26.370 105.505 ;
        RECT 26.735 105.335 26.905 106.695 ;
        RECT 27.075 105.785 27.425 106.405 ;
        RECT 27.595 106.185 27.950 106.405 ;
        RECT 27.595 105.595 27.765 106.185 ;
        RECT 28.120 105.985 28.290 106.695 ;
        RECT 29.165 106.625 29.495 107.085 ;
        RECT 29.705 106.725 30.055 106.895 ;
        RECT 28.495 106.155 29.285 106.405 ;
        RECT 29.705 106.335 29.965 106.725 ;
        RECT 30.275 106.635 31.225 106.915 ;
        RECT 31.395 106.645 31.585 107.085 ;
        RECT 31.755 106.705 32.825 106.875 ;
        RECT 29.455 105.985 29.625 106.165 ;
        RECT 26.735 105.165 27.130 105.335 ;
        RECT 27.300 105.205 27.765 105.595 ;
        RECT 27.935 105.815 29.625 105.985 ;
        RECT 26.960 105.035 27.130 105.165 ;
        RECT 27.935 105.035 28.105 105.815 ;
        RECT 29.795 105.645 29.965 106.335 ;
        RECT 28.465 105.475 29.965 105.645 ;
        RECT 30.155 105.675 30.365 106.465 ;
        RECT 30.535 105.845 30.885 106.465 ;
        RECT 31.055 105.855 31.225 106.635 ;
        RECT 31.755 106.475 31.925 106.705 ;
        RECT 31.395 106.305 31.925 106.475 ;
        RECT 31.395 106.025 31.615 106.305 ;
        RECT 32.095 106.135 32.335 106.535 ;
        RECT 31.055 105.685 31.460 105.855 ;
        RECT 31.795 105.765 32.335 106.135 ;
        RECT 32.505 106.350 32.825 106.705 ;
        RECT 32.505 106.095 32.830 106.350 ;
        RECT 33.025 106.275 33.195 107.085 ;
        RECT 33.365 106.435 33.695 106.915 ;
        RECT 33.865 106.615 34.035 107.085 ;
        RECT 34.205 106.435 34.535 106.915 ;
        RECT 34.705 106.615 34.875 107.085 ;
        RECT 33.365 106.265 35.130 106.435 ;
        RECT 35.355 106.360 35.645 107.085 ;
        RECT 36.335 106.265 36.545 107.085 ;
        RECT 36.715 106.285 37.045 106.915 ;
        RECT 32.505 105.885 34.535 106.095 ;
        RECT 32.505 105.875 32.850 105.885 ;
        RECT 30.155 105.515 30.830 105.675 ;
        RECT 31.290 105.595 31.460 105.685 ;
        RECT 30.155 105.505 31.120 105.515 ;
        RECT 29.795 105.335 29.965 105.475 ;
        RECT 26.540 104.535 26.790 104.995 ;
        RECT 26.960 104.705 27.210 105.035 ;
        RECT 27.425 104.705 28.105 105.035 ;
        RECT 28.275 105.135 29.350 105.305 ;
        RECT 29.795 105.165 30.355 105.335 ;
        RECT 30.660 105.215 31.120 105.505 ;
        RECT 31.290 105.425 32.510 105.595 ;
        RECT 28.275 104.795 28.445 105.135 ;
        RECT 28.680 104.535 29.010 104.965 ;
        RECT 29.180 104.795 29.350 105.135 ;
        RECT 29.645 104.535 30.015 104.995 ;
        RECT 30.185 104.705 30.355 105.165 ;
        RECT 31.290 105.045 31.460 105.425 ;
        RECT 32.680 105.255 32.850 105.875 ;
        RECT 34.720 105.715 35.130 106.265 ;
        RECT 30.590 104.705 31.460 105.045 ;
        RECT 32.050 105.085 32.850 105.255 ;
        RECT 31.630 104.535 31.880 104.995 ;
        RECT 32.050 104.795 32.220 105.085 ;
        RECT 32.400 104.535 32.730 104.915 ;
        RECT 33.025 104.535 33.195 105.595 ;
        RECT 33.405 105.545 35.130 105.715 ;
        RECT 33.405 104.705 33.695 105.545 ;
        RECT 33.865 104.535 34.035 105.375 ;
        RECT 34.245 104.705 34.495 105.545 ;
        RECT 34.705 104.535 34.875 105.375 ;
        RECT 35.355 104.535 35.645 105.700 ;
        RECT 36.715 105.685 36.965 106.285 ;
        RECT 37.215 106.265 37.445 107.085 ;
        RECT 38.115 106.315 39.785 107.085 ;
        RECT 39.960 106.535 40.215 106.825 ;
        RECT 40.385 106.705 40.715 107.085 ;
        RECT 39.960 106.365 40.710 106.535 ;
        RECT 37.135 105.845 37.465 106.095 ;
        RECT 36.335 104.535 36.545 105.675 ;
        RECT 36.715 104.705 37.045 105.685 ;
        RECT 37.215 104.535 37.445 105.675 ;
        RECT 38.115 105.625 38.865 106.145 ;
        RECT 39.035 105.795 39.785 106.315 ;
        RECT 38.115 104.535 39.785 105.625 ;
        RECT 39.960 105.545 40.310 106.195 ;
        RECT 40.480 105.375 40.710 106.365 ;
        RECT 39.960 105.205 40.710 105.375 ;
        RECT 39.960 104.705 40.215 105.205 ;
        RECT 40.385 104.535 40.715 105.035 ;
        RECT 40.885 104.705 41.055 106.825 ;
        RECT 41.415 106.725 41.745 107.085 ;
        RECT 41.915 106.695 42.410 106.865 ;
        RECT 42.615 106.695 43.470 106.865 ;
        RECT 41.285 105.505 41.745 106.555 ;
        RECT 41.225 104.720 41.550 105.505 ;
        RECT 41.915 105.335 42.085 106.695 ;
        RECT 42.255 105.785 42.605 106.405 ;
        RECT 42.775 106.185 43.130 106.405 ;
        RECT 42.775 105.595 42.945 106.185 ;
        RECT 43.300 105.985 43.470 106.695 ;
        RECT 44.345 106.625 44.675 107.085 ;
        RECT 44.885 106.725 45.235 106.895 ;
        RECT 43.675 106.155 44.465 106.405 ;
        RECT 44.885 106.335 45.145 106.725 ;
        RECT 45.455 106.635 46.405 106.915 ;
        RECT 46.575 106.645 46.765 107.085 ;
        RECT 46.935 106.705 48.005 106.875 ;
        RECT 44.635 105.985 44.805 106.165 ;
        RECT 41.915 105.165 42.310 105.335 ;
        RECT 42.480 105.205 42.945 105.595 ;
        RECT 43.115 105.815 44.805 105.985 ;
        RECT 42.140 105.035 42.310 105.165 ;
        RECT 43.115 105.035 43.285 105.815 ;
        RECT 44.975 105.645 45.145 106.335 ;
        RECT 43.645 105.475 45.145 105.645 ;
        RECT 45.335 105.675 45.545 106.465 ;
        RECT 45.715 105.845 46.065 106.465 ;
        RECT 46.235 105.855 46.405 106.635 ;
        RECT 46.935 106.475 47.105 106.705 ;
        RECT 46.575 106.305 47.105 106.475 ;
        RECT 46.575 106.025 46.795 106.305 ;
        RECT 47.275 106.135 47.515 106.535 ;
        RECT 46.235 105.685 46.640 105.855 ;
        RECT 46.975 105.765 47.515 106.135 ;
        RECT 47.685 106.350 48.005 106.705 ;
        RECT 47.685 106.095 48.010 106.350 ;
        RECT 48.205 106.275 48.375 107.085 ;
        RECT 48.545 106.435 48.875 106.915 ;
        RECT 49.045 106.615 49.215 107.085 ;
        RECT 49.385 106.435 49.715 106.915 ;
        RECT 49.885 106.615 50.055 107.085 ;
        RECT 50.540 106.535 50.795 106.825 ;
        RECT 50.965 106.705 51.295 107.085 ;
        RECT 48.545 106.265 50.310 106.435 ;
        RECT 50.540 106.365 51.290 106.535 ;
        RECT 47.685 105.885 49.715 106.095 ;
        RECT 47.685 105.875 48.030 105.885 ;
        RECT 45.335 105.515 46.010 105.675 ;
        RECT 46.470 105.595 46.640 105.685 ;
        RECT 45.335 105.505 46.300 105.515 ;
        RECT 44.975 105.335 45.145 105.475 ;
        RECT 41.720 104.535 41.970 104.995 ;
        RECT 42.140 104.705 42.390 105.035 ;
        RECT 42.605 104.705 43.285 105.035 ;
        RECT 43.455 105.135 44.530 105.305 ;
        RECT 44.975 105.165 45.535 105.335 ;
        RECT 45.840 105.215 46.300 105.505 ;
        RECT 46.470 105.425 47.690 105.595 ;
        RECT 43.455 104.795 43.625 105.135 ;
        RECT 43.860 104.535 44.190 104.965 ;
        RECT 44.360 104.795 44.530 105.135 ;
        RECT 44.825 104.535 45.195 104.995 ;
        RECT 45.365 104.705 45.535 105.165 ;
        RECT 46.470 105.045 46.640 105.425 ;
        RECT 47.860 105.255 48.030 105.875 ;
        RECT 49.900 105.715 50.310 106.265 ;
        RECT 45.770 104.705 46.640 105.045 ;
        RECT 47.230 105.085 48.030 105.255 ;
        RECT 46.810 104.535 47.060 104.995 ;
        RECT 47.230 104.795 47.400 105.085 ;
        RECT 47.580 104.535 47.910 104.915 ;
        RECT 48.205 104.535 48.375 105.595 ;
        RECT 48.585 105.545 50.310 105.715 ;
        RECT 50.540 105.545 50.890 106.195 ;
        RECT 48.585 104.705 48.875 105.545 ;
        RECT 49.045 104.535 49.215 105.375 ;
        RECT 49.425 104.705 49.675 105.545 ;
        RECT 51.060 105.375 51.290 106.365 ;
        RECT 49.885 104.535 50.055 105.375 ;
        RECT 50.540 105.205 51.290 105.375 ;
        RECT 50.540 104.705 50.795 105.205 ;
        RECT 50.965 104.535 51.295 105.035 ;
        RECT 51.465 104.705 51.635 106.825 ;
        RECT 51.995 106.725 52.325 107.085 ;
        RECT 52.495 106.695 52.990 106.865 ;
        RECT 53.195 106.695 54.050 106.865 ;
        RECT 51.865 105.505 52.325 106.555 ;
        RECT 51.805 104.720 52.130 105.505 ;
        RECT 52.495 105.335 52.665 106.695 ;
        RECT 52.835 105.785 53.185 106.405 ;
        RECT 53.355 106.185 53.710 106.405 ;
        RECT 53.355 105.595 53.525 106.185 ;
        RECT 53.880 105.985 54.050 106.695 ;
        RECT 54.925 106.625 55.255 107.085 ;
        RECT 55.465 106.725 55.815 106.895 ;
        RECT 54.255 106.155 55.045 106.405 ;
        RECT 55.465 106.335 55.725 106.725 ;
        RECT 56.035 106.635 56.985 106.915 ;
        RECT 57.155 106.645 57.345 107.085 ;
        RECT 57.515 106.705 58.585 106.875 ;
        RECT 55.215 105.985 55.385 106.165 ;
        RECT 52.495 105.165 52.890 105.335 ;
        RECT 53.060 105.205 53.525 105.595 ;
        RECT 53.695 105.815 55.385 105.985 ;
        RECT 52.720 105.035 52.890 105.165 ;
        RECT 53.695 105.035 53.865 105.815 ;
        RECT 55.555 105.645 55.725 106.335 ;
        RECT 54.225 105.475 55.725 105.645 ;
        RECT 55.915 105.675 56.125 106.465 ;
        RECT 56.295 105.845 56.645 106.465 ;
        RECT 56.815 105.855 56.985 106.635 ;
        RECT 57.515 106.475 57.685 106.705 ;
        RECT 57.155 106.305 57.685 106.475 ;
        RECT 57.155 106.025 57.375 106.305 ;
        RECT 57.855 106.135 58.095 106.535 ;
        RECT 56.815 105.685 57.220 105.855 ;
        RECT 57.555 105.765 58.095 106.135 ;
        RECT 58.265 106.350 58.585 106.705 ;
        RECT 58.265 106.095 58.590 106.350 ;
        RECT 58.785 106.275 58.955 107.085 ;
        RECT 59.125 106.435 59.455 106.915 ;
        RECT 59.625 106.615 59.795 107.085 ;
        RECT 59.965 106.435 60.295 106.915 ;
        RECT 60.465 106.615 60.635 107.085 ;
        RECT 59.125 106.265 60.890 106.435 ;
        RECT 61.115 106.360 61.405 107.085 ;
        RECT 61.885 106.615 62.055 107.085 ;
        RECT 62.225 106.435 62.555 106.915 ;
        RECT 62.725 106.615 62.895 107.085 ;
        RECT 63.065 106.435 63.395 106.915 ;
        RECT 58.265 105.885 60.295 106.095 ;
        RECT 58.265 105.875 58.610 105.885 ;
        RECT 55.915 105.515 56.590 105.675 ;
        RECT 57.050 105.595 57.220 105.685 ;
        RECT 55.915 105.505 56.880 105.515 ;
        RECT 55.555 105.335 55.725 105.475 ;
        RECT 52.300 104.535 52.550 104.995 ;
        RECT 52.720 104.705 52.970 105.035 ;
        RECT 53.185 104.705 53.865 105.035 ;
        RECT 54.035 105.135 55.110 105.305 ;
        RECT 55.555 105.165 56.115 105.335 ;
        RECT 56.420 105.215 56.880 105.505 ;
        RECT 57.050 105.425 58.270 105.595 ;
        RECT 54.035 104.795 54.205 105.135 ;
        RECT 54.440 104.535 54.770 104.965 ;
        RECT 54.940 104.795 55.110 105.135 ;
        RECT 55.405 104.535 55.775 104.995 ;
        RECT 55.945 104.705 56.115 105.165 ;
        RECT 57.050 105.045 57.220 105.425 ;
        RECT 58.440 105.255 58.610 105.875 ;
        RECT 60.480 105.715 60.890 106.265 ;
        RECT 56.350 104.705 57.220 105.045 ;
        RECT 57.810 105.085 58.610 105.255 ;
        RECT 57.390 104.535 57.640 104.995 ;
        RECT 57.810 104.795 57.980 105.085 ;
        RECT 58.160 104.535 58.490 104.915 ;
        RECT 58.785 104.535 58.955 105.595 ;
        RECT 59.165 105.545 60.890 105.715 ;
        RECT 61.630 106.265 63.395 106.435 ;
        RECT 63.565 106.275 63.735 107.085 ;
        RECT 63.935 106.705 65.005 106.875 ;
        RECT 63.935 106.350 64.255 106.705 ;
        RECT 61.630 105.715 62.040 106.265 ;
        RECT 63.930 106.095 64.255 106.350 ;
        RECT 62.225 105.885 64.255 106.095 ;
        RECT 63.910 105.875 64.255 105.885 ;
        RECT 64.425 106.135 64.665 106.535 ;
        RECT 64.835 106.475 65.005 106.705 ;
        RECT 65.175 106.645 65.365 107.085 ;
        RECT 65.535 106.635 66.485 106.915 ;
        RECT 66.705 106.725 67.055 106.895 ;
        RECT 64.835 106.305 65.365 106.475 ;
        RECT 59.165 104.705 59.455 105.545 ;
        RECT 59.625 104.535 59.795 105.375 ;
        RECT 60.005 104.705 60.255 105.545 ;
        RECT 60.465 104.535 60.635 105.375 ;
        RECT 61.115 104.535 61.405 105.700 ;
        RECT 61.630 105.545 63.355 105.715 ;
        RECT 61.885 104.535 62.055 105.375 ;
        RECT 62.265 104.705 62.515 105.545 ;
        RECT 62.725 104.535 62.895 105.375 ;
        RECT 63.065 104.705 63.355 105.545 ;
        RECT 63.565 104.535 63.735 105.595 ;
        RECT 63.910 105.255 64.080 105.875 ;
        RECT 64.425 105.765 64.965 106.135 ;
        RECT 65.145 106.025 65.365 106.305 ;
        RECT 65.535 105.855 65.705 106.635 ;
        RECT 65.300 105.685 65.705 105.855 ;
        RECT 65.875 105.845 66.225 106.465 ;
        RECT 65.300 105.595 65.470 105.685 ;
        RECT 66.395 105.675 66.605 106.465 ;
        RECT 64.250 105.425 65.470 105.595 ;
        RECT 65.930 105.515 66.605 105.675 ;
        RECT 63.910 105.085 64.710 105.255 ;
        RECT 64.030 104.535 64.360 104.915 ;
        RECT 64.540 104.795 64.710 105.085 ;
        RECT 65.300 105.045 65.470 105.425 ;
        RECT 65.640 105.505 66.605 105.515 ;
        RECT 66.795 106.335 67.055 106.725 ;
        RECT 67.265 106.625 67.595 107.085 ;
        RECT 68.470 106.695 69.325 106.865 ;
        RECT 69.530 106.695 70.025 106.865 ;
        RECT 70.195 106.725 70.525 107.085 ;
        RECT 66.795 105.645 66.965 106.335 ;
        RECT 67.135 105.985 67.305 106.165 ;
        RECT 67.475 106.155 68.265 106.405 ;
        RECT 68.470 105.985 68.640 106.695 ;
        RECT 68.810 106.185 69.165 106.405 ;
        RECT 67.135 105.815 68.825 105.985 ;
        RECT 65.640 105.215 66.100 105.505 ;
        RECT 66.795 105.475 68.295 105.645 ;
        RECT 66.795 105.335 66.965 105.475 ;
        RECT 66.405 105.165 66.965 105.335 ;
        RECT 64.880 104.535 65.130 104.995 ;
        RECT 65.300 104.705 66.170 105.045 ;
        RECT 66.405 104.705 66.575 105.165 ;
        RECT 67.410 105.135 68.485 105.305 ;
        RECT 66.745 104.535 67.115 104.995 ;
        RECT 67.410 104.795 67.580 105.135 ;
        RECT 67.750 104.535 68.080 104.965 ;
        RECT 68.315 104.795 68.485 105.135 ;
        RECT 68.655 105.035 68.825 105.815 ;
        RECT 68.995 105.595 69.165 106.185 ;
        RECT 69.335 105.785 69.685 106.405 ;
        RECT 68.995 105.205 69.460 105.595 ;
        RECT 69.855 105.335 70.025 106.695 ;
        RECT 70.195 105.505 70.655 106.555 ;
        RECT 69.630 105.165 70.025 105.335 ;
        RECT 69.630 105.035 69.800 105.165 ;
        RECT 68.655 104.705 69.335 105.035 ;
        RECT 69.550 104.705 69.800 105.035 ;
        RECT 69.970 104.535 70.220 104.995 ;
        RECT 70.390 104.720 70.715 105.505 ;
        RECT 70.885 104.705 71.055 106.825 ;
        RECT 71.225 106.705 71.555 107.085 ;
        RECT 71.725 106.535 71.980 106.825 ;
        RECT 72.465 106.615 72.635 107.085 ;
        RECT 71.230 106.365 71.980 106.535 ;
        RECT 72.805 106.435 73.135 106.915 ;
        RECT 73.305 106.615 73.475 107.085 ;
        RECT 73.645 106.435 73.975 106.915 ;
        RECT 71.230 105.375 71.460 106.365 ;
        RECT 72.210 106.265 73.975 106.435 ;
        RECT 74.145 106.275 74.315 107.085 ;
        RECT 74.515 106.705 75.585 106.875 ;
        RECT 74.515 106.350 74.835 106.705 ;
        RECT 71.630 105.545 71.980 106.195 ;
        RECT 72.210 105.715 72.620 106.265 ;
        RECT 74.510 106.095 74.835 106.350 ;
        RECT 72.805 105.885 74.835 106.095 ;
        RECT 74.490 105.875 74.835 105.885 ;
        RECT 75.005 106.135 75.245 106.535 ;
        RECT 75.415 106.475 75.585 106.705 ;
        RECT 75.755 106.645 75.945 107.085 ;
        RECT 76.115 106.635 77.065 106.915 ;
        RECT 77.285 106.725 77.635 106.895 ;
        RECT 75.415 106.305 75.945 106.475 ;
        RECT 72.210 105.545 73.935 105.715 ;
        RECT 71.230 105.205 71.980 105.375 ;
        RECT 71.225 104.535 71.555 105.035 ;
        RECT 71.725 104.705 71.980 105.205 ;
        RECT 72.465 104.535 72.635 105.375 ;
        RECT 72.845 104.705 73.095 105.545 ;
        RECT 73.305 104.535 73.475 105.375 ;
        RECT 73.645 104.705 73.935 105.545 ;
        RECT 74.145 104.535 74.315 105.595 ;
        RECT 74.490 105.255 74.660 105.875 ;
        RECT 75.005 105.765 75.545 106.135 ;
        RECT 75.725 106.025 75.945 106.305 ;
        RECT 76.115 105.855 76.285 106.635 ;
        RECT 75.880 105.685 76.285 105.855 ;
        RECT 76.455 105.845 76.805 106.465 ;
        RECT 75.880 105.595 76.050 105.685 ;
        RECT 76.975 105.675 77.185 106.465 ;
        RECT 74.830 105.425 76.050 105.595 ;
        RECT 76.510 105.515 77.185 105.675 ;
        RECT 74.490 105.085 75.290 105.255 ;
        RECT 74.610 104.535 74.940 104.915 ;
        RECT 75.120 104.795 75.290 105.085 ;
        RECT 75.880 105.045 76.050 105.425 ;
        RECT 76.220 105.505 77.185 105.515 ;
        RECT 77.375 106.335 77.635 106.725 ;
        RECT 77.845 106.625 78.175 107.085 ;
        RECT 79.050 106.695 79.905 106.865 ;
        RECT 80.110 106.695 80.605 106.865 ;
        RECT 80.775 106.725 81.105 107.085 ;
        RECT 77.375 105.645 77.545 106.335 ;
        RECT 77.715 105.985 77.885 106.165 ;
        RECT 78.055 106.155 78.845 106.405 ;
        RECT 79.050 105.985 79.220 106.695 ;
        RECT 79.390 106.185 79.745 106.405 ;
        RECT 77.715 105.815 79.405 105.985 ;
        RECT 76.220 105.215 76.680 105.505 ;
        RECT 77.375 105.475 78.875 105.645 ;
        RECT 77.375 105.335 77.545 105.475 ;
        RECT 76.985 105.165 77.545 105.335 ;
        RECT 75.460 104.535 75.710 104.995 ;
        RECT 75.880 104.705 76.750 105.045 ;
        RECT 76.985 104.705 77.155 105.165 ;
        RECT 77.990 105.135 79.065 105.305 ;
        RECT 77.325 104.535 77.695 104.995 ;
        RECT 77.990 104.795 78.160 105.135 ;
        RECT 78.330 104.535 78.660 104.965 ;
        RECT 78.895 104.795 79.065 105.135 ;
        RECT 79.235 105.035 79.405 105.815 ;
        RECT 79.575 105.595 79.745 106.185 ;
        RECT 79.915 105.785 80.265 106.405 ;
        RECT 79.575 105.205 80.040 105.595 ;
        RECT 80.435 105.335 80.605 106.695 ;
        RECT 80.775 105.505 81.235 106.555 ;
        RECT 80.210 105.165 80.605 105.335 ;
        RECT 80.210 105.035 80.380 105.165 ;
        RECT 79.235 104.705 79.915 105.035 ;
        RECT 80.130 104.705 80.380 105.035 ;
        RECT 80.550 104.535 80.800 104.995 ;
        RECT 80.970 104.720 81.295 105.505 ;
        RECT 81.465 104.705 81.635 106.825 ;
        RECT 81.805 106.705 82.135 107.085 ;
        RECT 82.305 106.535 82.560 106.825 ;
        RECT 81.810 106.365 82.560 106.535 ;
        RECT 81.810 105.375 82.040 106.365 ;
        RECT 82.735 106.335 83.945 107.085 ;
        RECT 82.210 105.545 82.560 106.195 ;
        RECT 82.735 105.625 83.255 106.165 ;
        RECT 83.425 105.795 83.945 106.335 ;
        RECT 84.175 106.265 84.385 107.085 ;
        RECT 84.555 106.285 84.885 106.915 ;
        RECT 84.555 105.685 84.805 106.285 ;
        RECT 85.055 106.265 85.285 107.085 ;
        RECT 85.535 106.265 85.765 107.085 ;
        RECT 85.935 106.285 86.265 106.915 ;
        RECT 84.975 105.845 85.305 106.095 ;
        RECT 85.515 105.845 85.845 106.095 ;
        RECT 86.015 105.685 86.265 106.285 ;
        RECT 86.435 106.265 86.645 107.085 ;
        RECT 86.875 106.360 87.165 107.085 ;
        RECT 87.340 106.535 87.595 106.825 ;
        RECT 87.765 106.705 88.095 107.085 ;
        RECT 87.340 106.365 88.090 106.535 ;
        RECT 81.810 105.205 82.560 105.375 ;
        RECT 81.805 104.535 82.135 105.035 ;
        RECT 82.305 104.705 82.560 105.205 ;
        RECT 82.735 104.535 83.945 105.625 ;
        RECT 84.175 104.535 84.385 105.675 ;
        RECT 84.555 104.705 84.885 105.685 ;
        RECT 85.055 104.535 85.285 105.675 ;
        RECT 85.535 104.535 85.765 105.675 ;
        RECT 85.935 104.705 86.265 105.685 ;
        RECT 86.435 104.535 86.645 105.675 ;
        RECT 86.875 104.535 87.165 105.700 ;
        RECT 87.340 105.545 87.690 106.195 ;
        RECT 87.860 105.375 88.090 106.365 ;
        RECT 87.340 105.205 88.090 105.375 ;
        RECT 87.340 104.705 87.595 105.205 ;
        RECT 87.765 104.535 88.095 105.035 ;
        RECT 88.265 104.705 88.435 106.825 ;
        RECT 88.795 106.725 89.125 107.085 ;
        RECT 89.295 106.695 89.790 106.865 ;
        RECT 89.995 106.695 90.850 106.865 ;
        RECT 88.665 105.505 89.125 106.555 ;
        RECT 88.605 104.720 88.930 105.505 ;
        RECT 89.295 105.335 89.465 106.695 ;
        RECT 89.635 105.785 89.985 106.405 ;
        RECT 90.155 106.185 90.510 106.405 ;
        RECT 90.155 105.595 90.325 106.185 ;
        RECT 90.680 105.985 90.850 106.695 ;
        RECT 91.725 106.625 92.055 107.085 ;
        RECT 92.265 106.725 92.615 106.895 ;
        RECT 91.055 106.155 91.845 106.405 ;
        RECT 92.265 106.335 92.525 106.725 ;
        RECT 92.835 106.635 93.785 106.915 ;
        RECT 93.955 106.645 94.145 107.085 ;
        RECT 94.315 106.705 95.385 106.875 ;
        RECT 92.015 105.985 92.185 106.165 ;
        RECT 89.295 105.165 89.690 105.335 ;
        RECT 89.860 105.205 90.325 105.595 ;
        RECT 90.495 105.815 92.185 105.985 ;
        RECT 89.520 105.035 89.690 105.165 ;
        RECT 90.495 105.035 90.665 105.815 ;
        RECT 92.355 105.645 92.525 106.335 ;
        RECT 91.025 105.475 92.525 105.645 ;
        RECT 92.715 105.675 92.925 106.465 ;
        RECT 93.095 105.845 93.445 106.465 ;
        RECT 93.615 105.855 93.785 106.635 ;
        RECT 94.315 106.475 94.485 106.705 ;
        RECT 93.955 106.305 94.485 106.475 ;
        RECT 93.955 106.025 94.175 106.305 ;
        RECT 94.655 106.135 94.895 106.535 ;
        RECT 93.615 105.685 94.020 105.855 ;
        RECT 94.355 105.765 94.895 106.135 ;
        RECT 95.065 106.350 95.385 106.705 ;
        RECT 95.065 106.095 95.390 106.350 ;
        RECT 95.585 106.275 95.755 107.085 ;
        RECT 95.925 106.435 96.255 106.915 ;
        RECT 96.425 106.615 96.595 107.085 ;
        RECT 96.765 106.435 97.095 106.915 ;
        RECT 97.265 106.615 97.435 107.085 ;
        RECT 98.225 106.615 98.395 107.085 ;
        RECT 98.565 106.435 98.895 106.915 ;
        RECT 99.065 106.615 99.235 107.085 ;
        RECT 99.405 106.435 99.735 106.915 ;
        RECT 95.925 106.265 97.690 106.435 ;
        RECT 95.065 105.885 97.095 106.095 ;
        RECT 95.065 105.875 95.410 105.885 ;
        RECT 92.715 105.515 93.390 105.675 ;
        RECT 93.850 105.595 94.020 105.685 ;
        RECT 92.715 105.505 93.680 105.515 ;
        RECT 92.355 105.335 92.525 105.475 ;
        RECT 89.100 104.535 89.350 104.995 ;
        RECT 89.520 104.705 89.770 105.035 ;
        RECT 89.985 104.705 90.665 105.035 ;
        RECT 90.835 105.135 91.910 105.305 ;
        RECT 92.355 105.165 92.915 105.335 ;
        RECT 93.220 105.215 93.680 105.505 ;
        RECT 93.850 105.425 95.070 105.595 ;
        RECT 90.835 104.795 91.005 105.135 ;
        RECT 91.240 104.535 91.570 104.965 ;
        RECT 91.740 104.795 91.910 105.135 ;
        RECT 92.205 104.535 92.575 104.995 ;
        RECT 92.745 104.705 92.915 105.165 ;
        RECT 93.850 105.045 94.020 105.425 ;
        RECT 95.240 105.255 95.410 105.875 ;
        RECT 97.280 105.715 97.690 106.265 ;
        RECT 93.150 104.705 94.020 105.045 ;
        RECT 94.610 105.085 95.410 105.255 ;
        RECT 94.190 104.535 94.440 104.995 ;
        RECT 94.610 104.795 94.780 105.085 ;
        RECT 94.960 104.535 95.290 104.915 ;
        RECT 95.585 104.535 95.755 105.595 ;
        RECT 95.965 105.545 97.690 105.715 ;
        RECT 97.970 106.265 99.735 106.435 ;
        RECT 99.905 106.275 100.075 107.085 ;
        RECT 100.275 106.705 101.345 106.875 ;
        RECT 100.275 106.350 100.595 106.705 ;
        RECT 97.970 105.715 98.380 106.265 ;
        RECT 100.270 106.095 100.595 106.350 ;
        RECT 98.565 105.885 100.595 106.095 ;
        RECT 100.250 105.875 100.595 105.885 ;
        RECT 100.765 106.135 101.005 106.535 ;
        RECT 101.175 106.475 101.345 106.705 ;
        RECT 101.515 106.645 101.705 107.085 ;
        RECT 101.875 106.635 102.825 106.915 ;
        RECT 103.045 106.725 103.395 106.895 ;
        RECT 101.175 106.305 101.705 106.475 ;
        RECT 97.970 105.545 99.695 105.715 ;
        RECT 95.965 104.705 96.255 105.545 ;
        RECT 96.425 104.535 96.595 105.375 ;
        RECT 96.805 104.705 97.055 105.545 ;
        RECT 97.265 104.535 97.435 105.375 ;
        RECT 98.225 104.535 98.395 105.375 ;
        RECT 98.605 104.705 98.855 105.545 ;
        RECT 99.065 104.535 99.235 105.375 ;
        RECT 99.405 104.705 99.695 105.545 ;
        RECT 99.905 104.535 100.075 105.595 ;
        RECT 100.250 105.255 100.420 105.875 ;
        RECT 100.765 105.765 101.305 106.135 ;
        RECT 101.485 106.025 101.705 106.305 ;
        RECT 101.875 105.855 102.045 106.635 ;
        RECT 101.640 105.685 102.045 105.855 ;
        RECT 102.215 105.845 102.565 106.465 ;
        RECT 101.640 105.595 101.810 105.685 ;
        RECT 102.735 105.675 102.945 106.465 ;
        RECT 100.590 105.425 101.810 105.595 ;
        RECT 102.270 105.515 102.945 105.675 ;
        RECT 100.250 105.085 101.050 105.255 ;
        RECT 100.370 104.535 100.700 104.915 ;
        RECT 100.880 104.795 101.050 105.085 ;
        RECT 101.640 105.045 101.810 105.425 ;
        RECT 101.980 105.505 102.945 105.515 ;
        RECT 103.135 106.335 103.395 106.725 ;
        RECT 103.605 106.625 103.935 107.085 ;
        RECT 104.810 106.695 105.665 106.865 ;
        RECT 105.870 106.695 106.365 106.865 ;
        RECT 106.535 106.725 106.865 107.085 ;
        RECT 103.135 105.645 103.305 106.335 ;
        RECT 103.475 105.985 103.645 106.165 ;
        RECT 103.815 106.155 104.605 106.405 ;
        RECT 104.810 105.985 104.980 106.695 ;
        RECT 105.150 106.185 105.505 106.405 ;
        RECT 103.475 105.815 105.165 105.985 ;
        RECT 101.980 105.215 102.440 105.505 ;
        RECT 103.135 105.475 104.635 105.645 ;
        RECT 103.135 105.335 103.305 105.475 ;
        RECT 102.745 105.165 103.305 105.335 ;
        RECT 101.220 104.535 101.470 104.995 ;
        RECT 101.640 104.705 102.510 105.045 ;
        RECT 102.745 104.705 102.915 105.165 ;
        RECT 103.750 105.135 104.825 105.305 ;
        RECT 103.085 104.535 103.455 104.995 ;
        RECT 103.750 104.795 103.920 105.135 ;
        RECT 104.090 104.535 104.420 104.965 ;
        RECT 104.655 104.795 104.825 105.135 ;
        RECT 104.995 105.035 105.165 105.815 ;
        RECT 105.335 105.595 105.505 106.185 ;
        RECT 105.675 105.785 106.025 106.405 ;
        RECT 105.335 105.205 105.800 105.595 ;
        RECT 106.195 105.335 106.365 106.695 ;
        RECT 106.535 105.505 106.995 106.555 ;
        RECT 105.970 105.165 106.365 105.335 ;
        RECT 105.970 105.035 106.140 105.165 ;
        RECT 104.995 104.705 105.675 105.035 ;
        RECT 105.890 104.705 106.140 105.035 ;
        RECT 106.310 104.535 106.560 104.995 ;
        RECT 106.730 104.720 107.055 105.505 ;
        RECT 107.225 104.705 107.395 106.825 ;
        RECT 107.565 106.705 107.895 107.085 ;
        RECT 108.065 106.535 108.320 106.825 ;
        RECT 107.570 106.365 108.320 106.535 ;
        RECT 107.570 105.375 107.800 106.365 ;
        RECT 108.955 106.315 112.465 107.085 ;
        RECT 112.635 106.360 112.925 107.085 ;
        RECT 113.405 106.615 113.575 107.085 ;
        RECT 113.745 106.435 114.075 106.915 ;
        RECT 114.245 106.615 114.415 107.085 ;
        RECT 114.585 106.435 114.915 106.915 ;
        RECT 107.970 105.545 108.320 106.195 ;
        RECT 108.955 105.625 110.645 106.145 ;
        RECT 110.815 105.795 112.465 106.315 ;
        RECT 113.150 106.265 114.915 106.435 ;
        RECT 115.085 106.275 115.255 107.085 ;
        RECT 115.455 106.705 116.525 106.875 ;
        RECT 115.455 106.350 115.775 106.705 ;
        RECT 113.150 105.715 113.560 106.265 ;
        RECT 115.450 106.095 115.775 106.350 ;
        RECT 113.745 105.885 115.775 106.095 ;
        RECT 115.430 105.875 115.775 105.885 ;
        RECT 115.945 106.135 116.185 106.535 ;
        RECT 116.355 106.475 116.525 106.705 ;
        RECT 116.695 106.645 116.885 107.085 ;
        RECT 117.055 106.635 118.005 106.915 ;
        RECT 118.225 106.725 118.575 106.895 ;
        RECT 116.355 106.305 116.885 106.475 ;
        RECT 107.570 105.205 108.320 105.375 ;
        RECT 107.565 104.535 107.895 105.035 ;
        RECT 108.065 104.705 108.320 105.205 ;
        RECT 108.955 104.535 112.465 105.625 ;
        RECT 112.635 104.535 112.925 105.700 ;
        RECT 113.150 105.545 114.875 105.715 ;
        RECT 113.405 104.535 113.575 105.375 ;
        RECT 113.785 104.705 114.035 105.545 ;
        RECT 114.245 104.535 114.415 105.375 ;
        RECT 114.585 104.705 114.875 105.545 ;
        RECT 115.085 104.535 115.255 105.595 ;
        RECT 115.430 105.255 115.600 105.875 ;
        RECT 115.945 105.765 116.485 106.135 ;
        RECT 116.665 106.025 116.885 106.305 ;
        RECT 117.055 105.855 117.225 106.635 ;
        RECT 116.820 105.685 117.225 105.855 ;
        RECT 117.395 105.845 117.745 106.465 ;
        RECT 116.820 105.595 116.990 105.685 ;
        RECT 117.915 105.675 118.125 106.465 ;
        RECT 115.770 105.425 116.990 105.595 ;
        RECT 117.450 105.515 118.125 105.675 ;
        RECT 115.430 105.085 116.230 105.255 ;
        RECT 115.550 104.535 115.880 104.915 ;
        RECT 116.060 104.795 116.230 105.085 ;
        RECT 116.820 105.045 116.990 105.425 ;
        RECT 117.160 105.505 118.125 105.515 ;
        RECT 118.315 106.335 118.575 106.725 ;
        RECT 118.785 106.625 119.115 107.085 ;
        RECT 119.990 106.695 120.845 106.865 ;
        RECT 121.050 106.695 121.545 106.865 ;
        RECT 121.715 106.725 122.045 107.085 ;
        RECT 118.315 105.645 118.485 106.335 ;
        RECT 118.655 105.985 118.825 106.165 ;
        RECT 118.995 106.155 119.785 106.405 ;
        RECT 119.990 105.985 120.160 106.695 ;
        RECT 120.330 106.185 120.685 106.405 ;
        RECT 118.655 105.815 120.345 105.985 ;
        RECT 117.160 105.215 117.620 105.505 ;
        RECT 118.315 105.475 119.815 105.645 ;
        RECT 118.315 105.335 118.485 105.475 ;
        RECT 117.925 105.165 118.485 105.335 ;
        RECT 116.400 104.535 116.650 104.995 ;
        RECT 116.820 104.705 117.690 105.045 ;
        RECT 117.925 104.705 118.095 105.165 ;
        RECT 118.930 105.135 120.005 105.305 ;
        RECT 118.265 104.535 118.635 104.995 ;
        RECT 118.930 104.795 119.100 105.135 ;
        RECT 119.270 104.535 119.600 104.965 ;
        RECT 119.835 104.795 120.005 105.135 ;
        RECT 120.175 105.035 120.345 105.815 ;
        RECT 120.515 105.595 120.685 106.185 ;
        RECT 120.855 105.785 121.205 106.405 ;
        RECT 120.515 105.205 120.980 105.595 ;
        RECT 121.375 105.335 121.545 106.695 ;
        RECT 121.715 105.505 122.175 106.555 ;
        RECT 121.150 105.165 121.545 105.335 ;
        RECT 121.150 105.035 121.320 105.165 ;
        RECT 120.175 104.705 120.855 105.035 ;
        RECT 121.070 104.705 121.320 105.035 ;
        RECT 121.490 104.535 121.740 104.995 ;
        RECT 121.910 104.720 122.235 105.505 ;
        RECT 122.405 104.705 122.575 106.825 ;
        RECT 122.745 106.705 123.075 107.085 ;
        RECT 123.245 106.535 123.500 106.825 ;
        RECT 122.750 106.365 123.500 106.535 ;
        RECT 122.750 105.375 122.980 106.365 ;
        RECT 124.595 106.335 125.805 107.085 ;
        RECT 123.150 105.545 123.500 106.195 ;
        RECT 124.595 105.625 125.115 106.165 ;
        RECT 125.285 105.795 125.805 106.335 ;
        RECT 122.750 105.205 123.500 105.375 ;
        RECT 122.745 104.535 123.075 105.035 ;
        RECT 123.245 104.705 123.500 105.205 ;
        RECT 124.595 104.535 125.805 105.625 ;
        RECT 11.810 104.365 125.890 104.535 ;
        RECT 11.895 103.275 13.105 104.365 ;
        RECT 11.895 102.565 12.415 103.105 ;
        RECT 12.585 102.735 13.105 103.275 ;
        RECT 13.275 103.275 16.785 104.365 ;
        RECT 16.960 103.930 22.305 104.365 ;
        RECT 13.275 102.755 14.965 103.275 ;
        RECT 15.135 102.585 16.785 103.105 ;
        RECT 18.550 102.680 18.900 103.930 ;
        RECT 22.475 103.200 22.765 104.365 ;
        RECT 23.245 103.525 23.415 104.365 ;
        RECT 23.625 103.355 23.875 104.195 ;
        RECT 24.085 103.525 24.255 104.365 ;
        RECT 24.425 103.355 24.715 104.195 ;
        RECT 11.895 101.815 13.105 102.565 ;
        RECT 13.275 101.815 16.785 102.585 ;
        RECT 20.380 102.360 20.720 103.190 ;
        RECT 22.990 103.185 24.715 103.355 ;
        RECT 24.925 103.305 25.095 104.365 ;
        RECT 25.390 103.985 25.720 104.365 ;
        RECT 25.900 103.815 26.070 104.105 ;
        RECT 26.240 103.905 26.490 104.365 ;
        RECT 25.270 103.645 26.070 103.815 ;
        RECT 26.660 103.855 27.530 104.195 ;
        RECT 22.990 102.635 23.400 103.185 ;
        RECT 25.270 103.025 25.440 103.645 ;
        RECT 26.660 103.475 26.830 103.855 ;
        RECT 27.765 103.735 27.935 104.195 ;
        RECT 28.105 103.905 28.475 104.365 ;
        RECT 28.770 103.765 28.940 104.105 ;
        RECT 29.110 103.935 29.440 104.365 ;
        RECT 29.675 103.765 29.845 104.105 ;
        RECT 25.610 103.305 26.830 103.475 ;
        RECT 27.000 103.395 27.460 103.685 ;
        RECT 27.765 103.565 28.325 103.735 ;
        RECT 28.770 103.595 29.845 103.765 ;
        RECT 30.015 103.865 30.695 104.195 ;
        RECT 30.910 103.865 31.160 104.195 ;
        RECT 31.330 103.905 31.580 104.365 ;
        RECT 28.155 103.425 28.325 103.565 ;
        RECT 27.000 103.385 27.965 103.395 ;
        RECT 26.660 103.215 26.830 103.305 ;
        RECT 27.290 103.225 27.965 103.385 ;
        RECT 25.270 103.015 25.615 103.025 ;
        RECT 23.585 102.805 25.615 103.015 ;
        RECT 16.960 101.815 22.305 102.360 ;
        RECT 22.475 101.815 22.765 102.540 ;
        RECT 22.990 102.465 24.755 102.635 ;
        RECT 23.245 101.815 23.415 102.285 ;
        RECT 23.585 101.985 23.915 102.465 ;
        RECT 24.085 101.815 24.255 102.285 ;
        RECT 24.425 101.985 24.755 102.465 ;
        RECT 24.925 101.815 25.095 102.625 ;
        RECT 25.290 102.550 25.615 102.805 ;
        RECT 25.295 102.195 25.615 102.550 ;
        RECT 25.785 102.765 26.325 103.135 ;
        RECT 26.660 103.045 27.065 103.215 ;
        RECT 25.785 102.365 26.025 102.765 ;
        RECT 26.505 102.595 26.725 102.875 ;
        RECT 26.195 102.425 26.725 102.595 ;
        RECT 26.195 102.195 26.365 102.425 ;
        RECT 26.895 102.265 27.065 103.045 ;
        RECT 27.235 102.435 27.585 103.055 ;
        RECT 27.755 102.435 27.965 103.225 ;
        RECT 28.155 103.255 29.655 103.425 ;
        RECT 28.155 102.565 28.325 103.255 ;
        RECT 30.015 103.085 30.185 103.865 ;
        RECT 30.990 103.735 31.160 103.865 ;
        RECT 28.495 102.915 30.185 103.085 ;
        RECT 30.355 103.305 30.820 103.695 ;
        RECT 30.990 103.565 31.385 103.735 ;
        RECT 28.495 102.735 28.665 102.915 ;
        RECT 25.295 102.025 26.365 102.195 ;
        RECT 26.535 101.815 26.725 102.255 ;
        RECT 26.895 101.985 27.845 102.265 ;
        RECT 28.155 102.175 28.415 102.565 ;
        RECT 28.835 102.495 29.625 102.745 ;
        RECT 28.065 102.005 28.415 102.175 ;
        RECT 28.625 101.815 28.955 102.275 ;
        RECT 29.830 102.205 30.000 102.915 ;
        RECT 30.355 102.715 30.525 103.305 ;
        RECT 30.170 102.495 30.525 102.715 ;
        RECT 30.695 102.495 31.045 103.115 ;
        RECT 31.215 102.205 31.385 103.565 ;
        RECT 31.750 103.395 32.075 104.180 ;
        RECT 31.555 102.345 32.015 103.395 ;
        RECT 29.830 102.035 30.685 102.205 ;
        RECT 30.890 102.035 31.385 102.205 ;
        RECT 31.555 101.815 31.885 102.175 ;
        RECT 32.245 102.075 32.415 104.195 ;
        RECT 32.585 103.865 32.915 104.365 ;
        RECT 33.085 103.695 33.340 104.195 ;
        RECT 32.590 103.525 33.340 103.695 ;
        RECT 32.590 102.535 32.820 103.525 ;
        RECT 32.990 102.705 33.340 103.355 ;
        RECT 33.515 103.275 35.185 104.365 ;
        RECT 33.515 102.755 34.265 103.275 ;
        RECT 35.355 103.200 35.645 104.365 ;
        RECT 35.820 103.930 41.165 104.365 ;
        RECT 41.340 103.930 46.685 104.365 ;
        RECT 34.435 102.585 35.185 103.105 ;
        RECT 37.410 102.680 37.760 103.930 ;
        RECT 32.590 102.365 33.340 102.535 ;
        RECT 32.585 101.815 32.915 102.195 ;
        RECT 33.085 102.075 33.340 102.365 ;
        RECT 33.515 101.815 35.185 102.585 ;
        RECT 35.355 101.815 35.645 102.540 ;
        RECT 39.240 102.360 39.580 103.190 ;
        RECT 42.930 102.680 43.280 103.930 ;
        RECT 46.915 103.225 47.125 104.365 ;
        RECT 47.295 103.215 47.625 104.195 ;
        RECT 47.795 103.225 48.025 104.365 ;
        RECT 44.760 102.360 45.100 103.190 ;
        RECT 35.820 101.815 41.165 102.360 ;
        RECT 41.340 101.815 46.685 102.360 ;
        RECT 46.915 101.815 47.125 102.635 ;
        RECT 47.295 102.615 47.545 103.215 ;
        RECT 48.235 103.200 48.525 104.365 ;
        RECT 48.700 103.930 54.045 104.365 ;
        RECT 54.220 103.930 59.565 104.365 ;
        RECT 47.715 102.805 48.045 103.055 ;
        RECT 50.290 102.680 50.640 103.930 ;
        RECT 47.295 101.985 47.625 102.615 ;
        RECT 47.795 101.815 48.025 102.635 ;
        RECT 48.235 101.815 48.525 102.540 ;
        RECT 52.120 102.360 52.460 103.190 ;
        RECT 55.810 102.680 56.160 103.930 ;
        RECT 59.775 103.225 60.005 104.365 ;
        RECT 60.175 103.215 60.505 104.195 ;
        RECT 60.675 103.225 60.885 104.365 ;
        RECT 57.640 102.360 57.980 103.190 ;
        RECT 59.755 102.805 60.085 103.055 ;
        RECT 48.700 101.815 54.045 102.360 ;
        RECT 54.220 101.815 59.565 102.360 ;
        RECT 59.775 101.815 60.005 102.635 ;
        RECT 60.255 102.615 60.505 103.215 ;
        RECT 61.115 103.200 61.405 104.365 ;
        RECT 62.075 103.225 62.305 104.365 ;
        RECT 62.475 103.215 62.805 104.195 ;
        RECT 62.975 103.225 63.185 104.365 ;
        RECT 63.415 103.275 66.925 104.365 ;
        RECT 67.100 103.930 72.445 104.365 ;
        RECT 62.055 102.805 62.385 103.055 ;
        RECT 60.175 101.985 60.505 102.615 ;
        RECT 60.675 101.815 60.885 102.635 ;
        RECT 61.115 101.815 61.405 102.540 ;
        RECT 62.075 101.815 62.305 102.635 ;
        RECT 62.555 102.615 62.805 103.215 ;
        RECT 63.415 102.755 65.105 103.275 ;
        RECT 62.475 101.985 62.805 102.615 ;
        RECT 62.975 101.815 63.185 102.635 ;
        RECT 65.275 102.585 66.925 103.105 ;
        RECT 68.690 102.680 69.040 103.930 ;
        RECT 72.675 103.225 72.885 104.365 ;
        RECT 73.055 103.215 73.385 104.195 ;
        RECT 73.555 103.225 73.785 104.365 ;
        RECT 63.415 101.815 66.925 102.585 ;
        RECT 70.520 102.360 70.860 103.190 ;
        RECT 67.100 101.815 72.445 102.360 ;
        RECT 72.675 101.815 72.885 102.635 ;
        RECT 73.055 102.615 73.305 103.215 ;
        RECT 73.995 103.200 74.285 104.365 ;
        RECT 74.955 103.225 75.185 104.365 ;
        RECT 75.355 103.215 75.685 104.195 ;
        RECT 75.855 103.225 76.065 104.365 ;
        RECT 76.605 103.525 76.775 104.365 ;
        RECT 76.985 103.355 77.235 104.195 ;
        RECT 77.445 103.525 77.615 104.365 ;
        RECT 77.785 103.355 78.075 104.195 ;
        RECT 73.475 102.805 73.805 103.055 ;
        RECT 74.935 102.805 75.265 103.055 ;
        RECT 73.055 101.985 73.385 102.615 ;
        RECT 73.555 101.815 73.785 102.635 ;
        RECT 73.995 101.815 74.285 102.540 ;
        RECT 74.955 101.815 75.185 102.635 ;
        RECT 75.435 102.615 75.685 103.215 ;
        RECT 76.350 103.185 78.075 103.355 ;
        RECT 78.285 103.305 78.455 104.365 ;
        RECT 78.750 103.985 79.080 104.365 ;
        RECT 79.260 103.815 79.430 104.105 ;
        RECT 79.600 103.905 79.850 104.365 ;
        RECT 78.630 103.645 79.430 103.815 ;
        RECT 80.020 103.855 80.890 104.195 ;
        RECT 76.350 102.635 76.760 103.185 ;
        RECT 78.630 103.025 78.800 103.645 ;
        RECT 80.020 103.475 80.190 103.855 ;
        RECT 81.125 103.735 81.295 104.195 ;
        RECT 81.465 103.905 81.835 104.365 ;
        RECT 82.130 103.765 82.300 104.105 ;
        RECT 82.470 103.935 82.800 104.365 ;
        RECT 83.035 103.765 83.205 104.105 ;
        RECT 78.970 103.305 80.190 103.475 ;
        RECT 80.360 103.395 80.820 103.685 ;
        RECT 81.125 103.565 81.685 103.735 ;
        RECT 82.130 103.595 83.205 103.765 ;
        RECT 83.375 103.865 84.055 104.195 ;
        RECT 84.270 103.865 84.520 104.195 ;
        RECT 84.690 103.905 84.940 104.365 ;
        RECT 81.515 103.425 81.685 103.565 ;
        RECT 80.360 103.385 81.325 103.395 ;
        RECT 80.020 103.215 80.190 103.305 ;
        RECT 80.650 103.225 81.325 103.385 ;
        RECT 78.630 103.015 78.975 103.025 ;
        RECT 76.945 102.805 78.975 103.015 ;
        RECT 75.355 101.985 75.685 102.615 ;
        RECT 75.855 101.815 76.065 102.635 ;
        RECT 76.350 102.465 78.115 102.635 ;
        RECT 76.605 101.815 76.775 102.285 ;
        RECT 76.945 101.985 77.275 102.465 ;
        RECT 77.445 101.815 77.615 102.285 ;
        RECT 77.785 101.985 78.115 102.465 ;
        RECT 78.285 101.815 78.455 102.625 ;
        RECT 78.650 102.550 78.975 102.805 ;
        RECT 78.655 102.195 78.975 102.550 ;
        RECT 79.145 102.765 79.685 103.135 ;
        RECT 80.020 103.045 80.425 103.215 ;
        RECT 79.145 102.365 79.385 102.765 ;
        RECT 79.865 102.595 80.085 102.875 ;
        RECT 79.555 102.425 80.085 102.595 ;
        RECT 79.555 102.195 79.725 102.425 ;
        RECT 80.255 102.265 80.425 103.045 ;
        RECT 80.595 102.435 80.945 103.055 ;
        RECT 81.115 102.435 81.325 103.225 ;
        RECT 81.515 103.255 83.015 103.425 ;
        RECT 81.515 102.565 81.685 103.255 ;
        RECT 83.375 103.085 83.545 103.865 ;
        RECT 84.350 103.735 84.520 103.865 ;
        RECT 81.855 102.915 83.545 103.085 ;
        RECT 83.715 103.305 84.180 103.695 ;
        RECT 84.350 103.565 84.745 103.735 ;
        RECT 81.855 102.735 82.025 102.915 ;
        RECT 78.655 102.025 79.725 102.195 ;
        RECT 79.895 101.815 80.085 102.255 ;
        RECT 80.255 101.985 81.205 102.265 ;
        RECT 81.515 102.175 81.775 102.565 ;
        RECT 82.195 102.495 82.985 102.745 ;
        RECT 81.425 102.005 81.775 102.175 ;
        RECT 81.985 101.815 82.315 102.275 ;
        RECT 83.190 102.205 83.360 102.915 ;
        RECT 83.715 102.715 83.885 103.305 ;
        RECT 83.530 102.495 83.885 102.715 ;
        RECT 84.055 102.495 84.405 103.115 ;
        RECT 84.575 102.205 84.745 103.565 ;
        RECT 85.110 103.395 85.435 104.180 ;
        RECT 84.915 102.345 85.375 103.395 ;
        RECT 83.190 102.035 84.045 102.205 ;
        RECT 84.250 102.035 84.745 102.205 ;
        RECT 84.915 101.815 85.245 102.175 ;
        RECT 85.605 102.075 85.775 104.195 ;
        RECT 85.945 103.865 86.275 104.365 ;
        RECT 86.445 103.695 86.700 104.195 ;
        RECT 85.950 103.525 86.700 103.695 ;
        RECT 85.950 102.535 86.180 103.525 ;
        RECT 86.350 102.705 86.700 103.355 ;
        RECT 86.875 103.200 87.165 104.365 ;
        RECT 87.335 103.275 89.005 104.365 ;
        RECT 89.180 103.930 94.525 104.365 ;
        RECT 87.335 102.755 88.085 103.275 ;
        RECT 88.255 102.585 89.005 103.105 ;
        RECT 90.770 102.680 91.120 103.930 ;
        RECT 94.755 103.225 94.965 104.365 ;
        RECT 95.135 103.215 95.465 104.195 ;
        RECT 95.635 103.225 95.865 104.365 ;
        RECT 96.075 103.275 99.585 104.365 ;
        RECT 85.950 102.365 86.700 102.535 ;
        RECT 85.945 101.815 86.275 102.195 ;
        RECT 86.445 102.075 86.700 102.365 ;
        RECT 86.875 101.815 87.165 102.540 ;
        RECT 87.335 101.815 89.005 102.585 ;
        RECT 92.600 102.360 92.940 103.190 ;
        RECT 89.180 101.815 94.525 102.360 ;
        RECT 94.755 101.815 94.965 102.635 ;
        RECT 95.135 102.615 95.385 103.215 ;
        RECT 95.555 102.805 95.885 103.055 ;
        RECT 96.075 102.755 97.765 103.275 ;
        RECT 99.755 103.200 100.045 104.365 ;
        RECT 100.215 103.275 101.425 104.365 ;
        RECT 101.600 103.930 106.945 104.365 ;
        RECT 107.120 103.930 112.465 104.365 ;
        RECT 95.135 101.985 95.465 102.615 ;
        RECT 95.635 101.815 95.865 102.635 ;
        RECT 97.935 102.585 99.585 103.105 ;
        RECT 100.215 102.735 100.735 103.275 ;
        RECT 96.075 101.815 99.585 102.585 ;
        RECT 100.905 102.565 101.425 103.105 ;
        RECT 103.190 102.680 103.540 103.930 ;
        RECT 99.755 101.815 100.045 102.540 ;
        RECT 100.215 101.815 101.425 102.565 ;
        RECT 105.020 102.360 105.360 103.190 ;
        RECT 108.710 102.680 109.060 103.930 ;
        RECT 112.635 103.200 112.925 104.365 ;
        RECT 113.095 103.275 116.605 104.365 ;
        RECT 110.540 102.360 110.880 103.190 ;
        RECT 113.095 102.755 114.785 103.275 ;
        RECT 116.815 103.225 117.045 104.365 ;
        RECT 117.215 103.215 117.545 104.195 ;
        RECT 117.715 103.225 117.925 104.365 ;
        RECT 119.080 103.930 124.425 104.365 ;
        RECT 114.955 102.585 116.605 103.105 ;
        RECT 116.795 102.805 117.125 103.055 ;
        RECT 101.600 101.815 106.945 102.360 ;
        RECT 107.120 101.815 112.465 102.360 ;
        RECT 112.635 101.815 112.925 102.540 ;
        RECT 113.095 101.815 116.605 102.585 ;
        RECT 116.815 101.815 117.045 102.635 ;
        RECT 117.295 102.615 117.545 103.215 ;
        RECT 120.670 102.680 121.020 103.930 ;
        RECT 124.595 103.275 125.805 104.365 ;
        RECT 117.215 101.985 117.545 102.615 ;
        RECT 117.715 101.815 117.925 102.635 ;
        RECT 122.500 102.360 122.840 103.190 ;
        RECT 124.595 102.735 125.115 103.275 ;
        RECT 125.285 102.565 125.805 103.105 ;
        RECT 119.080 101.815 124.425 102.360 ;
        RECT 124.595 101.815 125.805 102.565 ;
        RECT 11.810 101.645 125.890 101.815 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 11.010 215.730 125.890 216.210 ;
        RECT 11.810 213.010 125.890 213.490 ;
        RECT 11.010 210.290 125.890 210.770 ;
        RECT 11.810 207.570 125.890 208.050 ;
        RECT 11.010 204.850 125.890 205.330 ;
        RECT 11.810 202.130 125.890 202.610 ;
        RECT 11.010 199.410 125.890 199.890 ;
        RECT 64.435 198.870 64.725 198.915 ;
        RECT 65.240 198.870 65.560 198.930 ;
        RECT 67.675 198.870 68.325 198.915 ;
        RECT 64.435 198.730 68.325 198.870 ;
        RECT 64.435 198.685 65.025 198.730 ;
        RECT 64.735 198.370 65.025 198.685 ;
        RECT 65.240 198.670 65.560 198.730 ;
        RECT 67.675 198.685 68.325 198.730 ;
        RECT 65.815 198.530 66.105 198.575 ;
        RECT 69.395 198.530 69.685 198.575 ;
        RECT 71.230 198.530 71.520 198.575 ;
        RECT 65.815 198.390 71.520 198.530 ;
        RECT 65.815 198.345 66.105 198.390 ;
        RECT 69.395 198.345 69.685 198.390 ;
        RECT 71.230 198.345 71.520 198.390 ;
        RECT 71.680 197.990 72.000 198.250 ;
        RECT 65.815 197.850 66.105 197.895 ;
        RECT 68.935 197.850 69.225 197.895 ;
        RECT 70.825 197.850 71.115 197.895 ;
        RECT 65.815 197.710 71.115 197.850 ;
        RECT 65.815 197.665 66.105 197.710 ;
        RECT 68.935 197.665 69.225 197.710 ;
        RECT 70.825 197.665 71.115 197.710 ;
        RECT 62.955 197.510 63.245 197.555 ;
        RECT 64.780 197.510 65.100 197.570 ;
        RECT 62.955 197.370 65.100 197.510 ;
        RECT 62.955 197.325 63.245 197.370 ;
        RECT 64.780 197.310 65.100 197.370 ;
        RECT 70.410 197.510 70.700 197.555 ;
        RECT 71.220 197.510 71.540 197.570 ;
        RECT 70.410 197.370 71.540 197.510 ;
        RECT 70.410 197.325 70.700 197.370 ;
        RECT 71.220 197.310 71.540 197.370 ;
        RECT 11.810 196.690 125.890 197.170 ;
        RECT 65.240 196.490 65.560 196.550 ;
        RECT 69.395 196.490 69.685 196.535 ;
        RECT 65.240 196.350 69.685 196.490 ;
        RECT 65.240 196.290 65.560 196.350 ;
        RECT 69.395 196.305 69.685 196.350 ;
        RECT 78.210 196.350 84.330 196.490 ;
        RECT 59.225 196.150 59.515 196.195 ;
        RECT 61.115 196.150 61.405 196.195 ;
        RECT 64.235 196.150 64.525 196.195 ;
        RECT 59.225 196.010 64.525 196.150 ;
        RECT 59.225 195.965 59.515 196.010 ;
        RECT 61.115 195.965 61.405 196.010 ;
        RECT 64.235 195.965 64.525 196.010 ;
        RECT 71.680 196.150 72.000 196.210 ;
        RECT 78.210 196.150 78.350 196.350 ;
        RECT 71.680 196.010 78.350 196.150 ;
        RECT 78.695 196.150 78.985 196.195 ;
        RECT 81.815 196.150 82.105 196.195 ;
        RECT 83.705 196.150 83.995 196.195 ;
        RECT 78.695 196.010 83.995 196.150 ;
        RECT 71.680 195.950 72.000 196.010 ;
        RECT 78.695 195.965 78.985 196.010 ;
        RECT 81.815 195.965 82.105 196.010 ;
        RECT 83.705 195.965 83.995 196.010 ;
        RECT 62.940 195.810 63.260 195.870 ;
        RECT 79.500 195.810 79.820 195.870 ;
        RECT 83.195 195.810 83.485 195.855 ;
        RECT 62.940 195.670 66.620 195.810 ;
        RECT 62.940 195.610 63.260 195.670 ;
        RECT 57.420 195.470 57.740 195.530 ;
        RECT 58.355 195.470 58.645 195.515 ;
        RECT 57.420 195.330 58.645 195.470 ;
        RECT 57.420 195.270 57.740 195.330 ;
        RECT 58.355 195.285 58.645 195.330 ;
        RECT 58.820 195.470 59.110 195.515 ;
        RECT 60.655 195.470 60.945 195.515 ;
        RECT 64.235 195.470 64.525 195.515 ;
        RECT 58.820 195.330 64.525 195.470 ;
        RECT 58.820 195.285 59.110 195.330 ;
        RECT 60.655 195.285 60.945 195.330 ;
        RECT 64.235 195.285 64.525 195.330 ;
        RECT 59.720 194.930 60.040 195.190 ;
        RECT 62.015 195.130 62.665 195.175 ;
        RECT 63.400 195.130 63.720 195.190 ;
        RECT 65.315 195.175 65.605 195.490 ;
        RECT 66.480 195.470 66.620 195.670 ;
        RECT 79.500 195.670 83.485 195.810 ;
        RECT 84.190 195.810 84.330 196.350 ;
        RECT 84.560 195.810 84.880 195.870 ;
        RECT 84.190 195.670 84.880 195.810 ;
        RECT 79.500 195.610 79.820 195.670 ;
        RECT 83.195 195.625 83.485 195.670 ;
        RECT 84.560 195.610 84.880 195.670 ;
        RECT 69.855 195.470 70.145 195.515 ;
        RECT 74.455 195.470 74.745 195.515 ;
        RECT 66.480 195.330 74.745 195.470 ;
        RECT 69.855 195.285 70.145 195.330 ;
        RECT 74.455 195.285 74.745 195.330 ;
        RECT 65.315 195.130 65.905 195.175 ;
        RECT 62.015 194.990 65.905 195.130 ;
        RECT 62.015 194.945 62.665 194.990 ;
        RECT 63.400 194.930 63.720 194.990 ;
        RECT 65.615 194.945 65.905 194.990 ;
        RECT 68.475 194.945 68.765 195.175 ;
        RECT 74.530 195.130 74.670 195.285 ;
        RECT 77.615 195.175 77.905 195.490 ;
        RECT 78.695 195.470 78.985 195.515 ;
        RECT 82.275 195.470 82.565 195.515 ;
        RECT 84.110 195.470 84.400 195.515 ;
        RECT 78.695 195.330 84.400 195.470 ;
        RECT 78.695 195.285 78.985 195.330 ;
        RECT 82.275 195.285 82.565 195.330 ;
        RECT 84.110 195.285 84.400 195.330 ;
        RECT 80.880 195.175 81.200 195.190 ;
        RECT 77.315 195.130 77.905 195.175 ;
        RECT 80.555 195.130 81.205 195.175 ;
        RECT 74.530 194.990 76.970 195.130 ;
        RECT 68.550 194.790 68.690 194.945 ;
        RECT 69.840 194.790 70.160 194.850 ;
        RECT 68.550 194.650 70.160 194.790 ;
        RECT 69.840 194.590 70.160 194.650 ;
        RECT 74.915 194.790 75.205 194.835 ;
        RECT 75.360 194.790 75.680 194.850 ;
        RECT 74.915 194.650 75.680 194.790 ;
        RECT 74.915 194.605 75.205 194.650 ;
        RECT 75.360 194.590 75.680 194.650 ;
        RECT 75.820 194.590 76.140 194.850 ;
        RECT 76.830 194.790 76.970 194.990 ;
        RECT 77.315 194.990 81.205 195.130 ;
        RECT 77.315 194.945 77.605 194.990 ;
        RECT 80.555 194.945 81.205 194.990 ;
        RECT 80.880 194.930 81.200 194.945 ;
        RECT 85.020 194.790 85.340 194.850 ;
        RECT 76.830 194.650 85.340 194.790 ;
        RECT 85.020 194.590 85.340 194.650 ;
        RECT 11.010 193.970 125.890 194.450 ;
        RECT 63.400 193.770 63.720 193.830 ;
        RECT 63.875 193.770 64.165 193.815 ;
        RECT 63.400 193.630 64.165 193.770 ;
        RECT 63.400 193.570 63.720 193.630 ;
        RECT 63.875 193.585 64.165 193.630 ;
        RECT 71.220 193.770 71.540 193.830 ;
        RECT 71.695 193.770 71.985 193.815 ;
        RECT 71.220 193.630 71.985 193.770 ;
        RECT 71.220 193.570 71.540 193.630 ;
        RECT 71.695 193.585 71.985 193.630 ;
        RECT 80.880 193.770 81.200 193.830 ;
        RECT 84.575 193.770 84.865 193.815 ;
        RECT 80.880 193.630 84.865 193.770 ;
        RECT 80.880 193.570 81.200 193.630 ;
        RECT 84.575 193.585 84.865 193.630 ;
        RECT 75.360 193.430 75.680 193.490 ;
        RECT 76.395 193.430 76.685 193.475 ;
        RECT 79.635 193.430 80.285 193.475 ;
        RECT 75.360 193.290 80.285 193.430 ;
        RECT 75.360 193.230 75.680 193.290 ;
        RECT 76.395 193.245 76.985 193.290 ;
        RECT 79.635 193.245 80.285 193.290 ;
        RECT 98.015 193.430 98.305 193.475 ;
        RECT 98.820 193.430 99.140 193.490 ;
        RECT 101.255 193.430 101.905 193.475 ;
        RECT 98.015 193.290 101.905 193.430 ;
        RECT 98.015 193.245 98.605 193.290 ;
        RECT 62.940 193.090 63.260 193.150 ;
        RECT 63.415 193.090 63.705 193.135 ;
        RECT 62.940 192.950 63.705 193.090 ;
        RECT 62.940 192.890 63.260 192.950 ;
        RECT 63.415 192.905 63.705 192.950 ;
        RECT 64.780 193.090 65.100 193.150 ;
        RECT 65.715 193.090 66.005 193.135 ;
        RECT 64.780 192.950 66.005 193.090 ;
        RECT 64.780 192.890 65.100 192.950 ;
        RECT 65.715 192.905 66.005 192.950 ;
        RECT 67.080 193.090 67.400 193.150 ;
        RECT 68.935 193.090 69.225 193.135 ;
        RECT 67.080 192.950 69.225 193.090 ;
        RECT 67.080 192.890 67.400 192.950 ;
        RECT 68.935 192.905 69.225 192.950 ;
        RECT 69.840 192.890 70.160 193.150 ;
        RECT 73.535 192.905 73.825 193.135 ;
        RECT 76.695 192.930 76.985 193.245 ;
        RECT 77.775 193.090 78.065 193.135 ;
        RECT 81.355 193.090 81.645 193.135 ;
        RECT 83.190 193.090 83.480 193.135 ;
        RECT 77.775 192.950 83.480 193.090 ;
        RECT 77.775 192.905 78.065 192.950 ;
        RECT 81.355 192.905 81.645 192.950 ;
        RECT 83.190 192.905 83.480 192.950 ;
        RECT 83.655 193.090 83.945 193.135 ;
        RECT 84.560 193.090 84.880 193.150 ;
        RECT 83.655 192.950 84.880 193.090 ;
        RECT 83.655 192.905 83.945 192.950 ;
        RECT 68.475 192.565 68.765 192.795 ;
        RECT 66.635 192.410 66.925 192.455 ;
        RECT 68.550 192.410 68.690 192.565 ;
        RECT 69.380 192.550 69.700 192.810 ;
        RECT 69.840 192.410 70.160 192.470 ;
        RECT 73.610 192.410 73.750 192.905 ;
        RECT 84.560 192.890 84.880 192.950 ;
        RECT 85.020 193.090 85.340 193.150 ;
        RECT 91.000 193.090 91.320 193.150 ;
        RECT 85.020 192.950 91.320 193.090 ;
        RECT 85.020 192.890 85.340 192.950 ;
        RECT 91.000 192.890 91.320 192.950 ;
        RECT 98.315 192.930 98.605 193.245 ;
        RECT 98.820 193.230 99.140 193.290 ;
        RECT 101.255 193.245 101.905 193.290 ;
        RECT 103.420 193.430 103.740 193.490 ;
        RECT 103.420 193.290 105.950 193.430 ;
        RECT 103.420 193.230 103.740 193.290 ;
        RECT 105.810 193.135 105.950 193.290 ;
        RECT 99.395 193.090 99.685 193.135 ;
        RECT 102.975 193.090 103.265 193.135 ;
        RECT 104.810 193.090 105.100 193.135 ;
        RECT 99.395 192.950 105.100 193.090 ;
        RECT 99.395 192.905 99.685 192.950 ;
        RECT 102.975 192.905 103.265 192.950 ;
        RECT 104.810 192.905 105.100 192.950 ;
        RECT 105.735 192.905 106.025 193.135 ;
        RECT 107.560 192.890 107.880 193.150 ;
        RECT 73.980 192.550 74.300 192.810 ;
        RECT 81.800 192.750 82.120 192.810 ;
        RECT 82.275 192.750 82.565 192.795 ;
        RECT 81.800 192.610 82.565 192.750 ;
        RECT 81.800 192.550 82.120 192.610 ;
        RECT 82.275 192.565 82.565 192.610 ;
        RECT 103.880 192.550 104.200 192.810 ;
        RECT 105.275 192.750 105.565 192.795 ;
        RECT 109.860 192.750 110.180 192.810 ;
        RECT 105.275 192.610 110.180 192.750 ;
        RECT 105.275 192.565 105.565 192.610 ;
        RECT 109.860 192.550 110.180 192.610 ;
        RECT 66.635 192.270 73.750 192.410 ;
        RECT 77.775 192.410 78.065 192.455 ;
        RECT 80.895 192.410 81.185 192.455 ;
        RECT 82.785 192.410 83.075 192.455 ;
        RECT 77.775 192.270 83.075 192.410 ;
        RECT 66.635 192.225 66.925 192.270 ;
        RECT 69.840 192.210 70.160 192.270 ;
        RECT 77.775 192.225 78.065 192.270 ;
        RECT 80.895 192.225 81.185 192.270 ;
        RECT 82.785 192.225 83.075 192.270 ;
        RECT 99.395 192.410 99.685 192.455 ;
        RECT 102.515 192.410 102.805 192.455 ;
        RECT 104.405 192.410 104.695 192.455 ;
        RECT 99.395 192.270 104.695 192.410 ;
        RECT 99.395 192.225 99.685 192.270 ;
        RECT 102.515 192.225 102.805 192.270 ;
        RECT 104.405 192.225 104.695 192.270 ;
        RECT 67.540 191.870 67.860 192.130 ;
        RECT 72.140 192.070 72.460 192.130 ;
        RECT 74.915 192.070 75.205 192.115 ;
        RECT 72.140 191.930 75.205 192.070 ;
        RECT 72.140 191.870 72.460 191.930 ;
        RECT 74.915 191.885 75.205 191.930 ;
        RECT 96.535 192.070 96.825 192.115 ;
        RECT 100.200 192.070 100.520 192.130 ;
        RECT 96.535 191.930 100.520 192.070 ;
        RECT 96.535 191.885 96.825 191.930 ;
        RECT 100.200 191.870 100.520 191.930 ;
        RECT 106.180 191.870 106.500 192.130 ;
        RECT 108.495 192.070 108.785 192.115 ;
        RECT 109.400 192.070 109.720 192.130 ;
        RECT 108.495 191.930 109.720 192.070 ;
        RECT 108.495 191.885 108.785 191.930 ;
        RECT 109.400 191.870 109.720 191.930 ;
        RECT 11.810 191.250 125.890 191.730 ;
        RECT 68.935 191.050 69.225 191.095 ;
        RECT 70.760 191.050 71.080 191.110 ;
        RECT 68.935 190.910 71.080 191.050 ;
        RECT 68.935 190.865 69.225 190.910 ;
        RECT 70.760 190.850 71.080 190.910 ;
        RECT 79.500 190.850 79.820 191.110 ;
        RECT 81.355 191.050 81.645 191.095 ;
        RECT 81.800 191.050 82.120 191.110 ;
        RECT 81.355 190.910 82.120 191.050 ;
        RECT 81.355 190.865 81.645 190.910 ;
        RECT 81.800 190.850 82.120 190.910 ;
        RECT 98.820 190.850 99.140 191.110 ;
        RECT 109.860 191.050 110.180 191.110 ;
        RECT 109.860 190.910 111.470 191.050 ;
        RECT 109.860 190.850 110.180 190.910 ;
        RECT 65.255 190.710 65.545 190.755 ;
        RECT 69.380 190.710 69.700 190.770 ;
        RECT 65.255 190.570 69.700 190.710 ;
        RECT 65.255 190.525 65.545 190.570 ;
        RECT 69.380 190.510 69.700 190.570 ;
        RECT 69.840 190.510 70.160 190.770 ;
        RECT 105.375 190.710 105.665 190.755 ;
        RECT 108.495 190.710 108.785 190.755 ;
        RECT 110.385 190.710 110.675 190.755 ;
        RECT 105.375 190.570 110.675 190.710 ;
        RECT 105.375 190.525 105.665 190.570 ;
        RECT 108.495 190.525 108.785 190.570 ;
        RECT 110.385 190.525 110.675 190.570 ;
        RECT 65.700 190.170 66.020 190.430 ;
        RECT 68.140 190.370 68.430 190.415 ;
        RECT 72.140 190.370 72.460 190.430 ;
        RECT 103.420 190.370 103.740 190.430 ;
        RECT 68.090 190.230 72.460 190.370 ;
        RECT 68.090 190.185 68.430 190.230 ;
        RECT 64.780 190.030 65.100 190.090 ;
        RECT 67.095 190.030 67.385 190.075 ;
        RECT 64.780 189.890 67.385 190.030 ;
        RECT 64.780 189.830 65.100 189.890 ;
        RECT 67.095 189.845 67.385 189.890 ;
        RECT 64.335 189.690 64.625 189.735 ;
        RECT 68.090 189.690 68.230 190.185 ;
        RECT 72.140 190.170 72.460 190.230 ;
        RECT 91.090 190.230 103.740 190.370 ;
        RECT 91.090 190.090 91.230 190.230 ;
        RECT 69.380 190.030 69.700 190.090 ;
        RECT 71.220 190.030 71.540 190.090 ;
        RECT 75.360 190.030 75.680 190.090 ;
        RECT 69.380 189.890 75.680 190.030 ;
        RECT 69.380 189.830 69.700 189.890 ;
        RECT 71.220 189.830 71.540 189.890 ;
        RECT 75.360 189.830 75.680 189.890 ;
        RECT 76.280 190.030 76.600 190.090 ;
        RECT 78.135 190.030 78.425 190.075 ;
        RECT 79.055 190.030 79.345 190.075 ;
        RECT 76.280 189.890 79.345 190.030 ;
        RECT 76.280 189.830 76.600 189.890 ;
        RECT 78.135 189.845 78.425 189.890 ;
        RECT 79.055 189.845 79.345 189.890 ;
        RECT 80.420 189.830 80.740 190.090 ;
        RECT 91.000 189.830 91.320 190.090 ;
        RECT 91.920 190.030 92.240 190.090 ;
        RECT 98.450 190.075 98.590 190.230 ;
        RECT 103.420 190.170 103.740 190.230 ;
        RECT 109.400 190.370 109.720 190.430 ;
        RECT 111.330 190.415 111.470 190.910 ;
        RECT 109.875 190.370 110.165 190.415 ;
        RECT 109.400 190.230 110.165 190.370 ;
        RECT 109.400 190.170 109.720 190.230 ;
        RECT 109.875 190.185 110.165 190.230 ;
        RECT 111.255 190.370 111.545 190.415 ;
        RECT 114.000 190.370 114.320 190.430 ;
        RECT 111.255 190.230 114.320 190.370 ;
        RECT 111.255 190.185 111.545 190.230 ;
        RECT 114.000 190.170 114.320 190.230 ;
        RECT 92.395 190.030 92.685 190.075 ;
        RECT 91.920 189.890 92.685 190.030 ;
        RECT 91.920 189.830 92.240 189.890 ;
        RECT 92.395 189.845 92.685 189.890 ;
        RECT 98.375 189.845 98.665 190.075 ;
        RECT 64.335 189.550 68.230 189.690 ;
        RECT 69.855 189.690 70.145 189.735 ;
        RECT 70.300 189.690 70.620 189.750 ;
        RECT 75.820 189.690 76.140 189.750 ;
        RECT 104.295 189.735 104.585 190.050 ;
        RECT 105.375 190.030 105.665 190.075 ;
        RECT 108.955 190.030 109.245 190.075 ;
        RECT 110.790 190.030 111.080 190.075 ;
        RECT 105.375 189.890 111.080 190.030 ;
        RECT 105.375 189.845 105.665 189.890 ;
        RECT 108.955 189.845 109.245 189.890 ;
        RECT 110.790 189.845 111.080 189.890 ;
        RECT 77.215 189.690 77.505 189.735 ;
        RECT 69.855 189.550 70.620 189.690 ;
        RECT 64.335 189.505 64.625 189.550 ;
        RECT 69.855 189.505 70.145 189.550 ;
        RECT 70.300 189.490 70.620 189.550 ;
        RECT 72.690 189.550 77.505 189.690 ;
        RECT 72.690 189.395 72.830 189.550 ;
        RECT 75.820 189.490 76.140 189.550 ;
        RECT 77.215 189.505 77.505 189.550 ;
        RECT 103.995 189.690 104.585 189.735 ;
        RECT 106.180 189.690 106.500 189.750 ;
        RECT 107.235 189.690 107.885 189.735 ;
        RECT 103.995 189.550 107.885 189.690 ;
        RECT 103.995 189.505 104.285 189.550 ;
        RECT 106.180 189.490 106.500 189.550 ;
        RECT 107.235 189.505 107.885 189.550 ;
        RECT 67.555 189.350 67.845 189.395 ;
        RECT 72.615 189.350 72.905 189.395 ;
        RECT 67.555 189.210 72.905 189.350 ;
        RECT 67.555 189.165 67.845 189.210 ;
        RECT 72.615 189.165 72.905 189.210 ;
        RECT 73.520 189.150 73.840 189.410 ;
        RECT 74.440 189.150 74.760 189.410 ;
        RECT 90.555 189.350 90.845 189.395 ;
        RECT 91.000 189.350 91.320 189.410 ;
        RECT 90.555 189.210 91.320 189.350 ;
        RECT 90.555 189.165 90.845 189.210 ;
        RECT 91.000 189.150 91.320 189.210 ;
        RECT 93.300 189.150 93.620 189.410 ;
        RECT 102.500 189.150 102.820 189.410 ;
        RECT 11.010 188.530 125.890 189.010 ;
        RECT 59.720 188.330 60.040 188.390 ;
        RECT 67.540 188.375 67.860 188.390 ;
        RECT 65.255 188.330 65.545 188.375 ;
        RECT 38.650 188.190 50.750 188.330 ;
        RECT 32.120 187.650 32.440 187.710 ;
        RECT 38.650 187.695 38.790 188.190 ;
        RECT 39.035 187.990 39.325 188.035 ;
        RECT 41.435 187.990 41.725 188.035 ;
        RECT 44.675 187.990 45.325 188.035 ;
        RECT 39.035 187.850 45.325 187.990 ;
        RECT 39.035 187.805 39.325 187.850 ;
        RECT 41.435 187.805 42.025 187.850 ;
        RECT 44.675 187.805 45.325 187.850 ;
        RECT 50.610 187.990 50.750 188.190 ;
        RECT 59.720 188.190 65.545 188.330 ;
        RECT 59.720 188.130 60.040 188.190 ;
        RECT 65.255 188.145 65.545 188.190 ;
        RECT 66.635 188.145 66.925 188.375 ;
        RECT 67.475 188.145 67.860 188.375 ;
        RECT 70.300 188.330 70.620 188.390 ;
        RECT 50.610 187.850 54.890 187.990 ;
        RECT 38.575 187.650 38.865 187.695 ;
        RECT 32.120 187.510 38.865 187.650 ;
        RECT 32.120 187.450 32.440 187.510 ;
        RECT 38.575 187.465 38.865 187.510 ;
        RECT 41.735 187.490 42.025 187.805 ;
        RECT 50.610 187.695 50.750 187.850 ;
        RECT 42.815 187.650 43.105 187.695 ;
        RECT 46.395 187.650 46.685 187.695 ;
        RECT 48.230 187.650 48.520 187.695 ;
        RECT 42.815 187.510 48.520 187.650 ;
        RECT 42.815 187.465 43.105 187.510 ;
        RECT 46.395 187.465 46.685 187.510 ;
        RECT 48.230 187.465 48.520 187.510 ;
        RECT 50.535 187.465 50.825 187.695 ;
        RECT 50.980 187.650 51.300 187.710 ;
        RECT 54.750 187.695 54.890 187.850 ;
        RECT 52.375 187.650 52.665 187.695 ;
        RECT 50.980 187.510 52.665 187.650 ;
        RECT 50.980 187.450 51.300 187.510 ;
        RECT 52.375 187.465 52.665 187.510 ;
        RECT 54.675 187.465 54.965 187.695 ;
        RECT 66.175 187.650 66.465 187.695 ;
        RECT 66.710 187.650 66.850 188.145 ;
        RECT 67.540 188.130 67.860 188.145 ;
        RECT 68.090 188.190 70.620 188.330 ;
        RECT 66.175 187.510 66.850 187.650 ;
        RECT 68.090 187.650 68.230 188.190 ;
        RECT 70.300 188.130 70.620 188.190 ;
        RECT 71.695 188.330 71.985 188.375 ;
        RECT 74.075 188.330 74.365 188.375 ;
        RECT 71.695 188.190 74.365 188.330 ;
        RECT 71.695 188.145 71.985 188.190 ;
        RECT 74.075 188.145 74.365 188.190 ;
        RECT 74.915 188.330 75.205 188.375 ;
        RECT 80.420 188.330 80.740 188.390 ;
        RECT 74.915 188.190 80.740 188.330 ;
        RECT 74.915 188.145 75.205 188.190 ;
        RECT 68.475 187.990 68.765 188.035 ;
        RECT 71.770 187.990 71.910 188.145 ;
        RECT 80.420 188.130 80.740 188.190 ;
        RECT 87.335 188.330 87.625 188.375 ;
        RECT 89.620 188.330 89.940 188.390 ;
        RECT 106.195 188.330 106.485 188.375 ;
        RECT 107.560 188.330 107.880 188.390 ;
        RECT 87.335 188.190 95.370 188.330 ;
        RECT 87.335 188.145 87.625 188.190 ;
        RECT 89.620 188.130 89.940 188.190 ;
        RECT 68.475 187.850 71.910 187.990 ;
        RECT 73.075 187.990 73.365 188.035 ;
        RECT 75.835 187.990 76.125 188.035 ;
        RECT 73.075 187.850 76.125 187.990 ;
        RECT 68.475 187.805 68.765 187.850 ;
        RECT 73.075 187.805 73.365 187.850 ;
        RECT 74.070 187.710 74.210 187.850 ;
        RECT 75.835 187.805 76.125 187.850 ;
        RECT 88.815 187.990 89.105 188.035 ;
        RECT 91.000 187.990 91.320 188.050 ;
        RECT 92.055 187.990 92.705 188.035 ;
        RECT 88.815 187.850 92.705 187.990 ;
        RECT 88.815 187.805 89.405 187.850 ;
        RECT 68.935 187.650 69.225 187.695 ;
        RECT 73.520 187.650 73.840 187.710 ;
        RECT 68.090 187.510 73.840 187.650 ;
        RECT 66.175 187.465 66.465 187.510 ;
        RECT 47.300 187.110 47.620 187.370 ;
        RECT 48.695 187.310 48.985 187.355 ;
        RECT 57.420 187.310 57.740 187.370 ;
        RECT 48.695 187.170 57.740 187.310 ;
        RECT 48.695 187.125 48.985 187.170 ;
        RECT 57.420 187.110 57.740 187.170 ;
        RECT 65.700 187.310 66.020 187.370 ;
        RECT 68.090 187.310 68.230 187.510 ;
        RECT 68.935 187.465 69.225 187.510 ;
        RECT 73.520 187.450 73.840 187.510 ;
        RECT 73.980 187.450 74.300 187.710 ;
        RECT 75.360 187.450 75.680 187.710 ;
        RECT 76.280 187.450 76.600 187.710 ;
        RECT 89.115 187.490 89.405 187.805 ;
        RECT 91.000 187.790 91.320 187.850 ;
        RECT 92.055 187.805 92.705 187.850 ;
        RECT 93.300 187.990 93.620 188.050 ;
        RECT 94.695 187.990 94.985 188.035 ;
        RECT 93.300 187.850 94.985 187.990 ;
        RECT 95.230 187.990 95.370 188.190 ;
        RECT 106.195 188.190 107.880 188.330 ;
        RECT 106.195 188.145 106.485 188.190 ;
        RECT 107.560 188.130 107.880 188.190 ;
        RECT 100.215 187.990 100.505 188.035 ;
        RECT 104.355 187.990 104.645 188.035 ;
        RECT 95.230 187.850 100.505 187.990 ;
        RECT 93.300 187.790 93.620 187.850 ;
        RECT 94.695 187.805 94.985 187.850 ;
        RECT 100.215 187.805 100.505 187.850 ;
        RECT 101.670 187.850 104.645 187.990 ;
        RECT 90.195 187.650 90.485 187.695 ;
        RECT 93.775 187.650 94.065 187.695 ;
        RECT 95.610 187.650 95.900 187.695 ;
        RECT 90.195 187.510 95.900 187.650 ;
        RECT 90.195 187.465 90.485 187.510 ;
        RECT 93.775 187.465 94.065 187.510 ;
        RECT 95.610 187.465 95.900 187.510 ;
        RECT 101.670 187.370 101.810 187.850 ;
        RECT 104.355 187.805 104.645 187.850 ;
        RECT 102.500 187.650 102.820 187.710 ;
        RECT 102.500 187.510 104.110 187.650 ;
        RECT 102.500 187.450 102.820 187.510 ;
        RECT 65.700 187.170 68.230 187.310 ;
        RECT 65.700 187.110 66.020 187.170 ;
        RECT 69.840 187.110 70.160 187.370 ;
        RECT 70.300 187.110 70.620 187.370 ;
        RECT 87.780 187.310 88.100 187.370 ;
        RECT 96.075 187.310 96.365 187.355 ;
        RECT 98.835 187.310 99.125 187.355 ;
        RECT 87.780 187.170 96.365 187.310 ;
        RECT 87.780 187.110 88.100 187.170 ;
        RECT 96.075 187.125 96.365 187.170 ;
        RECT 96.610 187.170 99.125 187.310 ;
        RECT 42.815 186.970 43.105 187.015 ;
        RECT 45.935 186.970 46.225 187.015 ;
        RECT 47.825 186.970 48.115 187.015 ;
        RECT 42.815 186.830 48.115 186.970 ;
        RECT 69.930 186.970 70.070 187.110 ;
        RECT 90.195 186.970 90.485 187.015 ;
        RECT 93.315 186.970 93.605 187.015 ;
        RECT 95.205 186.970 95.495 187.015 ;
        RECT 69.930 186.830 70.530 186.970 ;
        RECT 42.815 186.785 43.105 186.830 ;
        RECT 45.935 186.785 46.225 186.830 ;
        RECT 47.825 186.785 48.115 186.830 ;
        RECT 39.955 186.630 40.245 186.675 ;
        RECT 43.620 186.630 43.940 186.690 ;
        RECT 39.955 186.490 43.940 186.630 ;
        RECT 39.955 186.445 40.245 186.490 ;
        RECT 43.620 186.430 43.940 186.490 ;
        RECT 50.980 186.430 51.300 186.690 ;
        RECT 53.280 186.430 53.600 186.690 ;
        RECT 54.215 186.630 54.505 186.675 ;
        RECT 55.580 186.630 55.900 186.690 ;
        RECT 54.215 186.490 55.900 186.630 ;
        RECT 54.215 186.445 54.505 186.490 ;
        RECT 55.580 186.430 55.900 186.490 ;
        RECT 67.555 186.630 67.845 186.675 ;
        RECT 69.840 186.630 70.160 186.690 ;
        RECT 70.390 186.675 70.530 186.830 ;
        RECT 90.195 186.830 95.495 186.970 ;
        RECT 90.195 186.785 90.485 186.830 ;
        RECT 93.315 186.785 93.605 186.830 ;
        RECT 95.205 186.785 95.495 186.830 ;
        RECT 67.555 186.490 70.160 186.630 ;
        RECT 67.555 186.445 67.845 186.490 ;
        RECT 69.840 186.430 70.160 186.490 ;
        RECT 70.315 186.630 70.605 186.675 ;
        RECT 72.600 186.630 72.920 186.690 ;
        RECT 70.315 186.490 72.920 186.630 ;
        RECT 70.315 186.445 70.605 186.490 ;
        RECT 72.600 186.430 72.920 186.490 ;
        RECT 73.995 186.630 74.285 186.675 ;
        RECT 74.440 186.630 74.760 186.690 ;
        RECT 73.995 186.490 74.760 186.630 ;
        RECT 73.995 186.445 74.285 186.490 ;
        RECT 74.440 186.430 74.760 186.490 ;
        RECT 89.160 186.630 89.480 186.690 ;
        RECT 96.610 186.630 96.750 187.170 ;
        RECT 98.835 187.125 99.125 187.170 ;
        RECT 99.755 187.310 100.045 187.355 ;
        RECT 100.200 187.310 100.520 187.370 ;
        RECT 101.580 187.310 101.900 187.370 ;
        RECT 103.970 187.355 104.110 187.510 ;
        RECT 109.860 187.450 110.180 187.710 ;
        RECT 99.755 187.170 101.900 187.310 ;
        RECT 99.755 187.125 100.045 187.170 ;
        RECT 98.910 186.970 99.050 187.125 ;
        RECT 100.200 187.110 100.520 187.170 ;
        RECT 101.580 187.110 101.900 187.170 ;
        RECT 103.435 187.125 103.725 187.355 ;
        RECT 103.895 187.310 104.185 187.355 ;
        RECT 106.180 187.310 106.500 187.370 ;
        RECT 103.895 187.170 106.500 187.310 ;
        RECT 103.895 187.125 104.185 187.170 ;
        RECT 98.910 186.830 102.730 186.970 ;
        RECT 89.160 186.490 96.750 186.630 ;
        RECT 89.160 186.430 89.480 186.490 ;
        RECT 102.040 186.430 102.360 186.690 ;
        RECT 102.590 186.630 102.730 186.830 ;
        RECT 103.510 186.630 103.650 187.125 ;
        RECT 106.180 187.110 106.500 187.170 ;
        RECT 104.340 186.630 104.660 186.690 ;
        RECT 102.590 186.490 104.660 186.630 ;
        RECT 104.340 186.430 104.660 186.490 ;
        RECT 110.795 186.630 111.085 186.675 ;
        RECT 112.620 186.630 112.940 186.690 ;
        RECT 110.795 186.490 112.940 186.630 ;
        RECT 110.795 186.445 111.085 186.490 ;
        RECT 112.620 186.430 112.940 186.490 ;
        RECT 11.810 185.810 125.890 186.290 ;
        RECT 68.475 185.425 68.765 185.655 ;
        RECT 70.300 185.610 70.620 185.670 ;
        RECT 70.775 185.610 71.065 185.655 ;
        RECT 70.300 185.470 71.065 185.610 ;
        RECT 34.845 185.270 35.135 185.315 ;
        RECT 36.735 185.270 37.025 185.315 ;
        RECT 39.855 185.270 40.145 185.315 ;
        RECT 34.845 185.130 40.145 185.270 ;
        RECT 34.845 185.085 35.135 185.130 ;
        RECT 36.735 185.085 37.025 185.130 ;
        RECT 39.855 185.085 40.145 185.130 ;
        RECT 51.555 185.270 51.845 185.315 ;
        RECT 54.675 185.270 54.965 185.315 ;
        RECT 56.565 185.270 56.855 185.315 ;
        RECT 68.550 185.270 68.690 185.425 ;
        RECT 70.300 185.410 70.620 185.470 ;
        RECT 70.775 185.425 71.065 185.470 ;
        RECT 91.920 185.410 92.240 185.670 ;
        RECT 103.435 185.610 103.725 185.655 ;
        RECT 103.880 185.610 104.200 185.670 ;
        RECT 103.435 185.470 104.200 185.610 ;
        RECT 103.435 185.425 103.725 185.470 ;
        RECT 103.880 185.410 104.200 185.470 ;
        RECT 51.555 185.130 56.855 185.270 ;
        RECT 51.555 185.085 51.845 185.130 ;
        RECT 54.675 185.085 54.965 185.130 ;
        RECT 56.565 185.085 56.855 185.130 ;
        RECT 66.480 185.130 68.690 185.270 ;
        RECT 69.840 185.270 70.160 185.330 ;
        RECT 71.695 185.270 71.985 185.315 ;
        RECT 72.140 185.270 72.460 185.330 ;
        RECT 94.680 185.270 95.000 185.330 ;
        RECT 69.840 185.130 72.460 185.270 ;
        RECT 66.480 184.990 66.620 185.130 ;
        RECT 69.840 185.070 70.160 185.130 ;
        RECT 71.695 185.085 71.985 185.130 ;
        RECT 72.140 185.070 72.460 185.130 ;
        RECT 85.110 185.130 95.000 185.270 ;
        RECT 35.340 184.730 35.660 184.990 ;
        RECT 43.620 184.930 43.940 184.990 ;
        RECT 46.395 184.930 46.685 184.975 ;
        RECT 43.620 184.790 46.685 184.930 ;
        RECT 43.620 184.730 43.940 184.790 ;
        RECT 46.395 184.745 46.685 184.790 ;
        RECT 47.315 184.930 47.605 184.975 ;
        RECT 47.760 184.930 48.080 184.990 ;
        RECT 47.315 184.790 48.080 184.930 ;
        RECT 47.315 184.745 47.605 184.790 ;
        RECT 47.760 184.730 48.080 184.790 ;
        RECT 53.280 184.930 53.600 184.990 ;
        RECT 56.055 184.930 56.345 184.975 ;
        RECT 53.280 184.790 56.345 184.930 ;
        RECT 53.280 184.730 53.600 184.790 ;
        RECT 56.055 184.745 56.345 184.790 ;
        RECT 63.875 184.930 64.165 184.975 ;
        RECT 66.160 184.930 66.620 184.990 ;
        RECT 63.875 184.790 66.620 184.930 ;
        RECT 69.395 184.930 69.685 184.975 ;
        RECT 71.220 184.930 71.540 184.990 ;
        RECT 69.395 184.790 71.540 184.930 ;
        RECT 63.875 184.745 64.165 184.790 ;
        RECT 66.160 184.730 66.480 184.790 ;
        RECT 69.395 184.745 69.685 184.790 ;
        RECT 71.220 184.730 71.540 184.790 ;
        RECT 82.720 184.930 83.040 184.990 ;
        RECT 84.575 184.930 84.865 184.975 ;
        RECT 82.720 184.790 84.865 184.930 ;
        RECT 82.720 184.730 83.040 184.790 ;
        RECT 84.575 184.745 84.865 184.790 ;
        RECT 32.120 184.590 32.440 184.650 ;
        RECT 32.595 184.590 32.885 184.635 ;
        RECT 32.120 184.450 32.885 184.590 ;
        RECT 32.120 184.390 32.440 184.450 ;
        RECT 32.595 184.405 32.885 184.450 ;
        RECT 33.055 184.590 33.345 184.635 ;
        RECT 33.055 184.450 33.730 184.590 ;
        RECT 33.055 184.405 33.345 184.450 ;
        RECT 33.590 184.250 33.730 184.450 ;
        RECT 33.960 184.390 34.280 184.650 ;
        RECT 34.440 184.590 34.730 184.635 ;
        RECT 36.275 184.590 36.565 184.635 ;
        RECT 39.855 184.590 40.145 184.635 ;
        RECT 34.440 184.450 40.145 184.590 ;
        RECT 34.440 184.405 34.730 184.450 ;
        RECT 36.275 184.405 36.565 184.450 ;
        RECT 39.855 184.405 40.145 184.450 ;
        RECT 40.935 184.295 41.225 184.610 ;
        RECT 50.475 184.590 50.765 184.610 ;
        RECT 50.980 184.590 51.300 184.650 ;
        RECT 50.475 184.450 51.300 184.590 ;
        RECT 50.475 184.295 50.765 184.450 ;
        RECT 50.980 184.390 51.300 184.450 ;
        RECT 51.555 184.590 51.845 184.635 ;
        RECT 55.135 184.590 55.425 184.635 ;
        RECT 56.970 184.590 57.260 184.635 ;
        RECT 51.555 184.450 57.260 184.590 ;
        RECT 51.555 184.405 51.845 184.450 ;
        RECT 55.135 184.405 55.425 184.450 ;
        RECT 56.970 184.405 57.260 184.450 ;
        RECT 57.420 184.590 57.740 184.650 ;
        RECT 60.640 184.590 60.960 184.650 ;
        RECT 57.420 184.450 60.960 184.590 ;
        RECT 57.420 184.390 57.740 184.450 ;
        RECT 60.640 184.390 60.960 184.450 ;
        RECT 62.480 184.390 62.800 184.650 ;
        RECT 62.940 184.390 63.260 184.650 ;
        RECT 67.080 184.590 67.400 184.650 ;
        RECT 68.015 184.590 68.305 184.635 ;
        RECT 67.080 184.450 68.305 184.590 ;
        RECT 67.080 184.390 67.400 184.450 ;
        RECT 68.015 184.405 68.305 184.450 ;
        RECT 37.635 184.250 38.285 184.295 ;
        RECT 40.935 184.250 41.525 184.295 ;
        RECT 45.935 184.250 46.225 184.295 ;
        RECT 33.590 184.110 41.525 184.250 ;
        RECT 37.635 184.065 38.285 184.110 ;
        RECT 41.235 184.065 41.525 184.110 ;
        RECT 42.330 184.110 46.225 184.250 ;
        RECT 38.560 183.910 38.880 183.970 ;
        RECT 42.330 183.910 42.470 184.110 ;
        RECT 45.935 184.065 46.225 184.110 ;
        RECT 50.175 184.250 50.765 184.295 ;
        RECT 53.415 184.250 54.065 184.295 ;
        RECT 50.175 184.110 54.065 184.250 ;
        RECT 68.090 184.250 68.230 184.405 ;
        RECT 72.600 184.390 72.920 184.650 ;
        RECT 73.075 184.590 73.365 184.635 ;
        RECT 73.520 184.590 73.840 184.650 ;
        RECT 85.110 184.635 85.250 185.130 ;
        RECT 94.680 185.070 95.000 185.130 ;
        RECT 108.135 185.270 108.425 185.315 ;
        RECT 111.255 185.270 111.545 185.315 ;
        RECT 113.145 185.270 113.435 185.315 ;
        RECT 108.135 185.130 113.435 185.270 ;
        RECT 108.135 185.085 108.425 185.130 ;
        RECT 111.255 185.085 111.545 185.130 ;
        RECT 113.145 185.085 113.435 185.130 ;
        RECT 89.160 184.730 89.480 184.990 ;
        RECT 89.620 184.730 89.940 184.990 ;
        RECT 112.620 184.730 112.940 184.990 ;
        RECT 114.000 184.730 114.320 184.990 ;
        RECT 73.075 184.450 73.840 184.590 ;
        RECT 73.075 184.405 73.365 184.450 ;
        RECT 73.520 184.390 73.840 184.450 ;
        RECT 83.195 184.590 83.485 184.635 ;
        RECT 85.035 184.590 85.325 184.635 ;
        RECT 83.195 184.450 85.325 184.590 ;
        RECT 83.195 184.405 83.485 184.450 ;
        RECT 85.035 184.405 85.325 184.450 ;
        RECT 102.040 184.590 102.360 184.650 ;
        RECT 102.515 184.590 102.805 184.635 ;
        RECT 102.040 184.450 102.805 184.590 ;
        RECT 102.040 184.390 102.360 184.450 ;
        RECT 102.515 184.405 102.805 184.450 ;
        RECT 103.420 184.590 103.740 184.650 ;
        RECT 103.895 184.590 104.185 184.635 ;
        RECT 103.420 184.450 104.185 184.590 ;
        RECT 103.420 184.390 103.740 184.450 ;
        RECT 103.895 184.405 104.185 184.450 ;
        RECT 104.355 184.590 104.645 184.635 ;
        RECT 107.055 184.590 107.345 184.610 ;
        RECT 104.355 184.450 107.345 184.590 ;
        RECT 104.355 184.405 104.645 184.450 ;
        RECT 75.820 184.250 76.140 184.310 ;
        RECT 107.055 184.295 107.345 184.450 ;
        RECT 108.135 184.590 108.425 184.635 ;
        RECT 111.715 184.590 112.005 184.635 ;
        RECT 113.550 184.590 113.840 184.635 ;
        RECT 108.135 184.450 113.840 184.590 ;
        RECT 108.135 184.405 108.425 184.450 ;
        RECT 111.715 184.405 112.005 184.450 ;
        RECT 113.550 184.405 113.840 184.450 ;
        RECT 90.095 184.250 90.385 184.295 ;
        RECT 68.090 184.110 72.370 184.250 ;
        RECT 50.175 184.065 50.465 184.110 ;
        RECT 53.415 184.065 54.065 184.110 ;
        RECT 38.560 183.770 42.470 183.910 ;
        RECT 38.560 183.710 38.880 183.770 ;
        RECT 42.700 183.710 43.020 183.970 ;
        RECT 44.095 183.910 44.385 183.955 ;
        RECT 45.460 183.910 45.780 183.970 ;
        RECT 44.095 183.770 45.780 183.910 ;
        RECT 46.010 183.910 46.150 184.065 ;
        RECT 48.220 183.910 48.540 183.970 ;
        RECT 48.695 183.910 48.985 183.955 ;
        RECT 46.010 183.770 48.985 183.910 ;
        RECT 44.095 183.725 44.385 183.770 ;
        RECT 45.460 183.710 45.780 183.770 ;
        RECT 48.220 183.710 48.540 183.770 ;
        RECT 48.695 183.725 48.985 183.770 ;
        RECT 66.635 183.910 66.925 183.955 ;
        RECT 71.220 183.910 71.540 183.970 ;
        RECT 72.230 183.955 72.370 184.110 ;
        RECT 75.820 184.110 90.385 184.250 ;
        RECT 75.820 184.050 76.140 184.110 ;
        RECT 90.095 184.065 90.385 184.110 ;
        RECT 106.755 184.250 107.345 184.295 ;
        RECT 109.995 184.250 110.645 184.295 ;
        RECT 106.755 184.110 110.645 184.250 ;
        RECT 106.755 184.065 107.045 184.110 ;
        RECT 109.995 184.065 110.645 184.110 ;
        RECT 66.635 183.770 71.540 183.910 ;
        RECT 66.635 183.725 66.925 183.770 ;
        RECT 71.220 183.710 71.540 183.770 ;
        RECT 72.155 183.910 72.445 183.955 ;
        RECT 73.060 183.910 73.380 183.970 ;
        RECT 76.280 183.910 76.600 183.970 ;
        RECT 72.155 183.770 76.600 183.910 ;
        RECT 72.155 183.725 72.445 183.770 ;
        RECT 73.060 183.710 73.380 183.770 ;
        RECT 76.280 183.710 76.600 183.770 ;
        RECT 81.800 183.910 82.120 183.970 ;
        RECT 82.735 183.910 83.025 183.955 ;
        RECT 81.800 183.770 83.025 183.910 ;
        RECT 81.800 183.710 82.120 183.770 ;
        RECT 82.735 183.725 83.025 183.770 ;
        RECT 105.260 183.710 105.580 183.970 ;
        RECT 11.010 183.090 125.890 183.570 ;
        RECT 35.340 182.890 35.660 182.950 ;
        RECT 39.495 182.890 39.785 182.935 ;
        RECT 35.340 182.750 39.785 182.890 ;
        RECT 35.340 182.690 35.660 182.750 ;
        RECT 39.495 182.705 39.785 182.750 ;
        RECT 46.395 182.890 46.685 182.935 ;
        RECT 47.300 182.890 47.620 182.950 ;
        RECT 46.395 182.750 47.620 182.890 ;
        RECT 46.395 182.705 46.685 182.750 ;
        RECT 47.300 182.690 47.620 182.750 ;
        RECT 48.220 182.690 48.540 182.950 ;
        RECT 50.520 182.690 50.840 182.950 ;
        RECT 70.775 182.890 71.065 182.935 ;
        RECT 69.010 182.750 71.065 182.890 ;
        RECT 42.715 182.550 43.005 182.595 ;
        RECT 43.620 182.550 43.940 182.610 ;
        RECT 55.580 182.595 55.900 182.610 ;
        RECT 42.715 182.410 43.940 182.550 ;
        RECT 42.715 182.365 43.005 182.410 ;
        RECT 43.620 182.350 43.940 182.410 ;
        RECT 52.475 182.550 52.765 182.595 ;
        RECT 55.580 182.550 56.365 182.595 ;
        RECT 52.475 182.410 56.365 182.550 ;
        RECT 52.475 182.365 53.065 182.410 ;
        RECT 40.415 182.210 40.705 182.255 ;
        RECT 40.415 182.070 41.090 182.210 ;
        RECT 40.415 182.025 40.705 182.070 ;
        RECT 40.950 181.575 41.090 182.070 ;
        RECT 45.460 182.010 45.780 182.270 ;
        RECT 47.300 182.210 47.620 182.270 ;
        RECT 48.695 182.210 48.985 182.255 ;
        RECT 47.300 182.070 51.210 182.210 ;
        RECT 47.300 182.010 47.620 182.070 ;
        RECT 48.695 182.025 48.985 182.070 ;
        RECT 41.320 181.870 41.640 181.930 ;
        RECT 42.700 181.870 43.020 181.930 ;
        RECT 43.175 181.870 43.465 181.915 ;
        RECT 41.320 181.730 43.465 181.870 ;
        RECT 41.320 181.670 41.640 181.730 ;
        RECT 42.700 181.670 43.020 181.730 ;
        RECT 43.175 181.685 43.465 181.730 ;
        RECT 44.095 181.870 44.385 181.915 ;
        RECT 47.760 181.870 48.080 181.930 ;
        RECT 51.070 181.915 51.210 182.070 ;
        RECT 52.775 182.050 53.065 182.365 ;
        RECT 55.580 182.365 56.365 182.410 ;
        RECT 62.480 182.550 62.800 182.610 ;
        RECT 69.010 182.595 69.150 182.750 ;
        RECT 70.775 182.705 71.065 182.750 ;
        RECT 87.335 182.705 87.625 182.935 ;
        RECT 109.860 182.890 110.180 182.950 ;
        RECT 111.255 182.890 111.545 182.935 ;
        RECT 109.860 182.750 111.545 182.890 ;
        RECT 63.055 182.550 63.345 182.595 ;
        RECT 66.295 182.550 66.945 182.595 ;
        RECT 62.480 182.410 66.945 182.550 ;
        RECT 55.580 182.350 55.900 182.365 ;
        RECT 62.480 182.350 62.800 182.410 ;
        RECT 63.055 182.365 63.645 182.410 ;
        RECT 66.295 182.365 66.945 182.410 ;
        RECT 68.935 182.365 69.225 182.595 ;
        RECT 71.220 182.550 71.540 182.610 ;
        RECT 82.720 182.595 83.040 182.610 ;
        RECT 79.450 182.550 79.740 182.595 ;
        RECT 82.710 182.550 83.040 182.595 ;
        RECT 71.220 182.410 72.830 182.550 ;
        RECT 53.855 182.210 54.145 182.255 ;
        RECT 57.435 182.210 57.725 182.255 ;
        RECT 59.270 182.210 59.560 182.255 ;
        RECT 53.855 182.070 59.560 182.210 ;
        RECT 53.855 182.025 54.145 182.070 ;
        RECT 57.435 182.025 57.725 182.070 ;
        RECT 59.270 182.025 59.560 182.070 ;
        RECT 63.355 182.050 63.645 182.365 ;
        RECT 71.220 182.350 71.540 182.410 ;
        RECT 64.435 182.210 64.725 182.255 ;
        RECT 68.015 182.210 68.305 182.255 ;
        RECT 69.850 182.210 70.140 182.255 ;
        RECT 64.435 182.070 70.140 182.210 ;
        RECT 64.435 182.025 64.725 182.070 ;
        RECT 68.015 182.025 68.305 182.070 ;
        RECT 69.850 182.025 70.140 182.070 ;
        RECT 70.315 182.210 70.605 182.255 ;
        RECT 71.680 182.210 72.000 182.270 ;
        RECT 72.690 182.255 72.830 182.410 ;
        RECT 79.450 182.410 83.040 182.550 ;
        RECT 79.450 182.365 79.740 182.410 ;
        RECT 82.710 182.365 83.040 182.410 ;
        RECT 82.720 182.350 83.040 182.365 ;
        RECT 83.630 182.550 83.920 182.595 ;
        RECT 85.490 182.550 85.780 182.595 ;
        RECT 83.630 182.410 85.780 182.550 ;
        RECT 83.630 182.365 83.920 182.410 ;
        RECT 85.490 182.365 85.780 182.410 ;
        RECT 70.315 182.070 72.000 182.210 ;
        RECT 70.315 182.025 70.605 182.070 ;
        RECT 71.680 182.010 72.000 182.070 ;
        RECT 72.615 182.025 72.905 182.255 ;
        RECT 81.310 182.210 81.600 182.255 ;
        RECT 83.630 182.210 83.845 182.365 ;
        RECT 81.310 182.070 83.845 182.210 ;
        RECT 84.575 182.210 84.865 182.255 ;
        RECT 87.410 182.210 87.550 182.705 ;
        RECT 109.860 182.690 110.180 182.750 ;
        RECT 111.255 182.705 111.545 182.750 ;
        RECT 106.180 182.550 106.500 182.610 ;
        RECT 109.415 182.550 109.705 182.595 ;
        RECT 106.180 182.410 109.705 182.550 ;
        RECT 106.180 182.350 106.500 182.410 ;
        RECT 109.415 182.365 109.705 182.410 ;
        RECT 84.575 182.070 87.550 182.210 ;
        RECT 81.310 182.025 81.600 182.070 ;
        RECT 84.575 182.025 84.865 182.070 ;
        RECT 88.255 182.025 88.545 182.255 ;
        RECT 94.680 182.210 95.000 182.270 ;
        RECT 98.375 182.210 98.665 182.255 ;
        RECT 94.680 182.070 98.665 182.210 ;
        RECT 44.095 181.730 48.080 181.870 ;
        RECT 44.095 181.685 44.385 181.730 ;
        RECT 47.760 181.670 48.080 181.730 ;
        RECT 50.995 181.685 51.285 181.915 ;
        RECT 58.340 181.670 58.660 181.930 ;
        RECT 59.735 181.870 60.025 181.915 ;
        RECT 60.640 181.870 60.960 181.930 ;
        RECT 59.735 181.730 60.960 181.870 ;
        RECT 59.735 181.685 60.025 181.730 ;
        RECT 60.640 181.670 60.960 181.730 ;
        RECT 40.875 181.345 41.165 181.575 ;
        RECT 53.855 181.530 54.145 181.575 ;
        RECT 56.975 181.530 57.265 181.575 ;
        RECT 58.865 181.530 59.155 181.575 ;
        RECT 53.855 181.390 59.155 181.530 ;
        RECT 53.855 181.345 54.145 181.390 ;
        RECT 56.975 181.345 57.265 181.390 ;
        RECT 58.865 181.345 59.155 181.390 ;
        RECT 64.435 181.530 64.725 181.575 ;
        RECT 67.555 181.530 67.845 181.575 ;
        RECT 69.445 181.530 69.735 181.575 ;
        RECT 64.435 181.390 69.735 181.530 ;
        RECT 71.770 181.530 71.910 182.010 ;
        RECT 72.140 181.670 72.460 181.930 ;
        RECT 86.415 181.870 86.705 181.915 ;
        RECT 87.780 181.870 88.100 181.930 ;
        RECT 80.970 181.730 88.100 181.870 ;
        RECT 80.970 181.530 81.110 181.730 ;
        RECT 86.415 181.685 86.705 181.730 ;
        RECT 87.780 181.670 88.100 181.730 ;
        RECT 71.770 181.390 81.110 181.530 ;
        RECT 81.310 181.530 81.600 181.575 ;
        RECT 84.090 181.530 84.380 181.575 ;
        RECT 85.950 181.530 86.240 181.575 ;
        RECT 81.310 181.390 86.240 181.530 ;
        RECT 64.435 181.345 64.725 181.390 ;
        RECT 67.555 181.345 67.845 181.390 ;
        RECT 69.445 181.345 69.735 181.390 ;
        RECT 81.310 181.345 81.600 181.390 ;
        RECT 84.090 181.345 84.380 181.390 ;
        RECT 85.950 181.345 86.240 181.390 ;
        RECT 61.575 181.190 61.865 181.235 ;
        RECT 66.160 181.190 66.480 181.250 ;
        RECT 61.575 181.050 66.480 181.190 ;
        RECT 61.575 181.005 61.865 181.050 ;
        RECT 66.160 180.990 66.480 181.050 ;
        RECT 67.080 181.190 67.400 181.250 ;
        RECT 75.820 181.190 76.140 181.250 ;
        RECT 77.445 181.190 77.735 181.235 ;
        RECT 67.080 181.050 77.735 181.190 ;
        RECT 67.080 180.990 67.400 181.050 ;
        RECT 75.820 180.990 76.140 181.050 ;
        RECT 77.445 181.005 77.735 181.050 ;
        RECT 78.120 181.190 78.440 181.250 ;
        RECT 88.330 181.190 88.470 182.025 ;
        RECT 94.680 182.010 95.000 182.070 ;
        RECT 98.375 182.025 98.665 182.070 ;
        RECT 102.055 182.210 102.345 182.255 ;
        RECT 103.420 182.210 103.740 182.270 ;
        RECT 102.055 182.070 103.740 182.210 ;
        RECT 102.055 182.025 102.345 182.070 ;
        RECT 103.420 182.010 103.740 182.070 ;
        RECT 105.260 182.210 105.580 182.270 ;
        RECT 107.560 182.210 107.880 182.270 ;
        RECT 108.955 182.210 109.245 182.255 ;
        RECT 105.260 182.070 109.245 182.210 ;
        RECT 105.260 182.010 105.580 182.070 ;
        RECT 107.560 182.010 107.880 182.070 ;
        RECT 108.955 182.025 109.245 182.070 ;
        RECT 104.340 181.670 104.660 181.930 ;
        RECT 104.815 181.870 105.105 181.915 ;
        RECT 106.640 181.870 106.960 181.930 ;
        RECT 104.815 181.730 106.960 181.870 ;
        RECT 104.815 181.685 105.105 181.730 ;
        RECT 106.640 181.670 106.960 181.730 ;
        RECT 108.035 181.685 108.325 181.915 ;
        RECT 104.430 181.530 104.570 181.670 ;
        RECT 108.110 181.530 108.250 181.685 ;
        RECT 104.430 181.390 108.250 181.530 ;
        RECT 78.120 181.050 88.470 181.190 ;
        RECT 97.440 181.190 97.760 181.250 ;
        RECT 97.915 181.190 98.205 181.235 ;
        RECT 97.440 181.050 98.205 181.190 ;
        RECT 78.120 180.990 78.440 181.050 ;
        RECT 97.440 180.990 97.760 181.050 ;
        RECT 97.915 181.005 98.205 181.050 ;
        RECT 102.500 180.990 102.820 181.250 ;
        RECT 107.100 180.990 107.420 181.250 ;
        RECT 11.810 180.370 125.890 180.850 ;
        RECT 57.435 180.170 57.725 180.215 ;
        RECT 58.340 180.170 58.660 180.230 ;
        RECT 57.435 180.030 58.660 180.170 ;
        RECT 57.435 179.985 57.725 180.030 ;
        RECT 58.340 179.970 58.660 180.030 ;
        RECT 78.120 179.970 78.440 180.230 ;
        RECT 82.690 179.830 82.980 179.875 ;
        RECT 85.470 179.830 85.760 179.875 ;
        RECT 87.330 179.830 87.620 179.875 ;
        RECT 82.690 179.690 87.620 179.830 ;
        RECT 82.690 179.645 82.980 179.690 ;
        RECT 85.470 179.645 85.760 179.690 ;
        RECT 87.330 179.645 87.620 179.690 ;
        RECT 91.425 179.830 91.715 179.875 ;
        RECT 93.315 179.830 93.605 179.875 ;
        RECT 96.435 179.830 96.725 179.875 ;
        RECT 91.425 179.690 96.725 179.830 ;
        RECT 91.425 179.645 91.715 179.690 ;
        RECT 93.315 179.645 93.605 179.690 ;
        RECT 96.435 179.645 96.725 179.690 ;
        RECT 106.295 179.830 106.585 179.875 ;
        RECT 109.415 179.830 109.705 179.875 ;
        RECT 111.305 179.830 111.595 179.875 ;
        RECT 106.295 179.690 111.595 179.830 ;
        RECT 106.295 179.645 106.585 179.690 ;
        RECT 109.415 179.645 109.705 179.690 ;
        RECT 111.305 179.645 111.595 179.690 ;
        RECT 43.635 179.490 43.925 179.535 ;
        RECT 47.760 179.490 48.080 179.550 ;
        RECT 52.835 179.490 53.125 179.535 ;
        RECT 58.340 179.490 58.660 179.550 ;
        RECT 43.635 179.350 58.660 179.490 ;
        RECT 43.635 179.305 43.925 179.350 ;
        RECT 47.760 179.290 48.080 179.350 ;
        RECT 52.835 179.305 53.125 179.350 ;
        RECT 58.340 179.290 58.660 179.350 ;
        RECT 62.940 179.490 63.260 179.550 ;
        RECT 67.095 179.490 67.385 179.535 ;
        RECT 62.940 179.350 67.385 179.490 ;
        RECT 62.940 179.290 63.260 179.350 ;
        RECT 67.095 179.305 67.385 179.350 ;
        RECT 75.375 179.305 75.665 179.535 ;
        RECT 39.495 179.150 39.785 179.195 ;
        RECT 41.320 179.150 41.640 179.210 ;
        RECT 39.495 179.010 41.640 179.150 ;
        RECT 39.495 178.965 39.785 179.010 ;
        RECT 41.320 178.950 41.640 179.010 ;
        RECT 42.255 179.150 42.545 179.195 ;
        RECT 44.555 179.150 44.845 179.195 ;
        RECT 42.255 179.010 44.845 179.150 ;
        RECT 42.255 178.965 42.545 179.010 ;
        RECT 44.555 178.965 44.845 179.010 ;
        RECT 47.300 179.150 47.620 179.210 ;
        RECT 53.295 179.150 53.585 179.195 ;
        RECT 56.515 179.150 56.805 179.195 ;
        RECT 47.300 179.010 53.585 179.150 ;
        RECT 47.300 178.950 47.620 179.010 ;
        RECT 53.295 178.965 53.585 179.010 ;
        RECT 55.670 179.010 56.805 179.150 ;
        RECT 44.095 178.470 44.385 178.515 ;
        RECT 45.460 178.470 45.780 178.530 ;
        RECT 44.095 178.330 45.780 178.470 ;
        RECT 44.095 178.285 44.385 178.330 ;
        RECT 45.460 178.270 45.780 178.330 ;
        RECT 45.920 178.470 46.240 178.530 ;
        RECT 46.395 178.470 46.685 178.515 ;
        RECT 45.920 178.330 46.685 178.470 ;
        RECT 45.920 178.270 46.240 178.330 ;
        RECT 46.395 178.285 46.685 178.330 ;
        RECT 53.280 178.470 53.600 178.530 ;
        RECT 55.670 178.515 55.810 179.010 ;
        RECT 56.515 178.965 56.805 179.010 ;
        RECT 64.320 179.150 64.640 179.210 ;
        RECT 66.175 179.150 66.465 179.195 ;
        RECT 64.320 179.010 66.465 179.150 ;
        RECT 75.450 179.150 75.590 179.305 ;
        RECT 75.820 179.290 76.140 179.550 ;
        RECT 87.780 179.490 88.100 179.550 ;
        RECT 90.555 179.490 90.845 179.535 ;
        RECT 87.780 179.350 90.845 179.490 ;
        RECT 87.780 179.290 88.100 179.350 ;
        RECT 90.555 179.305 90.845 179.350 ;
        RECT 91.935 179.490 92.225 179.535 ;
        RECT 98.360 179.490 98.680 179.550 ;
        RECT 91.935 179.350 98.680 179.490 ;
        RECT 91.935 179.305 92.225 179.350 ;
        RECT 98.360 179.290 98.680 179.350 ;
        RECT 112.175 179.490 112.465 179.535 ;
        RECT 114.000 179.490 114.320 179.550 ;
        RECT 112.175 179.350 114.320 179.490 ;
        RECT 112.175 179.305 112.465 179.350 ;
        RECT 114.000 179.290 114.320 179.350 ;
        RECT 82.690 179.150 82.980 179.195 ;
        RECT 85.955 179.150 86.245 179.195 ;
        RECT 86.400 179.150 86.720 179.210 ;
        RECT 75.450 179.010 76.050 179.150 ;
        RECT 64.320 178.950 64.640 179.010 ;
        RECT 66.175 178.965 66.465 179.010 ;
        RECT 75.910 178.870 76.050 179.010 ;
        RECT 82.690 179.010 85.225 179.150 ;
        RECT 82.690 178.965 82.980 179.010 ;
        RECT 75.820 178.610 76.140 178.870 ;
        RECT 80.830 178.810 81.120 178.855 ;
        RECT 81.800 178.810 82.120 178.870 ;
        RECT 85.010 178.855 85.225 179.010 ;
        RECT 85.955 179.010 86.720 179.150 ;
        RECT 85.955 178.965 86.245 179.010 ;
        RECT 86.400 178.950 86.720 179.010 ;
        RECT 91.020 179.150 91.310 179.195 ;
        RECT 92.855 179.150 93.145 179.195 ;
        RECT 96.435 179.150 96.725 179.195 ;
        RECT 91.020 179.010 96.725 179.150 ;
        RECT 91.020 178.965 91.310 179.010 ;
        RECT 92.855 178.965 93.145 179.010 ;
        RECT 96.435 178.965 96.725 179.010 ;
        RECT 97.440 179.170 97.760 179.210 ;
        RECT 97.440 178.950 97.805 179.170 ;
        RECT 97.515 178.855 97.805 178.950 ;
        RECT 84.090 178.810 84.380 178.855 ;
        RECT 80.830 178.670 84.380 178.810 ;
        RECT 80.830 178.625 81.120 178.670 ;
        RECT 81.800 178.610 82.120 178.670 ;
        RECT 84.090 178.625 84.380 178.670 ;
        RECT 85.010 178.810 85.300 178.855 ;
        RECT 86.870 178.810 87.160 178.855 ;
        RECT 85.010 178.670 87.160 178.810 ;
        RECT 85.010 178.625 85.300 178.670 ;
        RECT 86.870 178.625 87.160 178.670 ;
        RECT 94.215 178.810 94.865 178.855 ;
        RECT 97.515 178.810 98.105 178.855 ;
        RECT 94.215 178.670 98.105 178.810 ;
        RECT 94.215 178.625 94.865 178.670 ;
        RECT 97.815 178.625 98.105 178.670 ;
        RECT 102.500 178.810 102.820 178.870 ;
        RECT 105.215 178.855 105.505 179.170 ;
        RECT 106.295 179.150 106.585 179.195 ;
        RECT 109.875 179.150 110.165 179.195 ;
        RECT 111.710 179.150 112.000 179.195 ;
        RECT 106.295 179.010 112.000 179.150 ;
        RECT 106.295 178.965 106.585 179.010 ;
        RECT 109.875 178.965 110.165 179.010 ;
        RECT 111.710 178.965 112.000 179.010 ;
        RECT 104.915 178.810 105.505 178.855 ;
        RECT 108.155 178.810 108.805 178.855 ;
        RECT 102.500 178.670 108.805 178.810 ;
        RECT 102.500 178.610 102.820 178.670 ;
        RECT 104.915 178.625 105.205 178.670 ;
        RECT 108.155 178.625 108.805 178.670 ;
        RECT 109.400 178.810 109.720 178.870 ;
        RECT 110.795 178.810 111.085 178.855 ;
        RECT 109.400 178.670 111.085 178.810 ;
        RECT 109.400 178.610 109.720 178.670 ;
        RECT 110.795 178.625 111.085 178.670 ;
        RECT 53.755 178.470 54.045 178.515 ;
        RECT 53.280 178.330 54.045 178.470 ;
        RECT 53.280 178.270 53.600 178.330 ;
        RECT 53.755 178.285 54.045 178.330 ;
        RECT 55.595 178.285 55.885 178.515 ;
        RECT 76.295 178.470 76.585 178.515 ;
        RECT 78.120 178.470 78.440 178.530 ;
        RECT 78.825 178.470 79.115 178.515 ;
        RECT 76.295 178.330 79.115 178.470 ;
        RECT 76.295 178.285 76.585 178.330 ;
        RECT 78.120 178.270 78.440 178.330 ;
        RECT 78.825 178.285 79.115 178.330 ;
        RECT 99.295 178.470 99.585 178.515 ;
        RECT 100.660 178.470 100.980 178.530 ;
        RECT 99.295 178.330 100.980 178.470 ;
        RECT 99.295 178.285 99.585 178.330 ;
        RECT 100.660 178.270 100.980 178.330 ;
        RECT 103.435 178.470 103.725 178.515 ;
        RECT 106.640 178.470 106.960 178.530 ;
        RECT 103.435 178.330 106.960 178.470 ;
        RECT 103.435 178.285 103.725 178.330 ;
        RECT 106.640 178.270 106.960 178.330 ;
        RECT 11.010 177.650 125.890 178.130 ;
        RECT 39.495 177.450 39.785 177.495 ;
        RECT 45.460 177.450 45.780 177.510 ;
        RECT 73.520 177.450 73.840 177.510 ;
        RECT 39.495 177.310 45.780 177.450 ;
        RECT 39.495 177.265 39.785 177.310 ;
        RECT 45.460 177.250 45.780 177.310 ;
        RECT 69.930 177.310 73.840 177.450 ;
        RECT 38.575 177.110 38.865 177.155 ;
        RECT 40.975 177.110 41.265 177.155 ;
        RECT 44.215 177.110 44.865 177.155 ;
        RECT 38.575 176.970 44.865 177.110 ;
        RECT 38.575 176.925 38.865 176.970 ;
        RECT 40.975 176.925 41.565 176.970 ;
        RECT 44.215 176.925 44.865 176.970 ;
        RECT 30.295 176.770 30.585 176.815 ;
        RECT 32.120 176.770 32.440 176.830 ;
        RECT 36.720 176.770 37.040 176.830 ;
        RECT 38.115 176.770 38.405 176.815 ;
        RECT 30.295 176.630 38.405 176.770 ;
        RECT 30.295 176.585 30.585 176.630 ;
        RECT 32.120 176.570 32.440 176.630 ;
        RECT 36.720 176.570 37.040 176.630 ;
        RECT 38.115 176.585 38.405 176.630 ;
        RECT 41.275 176.610 41.565 176.925 ;
        RECT 42.355 176.770 42.645 176.815 ;
        RECT 45.935 176.770 46.225 176.815 ;
        RECT 47.770 176.770 48.060 176.815 ;
        RECT 42.355 176.630 48.060 176.770 ;
        RECT 42.355 176.585 42.645 176.630 ;
        RECT 45.935 176.585 46.225 176.630 ;
        RECT 47.770 176.585 48.060 176.630 ;
        RECT 56.040 176.770 56.360 176.830 ;
        RECT 56.515 176.770 56.805 176.815 ;
        RECT 56.040 176.630 56.805 176.770 ;
        RECT 56.040 176.570 56.360 176.630 ;
        RECT 56.515 176.585 56.805 176.630 ;
        RECT 67.540 176.770 67.860 176.830 ;
        RECT 69.930 176.770 70.070 177.310 ;
        RECT 73.520 177.250 73.840 177.310 ;
        RECT 86.400 177.250 86.720 177.510 ;
        RECT 94.220 177.450 94.540 177.510 ;
        RECT 88.790 177.310 94.540 177.450 ;
        RECT 73.060 177.110 73.380 177.170 ;
        RECT 75.360 177.110 75.680 177.170 ;
        RECT 76.280 177.110 76.600 177.170 ;
        RECT 71.770 176.970 73.380 177.110 ;
        RECT 71.770 176.815 71.910 176.970 ;
        RECT 73.060 176.910 73.380 176.970 ;
        RECT 73.610 176.970 76.600 177.110 ;
        RECT 70.775 176.770 71.065 176.815 ;
        RECT 67.540 176.630 71.065 176.770 ;
        RECT 67.540 176.570 67.860 176.630 ;
        RECT 70.775 176.585 71.065 176.630 ;
        RECT 71.695 176.585 71.985 176.815 ;
        RECT 72.140 176.770 72.460 176.830 ;
        RECT 73.610 176.770 73.750 176.970 ;
        RECT 75.360 176.910 75.680 176.970 ;
        RECT 76.280 176.910 76.600 176.970 ;
        RECT 78.120 177.110 78.440 177.170 ;
        RECT 78.595 177.110 78.885 177.155 ;
        RECT 82.735 177.110 83.025 177.155 ;
        RECT 78.120 176.970 78.885 177.110 ;
        RECT 78.120 176.910 78.440 176.970 ;
        RECT 78.595 176.925 78.885 176.970 ;
        RECT 79.590 176.970 83.025 177.110 ;
        RECT 79.590 176.830 79.730 176.970 ;
        RECT 82.735 176.925 83.025 176.970 ;
        RECT 83.195 177.110 83.485 177.155 ;
        RECT 84.560 177.110 84.880 177.170 ;
        RECT 83.195 176.970 84.880 177.110 ;
        RECT 83.195 176.925 83.485 176.970 ;
        RECT 84.560 176.910 84.880 176.970 ;
        RECT 72.140 176.630 73.750 176.770 ;
        RECT 72.140 176.570 72.460 176.630 ;
        RECT 74.455 176.585 74.745 176.815 ;
        RECT 79.055 176.770 79.345 176.815 ;
        RECT 79.500 176.770 79.820 176.830 ;
        RECT 88.790 176.815 88.930 177.310 ;
        RECT 94.220 177.250 94.540 177.310 ;
        RECT 109.400 177.250 109.720 177.510 ;
        RECT 89.175 177.110 89.465 177.155 ;
        RECT 91.575 177.110 91.865 177.155 ;
        RECT 94.815 177.110 95.465 177.155 ;
        RECT 89.175 176.970 95.465 177.110 ;
        RECT 89.175 176.925 89.465 176.970 ;
        RECT 91.575 176.925 92.165 176.970 ;
        RECT 94.815 176.925 95.465 176.970 ;
        RECT 85.495 176.770 85.785 176.815 ;
        RECT 88.715 176.770 89.005 176.815 ;
        RECT 79.055 176.630 79.820 176.770 ;
        RECT 79.055 176.585 79.345 176.630 ;
        RECT 46.840 176.230 47.160 176.490 ;
        RECT 48.235 176.430 48.525 176.475 ;
        RECT 60.640 176.430 60.960 176.490 ;
        RECT 48.235 176.290 60.960 176.430 ;
        RECT 48.235 176.245 48.525 176.290 ;
        RECT 60.640 176.230 60.960 176.290 ;
        RECT 71.235 176.430 71.525 176.475 ;
        RECT 72.600 176.430 72.920 176.490 ;
        RECT 71.235 176.290 72.920 176.430 ;
        RECT 71.235 176.245 71.525 176.290 ;
        RECT 72.600 176.230 72.920 176.290 ;
        RECT 42.355 176.090 42.645 176.135 ;
        RECT 45.475 176.090 45.765 176.135 ;
        RECT 47.365 176.090 47.655 176.135 ;
        RECT 42.355 175.950 47.655 176.090 ;
        RECT 42.355 175.905 42.645 175.950 ;
        RECT 45.475 175.905 45.765 175.950 ;
        RECT 47.365 175.905 47.655 175.950 ;
        RECT 64.320 176.090 64.640 176.150 ;
        RECT 74.530 176.090 74.670 176.585 ;
        RECT 79.500 176.570 79.820 176.630 ;
        RECT 80.970 176.630 85.785 176.770 ;
        RECT 75.375 176.245 75.665 176.475 ;
        RECT 75.820 176.430 76.140 176.490 ;
        RECT 77.675 176.430 77.965 176.475 ;
        RECT 75.820 176.290 77.965 176.430 ;
        RECT 64.320 175.950 74.670 176.090 ;
        RECT 75.450 176.090 75.590 176.245 ;
        RECT 75.820 176.230 76.140 176.290 ;
        RECT 77.675 176.245 77.965 176.290 ;
        RECT 77.200 176.090 77.520 176.150 ;
        RECT 75.450 175.950 77.520 176.090 ;
        RECT 64.320 175.890 64.640 175.950 ;
        RECT 77.200 175.890 77.520 175.950 ;
        RECT 30.280 175.750 30.600 175.810 ;
        RECT 30.755 175.750 31.045 175.795 ;
        RECT 30.280 175.610 31.045 175.750 ;
        RECT 30.280 175.550 30.600 175.610 ;
        RECT 30.755 175.565 31.045 175.610 ;
        RECT 56.055 175.750 56.345 175.795 ;
        RECT 56.500 175.750 56.820 175.810 ;
        RECT 56.055 175.610 56.820 175.750 ;
        RECT 56.055 175.565 56.345 175.610 ;
        RECT 56.500 175.550 56.820 175.610 ;
        RECT 69.855 175.750 70.145 175.795 ;
        RECT 70.300 175.750 70.620 175.810 ;
        RECT 69.855 175.610 70.620 175.750 ;
        RECT 77.750 175.750 77.890 176.245 ;
        RECT 80.970 176.135 81.110 176.630 ;
        RECT 85.495 176.585 85.785 176.630 ;
        RECT 86.030 176.630 89.005 176.770 ;
        RECT 81.815 176.430 82.105 176.475 ;
        RECT 81.430 176.290 82.105 176.430 ;
        RECT 80.895 175.905 81.185 176.135 ;
        RECT 79.960 175.750 80.280 175.810 ;
        RECT 81.430 175.750 81.570 176.290 ;
        RECT 81.815 176.245 82.105 176.290 ;
        RECT 84.100 176.430 84.420 176.490 ;
        RECT 86.030 176.430 86.170 176.630 ;
        RECT 88.715 176.585 89.005 176.630 ;
        RECT 91.875 176.610 92.165 176.925 ;
        RECT 97.440 176.910 97.760 177.170 ;
        RECT 101.135 177.110 101.425 177.155 ;
        RECT 103.435 177.110 103.725 177.155 ;
        RECT 101.135 176.970 103.725 177.110 ;
        RECT 101.135 176.925 101.425 176.970 ;
        RECT 103.435 176.925 103.725 176.970 ;
        RECT 115.495 177.110 115.785 177.155 ;
        RECT 118.735 177.110 119.385 177.155 ;
        RECT 115.495 176.970 119.385 177.110 ;
        RECT 115.495 176.925 116.085 176.970 ;
        RECT 118.735 176.925 119.385 176.970 ;
        RECT 119.980 177.110 120.300 177.170 ;
        RECT 121.375 177.110 121.665 177.155 ;
        RECT 119.980 176.970 121.665 177.110 ;
        RECT 92.955 176.770 93.245 176.815 ;
        RECT 96.535 176.770 96.825 176.815 ;
        RECT 98.370 176.770 98.660 176.815 ;
        RECT 92.955 176.630 98.660 176.770 ;
        RECT 92.955 176.585 93.245 176.630 ;
        RECT 96.535 176.585 96.825 176.630 ;
        RECT 98.370 176.585 98.660 176.630 ;
        RECT 107.100 176.770 107.420 176.830 ;
        RECT 108.495 176.770 108.785 176.815 ;
        RECT 107.100 176.630 108.785 176.770 ;
        RECT 107.100 176.570 107.420 176.630 ;
        RECT 108.495 176.585 108.785 176.630 ;
        RECT 110.320 176.770 110.640 176.830 ;
        RECT 111.255 176.770 111.545 176.815 ;
        RECT 110.320 176.630 111.545 176.770 ;
        RECT 110.320 176.570 110.640 176.630 ;
        RECT 111.255 176.585 111.545 176.630 ;
        RECT 114.920 176.770 115.240 176.830 ;
        RECT 115.795 176.770 116.085 176.925 ;
        RECT 119.980 176.910 120.300 176.970 ;
        RECT 121.375 176.925 121.665 176.970 ;
        RECT 114.920 176.630 116.085 176.770 ;
        RECT 114.920 176.570 115.240 176.630 ;
        RECT 115.795 176.610 116.085 176.630 ;
        RECT 116.875 176.770 117.165 176.815 ;
        RECT 120.455 176.770 120.745 176.815 ;
        RECT 122.290 176.770 122.580 176.815 ;
        RECT 116.875 176.630 122.580 176.770 ;
        RECT 116.875 176.585 117.165 176.630 ;
        RECT 120.455 176.585 120.745 176.630 ;
        RECT 122.290 176.585 122.580 176.630 ;
        RECT 84.100 176.290 86.170 176.430 ;
        RECT 88.240 176.430 88.560 176.490 ;
        RECT 98.835 176.430 99.125 176.475 ;
        RECT 88.240 176.290 99.125 176.430 ;
        RECT 84.100 176.230 84.420 176.290 ;
        RECT 88.240 176.230 88.560 176.290 ;
        RECT 98.835 176.245 99.125 176.290 ;
        RECT 99.755 176.245 100.045 176.475 ;
        RECT 100.675 176.430 100.965 176.475 ;
        RECT 101.120 176.430 101.440 176.490 ;
        RECT 100.675 176.290 101.440 176.430 ;
        RECT 100.675 176.245 100.965 176.290 ;
        RECT 84.560 176.090 84.880 176.150 ;
        RECT 90.095 176.090 90.385 176.135 ;
        RECT 84.560 175.950 90.385 176.090 ;
        RECT 84.560 175.890 84.880 175.950 ;
        RECT 90.095 175.905 90.385 175.950 ;
        RECT 92.955 176.090 93.245 176.135 ;
        RECT 96.075 176.090 96.365 176.135 ;
        RECT 97.965 176.090 98.255 176.135 ;
        RECT 92.955 175.950 98.255 176.090 ;
        RECT 92.955 175.905 93.245 175.950 ;
        RECT 96.075 175.905 96.365 175.950 ;
        RECT 97.965 175.905 98.255 175.950 ;
        RECT 77.750 175.610 81.570 175.750 ;
        RECT 69.855 175.565 70.145 175.610 ;
        RECT 70.300 175.550 70.620 175.610 ;
        RECT 79.960 175.550 80.280 175.610 ;
        RECT 85.020 175.550 85.340 175.810 ;
        RECT 89.160 175.750 89.480 175.810 ;
        RECT 99.830 175.750 99.970 176.245 ;
        RECT 101.120 176.230 101.440 176.290 ;
        RECT 106.640 176.230 106.960 176.490 ;
        RECT 114.000 176.430 114.320 176.490 ;
        RECT 121.360 176.430 121.680 176.490 ;
        RECT 122.755 176.430 123.045 176.475 ;
        RECT 114.000 176.290 123.045 176.430 ;
        RECT 114.000 176.230 114.320 176.290 ;
        RECT 121.360 176.230 121.680 176.290 ;
        RECT 122.755 176.245 123.045 176.290 ;
        RECT 116.875 176.090 117.165 176.135 ;
        RECT 119.995 176.090 120.285 176.135 ;
        RECT 121.885 176.090 122.175 176.135 ;
        RECT 116.875 175.950 122.175 176.090 ;
        RECT 116.875 175.905 117.165 175.950 ;
        RECT 119.995 175.905 120.285 175.950 ;
        RECT 121.885 175.905 122.175 175.950 ;
        RECT 89.160 175.610 99.970 175.750 ;
        RECT 89.160 175.550 89.480 175.610 ;
        RECT 102.960 175.550 103.280 175.810 ;
        RECT 111.715 175.750 112.005 175.795 ;
        RECT 112.620 175.750 112.940 175.810 ;
        RECT 111.715 175.610 112.940 175.750 ;
        RECT 111.715 175.565 112.005 175.610 ;
        RECT 112.620 175.550 112.940 175.610 ;
        RECT 114.015 175.750 114.305 175.795 ;
        RECT 114.460 175.750 114.780 175.810 ;
        RECT 114.015 175.610 114.780 175.750 ;
        RECT 114.015 175.565 114.305 175.610 ;
        RECT 114.460 175.550 114.780 175.610 ;
        RECT 11.810 174.930 125.890 175.410 ;
        RECT 46.840 174.530 47.160 174.790 ;
        RECT 73.520 174.530 73.840 174.790 ;
        RECT 73.980 174.730 74.300 174.790 ;
        RECT 77.200 174.730 77.520 174.790 ;
        RECT 84.100 174.730 84.420 174.790 ;
        RECT 73.980 174.590 75.590 174.730 ;
        RECT 73.980 174.530 74.300 174.590 ;
        RECT 30.855 174.390 31.145 174.435 ;
        RECT 33.975 174.390 34.265 174.435 ;
        RECT 35.865 174.390 36.155 174.435 ;
        RECT 30.855 174.250 36.155 174.390 ;
        RECT 30.855 174.205 31.145 174.250 ;
        RECT 33.975 174.205 34.265 174.250 ;
        RECT 35.865 174.205 36.155 174.250 ;
        RECT 37.195 174.205 37.485 174.435 ;
        RECT 56.010 174.390 56.300 174.435 ;
        RECT 58.790 174.390 59.080 174.435 ;
        RECT 60.650 174.390 60.940 174.435 ;
        RECT 56.010 174.250 60.940 174.390 ;
        RECT 56.010 174.205 56.300 174.250 ;
        RECT 58.790 174.205 59.080 174.250 ;
        RECT 60.650 174.205 60.940 174.250 ;
        RECT 61.560 174.390 61.880 174.450 ;
        RECT 66.175 174.390 66.465 174.435 ;
        RECT 61.560 174.250 66.465 174.390 ;
        RECT 32.120 174.050 32.440 174.110 ;
        RECT 25.310 173.910 32.440 174.050 ;
        RECT 23.380 173.710 23.700 173.770 ;
        RECT 25.310 173.755 25.450 173.910 ;
        RECT 32.120 173.850 32.440 173.910 ;
        RECT 35.355 174.050 35.645 174.095 ;
        RECT 37.270 174.050 37.410 174.205 ;
        RECT 61.560 174.190 61.880 174.250 ;
        RECT 66.175 174.205 66.465 174.250 ;
        RECT 69.855 174.390 70.145 174.435 ;
        RECT 73.060 174.390 73.380 174.450 ;
        RECT 69.855 174.250 73.380 174.390 ;
        RECT 69.855 174.205 70.145 174.250 ;
        RECT 73.060 174.190 73.380 174.250 ;
        RECT 35.355 173.910 37.410 174.050 ;
        RECT 35.355 173.865 35.645 173.910 ;
        RECT 55.580 173.850 55.900 174.110 ;
        RECT 67.540 173.850 67.860 174.110 ;
        RECT 68.015 174.050 68.305 174.095 ;
        RECT 71.220 174.050 71.540 174.110 ;
        RECT 72.140 174.050 72.460 174.110 ;
        RECT 75.450 174.095 75.590 174.590 ;
        RECT 77.200 174.590 84.420 174.730 ;
        RECT 77.200 174.530 77.520 174.590 ;
        RECT 84.100 174.530 84.420 174.590 ;
        RECT 84.560 174.730 84.880 174.790 ;
        RECT 97.440 174.730 97.760 174.790 ;
        RECT 97.915 174.730 98.205 174.775 ;
        RECT 84.560 174.590 93.990 174.730 ;
        RECT 84.560 174.530 84.880 174.590 ;
        RECT 82.375 174.390 82.665 174.435 ;
        RECT 85.495 174.390 85.785 174.435 ;
        RECT 87.385 174.390 87.675 174.435 ;
        RECT 89.160 174.390 89.480 174.450 ;
        RECT 93.850 174.390 93.990 174.590 ;
        RECT 97.440 174.590 98.205 174.730 ;
        RECT 97.440 174.530 97.760 174.590 ;
        RECT 97.915 174.545 98.205 174.590 ;
        RECT 98.360 174.730 98.680 174.790 ;
        RECT 103.435 174.730 103.725 174.775 ;
        RECT 98.360 174.590 103.725 174.730 ;
        RECT 98.360 174.530 98.680 174.590 ;
        RECT 103.435 174.545 103.725 174.590 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 111.715 174.390 112.005 174.435 ;
        RECT 114.920 174.390 115.240 174.450 ;
        RECT 82.375 174.250 87.675 174.390 ;
        RECT 82.375 174.205 82.665 174.250 ;
        RECT 85.495 174.205 85.785 174.250 ;
        RECT 87.385 174.205 87.675 174.250 ;
        RECT 87.870 174.250 93.530 174.390 ;
        RECT 93.850 174.250 94.450 174.390 ;
        RECT 72.615 174.050 72.905 174.095 ;
        RECT 68.015 173.910 72.905 174.050 ;
        RECT 68.015 173.865 68.305 173.910 ;
        RECT 71.220 173.850 71.540 173.910 ;
        RECT 72.140 173.850 72.460 173.910 ;
        RECT 72.615 173.865 72.905 173.910 ;
        RECT 75.375 173.865 75.665 174.095 ;
        RECT 76.280 173.850 76.600 174.110 ;
        RECT 79.960 174.050 80.280 174.110 ;
        RECT 87.870 174.050 88.010 174.250 ;
        RECT 89.160 174.190 89.480 174.250 ;
        RECT 79.960 173.910 88.010 174.050 ;
        RECT 79.960 173.850 80.280 173.910 ;
        RECT 88.240 173.850 88.560 174.110 ;
        RECT 93.390 174.095 93.530 174.250 ;
        RECT 94.310 174.095 94.450 174.250 ;
        RECT 111.715 174.250 115.240 174.390 ;
        RECT 111.715 174.205 112.005 174.250 ;
        RECT 114.920 174.190 115.240 174.250 ;
        RECT 115.495 174.390 115.785 174.435 ;
        RECT 118.615 174.390 118.905 174.435 ;
        RECT 120.505 174.390 120.795 174.435 ;
        RECT 115.495 174.250 120.795 174.390 ;
        RECT 115.495 174.205 115.785 174.250 ;
        RECT 118.615 174.205 118.905 174.250 ;
        RECT 120.505 174.205 120.795 174.250 ;
        RECT 93.315 173.865 93.605 174.095 ;
        RECT 94.235 173.865 94.525 174.095 ;
        RECT 101.120 174.050 101.440 174.110 ;
        RECT 94.770 173.910 101.440 174.050 ;
        RECT 23.855 173.710 24.145 173.755 ;
        RECT 25.235 173.710 25.525 173.755 ;
        RECT 23.380 173.570 25.525 173.710 ;
        RECT 23.380 173.510 23.700 173.570 ;
        RECT 23.855 173.525 24.145 173.570 ;
        RECT 25.235 173.525 25.525 173.570 ;
        RECT 26.615 173.525 26.905 173.755 ;
        RECT 22.000 173.370 22.320 173.430 ;
        RECT 26.690 173.370 26.830 173.525 ;
        RECT 29.775 173.415 30.065 173.730 ;
        RECT 30.855 173.710 31.145 173.755 ;
        RECT 34.435 173.710 34.725 173.755 ;
        RECT 36.270 173.710 36.560 173.755 ;
        RECT 30.855 173.570 36.560 173.710 ;
        RECT 30.855 173.525 31.145 173.570 ;
        RECT 34.435 173.525 34.725 173.570 ;
        RECT 36.270 173.525 36.560 173.570 ;
        RECT 36.735 173.525 37.025 173.755 ;
        RECT 38.115 173.525 38.405 173.755 ;
        RECT 22.000 173.230 26.830 173.370 ;
        RECT 29.475 173.370 30.065 173.415 ;
        RECT 30.280 173.370 30.600 173.430 ;
        RECT 32.715 173.370 33.365 173.415 ;
        RECT 29.475 173.230 33.365 173.370 ;
        RECT 22.000 173.170 22.320 173.230 ;
        RECT 29.475 173.185 29.765 173.230 ;
        RECT 30.280 173.170 30.600 173.230 ;
        RECT 32.715 173.185 33.365 173.230 ;
        RECT 33.960 173.370 34.280 173.430 ;
        RECT 36.810 173.370 36.950 173.525 ;
        RECT 33.960 173.230 36.950 173.370 ;
        RECT 33.960 173.170 34.280 173.230 ;
        RECT 24.315 173.030 24.605 173.075 ;
        RECT 24.760 173.030 25.080 173.090 ;
        RECT 24.315 172.890 25.080 173.030 ;
        RECT 24.315 172.845 24.605 172.890 ;
        RECT 24.760 172.830 25.080 172.890 ;
        RECT 25.695 173.030 25.985 173.075 ;
        RECT 27.060 173.030 27.380 173.090 ;
        RECT 25.695 172.890 27.380 173.030 ;
        RECT 25.695 172.845 25.985 172.890 ;
        RECT 27.060 172.830 27.380 172.890 ;
        RECT 27.520 172.830 27.840 173.090 ;
        RECT 27.995 173.030 28.285 173.075 ;
        RECT 33.500 173.030 33.820 173.090 ;
        RECT 27.995 172.890 33.820 173.030 ;
        RECT 27.995 172.845 28.285 172.890 ;
        RECT 33.500 172.830 33.820 172.890 ;
        RECT 34.880 173.030 35.200 173.090 ;
        RECT 38.190 173.030 38.330 173.525 ;
        RECT 45.920 173.510 46.240 173.770 ;
        RECT 51.455 173.710 51.745 173.755 ;
        RECT 55.670 173.710 55.810 173.850 ;
        RECT 51.455 173.570 55.810 173.710 ;
        RECT 56.010 173.710 56.300 173.755 ;
        RECT 59.275 173.710 59.565 173.755 ;
        RECT 59.720 173.710 60.040 173.770 ;
        RECT 56.010 173.570 58.545 173.710 ;
        RECT 51.455 173.525 51.745 173.570 ;
        RECT 56.010 173.525 56.300 173.570 ;
        RECT 54.150 173.370 54.440 173.415 ;
        RECT 56.500 173.370 56.820 173.430 ;
        RECT 58.330 173.415 58.545 173.570 ;
        RECT 59.275 173.570 60.040 173.710 ;
        RECT 59.275 173.525 59.565 173.570 ;
        RECT 59.720 173.510 60.040 173.570 ;
        RECT 60.640 173.710 60.960 173.770 ;
        RECT 61.115 173.710 61.405 173.755 ;
        RECT 60.640 173.570 61.405 173.710 ;
        RECT 60.640 173.510 60.960 173.570 ;
        RECT 61.115 173.525 61.405 173.570 ;
        RECT 66.160 173.710 66.480 173.770 ;
        RECT 67.095 173.710 67.385 173.755 ;
        RECT 66.160 173.570 67.385 173.710 ;
        RECT 66.160 173.510 66.480 173.570 ;
        RECT 67.095 173.525 67.385 173.570 ;
        RECT 57.410 173.370 57.700 173.415 ;
        RECT 54.150 173.230 57.700 173.370 ;
        RECT 54.150 173.185 54.440 173.230 ;
        RECT 56.500 173.170 56.820 173.230 ;
        RECT 57.410 173.185 57.700 173.230 ;
        RECT 58.330 173.370 58.620 173.415 ;
        RECT 60.190 173.370 60.480 173.415 ;
        RECT 58.330 173.230 60.480 173.370 ;
        RECT 67.630 173.370 67.770 173.850 ;
        RECT 68.475 173.710 68.765 173.755 ;
        RECT 75.835 173.710 76.125 173.755 ;
        RECT 76.755 173.710 77.045 173.755 ;
        RECT 68.475 173.570 76.125 173.710 ;
        RECT 68.475 173.525 68.765 173.570 ;
        RECT 69.840 173.370 70.160 173.430 ;
        RECT 72.230 173.415 72.370 173.570 ;
        RECT 75.835 173.525 76.125 173.570 ;
        RECT 76.370 173.570 77.045 173.710 ;
        RECT 67.630 173.230 70.160 173.370 ;
        RECT 58.330 173.185 58.620 173.230 ;
        RECT 60.190 173.185 60.480 173.230 ;
        RECT 69.840 173.170 70.160 173.230 ;
        RECT 72.155 173.370 72.445 173.415 ;
        RECT 72.600 173.370 72.920 173.430 ;
        RECT 72.155 173.230 72.920 173.370 ;
        RECT 72.155 173.185 72.445 173.230 ;
        RECT 72.600 173.170 72.920 173.230 ;
        RECT 73.980 173.370 74.300 173.430 ;
        RECT 74.455 173.370 74.745 173.415 ;
        RECT 73.980 173.230 74.745 173.370 ;
        RECT 73.980 173.170 74.300 173.230 ;
        RECT 74.455 173.185 74.745 173.230 ;
        RECT 34.880 172.890 38.330 173.030 ;
        RECT 50.995 173.030 51.285 173.075 ;
        RECT 51.440 173.030 51.760 173.090 ;
        RECT 50.995 172.890 51.760 173.030 ;
        RECT 34.880 172.830 35.200 172.890 ;
        RECT 50.995 172.845 51.285 172.890 ;
        RECT 51.440 172.830 51.760 172.890 ;
        RECT 52.145 173.030 52.435 173.075 ;
        RECT 53.280 173.030 53.600 173.090 ;
        RECT 52.145 172.890 53.600 173.030 ;
        RECT 52.145 172.845 52.435 172.890 ;
        RECT 53.280 172.830 53.600 172.890 ;
        RECT 73.060 173.030 73.380 173.090 ;
        RECT 76.370 173.030 76.510 173.570 ;
        RECT 76.755 173.525 77.045 173.570 ;
        RECT 77.200 173.710 77.520 173.770 ;
        RECT 94.770 173.755 94.910 173.910 ;
        RECT 101.120 173.850 101.440 173.910 ;
        RECT 112.160 174.050 112.480 174.110 ;
        RECT 112.635 174.050 112.925 174.095 ;
        RECT 112.160 173.910 112.925 174.050 ;
        RECT 112.160 173.850 112.480 173.910 ;
        RECT 112.635 173.865 112.925 173.910 ;
        RECT 78.135 173.710 78.425 173.755 ;
        RECT 77.200 173.570 78.425 173.710 ;
        RECT 77.200 173.510 77.520 173.570 ;
        RECT 78.135 173.525 78.425 173.570 ;
        RECT 81.295 173.415 81.585 173.730 ;
        RECT 82.375 173.710 82.665 173.755 ;
        RECT 85.955 173.710 86.245 173.755 ;
        RECT 87.790 173.710 88.080 173.755 ;
        RECT 82.375 173.570 88.080 173.710 ;
        RECT 82.375 173.525 82.665 173.570 ;
        RECT 85.955 173.525 86.245 173.570 ;
        RECT 87.790 173.525 88.080 173.570 ;
        RECT 94.695 173.525 94.985 173.755 ;
        RECT 96.995 173.710 97.285 173.755 ;
        RECT 96.610 173.570 97.285 173.710 ;
        RECT 78.595 173.370 78.885 173.415 ;
        RECT 80.995 173.370 81.585 173.415 ;
        RECT 84.235 173.370 84.885 173.415 ;
        RECT 78.595 173.230 84.885 173.370 ;
        RECT 78.595 173.185 78.885 173.230 ;
        RECT 80.995 173.185 81.285 173.230 ;
        RECT 84.235 173.185 84.885 173.230 ;
        RECT 86.860 173.170 87.180 173.430 ;
        RECT 73.060 172.890 76.510 173.030 ;
        RECT 73.060 172.830 73.380 172.890 ;
        RECT 79.500 172.830 79.820 173.090 ;
        RECT 96.610 173.075 96.750 173.570 ;
        RECT 96.995 173.525 97.285 173.570 ;
        RECT 102.960 173.710 103.280 173.770 ;
        RECT 104.355 173.710 104.645 173.755 ;
        RECT 102.960 173.570 104.645 173.710 ;
        RECT 102.960 173.510 103.280 173.570 ;
        RECT 104.355 173.525 104.645 173.570 ;
        RECT 108.020 173.710 108.340 173.770 ;
        RECT 110.320 173.710 110.640 173.770 ;
        RECT 111.255 173.710 111.545 173.755 ;
        RECT 108.020 173.570 111.545 173.710 ;
        RECT 108.020 173.510 108.340 173.570 ;
        RECT 110.320 173.510 110.640 173.570 ;
        RECT 111.255 173.525 111.545 173.570 ;
        RECT 112.620 173.370 112.940 173.430 ;
        RECT 114.415 173.415 114.705 173.730 ;
        RECT 115.495 173.710 115.785 173.755 ;
        RECT 119.075 173.710 119.365 173.755 ;
        RECT 120.910 173.710 121.200 173.755 ;
        RECT 115.495 173.570 121.200 173.710 ;
        RECT 115.495 173.525 115.785 173.570 ;
        RECT 119.075 173.525 119.365 173.570 ;
        RECT 120.910 173.525 121.200 173.570 ;
        RECT 121.360 173.510 121.680 173.770 ;
        RECT 122.740 173.510 123.060 173.770 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 114.115 173.370 114.705 173.415 ;
        RECT 117.355 173.370 118.005 173.415 ;
        RECT 112.620 173.230 118.005 173.370 ;
        RECT 112.620 173.170 112.940 173.230 ;
        RECT 114.115 173.185 114.405 173.230 ;
        RECT 117.355 173.185 118.005 173.230 ;
        RECT 119.520 173.370 119.840 173.430 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 119.995 173.370 120.285 173.415 ;
        RECT 119.520 173.230 120.285 173.370 ;
        RECT 119.520 173.170 119.840 173.230 ;
        RECT 119.995 173.185 120.285 173.230 ;
        RECT 96.535 172.845 96.825 173.075 ;
        RECT 116.760 173.030 117.080 173.090 ;
        RECT 122.295 173.030 122.585 173.075 ;
        RECT 116.760 172.890 122.585 173.030 ;
        RECT 116.760 172.830 117.080 172.890 ;
        RECT 122.295 172.845 122.585 172.890 ;
        RECT 11.010 172.210 125.890 172.690 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 34.880 171.810 35.200 172.070 ;
        RECT 53.280 172.010 53.600 172.070 ;
        RECT 56.975 172.010 57.265 172.055 ;
        RECT 53.280 171.870 57.265 172.010 ;
        RECT 53.280 171.810 53.600 171.870 ;
        RECT 56.975 171.825 57.265 171.870 ;
        RECT 59.720 171.810 60.040 172.070 ;
        RECT 60.640 171.810 60.960 172.070 ;
        RECT 85.955 172.010 86.245 172.055 ;
        RECT 86.860 172.010 87.180 172.070 ;
        RECT 85.955 171.870 87.180 172.010 ;
        RECT 85.955 171.825 86.245 171.870 ;
        RECT 86.860 171.810 87.180 171.870 ;
        RECT 114.460 171.810 114.780 172.070 ;
        RECT 118.155 172.010 118.445 172.055 ;
        RECT 119.520 172.010 119.840 172.070 ;
        RECT 118.155 171.870 119.840 172.010 ;
        RECT 118.155 171.825 118.445 171.870 ;
        RECT 119.520 171.810 119.840 171.870 ;
        RECT 119.980 171.810 120.300 172.070 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 19.650 171.670 19.940 171.715 ;
        RECT 22.910 171.670 23.200 171.715 ;
        RECT 19.650 171.530 23.200 171.670 ;
        RECT 19.650 171.485 19.940 171.530 ;
        RECT 22.910 171.485 23.200 171.530 ;
        RECT 23.830 171.670 24.120 171.715 ;
        RECT 25.690 171.670 25.980 171.715 ;
        RECT 23.830 171.530 25.980 171.670 ;
        RECT 23.830 171.485 24.120 171.530 ;
        RECT 25.690 171.485 25.980 171.530 ;
        RECT 30.755 171.670 31.045 171.715 ;
        RECT 33.055 171.670 33.345 171.715 ;
        RECT 30.755 171.530 33.345 171.670 ;
        RECT 30.755 171.485 31.045 171.530 ;
        RECT 33.055 171.485 33.345 171.530 ;
        RECT 36.260 171.670 36.580 171.730 ;
        RECT 51.440 171.715 51.760 171.730 ;
        RECT 37.295 171.670 37.585 171.715 ;
        RECT 40.535 171.670 41.185 171.715 ;
        RECT 36.260 171.530 41.185 171.670 ;
        RECT 17.400 171.330 17.720 171.390 ;
        RECT 19.790 171.330 19.930 171.485 ;
        RECT 17.400 171.190 19.930 171.330 ;
        RECT 21.510 171.330 21.800 171.375 ;
        RECT 23.830 171.330 24.045 171.485 ;
        RECT 36.260 171.470 36.580 171.530 ;
        RECT 37.295 171.485 37.885 171.530 ;
        RECT 40.535 171.485 41.185 171.530 ;
        RECT 48.170 171.670 48.460 171.715 ;
        RECT 51.430 171.670 51.760 171.715 ;
        RECT 48.170 171.530 51.760 171.670 ;
        RECT 48.170 171.485 48.460 171.530 ;
        RECT 51.430 171.485 51.760 171.530 ;
        RECT 21.510 171.190 24.045 171.330 ;
        RECT 27.995 171.330 28.285 171.375 ;
        RECT 27.995 171.190 36.030 171.330 ;
        RECT 17.400 171.130 17.720 171.190 ;
        RECT 21.510 171.145 21.800 171.190 ;
        RECT 27.995 171.145 28.285 171.190 ;
        RECT 21.080 170.990 21.400 171.050 ;
        RECT 24.775 170.990 25.065 171.035 ;
        RECT 21.080 170.850 25.065 170.990 ;
        RECT 21.080 170.790 21.400 170.850 ;
        RECT 24.775 170.805 25.065 170.850 ;
        RECT 26.615 170.805 26.905 171.035 ;
        RECT 21.510 170.650 21.800 170.695 ;
        RECT 24.290 170.650 24.580 170.695 ;
        RECT 26.150 170.650 26.440 170.695 ;
        RECT 21.510 170.510 26.440 170.650 ;
        RECT 26.690 170.650 26.830 170.805 ;
        RECT 32.120 170.790 32.440 171.050 ;
        RECT 32.595 170.990 32.885 171.035 ;
        RECT 33.500 170.990 33.820 171.050 ;
        RECT 34.880 170.990 35.200 171.050 ;
        RECT 32.595 170.850 35.200 170.990 ;
        RECT 32.595 170.805 32.885 170.850 ;
        RECT 33.500 170.790 33.820 170.850 ;
        RECT 34.880 170.790 35.200 170.850 ;
        RECT 35.890 170.710 36.030 171.190 ;
        RECT 37.595 171.170 37.885 171.485 ;
        RECT 51.440 171.470 51.760 171.485 ;
        RECT 52.350 171.670 52.640 171.715 ;
        RECT 54.210 171.670 54.500 171.715 ;
        RECT 60.730 171.670 60.870 171.810 ;
        RECT 73.060 171.670 73.380 171.730 ;
        RECT 52.350 171.530 54.500 171.670 ;
        RECT 52.350 171.485 52.640 171.530 ;
        RECT 54.210 171.485 54.500 171.530 ;
        RECT 55.210 171.530 60.870 171.670 ;
        RECT 71.770 171.530 73.380 171.670 ;
        RECT 38.675 171.330 38.965 171.375 ;
        RECT 42.255 171.330 42.545 171.375 ;
        RECT 44.090 171.330 44.380 171.375 ;
        RECT 38.675 171.190 44.380 171.330 ;
        RECT 38.675 171.145 38.965 171.190 ;
        RECT 42.255 171.145 42.545 171.190 ;
        RECT 44.090 171.145 44.380 171.190 ;
        RECT 46.165 171.330 46.455 171.375 ;
        RECT 46.840 171.330 47.160 171.390 ;
        RECT 46.165 171.190 47.160 171.330 ;
        RECT 46.165 171.145 46.455 171.190 ;
        RECT 46.840 171.130 47.160 171.190 ;
        RECT 50.030 171.330 50.320 171.375 ;
        RECT 52.350 171.330 52.565 171.485 ;
        RECT 50.030 171.190 52.565 171.330 ;
        RECT 52.820 171.330 53.140 171.390 ;
        RECT 55.210 171.375 55.350 171.530 ;
        RECT 53.295 171.330 53.585 171.375 ;
        RECT 52.820 171.190 53.585 171.330 ;
        RECT 50.030 171.145 50.320 171.190 ;
        RECT 52.820 171.130 53.140 171.190 ;
        RECT 53.295 171.145 53.585 171.190 ;
        RECT 55.135 171.145 55.425 171.375 ;
        RECT 43.160 170.790 43.480 171.050 ;
        RECT 44.555 170.990 44.845 171.035 ;
        RECT 55.210 170.990 55.350 171.145 ;
        RECT 57.420 171.130 57.740 171.390 ;
        RECT 60.655 171.330 60.945 171.375 ;
        RECT 59.350 171.190 60.945 171.330 ;
        RECT 44.555 170.850 55.350 170.990 ;
        RECT 56.515 170.990 56.805 171.035 ;
        RECT 58.340 170.990 58.660 171.050 ;
        RECT 56.515 170.850 58.660 170.990 ;
        RECT 44.555 170.805 44.845 170.850 ;
        RECT 56.515 170.805 56.805 170.850 ;
        RECT 58.340 170.790 58.660 170.850 ;
        RECT 33.960 170.650 34.280 170.710 ;
        RECT 26.690 170.510 34.280 170.650 ;
        RECT 21.510 170.465 21.800 170.510 ;
        RECT 24.290 170.465 24.580 170.510 ;
        RECT 26.150 170.465 26.440 170.510 ;
        RECT 33.960 170.450 34.280 170.510 ;
        RECT 35.800 170.450 36.120 170.710 ;
        RECT 59.350 170.695 59.490 171.190 ;
        RECT 60.655 171.145 60.945 171.190 ;
        RECT 62.020 171.330 62.340 171.390 ;
        RECT 63.415 171.330 63.705 171.375 ;
        RECT 62.020 171.190 63.705 171.330 ;
        RECT 62.020 171.130 62.340 171.190 ;
        RECT 63.415 171.145 63.705 171.190 ;
        RECT 66.160 171.330 66.480 171.390 ;
        RECT 68.935 171.330 69.225 171.375 ;
        RECT 66.160 171.190 69.225 171.330 ;
        RECT 66.160 171.130 66.480 171.190 ;
        RECT 68.935 171.145 69.225 171.190 ;
        RECT 69.840 171.330 70.160 171.390 ;
        RECT 70.775 171.330 71.065 171.375 ;
        RECT 69.840 171.190 71.065 171.330 ;
        RECT 69.840 171.130 70.160 171.190 ;
        RECT 70.775 171.145 71.065 171.190 ;
        RECT 71.220 171.130 71.540 171.390 ;
        RECT 71.770 171.375 71.910 171.530 ;
        RECT 73.060 171.470 73.380 171.530 ;
        RECT 75.820 171.470 76.140 171.730 ;
        RECT 89.620 171.670 89.940 171.730 ;
        RECT 108.480 171.670 108.800 171.730 ;
        RECT 109.875 171.670 110.165 171.715 ;
        RECT 112.160 171.670 112.480 171.730 ;
        RECT 114.935 171.670 115.225 171.715 ;
        RECT 89.620 171.530 92.150 171.670 ;
        RECT 89.620 171.470 89.940 171.530 ;
        RECT 71.695 171.145 71.985 171.375 ;
        RECT 72.155 171.330 72.445 171.375 ;
        RECT 72.600 171.330 72.920 171.390 ;
        RECT 72.155 171.190 72.920 171.330 ;
        RECT 72.155 171.145 72.445 171.190 ;
        RECT 72.600 171.130 72.920 171.190 ;
        RECT 73.995 171.145 74.285 171.375 ;
        RECT 74.070 170.990 74.210 171.145 ;
        RECT 85.020 171.130 85.340 171.390 ;
        RECT 88.255 171.330 88.545 171.375 ;
        RECT 88.700 171.330 89.020 171.390 ;
        RECT 92.010 171.375 92.150 171.530 ;
        RECT 108.480 171.530 115.225 171.670 ;
        RECT 108.480 171.470 108.800 171.530 ;
        RECT 109.875 171.485 110.165 171.530 ;
        RECT 112.160 171.470 112.480 171.530 ;
        RECT 114.935 171.485 115.225 171.530 ;
        RECT 88.255 171.190 89.020 171.330 ;
        RECT 88.255 171.145 88.545 171.190 ;
        RECT 88.700 171.130 89.020 171.190 ;
        RECT 91.015 171.145 91.305 171.375 ;
        RECT 91.935 171.145 92.225 171.375 ;
        RECT 71.770 170.850 74.210 170.990 ;
        RECT 87.320 170.990 87.640 171.050 ;
        RECT 91.090 170.990 91.230 171.145 ;
        RECT 92.380 171.130 92.700 171.390 ;
        RECT 92.855 171.145 93.145 171.375 ;
        RECT 92.930 170.990 93.070 171.145 ;
        RECT 100.660 171.130 100.980 171.390 ;
        RECT 105.275 171.145 105.565 171.375 ;
        RECT 103.420 170.990 103.740 171.050 ;
        RECT 105.350 170.990 105.490 171.145 ;
        RECT 105.720 171.130 106.040 171.390 ;
        RECT 106.180 171.130 106.500 171.390 ;
        RECT 107.100 171.130 107.420 171.390 ;
        RECT 108.940 171.330 109.260 171.390 ;
        RECT 110.335 171.330 110.625 171.375 ;
        RECT 117.235 171.330 117.525 171.375 ;
        RECT 108.940 171.190 110.625 171.330 ;
        RECT 108.940 171.130 109.260 171.190 ;
        RECT 110.335 171.145 110.625 171.190 ;
        RECT 114.780 171.190 117.525 171.330 ;
        RECT 87.320 170.850 91.230 170.990 ;
        RECT 92.470 170.850 105.490 170.990 ;
        RECT 109.415 170.990 109.705 171.035 ;
        RECT 113.555 170.990 113.845 171.035 ;
        RECT 109.415 170.850 113.845 170.990 ;
        RECT 71.770 170.710 71.910 170.850 ;
        RECT 87.320 170.790 87.640 170.850 ;
        RECT 38.675 170.650 38.965 170.695 ;
        RECT 41.795 170.650 42.085 170.695 ;
        RECT 43.685 170.650 43.975 170.695 ;
        RECT 50.030 170.650 50.320 170.695 ;
        RECT 52.810 170.650 53.100 170.695 ;
        RECT 54.670 170.650 54.960 170.695 ;
        RECT 38.675 170.510 43.975 170.650 ;
        RECT 38.675 170.465 38.965 170.510 ;
        RECT 41.795 170.465 42.085 170.510 ;
        RECT 43.685 170.465 43.975 170.510 ;
        RECT 45.550 170.510 47.070 170.650 ;
        RECT 17.645 170.310 17.935 170.355 ;
        RECT 23.840 170.310 24.160 170.370 ;
        RECT 17.645 170.170 24.160 170.310 ;
        RECT 17.645 170.125 17.935 170.170 ;
        RECT 23.840 170.110 24.160 170.170 ;
        RECT 32.120 170.310 32.440 170.370 ;
        RECT 33.500 170.310 33.820 170.370 ;
        RECT 37.640 170.310 37.960 170.370 ;
        RECT 45.550 170.310 45.690 170.510 ;
        RECT 32.120 170.170 45.690 170.310 ;
        RECT 46.930 170.310 47.070 170.510 ;
        RECT 50.030 170.510 54.960 170.650 ;
        RECT 50.030 170.465 50.320 170.510 ;
        RECT 52.810 170.465 53.100 170.510 ;
        RECT 54.670 170.465 54.960 170.510 ;
        RECT 59.275 170.465 59.565 170.695 ;
        RECT 62.495 170.650 62.785 170.695 ;
        RECT 64.320 170.650 64.640 170.710 ;
        RECT 62.495 170.510 64.640 170.650 ;
        RECT 62.495 170.465 62.785 170.510 ;
        RECT 64.320 170.450 64.640 170.510 ;
        RECT 71.680 170.450 72.000 170.710 ;
        RECT 86.860 170.650 87.180 170.710 ;
        RECT 87.795 170.650 88.085 170.695 ;
        RECT 86.860 170.510 88.085 170.650 ;
        RECT 86.860 170.450 87.180 170.510 ;
        RECT 87.795 170.465 88.085 170.510 ;
        RECT 60.180 170.310 60.500 170.370 ;
        RECT 46.930 170.170 60.500 170.310 ;
        RECT 32.120 170.110 32.440 170.170 ;
        RECT 33.500 170.110 33.820 170.170 ;
        RECT 37.640 170.110 37.960 170.170 ;
        RECT 60.180 170.110 60.500 170.170 ;
        RECT 69.395 170.310 69.685 170.355 ;
        RECT 72.600 170.310 72.920 170.370 ;
        RECT 69.395 170.170 72.920 170.310 ;
        RECT 69.395 170.125 69.685 170.170 ;
        RECT 72.600 170.110 72.920 170.170 ;
        RECT 73.060 170.110 73.380 170.370 ;
        RECT 76.740 170.310 77.060 170.370 ;
        RECT 92.470 170.310 92.610 170.850 ;
        RECT 103.420 170.790 103.740 170.850 ;
        RECT 109.415 170.805 109.705 170.850 ;
        RECT 113.555 170.805 113.845 170.850 ;
        RECT 94.235 170.650 94.525 170.695 ;
        RECT 95.140 170.650 95.460 170.710 ;
        RECT 94.235 170.510 95.460 170.650 ;
        RECT 94.235 170.465 94.525 170.510 ;
        RECT 95.140 170.450 95.460 170.510 ;
        RECT 102.960 170.650 103.280 170.710 ;
        RECT 103.895 170.650 104.185 170.695 ;
        RECT 102.960 170.510 104.185 170.650 ;
        RECT 109.490 170.650 109.630 170.805 ;
        RECT 110.320 170.650 110.640 170.710 ;
        RECT 109.490 170.510 110.640 170.650 ;
        RECT 102.960 170.450 103.280 170.510 ;
        RECT 103.895 170.465 104.185 170.510 ;
        RECT 110.320 170.450 110.640 170.510 ;
        RECT 112.175 170.650 112.465 170.695 ;
        RECT 114.780 170.650 114.920 171.190 ;
        RECT 117.235 171.145 117.525 171.190 ;
        RECT 119.075 171.145 119.365 171.375 ;
        RECT 119.150 170.990 119.290 171.145 ;
        RECT 116.850 170.850 119.290 170.990 ;
        RECT 116.850 170.695 116.990 170.850 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 112.175 170.510 114.920 170.650 ;
        RECT 112.175 170.465 112.465 170.510 ;
        RECT 116.775 170.465 117.065 170.695 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 76.740 170.170 92.610 170.310 ;
        RECT 76.740 170.110 77.060 170.170 ;
        RECT 99.740 170.110 100.060 170.370 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 11.810 169.490 125.890 169.970 ;
        RECT 17.400 169.090 17.720 169.350 ;
        RECT 22.000 169.090 22.320 169.350 ;
        RECT 36.260 169.090 36.580 169.350 ;
        RECT 42.255 169.290 42.545 169.335 ;
        RECT 43.160 169.290 43.480 169.350 ;
        RECT 42.255 169.150 43.480 169.290 ;
        RECT 42.255 169.105 42.545 169.150 ;
        RECT 43.160 169.090 43.480 169.150 ;
        RECT 51.915 169.290 52.205 169.335 ;
        RECT 52.360 169.290 52.680 169.350 ;
        RECT 51.915 169.150 52.680 169.290 ;
        RECT 51.915 169.105 52.205 169.150 ;
        RECT 52.360 169.090 52.680 169.150 ;
        RECT 55.580 169.290 55.900 169.350 ;
        RECT 71.695 169.290 71.985 169.335 ;
        RECT 87.320 169.290 87.640 169.350 ;
        RECT 55.580 169.150 87.640 169.290 ;
        RECT 55.580 169.090 55.900 169.150 ;
        RECT 71.695 169.105 71.985 169.150 ;
        RECT 87.320 169.090 87.640 169.150 ;
        RECT 88.240 169.290 88.560 169.350 ;
        RECT 90.095 169.290 90.385 169.335 ;
        RECT 88.240 169.150 90.385 169.290 ;
        RECT 88.240 169.090 88.560 169.150 ;
        RECT 90.095 169.105 90.385 169.150 ;
        RECT 98.835 169.290 99.125 169.335 ;
        RECT 100.660 169.290 100.980 169.350 ;
        RECT 98.835 169.150 100.980 169.290 ;
        RECT 98.835 169.105 99.125 169.150 ;
        RECT 100.660 169.090 100.980 169.150 ;
        RECT 25.795 168.950 26.085 168.995 ;
        RECT 28.915 168.950 29.205 168.995 ;
        RECT 30.805 168.950 31.095 168.995 ;
        RECT 25.795 168.810 31.095 168.950 ;
        RECT 25.795 168.765 26.085 168.810 ;
        RECT 28.915 168.765 29.205 168.810 ;
        RECT 30.805 168.765 31.095 168.810 ;
        RECT 35.800 168.950 36.120 169.010 ;
        RECT 39.020 168.950 39.340 169.010 ;
        RECT 71.220 168.950 71.540 169.010 ;
        RECT 92.380 168.950 92.700 169.010 ;
        RECT 102.040 168.950 102.360 169.010 ;
        RECT 105.720 168.950 106.040 169.010 ;
        RECT 35.800 168.810 38.790 168.950 ;
        RECT 35.800 168.750 36.120 168.810 ;
        RECT 19.255 168.610 19.545 168.655 ;
        RECT 24.300 168.610 24.620 168.670 ;
        RECT 19.255 168.470 24.620 168.610 ;
        RECT 19.255 168.425 19.545 168.470 ;
        RECT 24.300 168.410 24.620 168.470 ;
        RECT 27.520 168.610 27.840 168.670 ;
        RECT 30.295 168.610 30.585 168.655 ;
        RECT 27.520 168.470 30.585 168.610 ;
        RECT 27.520 168.410 27.840 168.470 ;
        RECT 30.295 168.425 30.585 168.470 ;
        RECT 31.675 168.610 31.965 168.655 ;
        RECT 32.120 168.610 32.440 168.670 ;
        RECT 33.960 168.610 34.280 168.670 ;
        RECT 31.675 168.470 34.280 168.610 ;
        RECT 31.675 168.425 31.965 168.470 ;
        RECT 32.120 168.410 32.440 168.470 ;
        RECT 33.960 168.410 34.280 168.470 ;
        RECT 37.640 168.410 37.960 168.670 ;
        RECT 38.650 168.655 38.790 168.810 ;
        RECT 39.020 168.810 57.190 168.950 ;
        RECT 39.020 168.750 39.340 168.810 ;
        RECT 38.575 168.610 38.865 168.655 ;
        RECT 38.575 168.470 42.010 168.610 ;
        RECT 38.575 168.425 38.865 168.470 ;
        RECT 17.875 168.270 18.165 168.315 ;
        RECT 23.380 168.270 23.700 168.330 ;
        RECT 24.760 168.290 25.080 168.330 ;
        RECT 17.875 168.130 23.700 168.270 ;
        RECT 17.875 168.085 18.165 168.130 ;
        RECT 23.380 168.070 23.700 168.130 ;
        RECT 24.715 168.070 25.080 168.290 ;
        RECT 25.795 168.270 26.085 168.315 ;
        RECT 29.375 168.270 29.665 168.315 ;
        RECT 31.210 168.270 31.500 168.315 ;
        RECT 25.795 168.130 31.500 168.270 ;
        RECT 25.795 168.085 26.085 168.130 ;
        RECT 29.375 168.085 29.665 168.130 ;
        RECT 31.210 168.085 31.500 168.130 ;
        RECT 35.815 168.270 36.105 168.315 ;
        RECT 36.720 168.270 37.040 168.330 ;
        RECT 39.020 168.270 39.340 168.330 ;
        RECT 41.335 168.270 41.625 168.315 ;
        RECT 35.815 168.130 39.340 168.270 ;
        RECT 35.815 168.085 36.105 168.130 ;
        RECT 36.720 168.070 37.040 168.130 ;
        RECT 39.020 168.070 39.340 168.130 ;
        RECT 40.950 168.130 41.625 168.270 ;
        RECT 24.715 167.975 25.005 168.070 ;
        RECT 20.175 167.930 20.465 167.975 ;
        RECT 24.415 167.930 25.005 167.975 ;
        RECT 27.655 167.930 28.305 167.975 ;
        RECT 34.880 167.930 35.200 167.990 ;
        RECT 20.175 167.790 24.070 167.930 ;
        RECT 20.175 167.745 20.465 167.790 ;
        RECT 19.715 167.590 20.005 167.635 ;
        RECT 22.920 167.590 23.240 167.650 ;
        RECT 19.715 167.450 23.240 167.590 ;
        RECT 23.930 167.590 24.070 167.790 ;
        RECT 24.415 167.790 28.305 167.930 ;
        RECT 24.415 167.745 24.705 167.790 ;
        RECT 27.655 167.745 28.305 167.790 ;
        RECT 31.290 167.790 35.200 167.930 ;
        RECT 31.290 167.590 31.430 167.790 ;
        RECT 34.880 167.730 35.200 167.790 ;
        RECT 23.930 167.450 31.430 167.590 ;
        RECT 32.580 167.590 32.900 167.650 ;
        RECT 40.950 167.635 41.090 168.130 ;
        RECT 41.335 168.085 41.625 168.130 ;
        RECT 41.870 167.930 42.010 168.470 ;
        RECT 45.000 168.410 45.320 168.670 ;
        RECT 57.050 168.655 57.190 168.810 ;
        RECT 71.220 168.810 106.040 168.950 ;
        RECT 71.220 168.750 71.540 168.810 ;
        RECT 92.380 168.750 92.700 168.810 ;
        RECT 102.040 168.750 102.360 168.810 ;
        RECT 56.975 168.425 57.265 168.655 ;
        RECT 73.980 168.610 74.300 168.670 ;
        RECT 70.850 168.470 74.300 168.610 ;
        RECT 45.935 168.270 46.225 168.315 ;
        RECT 46.380 168.270 46.700 168.330 ;
        RECT 48.220 168.270 48.540 168.330 ;
        RECT 45.935 168.130 46.700 168.270 ;
        RECT 45.935 168.085 46.225 168.130 ;
        RECT 46.380 168.070 46.700 168.130 ;
        RECT 46.930 168.130 48.540 168.270 ;
        RECT 46.930 167.930 47.070 168.130 ;
        RECT 48.220 168.070 48.540 168.130 ;
        RECT 50.995 168.085 51.285 168.315 ;
        RECT 54.675 168.270 54.965 168.315 ;
        RECT 56.500 168.270 56.820 168.330 ;
        RECT 54.675 168.130 56.820 168.270 ;
        RECT 54.675 168.085 54.965 168.130 ;
        RECT 41.870 167.790 47.070 167.930 ;
        RECT 39.035 167.590 39.325 167.635 ;
        RECT 32.580 167.450 39.325 167.590 ;
        RECT 19.715 167.405 20.005 167.450 ;
        RECT 22.920 167.390 23.240 167.450 ;
        RECT 32.580 167.390 32.900 167.450 ;
        RECT 39.035 167.405 39.325 167.450 ;
        RECT 40.875 167.405 41.165 167.635 ;
        RECT 45.475 167.590 45.765 167.635 ;
        RECT 46.840 167.590 47.160 167.650 ;
        RECT 45.475 167.450 47.160 167.590 ;
        RECT 45.475 167.405 45.765 167.450 ;
        RECT 46.840 167.390 47.160 167.450 ;
        RECT 47.775 167.590 48.065 167.635 ;
        RECT 51.070 167.590 51.210 168.085 ;
        RECT 56.500 168.070 56.820 168.130 ;
        RECT 58.355 168.270 58.645 168.315 ;
        RECT 61.115 168.270 61.405 168.315 ;
        RECT 62.020 168.270 62.340 168.330 ;
        RECT 70.850 168.315 70.990 168.470 ;
        RECT 73.980 168.410 74.300 168.470 ;
        RECT 87.320 168.610 87.640 168.670 ;
        RECT 87.320 168.470 95.370 168.610 ;
        RECT 87.320 168.410 87.640 168.470 ;
        RECT 58.355 168.130 62.340 168.270 ;
        RECT 58.355 168.085 58.645 168.130 ;
        RECT 61.115 168.085 61.405 168.130 ;
        RECT 62.020 168.070 62.340 168.130 ;
        RECT 70.775 168.085 71.065 168.315 ;
        RECT 72.600 168.070 72.920 168.330 ;
        RECT 94.680 168.070 95.000 168.330 ;
        RECT 95.230 168.270 95.370 168.470 ;
        RECT 96.060 168.410 96.380 168.670 ;
        RECT 101.135 168.270 101.425 168.315 ;
        RECT 95.230 168.130 101.425 168.270 ;
        RECT 101.135 168.085 101.425 168.130 ;
        RECT 101.580 168.270 101.900 168.330 ;
        RECT 102.590 168.315 102.730 168.810 ;
        RECT 105.720 168.750 106.040 168.810 ;
        RECT 110.895 168.950 111.185 168.995 ;
        RECT 114.015 168.950 114.305 168.995 ;
        RECT 115.905 168.950 116.195 168.995 ;
        RECT 110.895 168.810 116.195 168.950 ;
        RECT 110.895 168.765 111.185 168.810 ;
        RECT 114.015 168.765 114.305 168.810 ;
        RECT 115.905 168.765 116.195 168.810 ;
        RECT 117.235 168.765 117.525 168.995 ;
        RECT 107.100 168.610 107.420 168.670 ;
        RECT 106.270 168.470 107.420 168.610 ;
        RECT 102.055 168.270 102.345 168.315 ;
        RECT 101.580 168.130 102.345 168.270 ;
        RECT 56.590 167.930 56.730 168.070 ;
        RECT 59.735 167.930 60.025 167.975 ;
        RECT 56.590 167.790 60.025 167.930 ;
        RECT 59.735 167.745 60.025 167.790 ;
        RECT 60.180 167.930 60.500 167.990 ;
        RECT 67.095 167.930 67.385 167.975 ;
        RECT 60.180 167.790 67.385 167.930 ;
        RECT 60.180 167.730 60.500 167.790 ;
        RECT 67.095 167.745 67.385 167.790 ;
        RECT 68.935 167.930 69.225 167.975 ;
        RECT 71.680 167.930 72.000 167.990 ;
        RECT 68.935 167.790 72.000 167.930 ;
        RECT 68.935 167.745 69.225 167.790 ;
        RECT 71.680 167.730 72.000 167.790 ;
        RECT 83.640 167.730 83.960 167.990 ;
        RECT 96.995 167.930 97.285 167.975 ;
        RECT 84.190 167.790 97.285 167.930 ;
        RECT 101.210 167.930 101.350 168.085 ;
        RECT 101.580 168.070 101.900 168.130 ;
        RECT 102.055 168.085 102.345 168.130 ;
        RECT 102.515 168.085 102.805 168.315 ;
        RECT 102.975 168.270 103.265 168.315 ;
        RECT 103.420 168.270 103.740 168.330 ;
        RECT 102.975 168.130 103.740 168.270 ;
        RECT 102.975 168.085 103.265 168.130 ;
        RECT 103.420 168.070 103.740 168.130 ;
        RECT 106.270 167.930 106.410 168.470 ;
        RECT 107.100 168.410 107.420 168.470 ;
        RECT 115.395 168.610 115.685 168.655 ;
        RECT 117.310 168.610 117.450 168.765 ;
        RECT 115.395 168.470 117.450 168.610 ;
        RECT 115.395 168.425 115.685 168.470 ;
        RECT 106.655 168.270 106.945 168.315 ;
        RECT 108.020 168.270 108.340 168.330 ;
        RECT 106.655 168.130 108.340 168.270 ;
        RECT 106.655 168.085 106.945 168.130 ;
        RECT 108.020 168.070 108.340 168.130 ;
        RECT 109.815 167.975 110.105 168.290 ;
        RECT 110.895 168.270 111.185 168.315 ;
        RECT 114.475 168.270 114.765 168.315 ;
        RECT 116.310 168.270 116.600 168.315 ;
        RECT 110.895 168.130 116.600 168.270 ;
        RECT 110.895 168.085 111.185 168.130 ;
        RECT 114.475 168.085 114.765 168.130 ;
        RECT 116.310 168.085 116.600 168.130 ;
        RECT 116.775 168.085 117.065 168.315 ;
        RECT 101.210 167.790 106.410 167.930 ;
        RECT 107.115 167.930 107.405 167.975 ;
        RECT 109.515 167.930 110.105 167.975 ;
        RECT 112.755 167.930 113.405 167.975 ;
        RECT 107.115 167.790 113.405 167.930 ;
        RECT 116.850 167.930 116.990 168.085 ;
        RECT 118.140 168.070 118.460 168.330 ;
        RECT 121.360 167.930 121.680 167.990 ;
        RECT 116.850 167.790 121.680 167.930 ;
        RECT 47.775 167.450 51.210 167.590 ;
        RECT 47.775 167.405 48.065 167.450 ;
        RECT 55.120 167.390 55.440 167.650 ;
        RECT 69.840 167.390 70.160 167.650 ;
        RECT 78.580 167.590 78.900 167.650 ;
        RECT 84.190 167.590 84.330 167.790 ;
        RECT 96.995 167.745 97.285 167.790 ;
        RECT 107.115 167.745 107.405 167.790 ;
        RECT 109.515 167.745 109.805 167.790 ;
        RECT 112.755 167.745 113.405 167.790 ;
        RECT 121.360 167.730 121.680 167.790 ;
        RECT 78.580 167.450 84.330 167.590 ;
        RECT 92.840 167.590 93.160 167.650 ;
        RECT 94.235 167.590 94.525 167.635 ;
        RECT 92.840 167.450 94.525 167.590 ;
        RECT 78.580 167.390 78.900 167.450 ;
        RECT 92.840 167.390 93.160 167.450 ;
        RECT 94.235 167.405 94.525 167.450 ;
        RECT 96.535 167.590 96.825 167.635 ;
        RECT 98.360 167.590 98.680 167.650 ;
        RECT 96.535 167.450 98.680 167.590 ;
        RECT 96.535 167.405 96.825 167.450 ;
        RECT 98.360 167.390 98.680 167.450 ;
        RECT 104.355 167.590 104.645 167.635 ;
        RECT 106.180 167.590 106.500 167.650 ;
        RECT 104.355 167.450 106.500 167.590 ;
        RECT 104.355 167.405 104.645 167.450 ;
        RECT 106.180 167.390 106.500 167.450 ;
        RECT 108.035 167.590 108.325 167.635 ;
        RECT 108.940 167.590 109.260 167.650 ;
        RECT 108.035 167.450 109.260 167.590 ;
        RECT 108.035 167.405 108.325 167.450 ;
        RECT 108.940 167.390 109.260 167.450 ;
        RECT 11.010 166.770 125.890 167.250 ;
        RECT 21.080 166.370 21.400 166.630 ;
        RECT 21.555 166.385 21.845 166.615 ;
        RECT 23.840 166.570 24.160 166.630 ;
        RECT 39.940 166.570 40.260 166.630 ;
        RECT 23.840 166.430 40.260 166.570 ;
        RECT 20.175 165.890 20.465 165.935 ;
        RECT 21.630 165.890 21.770 166.385 ;
        RECT 23.840 166.370 24.160 166.430 ;
        RECT 39.940 166.370 40.260 166.430 ;
        RECT 40.860 166.570 41.180 166.630 ;
        RECT 45.460 166.570 45.780 166.630 ;
        RECT 51.685 166.570 51.975 166.615 ;
        RECT 52.820 166.570 53.140 166.630 ;
        RECT 57.420 166.570 57.740 166.630 ;
        RECT 40.860 166.430 49.370 166.570 ;
        RECT 40.860 166.370 41.180 166.430 ;
        RECT 45.460 166.370 45.780 166.430 ;
        RECT 27.175 166.230 27.465 166.275 ;
        RECT 30.415 166.230 31.065 166.275 ;
        RECT 27.175 166.090 31.065 166.230 ;
        RECT 27.175 166.045 27.765 166.090 ;
        RECT 30.415 166.045 31.065 166.090 ;
        RECT 36.720 166.230 37.040 166.290 ;
        RECT 36.720 166.090 48.910 166.230 ;
        RECT 27.475 165.950 27.765 166.045 ;
        RECT 36.720 166.030 37.040 166.090 ;
        RECT 20.175 165.750 21.770 165.890 ;
        RECT 22.920 165.890 23.240 165.950 ;
        RECT 23.395 165.890 23.685 165.935 ;
        RECT 24.300 165.890 24.620 165.950 ;
        RECT 22.920 165.750 24.620 165.890 ;
        RECT 20.175 165.705 20.465 165.750 ;
        RECT 22.920 165.690 23.240 165.750 ;
        RECT 23.395 165.705 23.685 165.750 ;
        RECT 24.300 165.690 24.620 165.750 ;
        RECT 27.475 165.730 27.840 165.950 ;
        RECT 27.520 165.690 27.840 165.730 ;
        RECT 28.555 165.890 28.845 165.935 ;
        RECT 32.135 165.890 32.425 165.935 ;
        RECT 33.970 165.890 34.260 165.935 ;
        RECT 28.555 165.750 34.260 165.890 ;
        RECT 28.555 165.705 28.845 165.750 ;
        RECT 32.135 165.705 32.425 165.750 ;
        RECT 33.970 165.705 34.260 165.750 ;
        RECT 34.420 165.690 34.740 165.950 ;
        RECT 39.570 165.935 39.710 166.090 ;
        RECT 39.035 165.705 39.325 165.935 ;
        RECT 39.495 165.705 39.785 165.935 ;
        RECT 24.760 165.350 25.080 165.610 ;
        RECT 33.040 165.350 33.360 165.610 ;
        RECT 37.180 165.550 37.500 165.610 ;
        RECT 39.110 165.550 39.250 165.705 ;
        RECT 39.940 165.690 40.260 165.950 ;
        RECT 40.860 165.690 41.180 165.950 ;
        RECT 44.170 165.935 44.310 166.090 ;
        RECT 43.635 165.705 43.925 165.935 ;
        RECT 44.095 165.705 44.385 165.935 ;
        RECT 43.710 165.550 43.850 165.705 ;
        RECT 44.540 165.690 44.860 165.950 ;
        RECT 45.460 165.690 45.780 165.950 ;
        RECT 47.850 165.935 47.990 166.090 ;
        RECT 47.315 165.705 47.605 165.935 ;
        RECT 47.775 165.705 48.065 165.935 ;
        RECT 47.390 165.550 47.530 165.705 ;
        RECT 48.220 165.690 48.540 165.950 ;
        RECT 48.770 165.550 48.910 166.090 ;
        RECT 49.230 165.935 49.370 166.430 ;
        RECT 51.685 166.430 57.740 166.570 ;
        RECT 51.685 166.385 51.975 166.430 ;
        RECT 52.820 166.370 53.140 166.430 ;
        RECT 57.420 166.370 57.740 166.430 ;
        RECT 58.340 166.570 58.660 166.630 ;
        RECT 63.415 166.570 63.705 166.615 ;
        RECT 58.340 166.430 63.705 166.570 ;
        RECT 58.340 166.370 58.660 166.430 ;
        RECT 63.415 166.385 63.705 166.430 ;
        RECT 68.475 166.570 68.765 166.615 ;
        RECT 71.220 166.570 71.540 166.630 ;
        RECT 68.475 166.430 71.540 166.570 ;
        RECT 68.475 166.385 68.765 166.430 ;
        RECT 53.690 166.230 53.980 166.275 ;
        RECT 55.120 166.230 55.440 166.290 ;
        RECT 56.950 166.230 57.240 166.275 ;
        RECT 53.690 166.090 57.240 166.230 ;
        RECT 53.690 166.045 53.980 166.090 ;
        RECT 55.120 166.030 55.440 166.090 ;
        RECT 56.950 166.045 57.240 166.090 ;
        RECT 57.870 166.230 58.160 166.275 ;
        RECT 59.730 166.230 60.020 166.275 ;
        RECT 57.870 166.090 60.020 166.230 ;
        RECT 57.870 166.045 58.160 166.090 ;
        RECT 59.730 166.045 60.020 166.090 ;
        RECT 60.180 166.230 60.500 166.290 ;
        RECT 68.550 166.230 68.690 166.385 ;
        RECT 71.220 166.370 71.540 166.430 ;
        RECT 71.680 166.370 72.000 166.630 ;
        RECT 74.455 166.570 74.745 166.615 ;
        RECT 86.860 166.570 87.180 166.630 ;
        RECT 72.230 166.430 74.745 166.570 ;
        RECT 72.230 166.230 72.370 166.430 ;
        RECT 74.455 166.385 74.745 166.430 ;
        RECT 83.270 166.430 87.180 166.570 ;
        RECT 60.180 166.090 68.690 166.230 ;
        RECT 69.470 166.090 72.370 166.230 ;
        RECT 49.155 165.890 49.445 165.935 ;
        RECT 54.200 165.890 54.520 165.950 ;
        RECT 49.155 165.750 54.520 165.890 ;
        RECT 49.155 165.705 49.445 165.750 ;
        RECT 54.200 165.690 54.520 165.750 ;
        RECT 55.550 165.890 55.840 165.935 ;
        RECT 57.870 165.890 58.085 166.045 ;
        RECT 60.180 166.030 60.500 166.090 ;
        RECT 69.470 165.950 69.610 166.090 ;
        RECT 72.600 166.030 72.920 166.290 ;
        RECT 79.450 166.230 79.740 166.275 ;
        RECT 82.710 166.230 83.000 166.275 ;
        RECT 83.270 166.230 83.410 166.430 ;
        RECT 86.860 166.370 87.180 166.430 ;
        RECT 94.680 166.570 95.000 166.630 ;
        RECT 98.360 166.570 98.680 166.630 ;
        RECT 109.415 166.570 109.705 166.615 ;
        RECT 94.680 166.430 96.290 166.570 ;
        RECT 94.680 166.370 95.000 166.430 ;
        RECT 73.610 166.090 75.590 166.230 ;
        RECT 55.550 165.750 58.085 165.890 ;
        RECT 58.815 165.890 59.105 165.935 ;
        RECT 58.815 165.750 61.330 165.890 ;
        RECT 55.550 165.705 55.840 165.750 ;
        RECT 58.815 165.705 59.105 165.750 ;
        RECT 59.720 165.550 60.040 165.610 ;
        RECT 37.180 165.410 47.990 165.550 ;
        RECT 48.770 165.410 60.040 165.550 ;
        RECT 37.180 165.350 37.500 165.410 ;
        RECT 28.555 165.210 28.845 165.255 ;
        RECT 31.675 165.210 31.965 165.255 ;
        RECT 33.565 165.210 33.855 165.255 ;
        RECT 28.555 165.070 33.855 165.210 ;
        RECT 28.555 165.025 28.845 165.070 ;
        RECT 31.675 165.025 31.965 165.070 ;
        RECT 33.565 165.025 33.855 165.070 ;
        RECT 34.880 165.210 35.200 165.270 ;
        RECT 44.540 165.210 44.860 165.270 ;
        RECT 34.880 165.070 44.860 165.210 ;
        RECT 34.880 165.010 35.200 165.070 ;
        RECT 44.540 165.010 44.860 165.070 ;
        RECT 25.695 164.870 25.985 164.915 ;
        RECT 27.980 164.870 28.300 164.930 ;
        RECT 25.695 164.730 28.300 164.870 ;
        RECT 25.695 164.685 25.985 164.730 ;
        RECT 27.980 164.670 28.300 164.730 ;
        RECT 37.640 164.670 37.960 164.930 ;
        RECT 38.560 164.870 38.880 164.930 ;
        RECT 42.255 164.870 42.545 164.915 ;
        RECT 38.560 164.730 42.545 164.870 ;
        RECT 38.560 164.670 38.880 164.730 ;
        RECT 42.255 164.685 42.545 164.730 ;
        RECT 45.920 164.670 46.240 164.930 ;
        RECT 47.850 164.870 47.990 165.410 ;
        RECT 59.720 165.350 60.040 165.410 ;
        RECT 60.640 165.350 60.960 165.610 ;
        RECT 55.550 165.210 55.840 165.255 ;
        RECT 58.330 165.210 58.620 165.255 ;
        RECT 60.190 165.210 60.480 165.255 ;
        RECT 55.550 165.070 60.480 165.210 ;
        RECT 61.190 165.210 61.330 165.750 ;
        RECT 62.480 165.690 62.800 165.950 ;
        RECT 64.795 165.890 65.085 165.935 ;
        RECT 68.920 165.890 69.240 165.950 ;
        RECT 64.795 165.750 69.240 165.890 ;
        RECT 64.795 165.705 65.085 165.750 ;
        RECT 68.920 165.690 69.240 165.750 ;
        RECT 69.380 165.690 69.700 165.950 ;
        RECT 69.840 165.690 70.160 165.950 ;
        RECT 72.155 165.890 72.445 165.935 ;
        RECT 72.690 165.890 72.830 166.030 ;
        RECT 72.155 165.750 72.830 165.890 ;
        RECT 73.060 165.890 73.380 165.950 ;
        RECT 73.610 165.935 73.750 166.090 ;
        RECT 73.535 165.890 73.825 165.935 ;
        RECT 73.060 165.750 73.825 165.890 ;
        RECT 72.155 165.705 72.445 165.750 ;
        RECT 73.060 165.690 73.380 165.750 ;
        RECT 73.535 165.705 73.825 165.750 ;
        RECT 73.980 165.690 74.300 165.950 ;
        RECT 75.450 165.935 75.590 166.090 ;
        RECT 79.450 166.090 83.410 166.230 ;
        RECT 83.630 166.230 83.920 166.275 ;
        RECT 85.490 166.230 85.780 166.275 ;
        RECT 83.630 166.090 85.780 166.230 ;
        RECT 79.450 166.045 79.740 166.090 ;
        RECT 82.710 166.045 83.000 166.090 ;
        RECT 83.630 166.045 83.920 166.090 ;
        RECT 85.490 166.045 85.780 166.090 ;
        RECT 75.375 165.705 75.665 165.935 ;
        RECT 81.310 165.890 81.600 165.935 ;
        RECT 83.630 165.890 83.845 166.045 ;
        RECT 95.600 166.030 95.920 166.290 ;
        RECT 96.150 166.230 96.290 166.430 ;
        RECT 98.360 166.430 109.705 166.570 ;
        RECT 98.360 166.370 98.680 166.430 ;
        RECT 109.415 166.385 109.705 166.430 ;
        RECT 111.255 166.570 111.545 166.615 ;
        RECT 118.140 166.570 118.460 166.630 ;
        RECT 111.255 166.430 118.460 166.570 ;
        RECT 111.255 166.385 111.545 166.430 ;
        RECT 118.140 166.370 118.460 166.430 ;
        RECT 108.020 166.230 108.340 166.290 ;
        RECT 96.150 166.090 116.070 166.230 ;
        RECT 108.020 166.030 108.340 166.090 ;
        RECT 81.310 165.750 83.845 165.890 ;
        RECT 86.415 165.890 86.705 165.935 ;
        RECT 88.240 165.890 88.560 165.950 ;
        RECT 90.080 165.890 90.400 165.950 ;
        RECT 115.930 165.935 116.070 166.090 ;
        RECT 92.395 165.890 92.685 165.935 ;
        RECT 86.415 165.750 92.685 165.890 ;
        RECT 81.310 165.705 81.600 165.750 ;
        RECT 86.415 165.705 86.705 165.750 ;
        RECT 88.240 165.690 88.560 165.750 ;
        RECT 90.080 165.690 90.400 165.750 ;
        RECT 92.395 165.705 92.685 165.750 ;
        RECT 93.775 165.705 94.065 165.935 ;
        RECT 115.855 165.705 116.145 165.935 ;
        RECT 72.615 165.365 72.905 165.595 ;
        RECT 84.575 165.550 84.865 165.595 ;
        RECT 84.575 165.410 93.070 165.550 ;
        RECT 84.575 165.365 84.865 165.410 ;
        RECT 61.575 165.210 61.865 165.255 ;
        RECT 61.190 165.070 61.865 165.210 ;
        RECT 55.550 165.025 55.840 165.070 ;
        RECT 58.330 165.025 58.620 165.070 ;
        RECT 60.190 165.025 60.480 165.070 ;
        RECT 61.575 165.025 61.865 165.070 ;
        RECT 72.140 165.210 72.460 165.270 ;
        RECT 72.690 165.210 72.830 165.365 ;
        RECT 92.930 165.255 93.070 165.410 ;
        RECT 72.140 165.070 72.830 165.210 ;
        RECT 81.310 165.210 81.600 165.255 ;
        RECT 84.090 165.210 84.380 165.255 ;
        RECT 85.950 165.210 86.240 165.255 ;
        RECT 81.310 165.070 86.240 165.210 ;
        RECT 72.140 165.010 72.460 165.070 ;
        RECT 81.310 165.025 81.600 165.070 ;
        RECT 84.090 165.025 84.380 165.070 ;
        RECT 85.950 165.025 86.240 165.070 ;
        RECT 92.855 165.025 93.145 165.255 ;
        RECT 70.775 164.870 71.065 164.915 ;
        RECT 76.740 164.870 77.060 164.930 ;
        RECT 77.660 164.915 77.980 164.930 ;
        RECT 47.850 164.730 77.060 164.870 ;
        RECT 70.775 164.685 71.065 164.730 ;
        RECT 76.740 164.670 77.060 164.730 ;
        RECT 77.445 164.870 77.980 164.915 ;
        RECT 78.580 164.870 78.900 164.930 ;
        RECT 77.445 164.730 78.900 164.870 ;
        RECT 77.445 164.685 77.980 164.730 ;
        RECT 77.660 164.670 77.980 164.685 ;
        RECT 78.580 164.670 78.900 164.730 ;
        RECT 80.420 164.870 80.740 164.930 ;
        RECT 93.850 164.870 93.990 165.705 ;
        RECT 118.600 165.690 118.920 165.950 ;
        RECT 96.060 165.550 96.380 165.610 ;
        RECT 108.035 165.550 108.325 165.595 ;
        RECT 96.060 165.410 108.325 165.550 ;
        RECT 96.060 165.350 96.380 165.410 ;
        RECT 108.035 165.365 108.325 165.410 ;
        RECT 108.110 165.210 108.250 165.365 ;
        RECT 108.940 165.350 109.260 165.610 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 110.320 165.210 110.640 165.270 ;
        RECT 108.110 165.070 110.640 165.210 ;
        RECT 110.320 165.010 110.640 165.070 ;
        RECT 80.420 164.730 93.990 164.870 ;
        RECT 102.500 164.870 102.820 164.930 ;
        RECT 102.975 164.870 103.265 164.915 ;
        RECT 102.500 164.730 103.265 164.870 ;
        RECT 80.420 164.670 80.740 164.730 ;
        RECT 102.500 164.670 102.820 164.730 ;
        RECT 102.975 164.685 103.265 164.730 ;
        RECT 115.840 164.870 116.160 164.930 ;
        RECT 116.315 164.870 116.605 164.915 ;
        RECT 115.840 164.730 116.605 164.870 ;
        RECT 115.840 164.670 116.160 164.730 ;
        RECT 116.315 164.685 116.605 164.730 ;
        RECT 119.535 164.870 119.825 164.915 ;
        RECT 120.900 164.870 121.220 164.930 ;
        RECT 119.535 164.730 121.220 164.870 ;
        RECT 119.535 164.685 119.825 164.730 ;
        RECT 120.900 164.670 121.220 164.730 ;
        RECT 11.810 164.050 125.890 164.530 ;
        RECT 32.135 163.850 32.425 163.895 ;
        RECT 32.580 163.850 32.900 163.910 ;
        RECT 32.135 163.710 32.900 163.850 ;
        RECT 32.135 163.665 32.425 163.710 ;
        RECT 32.580 163.650 32.900 163.710 ;
        RECT 33.040 163.850 33.360 163.910 ;
        RECT 33.975 163.850 34.265 163.895 ;
        RECT 62.480 163.850 62.800 163.910 ;
        RECT 33.040 163.710 34.265 163.850 ;
        RECT 33.040 163.650 33.360 163.710 ;
        RECT 33.975 163.665 34.265 163.710 ;
        RECT 59.350 163.710 62.800 163.850 ;
        RECT 55.595 163.510 55.885 163.555 ;
        RECT 59.350 163.510 59.490 163.710 ;
        RECT 62.480 163.650 62.800 163.710 ;
        RECT 70.760 163.850 71.080 163.910 ;
        RECT 71.695 163.850 71.985 163.895 ;
        RECT 70.760 163.710 71.985 163.850 ;
        RECT 70.760 163.650 71.080 163.710 ;
        RECT 71.695 163.665 71.985 163.710 ;
        RECT 72.155 163.665 72.445 163.895 ;
        RECT 55.595 163.370 59.490 163.510 ;
        RECT 60.150 163.510 60.440 163.555 ;
        RECT 62.930 163.510 63.220 163.555 ;
        RECT 64.790 163.510 65.080 163.555 ;
        RECT 60.150 163.370 65.080 163.510 ;
        RECT 55.595 163.325 55.885 163.370 ;
        RECT 60.150 163.325 60.440 163.370 ;
        RECT 62.930 163.325 63.220 163.370 ;
        RECT 64.790 163.325 65.080 163.370 ;
        RECT 68.920 163.510 69.240 163.570 ;
        RECT 72.230 163.510 72.370 163.665 ;
        RECT 80.420 163.650 80.740 163.910 ;
        RECT 98.010 163.850 98.300 163.895 ;
        RECT 99.740 163.850 100.060 163.910 ;
        RECT 98.010 163.710 100.060 163.850 ;
        RECT 98.010 163.665 98.300 163.710 ;
        RECT 99.740 163.650 100.060 163.710 ;
        RECT 72.600 163.510 72.920 163.570 ;
        RECT 68.920 163.370 72.920 163.510 ;
        RECT 68.920 163.310 69.240 163.370 ;
        RECT 72.600 163.310 72.920 163.370 ;
        RECT 84.990 163.510 85.280 163.555 ;
        RECT 87.770 163.510 88.060 163.555 ;
        RECT 89.630 163.510 89.920 163.555 ;
        RECT 84.990 163.370 89.920 163.510 ;
        RECT 84.990 163.325 85.280 163.370 ;
        RECT 87.770 163.325 88.060 163.370 ;
        RECT 89.630 163.325 89.920 163.370 ;
        RECT 93.415 163.510 93.705 163.555 ;
        RECT 96.535 163.510 96.825 163.555 ;
        RECT 98.425 163.510 98.715 163.555 ;
        RECT 93.415 163.370 98.715 163.510 ;
        RECT 93.415 163.325 93.705 163.370 ;
        RECT 96.535 163.325 96.825 163.370 ;
        RECT 98.425 163.325 98.715 163.370 ;
        RECT 116.415 163.510 116.705 163.555 ;
        RECT 119.535 163.510 119.825 163.555 ;
        RECT 121.425 163.510 121.715 163.555 ;
        RECT 116.415 163.370 121.715 163.510 ;
        RECT 116.415 163.325 116.705 163.370 ;
        RECT 119.535 163.325 119.825 163.370 ;
        RECT 121.425 163.325 121.715 163.370 ;
        RECT 27.980 163.170 28.300 163.230 ;
        RECT 28.915 163.170 29.205 163.215 ;
        RECT 45.000 163.170 45.320 163.230 ;
        RECT 52.360 163.170 52.680 163.230 ;
        RECT 27.980 163.030 36.490 163.170 ;
        RECT 27.980 162.970 28.300 163.030 ;
        RECT 28.915 162.985 29.205 163.030 ;
        RECT 34.880 162.630 35.200 162.890 ;
        RECT 36.350 162.875 36.490 163.030 ;
        RECT 45.000 163.030 52.680 163.170 ;
        RECT 45.000 162.970 45.320 163.030 ;
        RECT 52.360 162.970 52.680 163.030 ;
        RECT 53.280 162.970 53.600 163.230 ;
        RECT 60.640 163.170 60.960 163.230 ;
        RECT 70.300 163.170 70.620 163.230 ;
        RECT 60.640 163.030 65.470 163.170 ;
        RECT 60.640 162.970 60.960 163.030 ;
        RECT 65.330 162.890 65.470 163.030 ;
        RECT 69.010 163.030 70.620 163.170 ;
        RECT 35.355 162.645 35.645 162.875 ;
        RECT 36.275 162.645 36.565 162.875 ;
        RECT 35.430 162.490 35.570 162.645 ;
        RECT 36.720 162.630 37.040 162.890 ;
        RECT 37.180 162.630 37.500 162.890 ;
        RECT 41.780 162.830 42.100 162.890 ;
        RECT 38.650 162.690 42.100 162.830 ;
        RECT 38.650 162.490 38.790 162.690 ;
        RECT 41.780 162.630 42.100 162.690 ;
        RECT 60.150 162.830 60.440 162.875 ;
        RECT 60.150 162.690 62.685 162.830 ;
        RECT 60.150 162.645 60.440 162.690 ;
        RECT 35.430 162.350 38.790 162.490 ;
        RECT 39.020 162.290 39.340 162.550 ;
        RECT 47.760 162.290 48.080 162.550 ;
        RECT 53.280 162.490 53.600 162.550 ;
        RECT 56.285 162.490 56.575 162.535 ;
        RECT 53.280 162.350 56.575 162.490 ;
        RECT 53.280 162.290 53.600 162.350 ;
        RECT 56.285 162.305 56.575 162.350 ;
        RECT 57.420 162.490 57.740 162.550 ;
        RECT 62.470 162.535 62.685 162.690 ;
        RECT 63.400 162.630 63.720 162.890 ;
        RECT 65.240 162.630 65.560 162.890 ;
        RECT 69.010 162.875 69.150 163.030 ;
        RECT 70.300 162.970 70.620 163.030 ;
        RECT 71.680 163.170 72.000 163.230 ;
        RECT 73.060 163.170 73.380 163.230 ;
        RECT 71.680 163.030 73.380 163.170 ;
        RECT 71.680 162.970 72.000 163.030 ;
        RECT 73.060 162.970 73.380 163.030 ;
        RECT 77.200 162.970 77.520 163.230 ;
        RECT 78.135 163.170 78.425 163.215 ;
        RECT 78.580 163.170 78.900 163.230 ;
        RECT 78.135 163.030 78.900 163.170 ;
        RECT 78.135 162.985 78.425 163.030 ;
        RECT 78.580 162.970 78.900 163.030 ;
        RECT 90.080 162.970 90.400 163.230 ;
        RECT 90.555 163.170 90.845 163.215 ;
        RECT 97.900 163.170 98.220 163.230 ;
        RECT 99.740 163.170 100.060 163.230 ;
        RECT 90.555 163.030 100.060 163.170 ;
        RECT 90.555 162.985 90.845 163.030 ;
        RECT 97.900 162.970 98.220 163.030 ;
        RECT 99.740 162.970 100.060 163.030 ;
        RECT 101.120 163.170 101.440 163.230 ;
        RECT 101.120 163.030 102.730 163.170 ;
        RECT 101.120 162.970 101.440 163.030 ;
        RECT 68.935 162.645 69.225 162.875 ;
        RECT 69.380 162.630 69.700 162.890 ;
        RECT 70.390 162.830 70.530 162.970 ;
        RECT 71.235 162.830 71.525 162.875 ;
        RECT 70.390 162.690 71.525 162.830 ;
        RECT 71.235 162.645 71.525 162.690 ;
        RECT 72.140 162.830 72.460 162.890 ;
        RECT 72.615 162.830 72.905 162.875 ;
        RECT 72.140 162.690 72.905 162.830 ;
        RECT 72.140 162.630 72.460 162.690 ;
        RECT 72.615 162.645 72.905 162.690 ;
        RECT 84.990 162.830 85.280 162.875 ;
        RECT 84.990 162.690 87.525 162.830 ;
        RECT 84.990 162.645 85.280 162.690 ;
        RECT 87.310 162.535 87.525 162.690 ;
        RECT 88.240 162.630 88.560 162.890 ;
        RECT 92.335 162.535 92.625 162.850 ;
        RECT 93.415 162.830 93.705 162.875 ;
        RECT 96.995 162.830 97.285 162.875 ;
        RECT 98.830 162.830 99.120 162.875 ;
        RECT 93.415 162.690 99.120 162.830 ;
        RECT 93.415 162.645 93.705 162.690 ;
        RECT 96.995 162.645 97.285 162.690 ;
        RECT 98.830 162.645 99.120 162.690 ;
        RECT 99.295 162.645 99.585 162.875 ;
        RECT 101.595 162.645 101.885 162.875 ;
        RECT 58.290 162.490 58.580 162.535 ;
        RECT 61.550 162.490 61.840 162.535 ;
        RECT 57.420 162.350 61.840 162.490 ;
        RECT 57.420 162.290 57.740 162.350 ;
        RECT 58.290 162.305 58.580 162.350 ;
        RECT 61.550 162.305 61.840 162.350 ;
        RECT 62.470 162.490 62.760 162.535 ;
        RECT 64.330 162.490 64.620 162.535 ;
        RECT 62.470 162.350 64.620 162.490 ;
        RECT 62.470 162.305 62.760 162.350 ;
        RECT 64.330 162.305 64.620 162.350 ;
        RECT 83.130 162.490 83.420 162.535 ;
        RECT 86.390 162.490 86.680 162.535 ;
        RECT 87.310 162.490 87.600 162.535 ;
        RECT 89.170 162.490 89.460 162.535 ;
        RECT 83.130 162.350 87.090 162.490 ;
        RECT 83.130 162.305 83.420 162.350 ;
        RECT 86.390 162.305 86.680 162.350 ;
        RECT 34.420 162.150 34.740 162.210 ;
        RECT 38.575 162.150 38.865 162.195 ;
        RECT 34.420 162.010 38.865 162.150 ;
        RECT 34.420 161.950 34.740 162.010 ;
        RECT 38.575 161.965 38.865 162.010 ;
        RECT 53.755 162.150 54.045 162.195 ;
        RECT 56.960 162.150 57.280 162.210 ;
        RECT 53.755 162.010 57.280 162.150 ;
        RECT 53.755 161.965 54.045 162.010 ;
        RECT 56.960 161.950 57.280 162.010 ;
        RECT 66.160 162.150 66.480 162.210 ;
        RECT 68.015 162.150 68.305 162.195 ;
        RECT 66.160 162.010 68.305 162.150 ;
        RECT 66.160 161.950 66.480 162.010 ;
        RECT 68.015 161.965 68.305 162.010 ;
        RECT 70.315 162.150 70.605 162.195 ;
        RECT 73.060 162.150 73.380 162.210 ;
        RECT 70.315 162.010 73.380 162.150 ;
        RECT 70.315 161.965 70.605 162.010 ;
        RECT 73.060 161.950 73.380 162.010 ;
        RECT 78.580 162.150 78.900 162.210 ;
        RECT 81.125 162.150 81.415 162.195 ;
        RECT 78.580 162.010 81.415 162.150 ;
        RECT 86.950 162.150 87.090 162.350 ;
        RECT 87.310 162.350 89.460 162.490 ;
        RECT 87.310 162.305 87.600 162.350 ;
        RECT 89.170 162.305 89.460 162.350 ;
        RECT 92.035 162.490 92.625 162.535 ;
        RECT 92.840 162.490 93.160 162.550 ;
        RECT 95.275 162.490 95.925 162.535 ;
        RECT 99.370 162.490 99.510 162.645 ;
        RECT 92.035 162.350 95.925 162.490 ;
        RECT 92.035 162.305 92.325 162.350 ;
        RECT 92.840 162.290 93.160 162.350 ;
        RECT 95.275 162.305 95.925 162.350 ;
        RECT 98.910 162.350 99.510 162.490 ;
        RECT 101.670 162.490 101.810 162.645 ;
        RECT 102.040 162.630 102.360 162.890 ;
        RECT 102.590 162.875 102.730 163.030 ;
        RECT 103.510 163.030 107.330 163.170 ;
        RECT 103.510 162.875 103.650 163.030 ;
        RECT 107.190 162.890 107.330 163.030 ;
        RECT 120.900 162.970 121.220 163.230 ;
        RECT 102.515 162.645 102.805 162.875 ;
        RECT 103.435 162.645 103.725 162.875 ;
        RECT 103.880 162.830 104.200 162.890 ;
        RECT 105.275 162.830 105.565 162.875 ;
        RECT 103.880 162.690 105.565 162.830 ;
        RECT 103.880 162.630 104.200 162.690 ;
        RECT 105.275 162.645 105.565 162.690 ;
        RECT 105.720 162.630 106.040 162.890 ;
        RECT 106.195 162.830 106.485 162.875 ;
        RECT 106.640 162.830 106.960 162.890 ;
        RECT 106.195 162.690 106.960 162.830 ;
        RECT 106.195 162.645 106.485 162.690 ;
        RECT 106.640 162.630 106.960 162.690 ;
        RECT 107.100 162.630 107.420 162.890 ;
        RECT 103.970 162.490 104.110 162.630 ;
        RECT 115.335 162.535 115.625 162.850 ;
        RECT 116.415 162.830 116.705 162.875 ;
        RECT 119.995 162.830 120.285 162.875 ;
        RECT 121.830 162.830 122.120 162.875 ;
        RECT 116.415 162.690 122.120 162.830 ;
        RECT 116.415 162.645 116.705 162.690 ;
        RECT 119.995 162.645 120.285 162.690 ;
        RECT 121.830 162.645 122.120 162.690 ;
        RECT 122.280 162.830 122.600 162.890 ;
        RECT 123.660 162.830 123.980 162.890 ;
        RECT 122.280 162.690 123.980 162.830 ;
        RECT 122.280 162.630 122.600 162.690 ;
        RECT 123.660 162.630 123.980 162.690 ;
        RECT 101.670 162.350 104.110 162.490 ;
        RECT 115.035 162.490 115.625 162.535 ;
        RECT 115.840 162.490 116.160 162.550 ;
        RECT 118.275 162.490 118.925 162.535 ;
        RECT 115.035 162.350 118.925 162.490 ;
        RECT 89.620 162.150 89.940 162.210 ;
        RECT 86.950 162.010 89.940 162.150 ;
        RECT 78.580 161.950 78.900 162.010 ;
        RECT 81.125 161.965 81.415 162.010 ;
        RECT 89.620 161.950 89.940 162.010 ;
        RECT 90.080 162.150 90.400 162.210 ;
        RECT 93.760 162.150 94.080 162.210 ;
        RECT 98.910 162.150 99.050 162.350 ;
        RECT 115.035 162.305 115.325 162.350 ;
        RECT 115.840 162.290 116.160 162.350 ;
        RECT 118.275 162.305 118.925 162.350 ;
        RECT 90.080 162.010 99.050 162.150 ;
        RECT 90.080 161.950 90.400 162.010 ;
        RECT 93.760 161.950 94.080 162.010 ;
        RECT 100.200 161.950 100.520 162.210 ;
        RECT 103.420 162.150 103.740 162.210 ;
        RECT 103.895 162.150 104.185 162.195 ;
        RECT 103.420 162.010 104.185 162.150 ;
        RECT 103.420 161.950 103.740 162.010 ;
        RECT 103.895 161.965 104.185 162.010 ;
        RECT 112.620 162.150 112.940 162.210 ;
        RECT 113.555 162.150 113.845 162.195 ;
        RECT 112.620 162.010 113.845 162.150 ;
        RECT 112.620 161.950 112.940 162.010 ;
        RECT 113.555 161.965 113.845 162.010 ;
        RECT 11.010 161.330 125.890 161.810 ;
        RECT 21.555 161.130 21.845 161.175 ;
        RECT 23.840 161.130 24.160 161.190 ;
        RECT 21.555 160.990 24.160 161.130 ;
        RECT 21.555 160.945 21.845 160.990 ;
        RECT 23.840 160.930 24.160 160.990 ;
        RECT 27.980 161.130 28.300 161.190 ;
        RECT 30.755 161.130 31.045 161.175 ;
        RECT 27.980 160.990 31.045 161.130 ;
        RECT 27.980 160.930 28.300 160.990 ;
        RECT 30.755 160.945 31.045 160.990 ;
        RECT 33.055 161.130 33.345 161.175 ;
        RECT 34.880 161.130 35.200 161.190 ;
        RECT 33.055 160.990 35.200 161.130 ;
        RECT 33.055 160.945 33.345 160.990 ;
        RECT 34.880 160.930 35.200 160.990 ;
        RECT 53.280 161.130 53.600 161.190 ;
        RECT 58.355 161.130 58.645 161.175 ;
        RECT 53.280 160.990 58.645 161.130 ;
        RECT 53.280 160.930 53.600 160.990 ;
        RECT 58.355 160.945 58.645 160.990 ;
        RECT 60.195 161.130 60.485 161.175 ;
        RECT 68.920 161.130 69.240 161.190 ;
        RECT 75.835 161.130 76.125 161.175 ;
        RECT 76.280 161.130 76.600 161.190 ;
        RECT 77.200 161.130 77.520 161.190 ;
        RECT 60.195 160.990 61.790 161.130 ;
        RECT 60.195 160.945 60.485 160.990 ;
        RECT 41.320 160.790 41.640 160.850 ;
        RECT 37.730 160.650 41.640 160.790 ;
        RECT 22.460 160.450 22.780 160.510 ;
        RECT 31.215 160.450 31.505 160.495 ;
        RECT 20.710 160.310 21.770 160.450 ;
        RECT 20.710 160.155 20.850 160.310 ;
        RECT 20.635 159.925 20.925 160.155 ;
        RECT 21.095 159.925 21.385 160.155 ;
        RECT 21.630 160.110 21.770 160.310 ;
        RECT 22.460 160.310 31.505 160.450 ;
        RECT 22.460 160.250 22.780 160.310 ;
        RECT 31.215 160.265 31.505 160.310 ;
        RECT 36.735 160.450 37.025 160.495 ;
        RECT 37.180 160.450 37.500 160.510 ;
        RECT 37.730 160.495 37.870 160.650 ;
        RECT 41.320 160.590 41.640 160.650 ;
        RECT 47.760 160.790 48.080 160.850 ;
        RECT 60.640 160.790 60.960 160.850 ;
        RECT 47.760 160.650 60.960 160.790 ;
        RECT 47.760 160.590 48.080 160.650 ;
        RECT 36.735 160.310 37.500 160.450 ;
        RECT 36.735 160.265 37.025 160.310 ;
        RECT 37.180 160.250 37.500 160.310 ;
        RECT 37.655 160.265 37.945 160.495 ;
        RECT 38.115 160.265 38.405 160.495 ;
        RECT 38.575 160.450 38.865 160.495 ;
        RECT 42.240 160.450 42.560 160.510 ;
        RECT 51.070 160.495 51.210 160.650 ;
        RECT 60.640 160.590 60.960 160.650 ;
        RECT 38.575 160.310 42.560 160.450 ;
        RECT 38.575 160.265 38.865 160.310 ;
        RECT 22.920 160.110 23.240 160.170 ;
        RECT 24.760 160.110 25.080 160.170 ;
        RECT 30.295 160.110 30.585 160.155 ;
        RECT 33.500 160.110 33.820 160.170 ;
        RECT 21.630 159.970 33.820 160.110 ;
        RECT 38.190 160.110 38.330 160.265 ;
        RECT 42.240 160.250 42.560 160.310 ;
        RECT 50.995 160.265 51.285 160.495 ;
        RECT 52.835 160.265 53.125 160.495 ;
        RECT 53.295 160.265 53.585 160.495 ;
        RECT 39.480 160.110 39.800 160.170 ;
        RECT 38.190 159.970 39.800 160.110 ;
        RECT 21.170 159.770 21.310 159.925 ;
        RECT 22.920 159.910 23.240 159.970 ;
        RECT 24.760 159.910 25.080 159.970 ;
        RECT 30.295 159.925 30.585 159.970 ;
        RECT 33.500 159.910 33.820 159.970 ;
        RECT 39.480 159.910 39.800 159.970 ;
        RECT 33.040 159.770 33.360 159.830 ;
        RECT 11.510 159.630 33.360 159.770 ;
        RECT 11.510 158.410 11.650 159.630 ;
        RECT 33.040 159.570 33.360 159.630 ;
        RECT 45.920 159.770 46.240 159.830 ;
        RECT 52.910 159.770 53.050 160.265 ;
        RECT 53.370 160.110 53.510 160.265 ;
        RECT 53.740 160.250 54.060 160.510 ;
        RECT 54.675 160.450 54.965 160.495 ;
        RECT 55.580 160.450 55.900 160.510 ;
        RECT 58.340 160.450 58.660 160.510 ;
        RECT 61.650 160.495 61.790 160.990 ;
        RECT 68.920 160.990 75.130 161.130 ;
        RECT 68.920 160.930 69.240 160.990 ;
        RECT 72.600 160.790 72.920 160.850 ;
        RECT 74.455 160.790 74.745 160.835 ;
        RECT 72.600 160.650 74.745 160.790 ;
        RECT 74.990 160.790 75.130 160.990 ;
        RECT 75.835 160.990 77.520 161.130 ;
        RECT 75.835 160.945 76.125 160.990 ;
        RECT 76.280 160.930 76.600 160.990 ;
        RECT 77.200 160.930 77.520 160.990 ;
        RECT 78.580 160.930 78.900 161.190 ;
        RECT 79.040 161.130 79.360 161.190 ;
        RECT 84.115 161.130 84.405 161.175 ;
        RECT 79.040 160.990 84.405 161.130 ;
        RECT 79.040 160.930 79.360 160.990 ;
        RECT 84.115 160.945 84.405 160.990 ;
        RECT 85.955 160.945 86.245 161.175 ;
        RECT 78.670 160.790 78.810 160.930 ;
        RECT 83.655 160.790 83.945 160.835 ;
        RECT 74.990 160.650 78.350 160.790 ;
        RECT 78.670 160.650 83.945 160.790 ;
        RECT 72.600 160.590 72.920 160.650 ;
        RECT 74.455 160.605 74.745 160.650 ;
        RECT 54.675 160.310 55.900 160.450 ;
        RECT 54.675 160.265 54.965 160.310 ;
        RECT 55.580 160.250 55.900 160.310 ;
        RECT 57.050 160.310 58.660 160.450 ;
        RECT 54.200 160.110 54.520 160.170 ;
        RECT 53.370 159.970 54.520 160.110 ;
        RECT 54.200 159.910 54.520 159.970 ;
        RECT 56.040 160.110 56.360 160.170 ;
        RECT 57.050 160.155 57.190 160.310 ;
        RECT 58.340 160.250 58.660 160.310 ;
        RECT 61.575 160.265 61.865 160.495 ;
        RECT 66.160 160.250 66.480 160.510 ;
        RECT 68.015 160.450 68.305 160.495 ;
        RECT 69.380 160.450 69.700 160.510 ;
        RECT 68.015 160.310 69.700 160.450 ;
        RECT 68.015 160.265 68.305 160.310 ;
        RECT 69.380 160.250 69.700 160.310 ;
        RECT 69.855 160.450 70.145 160.495 ;
        RECT 70.760 160.450 71.080 160.510 ;
        RECT 69.855 160.310 71.080 160.450 ;
        RECT 69.855 160.265 70.145 160.310 ;
        RECT 70.760 160.250 71.080 160.310 ;
        RECT 71.680 160.450 72.000 160.510 ;
        RECT 72.155 160.450 72.445 160.495 ;
        RECT 71.680 160.310 72.445 160.450 ;
        RECT 71.680 160.250 72.000 160.310 ;
        RECT 72.155 160.265 72.445 160.310 ;
        RECT 76.755 160.265 77.045 160.495 ;
        RECT 56.975 160.110 57.265 160.155 ;
        RECT 56.040 159.970 57.265 160.110 ;
        RECT 56.040 159.910 56.360 159.970 ;
        RECT 56.975 159.925 57.265 159.970 ;
        RECT 57.880 159.910 58.200 160.170 ;
        RECT 71.220 160.110 71.540 160.170 ;
        RECT 76.830 160.110 76.970 160.265 ;
        RECT 77.660 160.250 77.980 160.510 ;
        RECT 78.210 160.495 78.350 160.650 ;
        RECT 83.655 160.605 83.945 160.650 ;
        RECT 78.135 160.265 78.425 160.495 ;
        RECT 78.595 160.265 78.885 160.495 ;
        RECT 86.030 160.450 86.170 160.945 ;
        RECT 88.240 160.930 88.560 161.190 ;
        RECT 89.620 161.130 89.940 161.190 ;
        RECT 92.395 161.130 92.685 161.175 ;
        RECT 89.620 160.990 92.685 161.130 ;
        RECT 89.620 160.930 89.940 160.990 ;
        RECT 92.395 160.945 92.685 160.990 ;
        RECT 107.100 160.930 107.420 161.190 ;
        RECT 108.020 161.130 108.340 161.190 ;
        RECT 114.460 161.130 114.780 161.190 ;
        RECT 114.935 161.130 115.225 161.175 ;
        RECT 108.020 160.990 115.225 161.130 ;
        RECT 108.020 160.930 108.340 160.990 ;
        RECT 114.460 160.930 114.780 160.990 ;
        RECT 114.935 160.945 115.225 160.990 ;
        RECT 116.775 161.130 117.065 161.175 ;
        RECT 118.600 161.130 118.920 161.190 ;
        RECT 116.775 160.990 118.920 161.130 ;
        RECT 116.775 160.945 117.065 160.990 ;
        RECT 118.600 160.930 118.920 160.990 ;
        RECT 88.700 160.790 89.020 160.850 ;
        RECT 94.680 160.790 95.000 160.850 ;
        RECT 95.550 160.790 95.840 160.835 ;
        RECT 98.810 160.790 99.100 160.835 ;
        RECT 88.700 160.650 93.070 160.790 ;
        RECT 88.700 160.590 89.020 160.650 ;
        RECT 89.710 160.495 89.850 160.650 ;
        RECT 92.930 160.495 93.070 160.650 ;
        RECT 94.680 160.650 99.100 160.790 ;
        RECT 94.680 160.590 95.000 160.650 ;
        RECT 95.550 160.605 95.840 160.650 ;
        RECT 98.810 160.605 99.100 160.650 ;
        RECT 99.730 160.790 100.020 160.835 ;
        RECT 101.590 160.790 101.880 160.835 ;
        RECT 99.730 160.650 101.880 160.790 ;
        RECT 99.730 160.605 100.020 160.650 ;
        RECT 101.590 160.605 101.880 160.650 ;
        RECT 105.720 160.790 106.040 160.850 ;
        RECT 107.190 160.790 107.330 160.930 ;
        RECT 105.720 160.650 106.870 160.790 ;
        RECT 107.190 160.650 108.250 160.790 ;
        RECT 87.335 160.450 87.625 160.495 ;
        RECT 86.030 160.310 87.625 160.450 ;
        RECT 87.335 160.265 87.625 160.310 ;
        RECT 89.635 160.265 89.925 160.495 ;
        RECT 90.555 160.265 90.845 160.495 ;
        RECT 92.855 160.450 93.145 160.495 ;
        RECT 93.300 160.450 93.620 160.510 ;
        RECT 92.855 160.310 93.620 160.450 ;
        RECT 92.855 160.265 93.145 160.310 ;
        RECT 71.220 159.970 76.970 160.110 ;
        RECT 77.200 160.110 77.520 160.170 ;
        RECT 78.210 160.110 78.350 160.265 ;
        RECT 77.200 159.970 78.350 160.110 ;
        RECT 71.220 159.910 71.540 159.970 ;
        RECT 77.200 159.910 77.520 159.970 ;
        RECT 65.255 159.770 65.545 159.815 ;
        RECT 77.660 159.770 77.980 159.830 ;
        RECT 78.670 159.770 78.810 160.265 ;
        RECT 81.340 160.110 81.660 160.170 ;
        RECT 82.735 160.110 83.025 160.155 ;
        RECT 81.340 159.970 83.025 160.110 ;
        RECT 81.340 159.910 81.660 159.970 ;
        RECT 82.735 159.925 83.025 159.970 ;
        RECT 84.100 160.110 84.420 160.170 ;
        RECT 90.630 160.110 90.770 160.265 ;
        RECT 93.300 160.250 93.620 160.310 ;
        RECT 97.410 160.450 97.700 160.495 ;
        RECT 99.730 160.450 99.945 160.605 ;
        RECT 105.720 160.590 106.040 160.650 ;
        RECT 97.410 160.310 99.945 160.450 ;
        RECT 103.880 160.450 104.200 160.510 ;
        RECT 106.730 160.495 106.870 160.650 ;
        RECT 106.195 160.450 106.485 160.495 ;
        RECT 103.880 160.310 106.485 160.450 ;
        RECT 97.410 160.265 97.700 160.310 ;
        RECT 103.880 160.250 104.200 160.310 ;
        RECT 106.195 160.265 106.485 160.310 ;
        RECT 106.655 160.265 106.945 160.495 ;
        RECT 107.115 160.450 107.405 160.495 ;
        RECT 107.560 160.450 107.880 160.510 ;
        RECT 108.110 160.495 108.250 160.650 ;
        RECT 107.115 160.310 107.880 160.450 ;
        RECT 107.115 160.265 107.405 160.310 ;
        RECT 107.560 160.250 107.880 160.310 ;
        RECT 108.035 160.265 108.325 160.495 ;
        RECT 112.620 160.450 112.940 160.510 ;
        RECT 114.475 160.450 114.765 160.495 ;
        RECT 112.620 160.310 114.765 160.450 ;
        RECT 112.620 160.250 112.940 160.310 ;
        RECT 114.475 160.265 114.765 160.310 ;
        RECT 115.380 160.450 115.700 160.510 ;
        RECT 117.695 160.450 117.985 160.495 ;
        RECT 115.380 160.310 117.985 160.450 ;
        RECT 115.380 160.250 115.700 160.310 ;
        RECT 117.695 160.265 117.985 160.310 ;
        RECT 119.520 160.250 119.840 160.510 ;
        RECT 84.100 159.970 90.770 160.110 ;
        RECT 84.100 159.910 84.420 159.970 ;
        RECT 100.660 159.910 100.980 160.170 ;
        RECT 102.500 159.910 102.820 160.170 ;
        RECT 110.320 160.110 110.640 160.170 ;
        RECT 113.555 160.110 113.845 160.155 ;
        RECT 110.320 159.970 113.845 160.110 ;
        RECT 110.320 159.910 110.640 159.970 ;
        RECT 113.555 159.925 113.845 159.970 ;
        RECT 45.920 159.630 56.730 159.770 ;
        RECT 45.920 159.570 46.240 159.630 ;
        RECT 23.380 159.230 23.700 159.490 ;
        RECT 39.940 159.230 40.260 159.490 ;
        RECT 50.060 159.430 50.380 159.490 ;
        RECT 51.455 159.430 51.745 159.475 ;
        RECT 50.060 159.290 51.745 159.430 ;
        RECT 50.060 159.230 50.380 159.290 ;
        RECT 51.455 159.245 51.745 159.290 ;
        RECT 52.360 159.430 52.680 159.490 ;
        RECT 56.040 159.430 56.360 159.490 ;
        RECT 52.360 159.290 56.360 159.430 ;
        RECT 56.590 159.430 56.730 159.630 ;
        RECT 57.510 159.630 78.810 159.770 ;
        RECT 97.410 159.770 97.700 159.815 ;
        RECT 100.190 159.770 100.480 159.815 ;
        RECT 102.050 159.770 102.340 159.815 ;
        RECT 97.410 159.630 102.340 159.770 ;
        RECT 57.510 159.430 57.650 159.630 ;
        RECT 65.255 159.585 65.545 159.630 ;
        RECT 77.660 159.570 77.980 159.630 ;
        RECT 97.410 159.585 97.700 159.630 ;
        RECT 100.190 159.585 100.480 159.630 ;
        RECT 102.050 159.585 102.340 159.630 ;
        RECT 56.590 159.290 57.650 159.430 ;
        RECT 52.360 159.230 52.680 159.290 ;
        RECT 56.040 159.230 56.360 159.290 ;
        RECT 62.480 159.230 62.800 159.490 ;
        RECT 66.620 159.430 66.940 159.490 ;
        RECT 67.095 159.430 67.385 159.475 ;
        RECT 66.620 159.290 67.385 159.430 ;
        RECT 66.620 159.230 66.940 159.290 ;
        RECT 67.095 159.245 67.385 159.290 ;
        RECT 71.220 159.230 71.540 159.490 ;
        RECT 76.740 159.430 77.060 159.490 ;
        RECT 79.975 159.430 80.265 159.475 ;
        RECT 76.740 159.290 80.265 159.430 ;
        RECT 76.740 159.230 77.060 159.290 ;
        RECT 79.975 159.245 80.265 159.290 ;
        RECT 89.160 159.230 89.480 159.490 ;
        RECT 91.475 159.430 91.765 159.475 ;
        RECT 91.920 159.430 92.240 159.490 ;
        RECT 91.475 159.290 92.240 159.430 ;
        RECT 91.475 159.245 91.765 159.290 ;
        RECT 91.920 159.230 92.240 159.290 ;
        RECT 93.545 159.430 93.835 159.475 ;
        RECT 94.220 159.430 94.540 159.490 ;
        RECT 93.545 159.290 94.540 159.430 ;
        RECT 93.545 159.245 93.835 159.290 ;
        RECT 94.220 159.230 94.540 159.290 ;
        RECT 99.280 159.430 99.600 159.490 ;
        RECT 104.815 159.430 105.105 159.475 ;
        RECT 99.280 159.290 105.105 159.430 ;
        RECT 99.280 159.230 99.600 159.290 ;
        RECT 104.815 159.245 105.105 159.290 ;
        RECT 118.140 159.230 118.460 159.490 ;
        RECT 120.440 159.230 120.760 159.490 ;
        RECT 11.810 158.610 125.890 159.090 ;
        RECT 13.275 158.410 13.565 158.455 ;
        RECT 11.510 158.270 13.565 158.410 ;
        RECT 13.275 158.225 13.565 158.270 ;
        RECT 29.835 158.410 30.125 158.455 ;
        RECT 31.660 158.410 31.980 158.470 ;
        RECT 33.960 158.410 34.280 158.470 ;
        RECT 29.835 158.270 34.280 158.410 ;
        RECT 29.835 158.225 30.125 158.270 ;
        RECT 31.660 158.210 31.980 158.270 ;
        RECT 33.960 158.210 34.280 158.270 ;
        RECT 37.180 158.410 37.500 158.470 ;
        RECT 76.280 158.410 76.600 158.470 ;
        RECT 81.340 158.410 81.660 158.470 ;
        RECT 37.180 158.270 41.550 158.410 ;
        RECT 37.180 158.210 37.500 158.270 ;
        RECT 16.135 158.070 16.425 158.115 ;
        RECT 19.255 158.070 19.545 158.115 ;
        RECT 21.145 158.070 21.435 158.115 ;
        RECT 16.135 157.930 21.435 158.070 ;
        RECT 16.135 157.885 16.425 157.930 ;
        RECT 19.255 157.885 19.545 157.930 ;
        RECT 21.145 157.885 21.435 157.930 ;
        RECT 22.935 157.885 23.225 158.115 ;
        RECT 35.800 158.070 36.120 158.130 ;
        RECT 40.875 158.070 41.165 158.115 ;
        RECT 35.800 157.930 41.165 158.070 ;
        RECT 20.635 157.730 20.925 157.775 ;
        RECT 23.010 157.730 23.150 157.885 ;
        RECT 35.800 157.870 36.120 157.930 ;
        RECT 40.875 157.885 41.165 157.930 ;
        RECT 39.480 157.730 39.800 157.790 ;
        RECT 20.635 157.590 23.150 157.730 ;
        RECT 38.650 157.590 39.800 157.730 ;
        RECT 41.410 157.730 41.550 158.270 ;
        RECT 76.280 158.270 81.660 158.410 ;
        RECT 76.280 158.210 76.600 158.270 ;
        RECT 81.340 158.210 81.660 158.270 ;
        RECT 84.100 158.210 84.420 158.470 ;
        RECT 88.330 158.270 94.450 158.410 ;
        RECT 60.150 158.070 60.440 158.115 ;
        RECT 62.930 158.070 63.220 158.115 ;
        RECT 64.790 158.070 65.080 158.115 ;
        RECT 60.150 157.930 65.080 158.070 ;
        RECT 60.150 157.885 60.440 157.930 ;
        RECT 62.930 157.885 63.220 157.930 ;
        RECT 64.790 157.885 65.080 157.930 ;
        RECT 81.430 158.070 81.570 158.210 ;
        RECT 88.330 158.070 88.470 158.270 ;
        RECT 81.430 157.930 88.470 158.070 ;
        RECT 88.670 158.070 88.960 158.115 ;
        RECT 91.450 158.070 91.740 158.115 ;
        RECT 93.310 158.070 93.600 158.115 ;
        RECT 88.670 157.930 93.600 158.070 ;
        RECT 41.410 157.590 47.990 157.730 ;
        RECT 20.635 157.545 20.925 157.590 ;
        RECT 13.720 157.050 14.040 157.110 ;
        RECT 15.055 157.095 15.345 157.410 ;
        RECT 16.135 157.390 16.425 157.435 ;
        RECT 19.715 157.390 20.005 157.435 ;
        RECT 21.550 157.390 21.840 157.435 ;
        RECT 16.135 157.250 21.840 157.390 ;
        RECT 16.135 157.205 16.425 157.250 ;
        RECT 19.715 157.205 20.005 157.250 ;
        RECT 21.550 157.205 21.840 157.250 ;
        RECT 22.000 157.190 22.320 157.450 ;
        RECT 23.380 157.390 23.700 157.450 ;
        RECT 23.855 157.390 24.145 157.435 ;
        RECT 23.380 157.250 24.145 157.390 ;
        RECT 23.380 157.190 23.700 157.250 ;
        RECT 23.855 157.205 24.145 157.250 ;
        RECT 26.155 157.390 26.445 157.435 ;
        RECT 30.280 157.390 30.600 157.450 ;
        RECT 26.155 157.250 30.600 157.390 ;
        RECT 26.155 157.205 26.445 157.250 ;
        RECT 30.280 157.190 30.600 157.250 ;
        RECT 36.260 157.190 36.580 157.450 ;
        RECT 37.180 157.190 37.500 157.450 ;
        RECT 38.100 157.190 38.420 157.450 ;
        RECT 38.650 157.435 38.790 157.590 ;
        RECT 39.480 157.530 39.800 157.590 ;
        RECT 38.575 157.205 38.865 157.435 ;
        RECT 39.035 157.390 39.325 157.435 ;
        RECT 42.240 157.390 42.560 157.450 ;
        RECT 39.035 157.250 42.560 157.390 ;
        RECT 39.035 157.205 39.325 157.250 ;
        RECT 14.755 157.050 15.345 157.095 ;
        RECT 17.995 157.050 18.645 157.095 ;
        RECT 13.720 156.910 18.645 157.050 ;
        RECT 38.650 157.050 38.790 157.205 ;
        RECT 42.240 157.190 42.560 157.250 ;
        RECT 42.715 157.205 43.005 157.435 ;
        RECT 43.175 157.390 43.465 157.435 ;
        RECT 43.620 157.390 43.940 157.450 ;
        RECT 44.170 157.435 44.310 157.590 ;
        RECT 47.850 157.450 47.990 157.590 ;
        RECT 52.360 157.530 52.680 157.790 ;
        RECT 53.280 157.530 53.600 157.790 ;
        RECT 56.960 157.730 57.280 157.790 ;
        RECT 57.880 157.730 58.200 157.790 ;
        RECT 56.960 157.590 58.200 157.730 ;
        RECT 56.960 157.530 57.280 157.590 ;
        RECT 57.880 157.530 58.200 157.590 ;
        RECT 62.480 157.730 62.800 157.790 ;
        RECT 81.430 157.775 81.570 157.930 ;
        RECT 88.670 157.885 88.960 157.930 ;
        RECT 91.450 157.885 91.740 157.930 ;
        RECT 93.310 157.885 93.600 157.930 ;
        RECT 63.415 157.730 63.705 157.775 ;
        RECT 62.480 157.590 63.705 157.730 ;
        RECT 62.480 157.530 62.800 157.590 ;
        RECT 63.415 157.545 63.705 157.590 ;
        RECT 81.355 157.545 81.645 157.775 ;
        RECT 91.920 157.530 92.240 157.790 ;
        RECT 93.760 157.530 94.080 157.790 ;
        RECT 94.310 157.730 94.450 158.270 ;
        RECT 94.680 158.210 95.000 158.470 ;
        RECT 100.660 158.410 100.980 158.470 ;
        RECT 101.135 158.410 101.425 158.455 ;
        RECT 119.520 158.410 119.840 158.470 ;
        RECT 96.610 158.270 99.970 158.410 ;
        RECT 96.060 157.730 96.380 157.790 ;
        RECT 94.310 157.590 96.380 157.730 ;
        RECT 96.060 157.530 96.380 157.590 ;
        RECT 43.175 157.250 43.940 157.390 ;
        RECT 43.175 157.205 43.465 157.250 ;
        RECT 42.790 157.050 42.930 157.205 ;
        RECT 43.620 157.190 43.940 157.250 ;
        RECT 44.095 157.205 44.385 157.435 ;
        RECT 45.920 157.190 46.240 157.450 ;
        RECT 46.395 157.205 46.685 157.435 ;
        RECT 46.855 157.390 47.145 157.435 ;
        RECT 47.300 157.390 47.620 157.450 ;
        RECT 46.855 157.250 47.620 157.390 ;
        RECT 46.855 157.205 47.145 157.250 ;
        RECT 45.460 157.050 45.780 157.110 ;
        RECT 46.470 157.050 46.610 157.205 ;
        RECT 47.300 157.190 47.620 157.250 ;
        RECT 47.760 157.190 48.080 157.450 ;
        RECT 60.150 157.390 60.440 157.435 ;
        RECT 60.150 157.250 62.685 157.390 ;
        RECT 60.150 157.205 60.440 157.250 ;
        RECT 48.220 157.050 48.540 157.110 ;
        RECT 38.650 156.910 48.540 157.050 ;
        RECT 13.720 156.850 14.040 156.910 ;
        RECT 14.755 156.865 15.045 156.910 ;
        RECT 17.995 156.865 18.645 156.910 ;
        RECT 45.460 156.850 45.780 156.910 ;
        RECT 48.220 156.850 48.540 156.910 ;
        RECT 53.280 157.050 53.600 157.110 ;
        RECT 56.285 157.050 56.575 157.095 ;
        RECT 56.960 157.050 57.280 157.110 ;
        RECT 53.280 156.910 57.280 157.050 ;
        RECT 53.280 156.850 53.600 156.910 ;
        RECT 56.285 156.865 56.575 156.910 ;
        RECT 56.960 156.850 57.280 156.910 ;
        RECT 58.290 157.050 58.580 157.095 ;
        RECT 58.800 157.050 59.120 157.110 ;
        RECT 62.470 157.095 62.685 157.250 ;
        RECT 65.240 157.190 65.560 157.450 ;
        RECT 66.160 157.390 66.480 157.450 ;
        RECT 66.635 157.390 66.925 157.435 ;
        RECT 66.160 157.250 66.925 157.390 ;
        RECT 66.160 157.190 66.480 157.250 ;
        RECT 66.635 157.205 66.925 157.250 ;
        RECT 68.475 157.390 68.765 157.435 ;
        RECT 70.760 157.390 71.080 157.450 ;
        RECT 68.475 157.250 71.080 157.390 ;
        RECT 68.475 157.205 68.765 157.250 ;
        RECT 70.760 157.190 71.080 157.250 ;
        RECT 71.680 157.390 72.000 157.450 ;
        RECT 72.615 157.390 72.905 157.435 ;
        RECT 71.680 157.250 72.905 157.390 ;
        RECT 71.680 157.190 72.000 157.250 ;
        RECT 72.615 157.205 72.905 157.250 ;
        RECT 77.660 157.190 77.980 157.450 ;
        RECT 78.135 157.205 78.425 157.435 ;
        RECT 61.550 157.050 61.840 157.095 ;
        RECT 58.290 156.910 61.840 157.050 ;
        RECT 58.290 156.865 58.580 156.910 ;
        RECT 58.800 156.850 59.120 156.910 ;
        RECT 61.550 156.865 61.840 156.910 ;
        RECT 62.470 157.050 62.760 157.095 ;
        RECT 64.330 157.050 64.620 157.095 ;
        RECT 62.470 156.910 64.620 157.050 ;
        RECT 62.470 156.865 62.760 156.910 ;
        RECT 64.330 156.865 64.620 156.910 ;
        RECT 76.280 156.850 76.600 157.110 ;
        RECT 77.200 157.050 77.520 157.110 ;
        RECT 78.210 157.050 78.350 157.205 ;
        RECT 78.580 157.190 78.900 157.450 ;
        RECT 79.515 157.390 79.805 157.435 ;
        RECT 79.960 157.390 80.280 157.450 ;
        RECT 79.515 157.250 80.280 157.390 ;
        RECT 79.515 157.205 79.805 157.250 ;
        RECT 79.960 157.190 80.280 157.250 ;
        RECT 88.670 157.390 88.960 157.435 ;
        RECT 93.300 157.390 93.620 157.450 ;
        RECT 94.235 157.390 94.525 157.435 ;
        RECT 96.610 157.390 96.750 158.270 ;
        RECT 99.295 157.885 99.585 158.115 ;
        RECT 99.830 158.070 99.970 158.270 ;
        RECT 100.660 158.270 101.425 158.410 ;
        RECT 100.660 158.210 100.980 158.270 ;
        RECT 101.135 158.225 101.425 158.270 ;
        RECT 118.230 158.270 119.840 158.410 ;
        RECT 114.015 158.070 114.305 158.115 ;
        RECT 118.230 158.070 118.370 158.270 ;
        RECT 119.520 158.210 119.840 158.270 ;
        RECT 99.830 157.930 111.470 158.070 ;
        RECT 88.670 157.250 91.205 157.390 ;
        RECT 88.670 157.205 88.960 157.250 ;
        RECT 82.275 157.050 82.565 157.095 ;
        RECT 86.810 157.050 87.100 157.095 ;
        RECT 89.160 157.050 89.480 157.110 ;
        RECT 90.990 157.095 91.205 157.250 ;
        RECT 93.300 157.250 96.750 157.390 ;
        RECT 99.370 157.390 99.510 157.885 ;
        RECT 105.735 157.730 106.025 157.775 ;
        RECT 101.210 157.590 106.025 157.730 ;
        RECT 100.215 157.390 100.505 157.435 ;
        RECT 99.370 157.250 100.505 157.390 ;
        RECT 93.300 157.190 93.620 157.250 ;
        RECT 94.235 157.205 94.525 157.250 ;
        RECT 100.215 157.205 100.505 157.250 ;
        RECT 90.070 157.050 90.360 157.095 ;
        RECT 77.200 156.910 78.350 157.050 ;
        RECT 78.670 156.910 86.630 157.050 ;
        RECT 77.200 156.850 77.520 156.910 ;
        RECT 26.615 156.710 26.905 156.755 ;
        RECT 27.060 156.710 27.380 156.770 ;
        RECT 26.615 156.570 27.380 156.710 ;
        RECT 26.615 156.525 26.905 156.570 ;
        RECT 27.060 156.510 27.380 156.570 ;
        RECT 37.180 156.710 37.500 156.770 ;
        RECT 38.560 156.710 38.880 156.770 ;
        RECT 37.180 156.570 38.880 156.710 ;
        RECT 37.180 156.510 37.500 156.570 ;
        RECT 38.560 156.510 38.880 156.570 ;
        RECT 40.415 156.710 40.705 156.755 ;
        RECT 42.700 156.710 43.020 156.770 ;
        RECT 40.415 156.570 43.020 156.710 ;
        RECT 40.415 156.525 40.705 156.570 ;
        RECT 42.700 156.510 43.020 156.570 ;
        RECT 44.540 156.510 44.860 156.770 ;
        RECT 46.840 156.710 47.160 156.770 ;
        RECT 49.600 156.710 49.920 156.770 ;
        RECT 53.755 156.710 54.045 156.755 ;
        RECT 46.840 156.570 54.045 156.710 ;
        RECT 46.840 156.510 47.160 156.570 ;
        RECT 49.600 156.510 49.920 156.570 ;
        RECT 53.755 156.525 54.045 156.570 ;
        RECT 55.595 156.710 55.885 156.755 ;
        RECT 59.260 156.710 59.580 156.770 ;
        RECT 55.595 156.570 59.580 156.710 ;
        RECT 55.595 156.525 55.885 156.570 ;
        RECT 59.260 156.510 59.580 156.570 ;
        RECT 67.540 156.510 67.860 156.770 ;
        RECT 69.395 156.710 69.685 156.755 ;
        RECT 69.840 156.710 70.160 156.770 ;
        RECT 69.395 156.570 70.160 156.710 ;
        RECT 69.395 156.525 69.685 156.570 ;
        RECT 69.840 156.510 70.160 156.570 ;
        RECT 70.300 156.710 70.620 156.770 ;
        RECT 71.695 156.710 71.985 156.755 ;
        RECT 70.300 156.570 71.985 156.710 ;
        RECT 70.300 156.510 70.620 156.570 ;
        RECT 71.695 156.525 71.985 156.570 ;
        RECT 73.980 156.710 74.300 156.770 ;
        RECT 78.670 156.710 78.810 156.910 ;
        RECT 82.275 156.865 82.565 156.910 ;
        RECT 73.980 156.570 78.810 156.710 ;
        RECT 79.040 156.710 79.360 156.770 ;
        RECT 81.815 156.710 82.105 156.755 ;
        RECT 84.805 156.710 85.095 156.755 ;
        RECT 79.040 156.570 85.095 156.710 ;
        RECT 86.490 156.710 86.630 156.910 ;
        RECT 86.810 156.910 90.360 157.050 ;
        RECT 86.810 156.865 87.100 156.910 ;
        RECT 89.160 156.850 89.480 156.910 ;
        RECT 90.070 156.865 90.360 156.910 ;
        RECT 90.990 157.050 91.280 157.095 ;
        RECT 92.850 157.050 93.140 157.095 ;
        RECT 90.990 156.910 93.140 157.050 ;
        RECT 90.990 156.865 91.280 156.910 ;
        RECT 92.850 156.865 93.140 156.910 ;
        RECT 96.060 157.050 96.380 157.110 ;
        RECT 101.210 157.050 101.350 157.590 ;
        RECT 105.735 157.545 106.025 157.590 ;
        RECT 110.320 157.730 110.640 157.790 ;
        RECT 110.795 157.730 111.085 157.775 ;
        RECT 110.320 157.590 111.085 157.730 ;
        RECT 111.330 157.730 111.470 157.930 ;
        RECT 114.015 157.930 118.370 158.070 ;
        RECT 118.570 158.070 118.860 158.115 ;
        RECT 121.350 158.070 121.640 158.115 ;
        RECT 123.210 158.070 123.500 158.115 ;
        RECT 118.570 157.930 123.500 158.070 ;
        RECT 114.015 157.885 114.305 157.930 ;
        RECT 118.570 157.885 118.860 157.930 ;
        RECT 121.350 157.885 121.640 157.930 ;
        RECT 123.210 157.885 123.500 157.930 ;
        RECT 115.380 157.730 115.700 157.790 ;
        RECT 111.330 157.590 115.700 157.730 ;
        RECT 110.320 157.530 110.640 157.590 ;
        RECT 110.795 157.545 111.085 157.590 ;
        RECT 115.380 157.530 115.700 157.590 ;
        RECT 120.440 157.730 120.760 157.790 ;
        RECT 121.835 157.730 122.125 157.775 ;
        RECT 120.440 157.590 122.125 157.730 ;
        RECT 120.440 157.530 120.760 157.590 ;
        RECT 121.835 157.545 122.125 157.590 ;
        RECT 106.640 157.390 106.960 157.450 ;
        RECT 107.115 157.390 107.405 157.435 ;
        RECT 96.060 156.910 101.350 157.050 ;
        RECT 102.130 157.250 105.950 157.390 ;
        RECT 96.060 156.850 96.380 156.910 ;
        RECT 94.220 156.710 94.540 156.770 ;
        RECT 96.995 156.710 97.285 156.755 ;
        RECT 86.490 156.570 97.285 156.710 ;
        RECT 73.980 156.510 74.300 156.570 ;
        RECT 79.040 156.510 79.360 156.570 ;
        RECT 81.815 156.525 82.105 156.570 ;
        RECT 84.805 156.525 85.095 156.570 ;
        RECT 94.220 156.510 94.540 156.570 ;
        RECT 96.995 156.525 97.285 156.570 ;
        RECT 97.455 156.710 97.745 156.755 ;
        RECT 98.360 156.710 98.680 156.770 ;
        RECT 102.130 156.710 102.270 157.250 ;
        RECT 102.500 157.050 102.820 157.110 ;
        RECT 104.355 157.050 104.645 157.095 ;
        RECT 102.500 156.910 104.645 157.050 ;
        RECT 105.810 157.050 105.950 157.250 ;
        RECT 106.640 157.250 107.405 157.390 ;
        RECT 106.640 157.190 106.960 157.250 ;
        RECT 107.115 157.205 107.405 157.250 ;
        RECT 107.560 157.190 107.880 157.450 ;
        RECT 108.020 157.190 108.340 157.450 ;
        RECT 108.955 157.390 109.245 157.435 ;
        RECT 109.400 157.390 109.720 157.450 ;
        RECT 108.955 157.250 109.720 157.390 ;
        RECT 108.955 157.205 109.245 157.250 ;
        RECT 109.400 157.190 109.720 157.250 ;
        RECT 111.715 157.390 112.005 157.435 ;
        RECT 114.705 157.390 114.995 157.435 ;
        RECT 111.715 157.250 114.995 157.390 ;
        RECT 111.715 157.205 112.005 157.250 ;
        RECT 114.705 157.205 114.995 157.250 ;
        RECT 118.570 157.390 118.860 157.435 ;
        RECT 118.570 157.250 121.105 157.390 ;
        RECT 118.570 157.205 118.860 157.250 ;
        RECT 111.790 157.050 111.930 157.205 ;
        RECT 105.810 156.910 111.930 157.050 ;
        RECT 102.500 156.850 102.820 156.910 ;
        RECT 104.355 156.865 104.645 156.910 ;
        RECT 97.455 156.570 102.270 156.710 ;
        RECT 104.430 156.710 104.570 156.865 ;
        RECT 112.160 156.850 112.480 157.110 ;
        RECT 116.710 157.050 117.000 157.095 ;
        RECT 118.140 157.050 118.460 157.110 ;
        RECT 120.890 157.095 121.105 157.250 ;
        RECT 123.660 157.190 123.980 157.450 ;
        RECT 119.970 157.050 120.260 157.095 ;
        RECT 116.710 156.910 120.260 157.050 ;
        RECT 116.710 156.865 117.000 156.910 ;
        RECT 118.140 156.850 118.460 156.910 ;
        RECT 119.970 156.865 120.260 156.910 ;
        RECT 120.890 157.050 121.180 157.095 ;
        RECT 122.750 157.050 123.040 157.095 ;
        RECT 120.890 156.910 123.040 157.050 ;
        RECT 120.890 156.865 121.180 156.910 ;
        RECT 122.750 156.865 123.040 156.910 ;
        RECT 123.660 156.710 123.980 156.770 ;
        RECT 104.430 156.570 123.980 156.710 ;
        RECT 97.455 156.525 97.745 156.570 ;
        RECT 98.360 156.510 98.680 156.570 ;
        RECT 123.660 156.510 123.980 156.570 ;
        RECT 11.010 155.890 125.890 156.370 ;
        RECT 13.720 155.490 14.040 155.750 ;
        RECT 14.655 155.690 14.945 155.735 ;
        RECT 14.655 155.550 21.770 155.690 ;
        RECT 14.655 155.505 14.945 155.550 ;
        RECT 21.630 155.410 21.770 155.550 ;
        RECT 45.920 155.490 46.240 155.750 ;
        RECT 51.440 155.690 51.760 155.750 ;
        RECT 51.440 155.550 53.050 155.690 ;
        RECT 51.440 155.490 51.760 155.550 ;
        RECT 16.135 155.350 16.425 155.395 ;
        RECT 19.375 155.350 20.025 155.395 ;
        RECT 16.135 155.210 20.025 155.350 ;
        RECT 16.135 155.165 16.725 155.210 ;
        RECT 19.375 155.165 20.025 155.210 ;
        RECT 21.540 155.350 21.860 155.410 ;
        RECT 22.460 155.350 22.780 155.410 ;
        RECT 21.540 155.210 22.780 155.350 ;
        RECT 16.435 155.070 16.725 155.165 ;
        RECT 21.540 155.150 21.860 155.210 ;
        RECT 22.460 155.150 22.780 155.210 ;
        RECT 27.635 155.350 27.925 155.395 ;
        RECT 30.875 155.350 31.525 155.395 ;
        RECT 27.635 155.210 31.525 155.350 ;
        RECT 27.635 155.165 28.225 155.210 ;
        RECT 30.875 155.165 31.525 155.210 ;
        RECT 27.935 155.070 28.225 155.165 ;
        RECT 33.500 155.150 33.820 155.410 ;
        RECT 33.960 155.350 34.280 155.410 ;
        RECT 42.240 155.350 42.560 155.410 ;
        RECT 46.010 155.350 46.150 155.490 ;
        RECT 52.910 155.350 53.050 155.550 ;
        RECT 57.420 155.490 57.740 155.750 ;
        RECT 58.800 155.490 59.120 155.750 ;
        RECT 60.655 155.690 60.945 155.735 ;
        RECT 63.400 155.690 63.720 155.750 ;
        RECT 72.600 155.690 72.920 155.750 ;
        RECT 97.900 155.690 98.220 155.750 ;
        RECT 107.560 155.690 107.880 155.750 ;
        RECT 60.655 155.550 63.720 155.690 ;
        RECT 60.655 155.505 60.945 155.550 ;
        RECT 63.400 155.490 63.720 155.550 ;
        RECT 66.480 155.550 71.450 155.690 ;
        RECT 66.480 155.350 66.620 155.550 ;
        RECT 71.310 155.410 71.450 155.550 ;
        RECT 72.600 155.550 98.220 155.690 ;
        RECT 72.600 155.490 72.920 155.550 ;
        RECT 97.900 155.490 98.220 155.550 ;
        RECT 107.190 155.550 107.880 155.690 ;
        RECT 33.960 155.210 35.110 155.350 ;
        RECT 33.960 155.150 34.280 155.210 ;
        RECT 14.180 154.810 14.500 155.070 ;
        RECT 16.435 154.850 16.800 155.070 ;
        RECT 16.480 154.810 16.800 154.850 ;
        RECT 17.515 155.010 17.805 155.055 ;
        RECT 21.095 155.010 21.385 155.055 ;
        RECT 22.930 155.010 23.220 155.055 ;
        RECT 17.515 154.870 23.220 155.010 ;
        RECT 17.515 154.825 17.805 154.870 ;
        RECT 21.095 154.825 21.385 154.870 ;
        RECT 22.930 154.825 23.220 154.870 ;
        RECT 24.760 155.010 25.080 155.070 ;
        RECT 25.695 155.010 25.985 155.055 ;
        RECT 24.760 154.870 25.985 155.010 ;
        RECT 24.760 154.810 25.080 154.870 ;
        RECT 25.695 154.825 25.985 154.870 ;
        RECT 27.935 154.850 28.300 155.070 ;
        RECT 27.980 154.810 28.300 154.850 ;
        RECT 29.015 155.010 29.305 155.055 ;
        RECT 32.595 155.010 32.885 155.055 ;
        RECT 34.430 155.010 34.720 155.055 ;
        RECT 29.015 154.870 34.720 155.010 ;
        RECT 29.015 154.825 29.305 154.870 ;
        RECT 32.595 154.825 32.885 154.870 ;
        RECT 34.430 154.825 34.720 154.870 ;
        RECT 34.970 155.010 35.110 155.210 ;
        RECT 42.240 155.210 46.150 155.350 ;
        RECT 48.770 155.210 52.590 155.350 ;
        RECT 52.910 155.210 66.620 155.350 ;
        RECT 71.220 155.350 71.540 155.410 ;
        RECT 97.990 155.350 98.130 155.490 ;
        RECT 107.190 155.350 107.330 155.550 ;
        RECT 107.560 155.490 107.880 155.550 ;
        RECT 112.160 155.350 112.480 155.410 ;
        RECT 71.220 155.210 80.190 155.350 ;
        RECT 97.990 155.210 107.330 155.350 ;
        RECT 42.240 155.150 42.560 155.210 ;
        RECT 36.720 155.010 37.040 155.070 ;
        RECT 45.090 155.055 45.230 155.210 ;
        RECT 38.115 155.010 38.405 155.055 ;
        RECT 34.970 154.870 38.405 155.010 ;
        RECT 19.240 154.670 19.560 154.730 ;
        RECT 22.015 154.670 22.305 154.715 ;
        RECT 19.240 154.530 22.305 154.670 ;
        RECT 19.240 154.470 19.560 154.530 ;
        RECT 22.015 154.485 22.305 154.530 ;
        RECT 23.380 154.670 23.700 154.730 ;
        RECT 34.970 154.715 35.110 154.870 ;
        RECT 36.720 154.810 37.040 154.870 ;
        RECT 38.115 154.825 38.405 154.870 ;
        RECT 45.015 154.825 45.305 155.055 ;
        RECT 45.460 154.810 45.780 155.070 ;
        RECT 45.935 155.010 46.225 155.055 ;
        RECT 46.380 155.010 46.700 155.070 ;
        RECT 45.935 154.870 46.700 155.010 ;
        RECT 45.935 154.825 46.225 154.870 ;
        RECT 46.380 154.810 46.700 154.870 ;
        RECT 46.855 155.010 47.145 155.055 ;
        RECT 47.760 155.010 48.080 155.070 ;
        RECT 48.770 155.055 48.910 155.210 ;
        RECT 52.450 155.070 52.590 155.210 ;
        RECT 71.220 155.150 71.540 155.210 ;
        RECT 46.855 154.870 48.450 155.010 ;
        RECT 46.855 154.825 47.145 154.870 ;
        RECT 47.760 154.810 48.080 154.870 ;
        RECT 34.895 154.670 35.185 154.715 ;
        RECT 23.380 154.530 35.185 154.670 ;
        RECT 23.380 154.470 23.700 154.530 ;
        RECT 34.895 154.485 35.185 154.530 ;
        RECT 17.515 154.330 17.805 154.375 ;
        RECT 20.635 154.330 20.925 154.375 ;
        RECT 22.525 154.330 22.815 154.375 ;
        RECT 17.515 154.190 22.815 154.330 ;
        RECT 17.515 154.145 17.805 154.190 ;
        RECT 20.635 154.145 20.925 154.190 ;
        RECT 22.525 154.145 22.815 154.190 ;
        RECT 29.015 154.330 29.305 154.375 ;
        RECT 32.135 154.330 32.425 154.375 ;
        RECT 34.025 154.330 34.315 154.375 ;
        RECT 29.015 154.190 34.315 154.330 ;
        RECT 29.015 154.145 29.305 154.190 ;
        RECT 32.135 154.145 32.425 154.190 ;
        RECT 34.025 154.145 34.315 154.190 ;
        RECT 35.340 154.330 35.660 154.390 ;
        RECT 48.310 154.330 48.450 154.870 ;
        RECT 48.695 154.825 48.985 155.055 ;
        RECT 49.155 154.825 49.445 155.055 ;
        RECT 49.230 154.670 49.370 154.825 ;
        RECT 49.600 154.810 49.920 155.070 ;
        RECT 50.535 155.010 50.825 155.055 ;
        RECT 51.440 155.010 51.760 155.070 ;
        RECT 50.535 154.870 51.760 155.010 ;
        RECT 50.535 154.825 50.825 154.870 ;
        RECT 51.440 154.810 51.760 154.870 ;
        RECT 52.360 154.810 52.680 155.070 ;
        RECT 52.835 154.825 53.125 155.055 ;
        RECT 53.295 155.010 53.585 155.055 ;
        RECT 53.740 155.010 54.060 155.070 ;
        RECT 53.295 154.870 54.060 155.010 ;
        RECT 53.295 154.825 53.585 154.870 ;
        RECT 51.900 154.670 52.220 154.730 ;
        RECT 52.910 154.670 53.050 154.825 ;
        RECT 53.740 154.810 54.060 154.870 ;
        RECT 54.215 155.010 54.505 155.055 ;
        RECT 55.580 155.010 55.900 155.070 ;
        RECT 54.215 154.870 55.900 155.010 ;
        RECT 54.215 154.825 54.505 154.870 ;
        RECT 55.580 154.810 55.900 154.870 ;
        RECT 56.960 155.010 57.280 155.070 ;
        RECT 58.355 155.010 58.645 155.055 ;
        RECT 56.960 154.870 58.645 155.010 ;
        RECT 56.960 154.810 57.280 154.870 ;
        RECT 58.355 154.825 58.645 154.870 ;
        RECT 59.260 155.010 59.580 155.070 ;
        RECT 59.735 155.010 60.025 155.055 ;
        RECT 59.260 154.870 60.025 155.010 ;
        RECT 59.260 154.810 59.580 154.870 ;
        RECT 59.735 154.825 60.025 154.870 ;
        RECT 62.020 155.010 62.340 155.070 ;
        RECT 68.935 155.010 69.225 155.055 ;
        RECT 62.020 154.870 69.225 155.010 ;
        RECT 62.020 154.810 62.340 154.870 ;
        RECT 49.230 154.530 53.050 154.670 ;
        RECT 51.900 154.470 52.220 154.530 ;
        RECT 51.440 154.330 51.760 154.390 ;
        RECT 35.340 154.190 47.990 154.330 ;
        RECT 48.310 154.190 51.760 154.330 ;
        RECT 35.340 154.130 35.660 154.190 ;
        RECT 24.300 153.990 24.620 154.050 ;
        RECT 24.775 153.990 25.065 154.035 ;
        RECT 24.300 153.850 25.065 153.990 ;
        RECT 24.300 153.790 24.620 153.850 ;
        RECT 24.775 153.805 25.065 153.850 ;
        RECT 26.155 153.990 26.445 154.035 ;
        RECT 27.520 153.990 27.840 154.050 ;
        RECT 26.155 153.850 27.840 153.990 ;
        RECT 26.155 153.805 26.445 153.850 ;
        RECT 27.520 153.790 27.840 153.850 ;
        RECT 34.880 153.990 35.200 154.050 ;
        RECT 38.100 153.990 38.420 154.050 ;
        RECT 34.880 153.850 38.420 153.990 ;
        RECT 34.880 153.790 35.200 153.850 ;
        RECT 38.100 153.790 38.420 153.850 ;
        RECT 42.240 153.990 42.560 154.050 ;
        RECT 43.635 153.990 43.925 154.035 ;
        RECT 42.240 153.850 43.925 153.990 ;
        RECT 42.240 153.790 42.560 153.850 ;
        RECT 43.635 153.805 43.925 153.850 ;
        RECT 47.300 153.790 47.620 154.050 ;
        RECT 47.850 153.990 47.990 154.190 ;
        RECT 51.440 154.130 51.760 154.190 ;
        RECT 50.995 153.990 51.285 154.035 ;
        RECT 47.850 153.850 51.285 153.990 ;
        RECT 67.170 153.990 67.310 154.870 ;
        RECT 68.935 154.825 69.225 154.870 ;
        RECT 69.840 155.010 70.160 155.070 ;
        RECT 72.600 155.010 72.920 155.070 ;
        RECT 73.150 155.055 73.290 155.210 ;
        RECT 80.050 155.070 80.190 155.210 ;
        RECT 69.840 154.870 72.920 155.010 ;
        RECT 69.840 154.810 70.160 154.870 ;
        RECT 72.600 154.810 72.920 154.870 ;
        RECT 73.075 154.825 73.365 155.055 ;
        RECT 73.980 154.810 74.300 155.070 ;
        RECT 74.455 154.825 74.745 155.055 ;
        RECT 74.915 155.010 75.205 155.055 ;
        RECT 77.660 155.010 77.980 155.070 ;
        RECT 78.135 155.010 78.425 155.055 ;
        RECT 74.915 154.870 78.425 155.010 ;
        RECT 74.915 154.825 75.205 154.870 ;
        RECT 68.000 154.470 68.320 154.730 ;
        RECT 74.530 154.670 74.670 154.825 ;
        RECT 77.660 154.810 77.980 154.870 ;
        RECT 78.135 154.825 78.425 154.870 ;
        RECT 78.595 154.825 78.885 155.055 ;
        RECT 77.200 154.670 77.520 154.730 ;
        RECT 78.670 154.670 78.810 154.825 ;
        RECT 79.040 154.810 79.360 155.070 ;
        RECT 79.960 154.810 80.280 155.070 ;
        RECT 98.820 155.010 99.140 155.070 ;
        RECT 103.050 155.055 103.190 155.210 ;
        RECT 107.190 155.070 107.330 155.210 ;
        RECT 107.650 155.210 112.480 155.350 ;
        RECT 101.595 155.010 101.885 155.055 ;
        RECT 98.820 154.870 101.885 155.010 ;
        RECT 98.820 154.810 99.140 154.870 ;
        RECT 101.595 154.825 101.885 154.870 ;
        RECT 102.515 154.825 102.805 155.055 ;
        RECT 102.975 154.825 103.265 155.055 ;
        RECT 103.435 155.010 103.725 155.055 ;
        RECT 104.340 155.010 104.660 155.070 ;
        RECT 106.640 155.010 106.960 155.070 ;
        RECT 103.435 154.870 106.960 155.010 ;
        RECT 103.435 154.825 103.725 154.870 ;
        RECT 74.530 154.530 78.810 154.670 ;
        RECT 102.590 154.670 102.730 154.825 ;
        RECT 104.340 154.810 104.660 154.870 ;
        RECT 106.640 154.810 106.960 154.870 ;
        RECT 107.100 154.810 107.420 155.070 ;
        RECT 107.650 155.055 107.790 155.210 ;
        RECT 112.160 155.150 112.480 155.210 ;
        RECT 115.380 155.150 115.700 155.410 ;
        RECT 107.575 154.825 107.865 155.055 ;
        RECT 108.020 155.010 108.340 155.070 ;
        RECT 108.495 155.010 108.785 155.055 ;
        RECT 109.400 155.010 109.720 155.070 ;
        RECT 108.020 154.870 109.720 155.010 ;
        RECT 108.020 154.810 108.340 154.870 ;
        RECT 108.495 154.825 108.785 154.870 ;
        RECT 109.400 154.810 109.720 154.870 ;
        RECT 116.760 154.810 117.080 155.070 ;
        RECT 108.940 154.670 109.260 154.730 ;
        RECT 102.590 154.530 109.260 154.670 ;
        RECT 77.200 154.470 77.520 154.530 ;
        RECT 108.940 154.470 109.260 154.530 ;
        RECT 67.540 154.330 67.860 154.390 ;
        RECT 97.440 154.330 97.760 154.390 ;
        RECT 67.540 154.190 97.760 154.330 ;
        RECT 67.540 154.130 67.860 154.190 ;
        RECT 97.440 154.130 97.760 154.190 ;
        RECT 102.960 154.330 103.280 154.390 ;
        RECT 105.275 154.330 105.565 154.375 ;
        RECT 102.960 154.190 105.565 154.330 ;
        RECT 102.960 154.130 103.280 154.190 ;
        RECT 105.275 154.145 105.565 154.190 ;
        RECT 72.140 153.990 72.460 154.050 ;
        RECT 67.170 153.850 72.460 153.990 ;
        RECT 50.995 153.805 51.285 153.850 ;
        RECT 72.140 153.790 72.460 153.850 ;
        RECT 74.900 153.990 75.220 154.050 ;
        RECT 76.295 153.990 76.585 154.035 ;
        RECT 74.900 153.850 76.585 153.990 ;
        RECT 74.900 153.790 75.220 153.850 ;
        RECT 76.295 153.805 76.585 153.850 ;
        RECT 76.755 153.990 77.045 154.035 ;
        RECT 77.200 153.990 77.520 154.050 ;
        RECT 76.755 153.850 77.520 153.990 ;
        RECT 76.755 153.805 77.045 153.850 ;
        RECT 77.200 153.790 77.520 153.850 ;
        RECT 99.740 153.990 100.060 154.050 ;
        RECT 103.880 153.990 104.200 154.050 ;
        RECT 99.740 153.850 104.200 153.990 ;
        RECT 99.740 153.790 100.060 153.850 ;
        RECT 103.880 153.790 104.200 153.850 ;
        RECT 104.815 153.990 105.105 154.035 ;
        RECT 105.720 153.990 106.040 154.050 ;
        RECT 104.815 153.850 106.040 153.990 ;
        RECT 104.815 153.805 105.105 153.850 ;
        RECT 105.720 153.790 106.040 153.850 ;
        RECT 11.810 153.170 125.890 153.650 ;
        RECT 22.935 152.970 23.225 153.015 ;
        RECT 24.760 152.970 25.080 153.030 ;
        RECT 22.935 152.830 25.080 152.970 ;
        RECT 22.935 152.785 23.225 152.830 ;
        RECT 24.760 152.770 25.080 152.830 ;
        RECT 30.280 152.970 30.600 153.030 ;
        RECT 52.360 152.970 52.680 153.030 ;
        RECT 67.540 152.970 67.860 153.030 ;
        RECT 73.060 152.970 73.380 153.030 ;
        RECT 78.120 152.970 78.440 153.030 ;
        RECT 81.800 152.970 82.120 153.030 ;
        RECT 30.280 152.830 50.290 152.970 ;
        RECT 30.280 152.770 30.600 152.830 ;
        RECT 16.135 152.630 16.425 152.675 ;
        RECT 19.255 152.630 19.545 152.675 ;
        RECT 21.145 152.630 21.435 152.675 ;
        RECT 16.135 152.490 21.435 152.630 ;
        RECT 16.135 152.445 16.425 152.490 ;
        RECT 19.255 152.445 19.545 152.490 ;
        RECT 21.145 152.445 21.435 152.490 ;
        RECT 23.840 152.630 24.160 152.690 ;
        RECT 30.855 152.630 31.145 152.675 ;
        RECT 33.975 152.630 34.265 152.675 ;
        RECT 35.865 152.630 36.155 152.675 ;
        RECT 23.840 152.490 25.910 152.630 ;
        RECT 23.840 152.430 24.160 152.490 ;
        RECT 20.635 152.290 20.925 152.335 ;
        RECT 24.300 152.290 24.620 152.350 ;
        RECT 25.770 152.335 25.910 152.490 ;
        RECT 30.855 152.490 36.155 152.630 ;
        RECT 30.855 152.445 31.145 152.490 ;
        RECT 33.975 152.445 34.265 152.490 ;
        RECT 35.865 152.445 36.155 152.490 ;
        RECT 36.350 152.490 42.930 152.630 ;
        RECT 20.635 152.150 24.620 152.290 ;
        RECT 20.635 152.105 20.925 152.150 ;
        RECT 24.300 152.090 24.620 152.150 ;
        RECT 25.695 152.105 25.985 152.335 ;
        RECT 36.350 152.290 36.490 152.490 ;
        RECT 27.150 152.150 36.490 152.290 ;
        RECT 15.055 151.655 15.345 151.970 ;
        RECT 16.135 151.950 16.425 151.995 ;
        RECT 19.715 151.950 20.005 151.995 ;
        RECT 21.550 151.950 21.840 151.995 ;
        RECT 16.135 151.810 21.840 151.950 ;
        RECT 16.135 151.765 16.425 151.810 ;
        RECT 19.715 151.765 20.005 151.810 ;
        RECT 21.550 151.765 21.840 151.810 ;
        RECT 22.015 151.950 22.305 151.995 ;
        RECT 22.920 151.950 23.240 152.010 ;
        RECT 22.015 151.810 23.240 151.950 ;
        RECT 22.015 151.765 22.305 151.810 ;
        RECT 22.920 151.750 23.240 151.810 ;
        RECT 25.235 151.950 25.525 151.995 ;
        RECT 27.150 151.950 27.290 152.150 ;
        RECT 36.720 152.090 37.040 152.350 ;
        RECT 25.235 151.810 27.290 151.950 ;
        RECT 25.235 151.765 25.525 151.810 ;
        RECT 14.755 151.610 15.345 151.655 ;
        RECT 17.400 151.610 17.720 151.670 ;
        RECT 17.995 151.610 18.645 151.655 ;
        RECT 14.755 151.470 18.645 151.610 ;
        RECT 14.755 151.425 15.045 151.470 ;
        RECT 17.400 151.410 17.720 151.470 ;
        RECT 17.995 151.425 18.645 151.470 ;
        RECT 24.760 151.410 25.080 151.670 ;
        RECT 13.275 151.270 13.565 151.315 ;
        RECT 21.540 151.270 21.860 151.330 ;
        RECT 25.310 151.270 25.450 151.765 ;
        RECT 27.060 151.610 27.380 151.670 ;
        RECT 29.775 151.655 30.065 151.970 ;
        RECT 30.855 151.950 31.145 151.995 ;
        RECT 34.435 151.950 34.725 151.995 ;
        RECT 36.270 151.950 36.560 151.995 ;
        RECT 30.855 151.810 36.560 151.950 ;
        RECT 30.855 151.765 31.145 151.810 ;
        RECT 34.435 151.765 34.725 151.810 ;
        RECT 36.270 151.765 36.560 151.810 ;
        RECT 38.100 151.750 38.420 152.010 ;
        RECT 41.780 151.750 42.100 152.010 ;
        RECT 42.790 151.995 42.930 152.490 ;
        RECT 50.150 152.290 50.290 152.830 ;
        RECT 52.360 152.830 67.860 152.970 ;
        RECT 52.360 152.770 52.680 152.830 ;
        RECT 67.540 152.770 67.860 152.830 ;
        RECT 71.770 152.830 82.120 152.970 ;
        RECT 50.520 152.630 50.840 152.690 ;
        RECT 56.960 152.630 57.280 152.690 ;
        RECT 50.520 152.490 57.280 152.630 ;
        RECT 50.520 152.430 50.840 152.490 ;
        RECT 56.960 152.430 57.280 152.490 ;
        RECT 57.420 152.630 57.740 152.690 ;
        RECT 71.770 152.630 71.910 152.830 ;
        RECT 73.060 152.770 73.380 152.830 ;
        RECT 78.120 152.770 78.440 152.830 ;
        RECT 81.800 152.770 82.120 152.830 ;
        RECT 88.240 152.970 88.560 153.030 ;
        RECT 88.240 152.830 111.470 152.970 ;
        RECT 88.240 152.770 88.560 152.830 ;
        RECT 57.420 152.490 71.910 152.630 ;
        RECT 57.420 152.430 57.740 152.490 ;
        RECT 51.900 152.290 52.220 152.350 ;
        RECT 67.080 152.290 67.400 152.350 ;
        RECT 50.150 152.150 51.670 152.290 ;
        RECT 42.715 151.765 43.005 151.995 ;
        RECT 43.175 151.765 43.465 151.995 ;
        RECT 43.635 151.950 43.925 151.995 ;
        RECT 43.635 151.810 45.690 151.950 ;
        RECT 43.635 151.765 43.925 151.810 ;
        RECT 29.475 151.610 30.065 151.655 ;
        RECT 32.715 151.610 33.365 151.655 ;
        RECT 27.060 151.470 33.365 151.610 ;
        RECT 27.060 151.410 27.380 151.470 ;
        RECT 29.475 151.425 29.765 151.470 ;
        RECT 32.715 151.425 33.365 151.470 ;
        RECT 35.355 151.425 35.645 151.655 ;
        RECT 41.320 151.610 41.640 151.670 ;
        RECT 43.250 151.610 43.390 151.765 ;
        RECT 44.080 151.610 44.400 151.670 ;
        RECT 41.320 151.470 44.400 151.610 ;
        RECT 13.275 151.130 25.450 151.270 ;
        RECT 27.995 151.270 28.285 151.315 ;
        RECT 28.900 151.270 29.220 151.330 ;
        RECT 27.995 151.130 29.220 151.270 ;
        RECT 35.430 151.270 35.570 151.425 ;
        RECT 41.320 151.410 41.640 151.470 ;
        RECT 44.080 151.410 44.400 151.470 ;
        RECT 45.550 151.330 45.690 151.810 ;
        RECT 46.380 151.610 46.700 151.670 ;
        RECT 50.995 151.610 51.285 151.655 ;
        RECT 46.380 151.470 51.285 151.610 ;
        RECT 51.530 151.610 51.670 152.150 ;
        RECT 51.900 152.150 66.620 152.290 ;
        RECT 51.900 152.090 52.220 152.150 ;
        RECT 52.360 151.750 52.680 152.010 ;
        RECT 52.910 151.995 53.050 152.150 ;
        RECT 52.835 151.765 53.125 151.995 ;
        RECT 53.280 151.750 53.600 152.010 ;
        RECT 54.200 151.950 54.520 152.010 ;
        RECT 55.580 151.950 55.900 152.010 ;
        RECT 54.200 151.810 55.900 151.950 ;
        RECT 66.480 151.950 66.620 152.150 ;
        RECT 67.080 152.150 70.990 152.290 ;
        RECT 67.080 152.090 67.400 152.150 ;
        RECT 69.380 151.950 69.700 152.010 ;
        RECT 66.480 151.810 69.700 151.950 ;
        RECT 54.200 151.750 54.520 151.810 ;
        RECT 55.580 151.750 55.900 151.810 ;
        RECT 69.380 151.750 69.700 151.810 ;
        RECT 70.300 151.750 70.620 152.010 ;
        RECT 70.850 151.935 70.990 152.150 ;
        RECT 71.770 151.995 71.910 152.490 ;
        RECT 72.140 152.630 72.460 152.690 ;
        RECT 72.140 152.490 110.550 152.630 ;
        RECT 72.140 152.430 72.460 152.490 ;
        RECT 84.100 152.290 84.420 152.350 ;
        RECT 107.100 152.290 107.420 152.350 ;
        RECT 77.750 152.150 81.570 152.290 ;
        RECT 77.750 152.010 77.890 152.150 ;
        RECT 71.235 151.935 71.525 151.995 ;
        RECT 70.850 151.795 71.525 151.935 ;
        RECT 71.235 151.765 71.525 151.795 ;
        RECT 71.695 151.765 71.985 151.995 ;
        RECT 72.140 151.950 72.460 152.010 ;
        RECT 77.660 151.950 77.980 152.010 ;
        RECT 72.140 151.810 77.980 151.950 ;
        RECT 72.140 151.750 72.460 151.810 ;
        RECT 77.660 151.750 77.980 151.810 ;
        RECT 78.120 151.750 78.440 152.010 ;
        RECT 78.595 151.950 78.885 151.995 ;
        RECT 79.040 151.950 79.360 152.010 ;
        RECT 81.430 151.995 81.570 152.150 ;
        RECT 82.350 152.150 84.420 152.290 ;
        RECT 78.595 151.810 79.360 151.950 ;
        RECT 78.595 151.765 78.885 151.810 ;
        RECT 79.040 151.750 79.360 151.810 ;
        RECT 79.515 151.950 79.805 151.995 ;
        RECT 79.515 151.810 80.190 151.950 ;
        RECT 79.515 151.765 79.805 151.810 ;
        RECT 67.080 151.610 67.400 151.670 ;
        RECT 51.530 151.470 67.400 151.610 ;
        RECT 70.390 151.610 70.530 151.750 ;
        RECT 80.050 151.610 80.190 151.810 ;
        RECT 81.355 151.765 81.645 151.995 ;
        RECT 81.800 151.750 82.120 152.010 ;
        RECT 82.350 151.995 82.490 152.150 ;
        RECT 84.100 152.090 84.420 152.150 ;
        RECT 97.990 152.150 103.650 152.290 ;
        RECT 97.990 152.010 98.130 152.150 ;
        RECT 82.275 151.765 82.565 151.995 ;
        RECT 83.195 151.765 83.485 151.995 ;
        RECT 83.270 151.610 83.410 151.765 ;
        RECT 97.440 151.750 97.760 152.010 ;
        RECT 97.900 151.750 98.220 152.010 ;
        RECT 98.360 151.750 98.680 152.010 ;
        RECT 98.820 151.950 99.140 152.010 ;
        RECT 103.510 151.995 103.650 152.150 ;
        RECT 107.100 152.150 108.250 152.290 ;
        RECT 107.100 152.090 107.420 152.150 ;
        RECT 99.295 151.950 99.585 151.995 ;
        RECT 98.820 151.810 99.585 151.950 ;
        RECT 98.820 151.750 99.140 151.810 ;
        RECT 99.295 151.765 99.585 151.810 ;
        RECT 102.975 151.765 103.265 151.995 ;
        RECT 103.435 151.765 103.725 151.995 ;
        RECT 70.390 151.470 83.410 151.610 ;
        RECT 97.530 151.610 97.670 151.750 ;
        RECT 103.050 151.610 103.190 151.765 ;
        RECT 103.880 151.750 104.200 152.010 ;
        RECT 104.800 151.750 105.120 152.010 ;
        RECT 108.110 151.995 108.250 152.150 ;
        RECT 107.575 151.765 107.865 151.995 ;
        RECT 108.035 151.765 108.325 151.995 ;
        RECT 104.340 151.610 104.660 151.670 ;
        RECT 107.650 151.610 107.790 151.765 ;
        RECT 108.480 151.750 108.800 152.010 ;
        RECT 110.410 151.995 110.550 152.490 ;
        RECT 111.330 152.335 111.470 152.830 ;
        RECT 115.955 152.630 116.245 152.675 ;
        RECT 119.075 152.630 119.365 152.675 ;
        RECT 120.965 152.630 121.255 152.675 ;
        RECT 115.955 152.490 121.255 152.630 ;
        RECT 115.955 152.445 116.245 152.490 ;
        RECT 119.075 152.445 119.365 152.490 ;
        RECT 120.965 152.445 121.255 152.490 ;
        RECT 111.255 152.105 111.545 152.335 ;
        RECT 116.760 152.290 117.080 152.350 ;
        RECT 111.790 152.150 117.080 152.290 ;
        RECT 109.415 151.765 109.705 151.995 ;
        RECT 110.335 151.950 110.625 151.995 ;
        RECT 111.790 151.950 111.930 152.150 ;
        RECT 116.760 152.090 117.080 152.150 ;
        RECT 121.835 152.290 122.125 152.335 ;
        RECT 123.660 152.290 123.980 152.350 ;
        RECT 121.835 152.150 123.980 152.290 ;
        RECT 121.835 152.105 122.125 152.150 ;
        RECT 123.660 152.090 123.980 152.150 ;
        RECT 110.335 151.810 111.930 151.950 ;
        RECT 110.335 151.765 110.625 151.810 ;
        RECT 109.490 151.610 109.630 151.765 ;
        RECT 114.875 151.655 115.165 151.970 ;
        RECT 115.955 151.950 116.245 151.995 ;
        RECT 119.535 151.950 119.825 151.995 ;
        RECT 121.370 151.950 121.660 151.995 ;
        RECT 115.955 151.810 121.660 151.950 ;
        RECT 115.955 151.765 116.245 151.810 ;
        RECT 119.535 151.765 119.825 151.810 ;
        RECT 121.370 151.765 121.660 151.810 ;
        RECT 97.530 151.470 107.790 151.610 ;
        RECT 108.110 151.470 109.630 151.610 ;
        RECT 114.575 151.610 115.165 151.655 ;
        RECT 116.760 151.610 117.080 151.670 ;
        RECT 117.815 151.610 118.465 151.655 ;
        RECT 114.575 151.470 118.465 151.610 ;
        RECT 46.380 151.410 46.700 151.470 ;
        RECT 50.995 151.425 51.285 151.470 ;
        RECT 67.080 151.410 67.400 151.470 ;
        RECT 79.590 151.330 79.730 151.470 ;
        RECT 104.340 151.410 104.660 151.470 ;
        RECT 108.110 151.330 108.250 151.470 ;
        RECT 114.575 151.425 114.865 151.470 ;
        RECT 116.760 151.410 117.080 151.470 ;
        RECT 117.815 151.425 118.465 151.470 ;
        RECT 120.440 151.410 120.760 151.670 ;
        RECT 37.195 151.270 37.485 151.315 ;
        RECT 35.430 151.130 37.485 151.270 ;
        RECT 13.275 151.085 13.565 151.130 ;
        RECT 21.540 151.070 21.860 151.130 ;
        RECT 27.995 151.085 28.285 151.130 ;
        RECT 28.900 151.070 29.220 151.130 ;
        RECT 37.195 151.085 37.485 151.130 ;
        RECT 43.620 151.270 43.940 151.330 ;
        RECT 45.015 151.270 45.305 151.315 ;
        RECT 43.620 151.130 45.305 151.270 ;
        RECT 43.620 151.070 43.940 151.130 ;
        RECT 45.015 151.085 45.305 151.130 ;
        RECT 45.460 151.270 45.780 151.330 ;
        RECT 66.620 151.270 66.940 151.330 ;
        RECT 72.140 151.270 72.460 151.330 ;
        RECT 45.460 151.130 72.460 151.270 ;
        RECT 45.460 151.070 45.780 151.130 ;
        RECT 66.620 151.070 66.940 151.130 ;
        RECT 72.140 151.070 72.460 151.130 ;
        RECT 73.535 151.270 73.825 151.315 ;
        RECT 73.980 151.270 74.300 151.330 ;
        RECT 73.535 151.130 74.300 151.270 ;
        RECT 73.535 151.085 73.825 151.130 ;
        RECT 73.980 151.070 74.300 151.130 ;
        RECT 76.280 151.070 76.600 151.330 ;
        RECT 79.500 151.070 79.820 151.330 ;
        RECT 79.975 151.270 80.265 151.315 ;
        RECT 80.880 151.270 81.200 151.330 ;
        RECT 79.975 151.130 81.200 151.270 ;
        RECT 79.975 151.085 80.265 151.130 ;
        RECT 80.880 151.070 81.200 151.130 ;
        RECT 94.680 151.270 95.000 151.330 ;
        RECT 96.075 151.270 96.365 151.315 ;
        RECT 94.680 151.130 96.365 151.270 ;
        RECT 94.680 151.070 95.000 151.130 ;
        RECT 96.075 151.085 96.365 151.130 ;
        RECT 100.660 151.270 100.980 151.330 ;
        RECT 101.595 151.270 101.885 151.315 ;
        RECT 100.660 151.130 101.885 151.270 ;
        RECT 100.660 151.070 100.980 151.130 ;
        RECT 101.595 151.085 101.885 151.130 ;
        RECT 102.040 151.270 102.360 151.330 ;
        RECT 106.195 151.270 106.485 151.315 ;
        RECT 102.040 151.130 106.485 151.270 ;
        RECT 102.040 151.070 102.360 151.130 ;
        RECT 106.195 151.085 106.485 151.130 ;
        RECT 108.020 151.070 108.340 151.330 ;
        RECT 112.620 151.270 112.940 151.330 ;
        RECT 113.095 151.270 113.385 151.315 ;
        RECT 112.620 151.130 113.385 151.270 ;
        RECT 112.620 151.070 112.940 151.130 ;
        RECT 113.095 151.085 113.385 151.130 ;
        RECT 11.010 150.450 125.890 150.930 ;
        RECT 16.035 150.250 16.325 150.295 ;
        RECT 16.480 150.250 16.800 150.310 ;
        RECT 16.035 150.110 16.800 150.250 ;
        RECT 16.035 150.065 16.325 150.110 ;
        RECT 16.480 150.050 16.800 150.110 ;
        RECT 17.400 150.050 17.720 150.310 ;
        RECT 19.240 150.050 19.560 150.310 ;
        RECT 21.540 150.050 21.860 150.310 ;
        RECT 26.155 150.250 26.445 150.295 ;
        RECT 27.980 150.250 28.300 150.310 ;
        RECT 26.155 150.110 28.300 150.250 ;
        RECT 26.155 150.065 26.445 150.110 ;
        RECT 27.980 150.050 28.300 150.110 ;
        RECT 28.900 150.250 29.220 150.310 ;
        RECT 31.660 150.250 31.980 150.310 ;
        RECT 28.900 150.110 31.980 150.250 ;
        RECT 28.900 150.050 29.220 150.110 ;
        RECT 31.660 150.050 31.980 150.110 ;
        RECT 33.040 150.050 33.360 150.310 ;
        RECT 33.500 150.250 33.820 150.310 ;
        RECT 35.815 150.250 36.105 150.295 ;
        RECT 52.820 150.250 53.140 150.310 ;
        RECT 33.500 150.110 36.105 150.250 ;
        RECT 33.500 150.050 33.820 150.110 ;
        RECT 35.815 150.065 36.105 150.110 ;
        RECT 52.450 150.110 53.140 150.250 ;
        RECT 25.220 149.910 25.540 149.970 ;
        RECT 27.520 149.910 27.840 149.970 ;
        RECT 28.455 149.910 28.745 149.955 ;
        RECT 17.950 149.770 20.390 149.910 ;
        RECT 14.180 149.570 14.500 149.630 ;
        RECT 17.950 149.615 18.090 149.770 ;
        RECT 15.575 149.570 15.865 149.615 ;
        RECT 17.875 149.570 18.165 149.615 ;
        RECT 14.180 149.430 18.165 149.570 ;
        RECT 14.180 149.370 14.500 149.430 ;
        RECT 15.575 149.385 15.865 149.430 ;
        RECT 17.875 149.385 18.165 149.430 ;
        RECT 18.335 149.570 18.625 149.615 ;
        RECT 20.250 149.570 20.390 149.770 ;
        RECT 25.220 149.770 37.410 149.910 ;
        RECT 25.220 149.710 25.540 149.770 ;
        RECT 27.520 149.710 27.840 149.770 ;
        RECT 28.455 149.725 28.745 149.770 ;
        RECT 25.695 149.570 25.985 149.615 ;
        RECT 30.280 149.570 30.600 149.630 ;
        RECT 36.735 149.570 37.025 149.615 ;
        RECT 18.335 149.430 19.930 149.570 ;
        RECT 20.250 149.430 30.600 149.570 ;
        RECT 18.335 149.385 18.625 149.430 ;
        RECT 19.790 148.935 19.930 149.430 ;
        RECT 25.695 149.385 25.985 149.430 ;
        RECT 30.280 149.370 30.600 149.430 ;
        RECT 30.830 149.430 37.025 149.570 ;
        RECT 37.270 149.570 37.410 149.770 ;
        RECT 40.490 149.770 44.770 149.910 ;
        RECT 40.490 149.630 40.630 149.770 ;
        RECT 37.270 149.430 39.250 149.570 ;
        RECT 22.000 149.030 22.320 149.290 ;
        RECT 22.935 149.230 23.225 149.275 ;
        RECT 23.840 149.230 24.160 149.290 ;
        RECT 27.535 149.230 27.825 149.275 ;
        RECT 22.935 149.090 27.825 149.230 ;
        RECT 22.935 149.045 23.225 149.090 ;
        RECT 23.840 149.030 24.160 149.090 ;
        RECT 27.535 149.045 27.825 149.090 ;
        RECT 19.715 148.705 20.005 148.935 ;
        RECT 27.610 148.550 27.750 149.045 ;
        RECT 30.830 148.935 30.970 149.430 ;
        RECT 36.735 149.385 37.025 149.430 ;
        RECT 31.675 149.230 31.965 149.275 ;
        RECT 31.290 149.090 31.965 149.230 ;
        RECT 30.755 148.705 31.045 148.935 ;
        RECT 31.290 148.550 31.430 149.090 ;
        RECT 31.675 149.045 31.965 149.090 ;
        RECT 32.595 149.045 32.885 149.275 ;
        RECT 39.110 149.230 39.250 149.430 ;
        RECT 40.400 149.370 40.720 149.630 ;
        RECT 40.860 149.370 41.180 149.630 ;
        RECT 41.335 149.385 41.625 149.615 ;
        RECT 41.780 149.570 42.100 149.630 ;
        RECT 42.255 149.570 42.545 149.615 ;
        RECT 42.715 149.570 43.005 149.615 ;
        RECT 41.780 149.430 43.005 149.570 ;
        RECT 41.410 149.230 41.550 149.385 ;
        RECT 41.780 149.370 42.100 149.430 ;
        RECT 42.255 149.385 42.545 149.430 ;
        RECT 42.715 149.385 43.005 149.430 ;
        RECT 43.160 149.570 43.480 149.630 ;
        RECT 43.635 149.570 43.925 149.615 ;
        RECT 43.160 149.430 43.925 149.570 ;
        RECT 43.160 149.370 43.480 149.430 ;
        RECT 43.635 149.385 43.925 149.430 ;
        RECT 44.080 149.370 44.400 149.630 ;
        RECT 44.630 149.615 44.770 149.770 ;
        RECT 44.555 149.570 44.845 149.615 ;
        RECT 45.460 149.570 45.780 149.630 ;
        RECT 44.555 149.430 45.780 149.570 ;
        RECT 44.555 149.385 44.845 149.430 ;
        RECT 45.460 149.370 45.780 149.430 ;
        RECT 50.995 149.385 51.285 149.615 ;
        RECT 39.110 149.090 41.550 149.230 ;
        RECT 44.170 149.230 44.310 149.370 ;
        RECT 51.070 149.230 51.210 149.385 ;
        RECT 51.440 149.370 51.760 149.630 ;
        RECT 51.915 149.570 52.205 149.615 ;
        RECT 52.450 149.570 52.590 150.110 ;
        RECT 52.820 150.050 53.140 150.110 ;
        RECT 69.840 150.250 70.160 150.310 ;
        RECT 70.315 150.250 70.605 150.295 ;
        RECT 69.840 150.110 70.605 150.250 ;
        RECT 69.840 150.050 70.160 150.110 ;
        RECT 70.315 150.065 70.605 150.110 ;
        RECT 71.695 150.250 71.985 150.295 ;
        RECT 98.820 150.250 99.140 150.310 ;
        RECT 104.800 150.250 105.120 150.310 ;
        RECT 108.020 150.250 108.340 150.310 ;
        RECT 71.695 150.110 108.340 150.250 ;
        RECT 71.695 150.065 71.985 150.110 ;
        RECT 58.800 149.910 59.120 149.970 ;
        RECT 71.770 149.910 71.910 150.065 ;
        RECT 98.820 150.050 99.140 150.110 ;
        RECT 104.800 150.050 105.120 150.110 ;
        RECT 108.020 150.050 108.340 150.110 ;
        RECT 116.760 150.050 117.080 150.310 ;
        RECT 118.615 150.250 118.905 150.295 ;
        RECT 120.440 150.250 120.760 150.310 ;
        RECT 118.615 150.110 120.760 150.250 ;
        RECT 118.615 150.065 118.905 150.110 ;
        RECT 120.440 150.050 120.760 150.110 ;
        RECT 58.800 149.770 71.910 149.910 ;
        RECT 90.655 149.910 90.945 149.955 ;
        RECT 92.840 149.910 93.160 149.970 ;
        RECT 93.895 149.910 94.545 149.955 ;
        RECT 90.655 149.770 94.545 149.910 ;
        RECT 58.800 149.710 59.120 149.770 ;
        RECT 90.655 149.725 91.245 149.770 ;
        RECT 51.915 149.430 52.590 149.570 ;
        RECT 52.835 149.570 53.125 149.615 ;
        RECT 54.200 149.570 54.520 149.630 ;
        RECT 58.890 149.570 59.030 149.710 ;
        RECT 52.835 149.430 59.030 149.570 ;
        RECT 63.415 149.570 63.705 149.615 ;
        RECT 64.320 149.570 64.640 149.630 ;
        RECT 63.415 149.430 64.640 149.570 ;
        RECT 51.915 149.385 52.205 149.430 ;
        RECT 52.835 149.385 53.125 149.430 ;
        RECT 54.200 149.370 54.520 149.430 ;
        RECT 63.415 149.385 63.705 149.430 ;
        RECT 64.320 149.370 64.640 149.430 ;
        RECT 65.255 149.385 65.545 149.615 ;
        RECT 69.395 149.570 69.685 149.615 ;
        RECT 71.680 149.570 72.000 149.630 ;
        RECT 72.615 149.570 72.905 149.615 ;
        RECT 73.060 149.570 73.380 149.630 ;
        RECT 69.395 149.430 73.380 149.570 ;
        RECT 69.395 149.385 69.685 149.430 ;
        RECT 52.360 149.230 52.680 149.290 ;
        RECT 44.170 149.090 50.290 149.230 ;
        RECT 51.070 149.090 52.680 149.230 ;
        RECT 27.610 148.410 31.430 148.550 ;
        RECT 31.660 148.550 31.980 148.610 ;
        RECT 32.670 148.550 32.810 149.045 ;
        RECT 34.880 148.690 35.200 148.950 ;
        RECT 40.860 148.890 41.180 148.950 ;
        RECT 38.190 148.750 41.180 148.890 ;
        RECT 38.190 148.550 38.330 148.750 ;
        RECT 40.860 148.690 41.180 148.750 ;
        RECT 41.320 148.890 41.640 148.950 ;
        RECT 49.615 148.890 49.905 148.935 ;
        RECT 41.320 148.750 49.905 148.890 ;
        RECT 50.150 148.890 50.290 149.090 ;
        RECT 52.360 149.030 52.680 149.090 ;
        RECT 60.640 149.230 60.960 149.290 ;
        RECT 65.330 149.230 65.470 149.385 ;
        RECT 71.680 149.370 72.000 149.430 ;
        RECT 72.615 149.385 72.905 149.430 ;
        RECT 73.060 149.370 73.380 149.430 ;
        RECT 77.660 149.370 77.980 149.630 ;
        RECT 78.120 149.370 78.440 149.630 ;
        RECT 78.580 149.370 78.900 149.630 ;
        RECT 79.500 149.370 79.820 149.630 ;
        RECT 88.240 149.370 88.560 149.630 ;
        RECT 90.955 149.410 91.245 149.725 ;
        RECT 92.840 149.710 93.160 149.770 ;
        RECT 93.895 149.725 94.545 149.770 ;
        RECT 92.035 149.570 92.325 149.615 ;
        RECT 95.615 149.570 95.905 149.615 ;
        RECT 97.450 149.570 97.740 149.615 ;
        RECT 92.035 149.430 97.740 149.570 ;
        RECT 92.035 149.385 92.325 149.430 ;
        RECT 95.615 149.385 95.905 149.430 ;
        RECT 97.450 149.385 97.740 149.430 ;
        RECT 105.720 149.370 106.040 149.630 ;
        RECT 106.180 149.370 106.500 149.630 ;
        RECT 107.100 149.370 107.420 149.630 ;
        RECT 115.380 149.570 115.700 149.630 ;
        RECT 117.235 149.570 117.525 149.615 ;
        RECT 115.380 149.430 117.525 149.570 ;
        RECT 115.380 149.370 115.700 149.430 ;
        RECT 117.235 149.385 117.525 149.430 ;
        RECT 117.680 149.370 118.000 149.630 ;
        RECT 60.640 149.090 65.470 149.230 ;
        RECT 60.640 149.030 60.960 149.090 ;
        RECT 96.520 149.030 96.840 149.290 ;
        RECT 97.915 149.230 98.205 149.275 ;
        RECT 98.360 149.230 98.680 149.290 ;
        RECT 97.915 149.090 98.680 149.230 ;
        RECT 97.915 149.045 98.205 149.090 ;
        RECT 98.360 149.030 98.680 149.090 ;
        RECT 57.420 148.890 57.740 148.950 ;
        RECT 50.150 148.750 57.740 148.890 ;
        RECT 41.320 148.690 41.640 148.750 ;
        RECT 49.615 148.705 49.905 148.750 ;
        RECT 57.420 148.690 57.740 148.750 ;
        RECT 92.035 148.890 92.325 148.935 ;
        RECT 95.155 148.890 95.445 148.935 ;
        RECT 97.045 148.890 97.335 148.935 ;
        RECT 92.035 148.750 97.335 148.890 ;
        RECT 92.035 148.705 92.325 148.750 ;
        RECT 95.155 148.705 95.445 148.750 ;
        RECT 97.045 148.705 97.335 148.750 ;
        RECT 104.815 148.890 105.105 148.935 ;
        RECT 118.600 148.890 118.920 148.950 ;
        RECT 104.815 148.750 118.920 148.890 ;
        RECT 104.815 148.705 105.105 148.750 ;
        RECT 118.600 148.690 118.920 148.750 ;
        RECT 31.660 148.410 38.330 148.550 ;
        RECT 38.560 148.550 38.880 148.610 ;
        RECT 39.035 148.550 39.325 148.595 ;
        RECT 38.560 148.410 39.325 148.550 ;
        RECT 31.660 148.350 31.980 148.410 ;
        RECT 38.560 148.350 38.880 148.410 ;
        RECT 39.035 148.365 39.325 148.410 ;
        RECT 45.000 148.550 45.320 148.610 ;
        RECT 45.935 148.550 46.225 148.595 ;
        RECT 45.000 148.410 46.225 148.550 ;
        RECT 45.000 148.350 45.320 148.410 ;
        RECT 45.935 148.365 46.225 148.410 ;
        RECT 63.860 148.350 64.180 148.610 ;
        RECT 66.175 148.550 66.465 148.595 ;
        RECT 70.300 148.550 70.620 148.610 ;
        RECT 66.175 148.410 70.620 148.550 ;
        RECT 66.175 148.365 66.465 148.410 ;
        RECT 70.300 148.350 70.620 148.410 ;
        RECT 71.680 148.550 72.000 148.610 ;
        RECT 73.520 148.550 73.840 148.610 ;
        RECT 71.680 148.410 73.840 148.550 ;
        RECT 71.680 148.350 72.000 148.410 ;
        RECT 73.520 148.350 73.840 148.410 ;
        RECT 76.295 148.550 76.585 148.595 ;
        RECT 77.660 148.550 77.980 148.610 ;
        RECT 76.295 148.410 77.980 148.550 ;
        RECT 76.295 148.365 76.585 148.410 ;
        RECT 77.660 148.350 77.980 148.410 ;
        RECT 87.795 148.550 88.085 148.595 ;
        RECT 88.240 148.550 88.560 148.610 ;
        RECT 87.795 148.410 88.560 148.550 ;
        RECT 87.795 148.365 88.085 148.410 ;
        RECT 88.240 148.350 88.560 148.410 ;
        RECT 89.175 148.550 89.465 148.595 ;
        RECT 90.540 148.550 90.860 148.610 ;
        RECT 89.175 148.410 90.860 148.550 ;
        RECT 89.175 148.365 89.465 148.410 ;
        RECT 90.540 148.350 90.860 148.410 ;
        RECT 107.115 148.550 107.405 148.595 ;
        RECT 107.560 148.550 107.880 148.610 ;
        RECT 107.115 148.410 107.880 148.550 ;
        RECT 107.115 148.365 107.405 148.410 ;
        RECT 107.560 148.350 107.880 148.410 ;
        RECT 11.810 147.730 125.890 148.210 ;
        RECT 33.040 147.530 33.360 147.590 ;
        RECT 43.160 147.530 43.480 147.590 ;
        RECT 33.040 147.390 43.480 147.530 ;
        RECT 33.040 147.330 33.360 147.390 ;
        RECT 43.160 147.330 43.480 147.390 ;
        RECT 61.100 147.330 61.420 147.590 ;
        RECT 71.680 147.330 72.000 147.590 ;
        RECT 73.535 147.530 73.825 147.575 ;
        RECT 75.360 147.530 75.680 147.590 ;
        RECT 73.535 147.390 75.680 147.530 ;
        RECT 73.535 147.345 73.825 147.390 ;
        RECT 75.360 147.330 75.680 147.390 ;
        RECT 92.840 147.330 93.160 147.590 ;
        RECT 95.155 147.530 95.445 147.575 ;
        RECT 96.520 147.530 96.840 147.590 ;
        RECT 95.155 147.390 96.840 147.530 ;
        RECT 95.155 147.345 95.445 147.390 ;
        RECT 96.520 147.330 96.840 147.390 ;
        RECT 98.375 147.530 98.665 147.575 ;
        RECT 98.820 147.530 99.140 147.590 ;
        RECT 98.375 147.390 99.140 147.530 ;
        RECT 98.375 147.345 98.665 147.390 ;
        RECT 98.820 147.330 99.140 147.390 ;
        RECT 106.655 147.530 106.945 147.575 ;
        RECT 107.100 147.530 107.420 147.590 ;
        RECT 106.655 147.390 107.420 147.530 ;
        RECT 106.655 147.345 106.945 147.390 ;
        RECT 107.100 147.330 107.420 147.390 ;
        RECT 114.935 147.530 115.225 147.575 ;
        RECT 117.680 147.530 118.000 147.590 ;
        RECT 114.935 147.390 118.000 147.530 ;
        RECT 114.935 147.345 115.225 147.390 ;
        RECT 117.680 147.330 118.000 147.390 ;
        RECT 22.000 147.190 22.320 147.250 ;
        RECT 44.080 147.190 44.400 147.250 ;
        RECT 22.000 147.050 39.710 147.190 ;
        RECT 22.000 146.990 22.320 147.050 ;
        RECT 39.570 146.555 39.710 147.050 ;
        RECT 40.490 147.050 44.400 147.190 ;
        RECT 40.490 146.850 40.630 147.050 ;
        RECT 44.080 146.990 44.400 147.050 ;
        RECT 59.260 146.990 59.580 147.250 ;
        RECT 69.395 147.005 69.685 147.235 ;
        RECT 74.440 147.190 74.760 147.250 ;
        RECT 71.310 147.050 74.760 147.190 ;
        RECT 40.030 146.710 40.630 146.850 ;
        RECT 40.860 146.850 41.180 146.910 ;
        RECT 44.170 146.850 44.310 146.990 ;
        RECT 59.350 146.850 59.490 146.990 ;
        RECT 69.470 146.850 69.610 147.005 ;
        RECT 70.760 146.850 71.080 146.910 ;
        RECT 40.860 146.710 43.390 146.850 ;
        RECT 40.030 146.555 40.170 146.710 ;
        RECT 40.860 146.650 41.180 146.710 ;
        RECT 38.575 146.325 38.865 146.555 ;
        RECT 39.495 146.325 39.785 146.555 ;
        RECT 39.955 146.325 40.245 146.555 ;
        RECT 38.650 146.170 38.790 146.325 ;
        RECT 40.400 146.310 40.720 146.570 ;
        RECT 41.780 146.510 42.100 146.570 ;
        RECT 43.250 146.555 43.390 146.710 ;
        RECT 43.710 146.710 44.310 146.850 ;
        RECT 53.830 146.710 71.080 146.850 ;
        RECT 43.710 146.555 43.850 146.710 ;
        RECT 53.830 146.570 53.970 146.710 ;
        RECT 42.255 146.510 42.545 146.555 ;
        RECT 41.780 146.370 42.545 146.510 ;
        RECT 41.780 146.310 42.100 146.370 ;
        RECT 42.255 146.325 42.545 146.370 ;
        RECT 43.175 146.325 43.465 146.555 ;
        RECT 43.635 146.325 43.925 146.555 ;
        RECT 44.080 146.510 44.400 146.570 ;
        RECT 45.460 146.510 45.780 146.570 ;
        RECT 44.080 146.370 45.780 146.510 ;
        RECT 41.870 146.170 42.010 146.310 ;
        RECT 38.650 146.030 42.010 146.170 ;
        RECT 39.020 145.830 39.340 145.890 ;
        RECT 41.795 145.830 42.085 145.875 ;
        RECT 39.020 145.690 42.085 145.830 ;
        RECT 39.020 145.630 39.340 145.690 ;
        RECT 41.795 145.645 42.085 145.690 ;
        RECT 43.160 145.830 43.480 145.890 ;
        RECT 43.710 145.830 43.850 146.325 ;
        RECT 44.080 146.310 44.400 146.370 ;
        RECT 45.460 146.310 45.780 146.370 ;
        RECT 53.740 146.310 54.060 146.570 ;
        RECT 54.215 146.325 54.505 146.555 ;
        RECT 54.290 146.170 54.430 146.325 ;
        RECT 54.660 146.310 54.980 146.570 ;
        RECT 55.595 146.510 55.885 146.555 ;
        RECT 56.500 146.510 56.820 146.570 ;
        RECT 57.510 146.555 57.650 146.710 ;
        RECT 70.760 146.650 71.080 146.710 ;
        RECT 55.595 146.370 56.820 146.510 ;
        RECT 55.595 146.325 55.885 146.370 ;
        RECT 56.500 146.310 56.820 146.370 ;
        RECT 57.435 146.325 57.725 146.555 ;
        RECT 57.895 146.325 58.185 146.555 ;
        RECT 55.120 146.170 55.440 146.230 ;
        RECT 57.970 146.170 58.110 146.325 ;
        RECT 58.340 146.310 58.660 146.570 ;
        RECT 58.800 146.510 59.120 146.570 ;
        RECT 71.310 146.555 71.450 147.050 ;
        RECT 74.440 146.990 74.760 147.050 ;
        RECT 86.830 147.190 87.120 147.235 ;
        RECT 89.610 147.190 89.900 147.235 ;
        RECT 91.470 147.190 91.760 147.235 ;
        RECT 86.830 147.050 91.760 147.190 ;
        RECT 86.830 147.005 87.120 147.050 ;
        RECT 89.610 147.005 89.900 147.050 ;
        RECT 91.470 147.005 91.760 147.050 ;
        RECT 99.295 147.190 99.585 147.235 ;
        RECT 117.220 147.190 117.540 147.250 ;
        RECT 99.295 147.050 117.540 147.190 ;
        RECT 99.295 147.005 99.585 147.050 ;
        RECT 117.220 146.990 117.540 147.050 ;
        RECT 73.060 146.850 73.380 146.910 ;
        RECT 95.140 146.850 95.460 146.910 ;
        RECT 97.455 146.850 97.745 146.895 ;
        RECT 110.320 146.850 110.640 146.910 ;
        RECT 111.715 146.850 112.005 146.895 ;
        RECT 73.060 146.710 76.510 146.850 ;
        RECT 73.060 146.650 73.380 146.710 ;
        RECT 59.275 146.510 59.565 146.555 ;
        RECT 58.800 146.370 59.565 146.510 ;
        RECT 58.800 146.310 59.120 146.370 ;
        RECT 59.275 146.325 59.565 146.370 ;
        RECT 70.315 146.510 70.605 146.555 ;
        RECT 71.235 146.510 71.525 146.555 ;
        RECT 70.315 146.370 71.525 146.510 ;
        RECT 70.315 146.325 70.605 146.370 ;
        RECT 71.235 146.325 71.525 146.370 ;
        RECT 72.600 146.310 72.920 146.570 ;
        RECT 73.520 146.510 73.840 146.570 ;
        RECT 76.370 146.555 76.510 146.710 ;
        RECT 95.140 146.710 97.745 146.850 ;
        RECT 95.140 146.650 95.460 146.710 ;
        RECT 97.455 146.665 97.745 146.710 ;
        RECT 103.970 146.710 108.250 146.850 ;
        RECT 103.970 146.570 104.110 146.710 ;
        RECT 74.455 146.510 74.745 146.555 ;
        RECT 73.520 146.370 74.745 146.510 ;
        RECT 73.520 146.310 73.840 146.370 ;
        RECT 74.455 146.325 74.745 146.370 ;
        RECT 76.295 146.325 76.585 146.555 ;
        RECT 86.830 146.510 87.120 146.555 ;
        RECT 86.830 146.370 89.365 146.510 ;
        RECT 86.830 146.325 87.120 146.370 ;
        RECT 59.720 146.170 60.040 146.230 ;
        RECT 68.475 146.170 68.765 146.215 ;
        RECT 73.060 146.170 73.380 146.230 ;
        RECT 84.100 146.170 84.420 146.230 ;
        RECT 88.240 146.215 88.560 146.230 ;
        RECT 54.290 146.030 66.620 146.170 ;
        RECT 55.120 145.970 55.440 146.030 ;
        RECT 59.720 145.970 60.040 146.030 ;
        RECT 43.160 145.690 43.850 145.830 ;
        RECT 43.160 145.630 43.480 145.690 ;
        RECT 45.460 145.630 45.780 145.890 ;
        RECT 52.360 145.630 52.680 145.890 ;
        RECT 56.055 145.830 56.345 145.875 ;
        RECT 57.880 145.830 58.200 145.890 ;
        RECT 56.055 145.690 58.200 145.830 ;
        RECT 66.480 145.830 66.620 146.030 ;
        RECT 68.475 146.030 73.380 146.170 ;
        RECT 68.475 145.985 68.765 146.030 ;
        RECT 73.060 145.970 73.380 146.030 ;
        RECT 75.450 146.030 84.420 146.170 ;
        RECT 75.450 145.875 75.590 146.030 ;
        RECT 84.100 145.970 84.420 146.030 ;
        RECT 84.970 146.170 85.260 146.215 ;
        RECT 88.230 146.170 88.560 146.215 ;
        RECT 84.970 146.030 88.560 146.170 ;
        RECT 84.970 145.985 85.260 146.030 ;
        RECT 88.230 145.985 88.560 146.030 ;
        RECT 89.150 146.215 89.365 146.370 ;
        RECT 90.080 146.310 90.400 146.570 ;
        RECT 91.920 146.310 92.240 146.570 ;
        RECT 93.300 146.310 93.620 146.570 ;
        RECT 94.220 146.310 94.540 146.570 ;
        RECT 98.375 146.510 98.665 146.555 ;
        RECT 100.660 146.510 100.980 146.570 ;
        RECT 98.375 146.370 100.980 146.510 ;
        RECT 98.375 146.325 98.665 146.370 ;
        RECT 100.660 146.310 100.980 146.370 ;
        RECT 103.880 146.310 104.200 146.570 ;
        RECT 104.340 146.310 104.660 146.570 ;
        RECT 104.815 146.325 105.105 146.555 ;
        RECT 89.150 146.170 89.440 146.215 ;
        RECT 91.010 146.170 91.300 146.215 ;
        RECT 89.150 146.030 91.300 146.170 ;
        RECT 89.150 145.985 89.440 146.030 ;
        RECT 91.010 145.985 91.300 146.030 ;
        RECT 96.995 146.170 97.285 146.215 ;
        RECT 102.515 146.170 102.805 146.215 ;
        RECT 96.995 146.030 102.805 146.170 ;
        RECT 96.995 145.985 97.285 146.030 ;
        RECT 102.515 145.985 102.805 146.030 ;
        RECT 88.240 145.970 88.560 145.985 ;
        RECT 75.375 145.830 75.665 145.875 ;
        RECT 66.480 145.690 75.665 145.830 ;
        RECT 56.055 145.645 56.345 145.690 ;
        RECT 57.880 145.630 58.200 145.690 ;
        RECT 75.375 145.645 75.665 145.690 ;
        RECT 77.215 145.830 77.505 145.875 ;
        RECT 78.580 145.830 78.900 145.890 ;
        RECT 83.180 145.875 83.500 145.890 ;
        RECT 77.215 145.690 78.900 145.830 ;
        RECT 77.215 145.645 77.505 145.690 ;
        RECT 78.580 145.630 78.900 145.690 ;
        RECT 82.965 145.645 83.500 145.875 ;
        RECT 83.180 145.630 83.500 145.645 ;
        RECT 90.540 145.830 90.860 145.890 ;
        RECT 104.890 145.830 105.030 146.325 ;
        RECT 105.720 146.310 106.040 146.570 ;
        RECT 108.110 146.555 108.250 146.710 ;
        RECT 110.320 146.710 112.005 146.850 ;
        RECT 110.320 146.650 110.640 146.710 ;
        RECT 111.715 146.665 112.005 146.710 ;
        RECT 108.035 146.325 108.325 146.555 ;
        RECT 108.495 146.325 108.785 146.555 ;
        RECT 105.260 146.170 105.580 146.230 ;
        RECT 108.570 146.170 108.710 146.325 ;
        RECT 108.940 146.310 109.260 146.570 ;
        RECT 109.400 146.510 109.720 146.570 ;
        RECT 109.875 146.510 110.165 146.555 ;
        RECT 109.400 146.370 110.165 146.510 ;
        RECT 109.400 146.310 109.720 146.370 ;
        RECT 109.875 146.325 110.165 146.370 ;
        RECT 115.380 146.510 115.700 146.570 ;
        RECT 117.680 146.510 118.000 146.570 ;
        RECT 115.380 146.370 118.000 146.510 ;
        RECT 115.380 146.310 115.700 146.370 ;
        RECT 117.680 146.310 118.000 146.370 ;
        RECT 119.520 146.310 119.840 146.570 ;
        RECT 105.260 146.030 108.710 146.170 ;
        RECT 109.030 146.170 109.170 146.310 ;
        RECT 112.620 146.170 112.940 146.230 ;
        RECT 109.030 146.030 112.940 146.170 ;
        RECT 105.260 145.970 105.580 146.030 ;
        RECT 112.620 145.970 112.940 146.030 ;
        RECT 113.095 145.830 113.385 145.875 ;
        RECT 90.540 145.690 113.385 145.830 ;
        RECT 90.540 145.630 90.860 145.690 ;
        RECT 113.095 145.645 113.385 145.690 ;
        RECT 118.140 145.630 118.460 145.890 ;
        RECT 120.455 145.830 120.745 145.875 ;
        RECT 121.820 145.830 122.140 145.890 ;
        RECT 120.455 145.690 122.140 145.830 ;
        RECT 120.455 145.645 120.745 145.690 ;
        RECT 121.820 145.630 122.140 145.690 ;
        RECT 11.010 145.010 125.890 145.490 ;
        RECT 31.660 144.810 31.980 144.870 ;
        RECT 39.955 144.810 40.245 144.855 ;
        RECT 52.360 144.810 52.680 144.870 ;
        RECT 31.660 144.670 40.245 144.810 ;
        RECT 31.660 144.610 31.980 144.670 ;
        RECT 39.955 144.625 40.245 144.670 ;
        RECT 41.870 144.670 52.680 144.810 ;
        RECT 14.640 144.470 14.960 144.530 ;
        RECT 15.970 144.470 16.260 144.515 ;
        RECT 19.230 144.470 19.520 144.515 ;
        RECT 14.640 144.330 19.520 144.470 ;
        RECT 14.640 144.270 14.960 144.330 ;
        RECT 15.970 144.285 16.260 144.330 ;
        RECT 19.230 144.285 19.520 144.330 ;
        RECT 20.150 144.470 20.440 144.515 ;
        RECT 22.010 144.470 22.300 144.515 ;
        RECT 20.150 144.330 22.300 144.470 ;
        RECT 20.150 144.285 20.440 144.330 ;
        RECT 22.010 144.285 22.300 144.330 ;
        RECT 23.380 144.470 23.700 144.530 ;
        RECT 36.720 144.470 37.040 144.530 ;
        RECT 23.380 144.330 37.040 144.470 ;
        RECT 17.830 144.130 18.120 144.175 ;
        RECT 20.150 144.130 20.365 144.285 ;
        RECT 23.380 144.270 23.700 144.330 ;
        RECT 36.720 144.270 37.040 144.330 ;
        RECT 39.035 144.470 39.325 144.515 ;
        RECT 41.870 144.470 42.010 144.670 ;
        RECT 52.360 144.610 52.680 144.670 ;
        RECT 60.640 144.610 60.960 144.870 ;
        RECT 86.415 144.625 86.705 144.855 ;
        RECT 88.715 144.810 89.005 144.855 ;
        RECT 90.080 144.810 90.400 144.870 ;
        RECT 88.715 144.670 90.400 144.810 ;
        RECT 88.715 144.625 89.005 144.670 ;
        RECT 39.035 144.330 42.010 144.470 ;
        RECT 42.255 144.470 42.545 144.515 ;
        RECT 42.715 144.470 43.005 144.515 ;
        RECT 42.255 144.330 43.005 144.470 ;
        RECT 39.035 144.285 39.325 144.330 ;
        RECT 42.255 144.285 42.545 144.330 ;
        RECT 42.715 144.285 43.005 144.330 ;
        RECT 43.160 144.470 43.480 144.530 ;
        RECT 58.340 144.470 58.660 144.530 ;
        RECT 63.860 144.515 64.180 144.530 ;
        RECT 61.805 144.470 62.095 144.515 ;
        RECT 43.160 144.330 44.770 144.470 ;
        RECT 43.160 144.270 43.480 144.330 ;
        RECT 17.830 143.990 20.365 144.130 ;
        RECT 17.830 143.945 18.120 143.990 ;
        RECT 22.920 143.930 23.240 144.190 ;
        RECT 37.655 143.945 37.945 144.175 ;
        RECT 21.095 143.790 21.385 143.835 ;
        RECT 22.000 143.790 22.320 143.850 ;
        RECT 21.095 143.650 22.320 143.790 ;
        RECT 21.095 143.605 21.385 143.650 ;
        RECT 22.000 143.590 22.320 143.650 ;
        RECT 17.830 143.450 18.120 143.495 ;
        RECT 20.610 143.450 20.900 143.495 ;
        RECT 22.470 143.450 22.760 143.495 ;
        RECT 17.830 143.310 22.760 143.450 ;
        RECT 17.830 143.265 18.120 143.310 ;
        RECT 20.610 143.265 20.900 143.310 ;
        RECT 22.470 143.265 22.760 143.310 ;
        RECT 24.760 143.450 25.080 143.510 ;
        RECT 36.735 143.450 37.025 143.495 ;
        RECT 24.760 143.310 37.025 143.450 ;
        RECT 37.730 143.450 37.870 143.945 ;
        RECT 38.100 143.930 38.420 144.190 ;
        RECT 40.795 144.160 41.085 144.175 ;
        RECT 41.320 144.160 41.640 144.190 ;
        RECT 44.080 144.175 44.400 144.190 ;
        RECT 44.630 144.175 44.770 144.330 ;
        RECT 55.670 144.330 57.190 144.470 ;
        RECT 40.795 144.020 41.640 144.160 ;
        RECT 40.795 143.990 41.090 144.020 ;
        RECT 40.795 143.945 41.085 143.990 ;
        RECT 41.320 143.930 41.640 144.020 ;
        RECT 43.865 143.945 44.400 144.175 ;
        RECT 44.555 143.945 44.845 144.175 ;
        RECT 45.120 144.145 45.410 144.190 ;
        RECT 45.120 144.005 45.690 144.145 ;
        RECT 45.120 143.960 45.410 144.005 ;
        RECT 44.080 143.930 44.400 143.945 ;
        RECT 41.795 143.605 42.085 143.835 ;
        RECT 43.160 143.790 43.480 143.850 ;
        RECT 45.550 143.790 45.690 144.005 ;
        RECT 45.935 143.945 46.225 144.175 ;
        RECT 43.160 143.650 45.690 143.790 ;
        RECT 46.010 143.790 46.150 143.945 ;
        RECT 51.900 143.930 52.220 144.190 ;
        RECT 53.740 144.130 54.060 144.190 ;
        RECT 54.675 144.130 54.965 144.175 ;
        RECT 53.740 143.990 54.965 144.130 ;
        RECT 53.740 143.930 54.060 143.990 ;
        RECT 54.675 143.945 54.965 143.990 ;
        RECT 55.120 143.930 55.440 144.190 ;
        RECT 55.670 144.175 55.810 144.330 ;
        RECT 55.595 143.945 55.885 144.175 ;
        RECT 56.500 143.930 56.820 144.190 ;
        RECT 57.050 144.130 57.190 144.330 ;
        RECT 58.340 144.330 62.095 144.470 ;
        RECT 58.340 144.270 58.660 144.330 ;
        RECT 61.805 144.285 62.095 144.330 ;
        RECT 63.810 144.470 64.180 144.515 ;
        RECT 67.070 144.470 67.360 144.515 ;
        RECT 63.810 144.330 67.360 144.470 ;
        RECT 63.810 144.285 64.180 144.330 ;
        RECT 67.070 144.285 67.360 144.330 ;
        RECT 67.990 144.470 68.280 144.515 ;
        RECT 69.850 144.470 70.140 144.515 ;
        RECT 67.990 144.330 70.140 144.470 ;
        RECT 67.990 144.285 68.280 144.330 ;
        RECT 69.850 144.285 70.140 144.330 ;
        RECT 63.860 144.270 64.180 144.285 ;
        RECT 58.800 144.130 59.120 144.190 ;
        RECT 57.050 143.990 59.120 144.130 ;
        RECT 58.800 143.930 59.120 143.990 ;
        RECT 65.670 144.130 65.960 144.175 ;
        RECT 67.990 144.130 68.205 144.285 ;
        RECT 70.760 144.270 71.080 144.530 ;
        RECT 73.075 144.470 73.365 144.515 ;
        RECT 75.360 144.470 75.680 144.530 ;
        RECT 76.755 144.470 77.045 144.515 ;
        RECT 73.075 144.330 77.045 144.470 ;
        RECT 73.075 144.285 73.365 144.330 ;
        RECT 75.360 144.270 75.680 144.330 ;
        RECT 76.755 144.285 77.045 144.330 ;
        RECT 83.640 144.470 83.960 144.530 ;
        RECT 85.940 144.470 86.260 144.530 ;
        RECT 83.640 144.330 86.260 144.470 ;
        RECT 83.640 144.270 83.960 144.330 ;
        RECT 85.940 144.270 86.260 144.330 ;
        RECT 65.670 143.990 68.205 144.130 ;
        RECT 68.935 144.130 69.225 144.175 ;
        RECT 70.300 144.130 70.620 144.190 ;
        RECT 68.935 143.990 70.620 144.130 ;
        RECT 70.850 144.130 70.990 144.270 ;
        RECT 73.995 144.130 74.285 144.175 ;
        RECT 74.440 144.130 74.760 144.190 ;
        RECT 70.850 143.990 73.750 144.130 ;
        RECT 65.670 143.945 65.960 143.990 ;
        RECT 68.935 143.945 69.225 143.990 ;
        RECT 70.300 143.930 70.620 143.990 ;
        RECT 56.590 143.790 56.730 143.930 ;
        RECT 46.010 143.650 57.190 143.790 ;
        RECT 40.860 143.450 41.180 143.510 ;
        RECT 37.730 143.310 41.180 143.450 ;
        RECT 41.870 143.450 42.010 143.605 ;
        RECT 43.160 143.590 43.480 143.650 ;
        RECT 46.840 143.450 47.160 143.510 ;
        RECT 53.295 143.450 53.585 143.495 ;
        RECT 41.870 143.310 43.850 143.450 ;
        RECT 24.760 143.250 25.080 143.310 ;
        RECT 36.735 143.265 37.025 143.310 ;
        RECT 40.860 143.250 41.180 143.310 ;
        RECT 13.965 143.110 14.255 143.155 ;
        RECT 17.400 143.110 17.720 143.170 ;
        RECT 13.965 142.970 17.720 143.110 ;
        RECT 13.965 142.925 14.255 142.970 ;
        RECT 17.400 142.910 17.720 142.970 ;
        RECT 33.960 143.110 34.280 143.170 ;
        RECT 37.655 143.110 37.945 143.155 ;
        RECT 33.960 142.970 37.945 143.110 ;
        RECT 33.960 142.910 34.280 142.970 ;
        RECT 37.655 142.925 37.945 142.970 ;
        RECT 41.780 142.910 42.100 143.170 ;
        RECT 43.710 143.110 43.850 143.310 ;
        RECT 46.840 143.310 53.585 143.450 ;
        RECT 57.050 143.450 57.190 143.650 ;
        RECT 57.420 143.590 57.740 143.850 ;
        RECT 65.240 143.790 65.560 143.850 ;
        RECT 70.775 143.790 71.065 143.835 ;
        RECT 65.240 143.650 71.065 143.790 ;
        RECT 65.240 143.590 65.560 143.650 ;
        RECT 70.775 143.605 71.065 143.650 ;
        RECT 61.100 143.450 61.420 143.510 ;
        RECT 57.050 143.310 61.420 143.450 ;
        RECT 46.840 143.250 47.160 143.310 ;
        RECT 53.295 143.265 53.585 143.310 ;
        RECT 61.100 143.250 61.420 143.310 ;
        RECT 65.670 143.450 65.960 143.495 ;
        RECT 68.450 143.450 68.740 143.495 ;
        RECT 70.310 143.450 70.600 143.495 ;
        RECT 65.670 143.310 70.600 143.450 ;
        RECT 73.610 143.450 73.750 143.990 ;
        RECT 73.995 143.990 74.760 144.130 ;
        RECT 73.995 143.945 74.285 143.990 ;
        RECT 74.440 143.930 74.760 143.990 ;
        RECT 80.420 144.130 80.740 144.190 ;
        RECT 83.180 144.130 83.500 144.190 ;
        RECT 84.115 144.130 84.405 144.175 ;
        RECT 80.420 143.990 84.405 144.130 ;
        RECT 80.420 143.930 80.740 143.990 ;
        RECT 83.180 143.930 83.500 143.990 ;
        RECT 84.115 143.945 84.405 143.990 ;
        RECT 78.135 143.790 78.425 143.835 ;
        RECT 81.800 143.790 82.120 143.850 ;
        RECT 83.640 143.790 83.960 143.850 ;
        RECT 78.135 143.650 83.960 143.790 ;
        RECT 84.190 143.790 84.330 143.945 ;
        RECT 84.560 143.930 84.880 144.190 ;
        RECT 86.490 144.130 86.630 144.625 ;
        RECT 90.080 144.610 90.400 144.670 ;
        RECT 90.540 144.610 90.860 144.870 ;
        RECT 92.855 144.810 93.145 144.855 ;
        RECT 94.220 144.810 94.540 144.870 ;
        RECT 108.940 144.810 109.260 144.870 ;
        RECT 92.855 144.670 94.540 144.810 ;
        RECT 92.855 144.625 93.145 144.670 ;
        RECT 94.220 144.610 94.540 144.670 ;
        RECT 108.110 144.670 109.260 144.810 ;
        RECT 86.860 144.470 87.180 144.530 ;
        RECT 102.975 144.470 103.265 144.515 ;
        RECT 107.115 144.470 107.405 144.515 ;
        RECT 86.860 144.330 91.690 144.470 ;
        RECT 86.860 144.270 87.180 144.330 ;
        RECT 87.795 144.130 88.085 144.175 ;
        RECT 91.015 144.130 91.305 144.175 ;
        RECT 86.490 143.990 88.085 144.130 ;
        RECT 87.795 143.945 88.085 143.990 ;
        RECT 89.710 143.990 91.305 144.130 ;
        RECT 89.710 143.790 89.850 143.990 ;
        RECT 91.015 143.945 91.305 143.990 ;
        RECT 84.190 143.650 89.850 143.790 ;
        RECT 90.095 143.790 90.385 143.835 ;
        RECT 91.550 143.790 91.690 144.330 ;
        RECT 102.975 144.330 107.405 144.470 ;
        RECT 102.975 144.285 103.265 144.330 ;
        RECT 107.115 144.285 107.405 144.330 ;
        RECT 101.595 144.130 101.885 144.175 ;
        RECT 102.040 144.130 102.360 144.190 ;
        RECT 101.595 143.990 102.360 144.130 ;
        RECT 101.595 143.945 101.885 143.990 ;
        RECT 102.040 143.930 102.360 143.990 ;
        RECT 103.895 144.130 104.185 144.175 ;
        RECT 108.110 144.130 108.250 144.670 ;
        RECT 108.940 144.610 109.260 144.670 ;
        RECT 116.710 144.470 117.000 144.515 ;
        RECT 118.140 144.470 118.460 144.530 ;
        RECT 119.970 144.470 120.260 144.515 ;
        RECT 116.710 144.330 120.260 144.470 ;
        RECT 116.710 144.285 117.000 144.330 ;
        RECT 118.140 144.270 118.460 144.330 ;
        RECT 119.970 144.285 120.260 144.330 ;
        RECT 120.890 144.470 121.180 144.515 ;
        RECT 122.750 144.470 123.040 144.515 ;
        RECT 120.890 144.330 123.040 144.470 ;
        RECT 120.890 144.285 121.180 144.330 ;
        RECT 122.750 144.285 123.040 144.330 ;
        RECT 103.895 143.990 108.250 144.130 ;
        RECT 103.895 143.945 104.185 143.990 ;
        RECT 108.495 143.945 108.785 144.175 ;
        RECT 108.955 143.945 109.245 144.175 ;
        RECT 90.095 143.650 91.690 143.790 ;
        RECT 78.135 143.605 78.425 143.650 ;
        RECT 81.800 143.590 82.120 143.650 ;
        RECT 83.640 143.590 83.960 143.650 ;
        RECT 90.095 143.605 90.385 143.650 ;
        RECT 102.500 143.590 102.820 143.850 ;
        RECT 108.570 143.790 108.710 143.945 ;
        RECT 103.970 143.650 108.710 143.790 ;
        RECT 103.970 143.510 104.110 143.650 ;
        RECT 97.440 143.450 97.760 143.510 ;
        RECT 103.880 143.450 104.200 143.510 ;
        RECT 73.610 143.310 104.200 143.450 ;
        RECT 65.670 143.265 65.960 143.310 ;
        RECT 68.450 143.265 68.740 143.310 ;
        RECT 70.310 143.265 70.600 143.310 ;
        RECT 97.440 143.250 97.760 143.310 ;
        RECT 103.880 143.250 104.200 143.310 ;
        RECT 104.340 143.450 104.660 143.510 ;
        RECT 109.030 143.450 109.170 143.945 ;
        RECT 109.400 143.930 109.720 144.190 ;
        RECT 109.860 144.130 110.180 144.190 ;
        RECT 110.335 144.130 110.625 144.175 ;
        RECT 109.860 143.990 110.625 144.130 ;
        RECT 109.860 143.930 110.180 143.990 ;
        RECT 110.335 143.945 110.625 143.990 ;
        RECT 118.570 144.130 118.860 144.175 ;
        RECT 120.890 144.130 121.105 144.285 ;
        RECT 118.570 143.990 121.105 144.130 ;
        RECT 118.570 143.945 118.860 143.990 ;
        RECT 121.820 143.930 122.140 144.190 ;
        RECT 109.490 143.790 109.630 143.930 ;
        RECT 114.920 143.835 115.240 143.850 ;
        RECT 114.705 143.790 115.240 143.835 ;
        RECT 109.490 143.650 115.240 143.790 ;
        RECT 114.705 143.605 115.240 143.650 ;
        RECT 114.920 143.590 115.240 143.605 ;
        RECT 122.280 143.790 122.600 143.850 ;
        RECT 123.675 143.790 123.965 143.835 ;
        RECT 122.280 143.650 123.965 143.790 ;
        RECT 122.280 143.590 122.600 143.650 ;
        RECT 123.675 143.605 123.965 143.650 ;
        RECT 104.340 143.310 109.170 143.450 ;
        RECT 118.570 143.450 118.860 143.495 ;
        RECT 121.350 143.450 121.640 143.495 ;
        RECT 123.210 143.450 123.500 143.495 ;
        RECT 118.570 143.310 123.500 143.450 ;
        RECT 104.340 143.250 104.660 143.310 ;
        RECT 118.570 143.265 118.860 143.310 ;
        RECT 121.350 143.265 121.640 143.310 ;
        RECT 123.210 143.265 123.500 143.310 ;
        RECT 50.060 143.110 50.380 143.170 ;
        RECT 43.710 142.970 50.380 143.110 ;
        RECT 50.060 142.910 50.380 142.970 ;
        RECT 52.835 143.110 53.125 143.155 ;
        RECT 56.040 143.110 56.360 143.170 ;
        RECT 52.835 142.970 56.360 143.110 ;
        RECT 52.835 142.925 53.125 142.970 ;
        RECT 56.040 142.910 56.360 142.970 ;
        RECT 69.840 143.110 70.160 143.170 ;
        RECT 71.695 143.110 71.985 143.155 ;
        RECT 69.840 142.970 71.985 143.110 ;
        RECT 69.840 142.910 70.160 142.970 ;
        RECT 71.695 142.925 71.985 142.970 ;
        RECT 74.915 143.110 75.205 143.155 ;
        RECT 79.040 143.110 79.360 143.170 ;
        RECT 74.915 142.970 79.360 143.110 ;
        RECT 74.915 142.925 75.205 142.970 ;
        RECT 79.040 142.910 79.360 142.970 ;
        RECT 84.100 143.110 84.420 143.170 ;
        RECT 97.900 143.110 98.220 143.170 ;
        RECT 84.100 142.970 98.220 143.110 ;
        RECT 84.100 142.910 84.420 142.970 ;
        RECT 97.900 142.910 98.220 142.970 ;
        RECT 100.660 142.910 100.980 143.170 ;
        RECT 102.975 143.110 103.265 143.155 ;
        RECT 105.260 143.110 105.580 143.170 ;
        RECT 102.975 142.970 105.580 143.110 ;
        RECT 102.975 142.925 103.265 142.970 ;
        RECT 105.260 142.910 105.580 142.970 ;
        RECT 106.640 142.910 106.960 143.170 ;
        RECT 11.810 142.290 125.890 142.770 ;
        RECT 22.000 141.890 22.320 142.150 ;
        RECT 33.960 141.890 34.280 142.150 ;
        RECT 34.880 142.090 35.200 142.150 ;
        RECT 35.355 142.090 35.645 142.135 ;
        RECT 37.195 142.090 37.485 142.135 ;
        RECT 34.880 141.950 35.645 142.090 ;
        RECT 34.880 141.890 35.200 141.950 ;
        RECT 35.355 141.905 35.645 141.950 ;
        RECT 36.350 141.950 37.485 142.090 ;
        RECT 33.040 141.750 33.360 141.810 ;
        RECT 36.350 141.750 36.490 141.950 ;
        RECT 37.195 141.905 37.485 141.950 ;
        RECT 37.640 142.090 37.960 142.150 ;
        RECT 38.575 142.090 38.865 142.135 ;
        RECT 37.640 141.950 38.865 142.090 ;
        RECT 37.640 141.890 37.960 141.950 ;
        RECT 38.575 141.905 38.865 141.950 ;
        RECT 41.780 141.890 42.100 142.150 ;
        RECT 57.895 142.090 58.185 142.135 ;
        RECT 47.390 141.950 58.185 142.090 ;
        RECT 18.180 141.610 32.350 141.750 ;
        RECT 17.400 141.410 17.720 141.470 ;
        RECT 18.180 141.410 18.320 141.610 ;
        RECT 17.400 141.270 18.320 141.410 ;
        RECT 19.700 141.410 20.020 141.470 ;
        RECT 27.075 141.410 27.365 141.455 ;
        RECT 30.740 141.410 31.060 141.470 ;
        RECT 32.210 141.455 32.350 141.610 ;
        RECT 33.040 141.610 36.490 141.750 ;
        RECT 38.100 141.750 38.420 141.810 ;
        RECT 46.380 141.750 46.700 141.810 ;
        RECT 38.100 141.610 46.700 141.750 ;
        RECT 33.040 141.550 33.360 141.610 ;
        RECT 38.100 141.550 38.420 141.610 ;
        RECT 46.380 141.550 46.700 141.610 ;
        RECT 19.700 141.270 24.530 141.410 ;
        RECT 17.400 141.210 17.720 141.270 ;
        RECT 19.700 141.210 20.020 141.270 ;
        RECT 19.240 141.070 19.560 141.130 ;
        RECT 21.095 141.070 21.385 141.115 ;
        RECT 19.240 140.930 21.385 141.070 ;
        RECT 19.240 140.870 19.560 140.930 ;
        RECT 21.095 140.885 21.385 140.930 ;
        RECT 22.935 140.885 23.225 141.115 ;
        RECT 24.390 141.070 24.530 141.270 ;
        RECT 27.075 141.270 31.060 141.410 ;
        RECT 27.075 141.225 27.365 141.270 ;
        RECT 30.740 141.210 31.060 141.270 ;
        RECT 32.135 141.225 32.425 141.455 ;
        RECT 36.260 141.210 36.580 141.470 ;
        RECT 37.180 141.410 37.500 141.470 ;
        RECT 38.575 141.410 38.865 141.455 ;
        RECT 37.180 141.270 38.865 141.410 ;
        RECT 37.180 141.210 37.500 141.270 ;
        RECT 38.575 141.225 38.865 141.270 ;
        RECT 39.940 141.210 40.260 141.470 ;
        RECT 46.840 141.410 47.160 141.470 ;
        RECT 40.490 141.270 47.160 141.410 ;
        RECT 27.995 141.070 28.285 141.115 ;
        RECT 33.055 141.070 33.345 141.115 ;
        RECT 33.500 141.070 33.820 141.130 ;
        RECT 24.390 140.930 32.120 141.070 ;
        RECT 27.995 140.885 28.285 140.930 ;
        RECT 15.100 140.730 15.420 140.790 ;
        RECT 23.010 140.730 23.150 140.885 ;
        RECT 15.100 140.590 23.150 140.730 ;
        RECT 31.980 140.730 32.120 140.930 ;
        RECT 33.055 140.930 33.820 141.070 ;
        RECT 33.055 140.885 33.345 140.930 ;
        RECT 33.500 140.870 33.820 140.930 ;
        RECT 35.340 140.870 35.660 141.130 ;
        RECT 38.100 140.870 38.420 141.130 ;
        RECT 39.495 141.070 39.785 141.115 ;
        RECT 40.490 141.070 40.630 141.270 ;
        RECT 46.840 141.210 47.160 141.270 ;
        RECT 39.495 140.930 40.630 141.070 ;
        RECT 40.875 141.070 41.165 141.115 ;
        RECT 41.780 141.070 42.100 141.130 ;
        RECT 40.875 140.930 42.100 141.070 ;
        RECT 39.495 140.885 39.785 140.930 ;
        RECT 40.875 140.885 41.165 140.930 ;
        RECT 41.780 140.870 42.100 140.930 ;
        RECT 36.735 140.730 37.025 140.775 ;
        RECT 47.390 140.730 47.530 141.950 ;
        RECT 57.895 141.905 58.185 141.950 ;
        RECT 68.920 142.090 69.240 142.150 ;
        RECT 77.675 142.090 77.965 142.135 ;
        RECT 79.500 142.090 79.820 142.150 ;
        RECT 68.920 141.950 77.430 142.090 ;
        RECT 68.920 141.890 69.240 141.950 ;
        RECT 51.555 141.750 51.845 141.795 ;
        RECT 54.675 141.750 54.965 141.795 ;
        RECT 56.565 141.750 56.855 141.795 ;
        RECT 51.555 141.610 56.855 141.750 ;
        RECT 51.555 141.565 51.845 141.610 ;
        RECT 54.675 141.565 54.965 141.610 ;
        RECT 56.565 141.565 56.855 141.610 ;
        RECT 67.970 141.750 68.260 141.795 ;
        RECT 70.750 141.750 71.040 141.795 ;
        RECT 72.610 141.750 72.900 141.795 ;
        RECT 67.970 141.610 72.900 141.750 ;
        RECT 77.290 141.750 77.430 141.950 ;
        RECT 77.675 141.950 79.820 142.090 ;
        RECT 77.675 141.905 77.965 141.950 ;
        RECT 79.500 141.890 79.820 141.950 ;
        RECT 85.570 141.950 93.530 142.090 ;
        RECT 85.570 141.750 85.710 141.950 ;
        RECT 77.290 141.610 85.710 141.750 ;
        RECT 85.910 141.750 86.200 141.795 ;
        RECT 88.690 141.750 88.980 141.795 ;
        RECT 90.550 141.750 90.840 141.795 ;
        RECT 85.910 141.610 90.840 141.750 ;
        RECT 93.390 141.750 93.530 141.950 ;
        RECT 93.760 141.890 94.080 142.150 ;
        RECT 97.900 142.090 98.220 142.150 ;
        RECT 104.340 142.090 104.660 142.150 ;
        RECT 97.900 141.950 104.660 142.090 ;
        RECT 97.900 141.890 98.220 141.950 ;
        RECT 104.340 141.890 104.660 141.950 ;
        RECT 106.640 142.090 106.960 142.150 ;
        RECT 117.235 142.090 117.525 142.135 ;
        RECT 119.520 142.090 119.840 142.150 ;
        RECT 106.640 141.950 115.610 142.090 ;
        RECT 106.640 141.890 106.960 141.950 ;
        RECT 105.720 141.750 106.040 141.810 ;
        RECT 93.390 141.610 107.330 141.750 ;
        RECT 67.970 141.565 68.260 141.610 ;
        RECT 70.750 141.565 71.040 141.610 ;
        RECT 72.610 141.565 72.900 141.610 ;
        RECT 85.910 141.565 86.200 141.610 ;
        RECT 88.690 141.565 88.980 141.610 ;
        RECT 90.550 141.565 90.840 141.610 ;
        RECT 56.040 141.210 56.360 141.470 ;
        RECT 57.435 141.410 57.725 141.455 ;
        RECT 57.435 141.270 70.990 141.410 ;
        RECT 57.435 141.225 57.725 141.270 ;
        RECT 70.850 141.130 70.990 141.270 ;
        RECT 71.220 141.210 71.540 141.470 ;
        RECT 73.980 141.410 74.300 141.470 ;
        RECT 77.215 141.410 77.505 141.455 ;
        RECT 73.980 141.270 77.505 141.410 ;
        RECT 73.980 141.210 74.300 141.270 ;
        RECT 77.215 141.225 77.505 141.270 ;
        RECT 91.015 141.410 91.305 141.455 ;
        RECT 91.920 141.410 92.240 141.470 ;
        RECT 91.015 141.270 92.240 141.410 ;
        RECT 91.015 141.225 91.305 141.270 ;
        RECT 91.920 141.210 92.240 141.270 ;
        RECT 94.235 141.410 94.525 141.455 ;
        RECT 94.235 141.270 97.210 141.410 ;
        RECT 94.235 141.225 94.525 141.270 ;
        RECT 50.475 140.775 50.765 141.090 ;
        RECT 51.555 141.070 51.845 141.115 ;
        RECT 55.135 141.070 55.425 141.115 ;
        RECT 56.970 141.070 57.260 141.115 ;
        RECT 51.555 140.930 57.260 141.070 ;
        RECT 51.555 140.885 51.845 140.930 ;
        RECT 55.135 140.885 55.425 140.930 ;
        RECT 56.970 140.885 57.260 140.930 ;
        RECT 59.260 140.870 59.580 141.130 ;
        RECT 59.720 140.870 60.040 141.130 ;
        RECT 60.180 140.870 60.500 141.130 ;
        RECT 61.100 141.070 61.420 141.130 ;
        RECT 67.970 141.070 68.260 141.115 ;
        RECT 70.760 141.070 71.080 141.130 ;
        RECT 73.075 141.070 73.365 141.115 ;
        RECT 61.100 140.930 65.010 141.070 ;
        RECT 61.100 140.870 61.420 140.930 ;
        RECT 31.980 140.590 35.110 140.730 ;
        RECT 15.100 140.530 15.420 140.590 ;
        RECT 23.380 140.190 23.700 140.450 ;
        RECT 27.520 140.190 27.840 140.450 ;
        RECT 29.820 140.190 30.140 140.450 ;
        RECT 33.960 140.390 34.280 140.450 ;
        RECT 34.435 140.390 34.725 140.435 ;
        RECT 33.960 140.250 34.725 140.390 ;
        RECT 34.970 140.390 35.110 140.590 ;
        RECT 36.735 140.590 47.530 140.730 ;
        RECT 50.175 140.730 50.765 140.775 ;
        RECT 52.360 140.730 52.680 140.790 ;
        RECT 53.415 140.730 54.065 140.775 ;
        RECT 50.175 140.590 54.065 140.730 ;
        RECT 36.735 140.545 37.025 140.590 ;
        RECT 50.175 140.545 50.465 140.590 ;
        RECT 52.360 140.530 52.680 140.590 ;
        RECT 53.415 140.545 54.065 140.590 ;
        RECT 39.940 140.390 40.260 140.450 ;
        RECT 34.970 140.250 40.260 140.390 ;
        RECT 33.960 140.190 34.280 140.250 ;
        RECT 34.435 140.205 34.725 140.250 ;
        RECT 39.940 140.190 40.260 140.250 ;
        RECT 48.695 140.390 48.985 140.435 ;
        RECT 49.600 140.390 49.920 140.450 ;
        RECT 48.695 140.250 49.920 140.390 ;
        RECT 48.695 140.205 48.985 140.250 ;
        RECT 49.600 140.190 49.920 140.250 ;
        RECT 62.940 140.390 63.260 140.450 ;
        RECT 64.105 140.390 64.395 140.435 ;
        RECT 62.940 140.250 64.395 140.390 ;
        RECT 64.870 140.390 65.010 140.930 ;
        RECT 67.970 140.930 70.505 141.070 ;
        RECT 67.970 140.885 68.260 140.930 ;
        RECT 66.110 140.730 66.400 140.775 ;
        RECT 67.540 140.730 67.860 140.790 ;
        RECT 70.290 140.775 70.505 140.930 ;
        RECT 70.760 140.930 73.365 141.070 ;
        RECT 70.760 140.870 71.080 140.930 ;
        RECT 73.075 140.885 73.365 140.930 ;
        RECT 76.295 141.070 76.585 141.115 ;
        RECT 76.740 141.070 77.060 141.130 ;
        RECT 76.295 140.930 77.060 141.070 ;
        RECT 76.295 140.885 76.585 140.930 ;
        RECT 76.740 140.870 77.060 140.930 ;
        RECT 79.040 141.070 79.360 141.130 ;
        RECT 79.515 141.070 79.805 141.115 ;
        RECT 79.040 140.930 79.805 141.070 ;
        RECT 79.040 140.870 79.360 140.930 ;
        RECT 79.515 140.885 79.805 140.930 ;
        RECT 79.960 140.870 80.280 141.130 ;
        RECT 80.420 140.870 80.740 141.130 ;
        RECT 81.340 140.870 81.660 141.130 ;
        RECT 85.910 141.070 86.200 141.115 ;
        RECT 85.910 140.930 88.445 141.070 ;
        RECT 85.910 140.885 86.200 140.930 ;
        RECT 69.370 140.730 69.660 140.775 ;
        RECT 66.110 140.590 69.660 140.730 ;
        RECT 66.110 140.545 66.400 140.590 ;
        RECT 67.540 140.530 67.860 140.590 ;
        RECT 69.370 140.545 69.660 140.590 ;
        RECT 70.290 140.730 70.580 140.775 ;
        RECT 72.150 140.730 72.440 140.775 ;
        RECT 70.290 140.590 72.440 140.730 ;
        RECT 70.290 140.545 70.580 140.590 ;
        RECT 72.150 140.545 72.440 140.590 ;
        RECT 77.675 140.730 77.965 140.775 ;
        RECT 78.135 140.730 78.425 140.775 ;
        RECT 77.675 140.590 78.425 140.730 ;
        RECT 77.675 140.545 77.965 140.590 ;
        RECT 78.135 140.545 78.425 140.590 ;
        RECT 84.050 140.730 84.340 140.775 ;
        RECT 86.400 140.730 86.720 140.790 ;
        RECT 88.230 140.775 88.445 140.930 ;
        RECT 89.160 140.870 89.480 141.130 ;
        RECT 94.680 140.870 95.000 141.130 ;
        RECT 87.310 140.730 87.600 140.775 ;
        RECT 84.050 140.590 87.600 140.730 ;
        RECT 84.050 140.545 84.340 140.590 ;
        RECT 86.400 140.530 86.720 140.590 ;
        RECT 87.310 140.545 87.600 140.590 ;
        RECT 88.230 140.730 88.520 140.775 ;
        RECT 90.090 140.730 90.380 140.775 ;
        RECT 88.230 140.590 90.380 140.730 ;
        RECT 88.230 140.545 88.520 140.590 ;
        RECT 90.090 140.545 90.380 140.590 ;
        RECT 93.315 140.730 93.605 140.775 ;
        RECT 96.075 140.730 96.365 140.775 ;
        RECT 93.315 140.590 96.365 140.730 ;
        RECT 93.315 140.545 93.605 140.590 ;
        RECT 96.075 140.545 96.365 140.590 ;
        RECT 68.920 140.390 69.240 140.450 ;
        RECT 64.870 140.250 69.240 140.390 ;
        RECT 62.940 140.190 63.260 140.250 ;
        RECT 64.105 140.205 64.395 140.250 ;
        RECT 68.920 140.190 69.240 140.250 ;
        RECT 75.360 140.190 75.680 140.450 ;
        RECT 80.420 140.390 80.740 140.450 ;
        RECT 82.045 140.390 82.335 140.435 ;
        RECT 84.560 140.390 84.880 140.450 ;
        RECT 80.420 140.250 84.880 140.390 ;
        RECT 80.420 140.190 80.740 140.250 ;
        RECT 82.045 140.205 82.335 140.250 ;
        RECT 84.560 140.190 84.880 140.250 ;
        RECT 95.140 140.390 95.460 140.450 ;
        RECT 95.615 140.390 95.905 140.435 ;
        RECT 95.140 140.250 95.905 140.390 ;
        RECT 97.070 140.390 97.210 141.270 ;
        RECT 97.440 140.870 97.760 141.130 ;
        RECT 97.900 140.870 98.220 141.130 ;
        RECT 99.370 141.115 99.510 141.610 ;
        RECT 105.720 141.550 106.040 141.610 ;
        RECT 104.340 141.410 104.660 141.470 ;
        RECT 106.640 141.410 106.960 141.470 ;
        RECT 104.340 141.270 106.960 141.410 ;
        RECT 104.340 141.210 104.660 141.270 ;
        RECT 98.375 140.885 98.665 141.115 ;
        RECT 99.295 140.885 99.585 141.115 ;
        RECT 103.880 141.070 104.200 141.130 ;
        RECT 104.800 141.070 105.120 141.130 ;
        RECT 105.810 141.115 105.950 141.270 ;
        RECT 106.640 141.210 106.960 141.270 ;
        RECT 107.190 141.115 107.330 141.610 ;
        RECT 108.940 141.410 109.260 141.470 ;
        RECT 109.875 141.410 110.165 141.455 ;
        RECT 110.320 141.410 110.640 141.470 ;
        RECT 114.015 141.410 114.305 141.455 ;
        RECT 108.940 141.270 114.305 141.410 ;
        RECT 108.940 141.210 109.260 141.270 ;
        RECT 109.875 141.225 110.165 141.270 ;
        RECT 110.320 141.210 110.640 141.270 ;
        RECT 114.015 141.225 114.305 141.270 ;
        RECT 114.920 141.210 115.240 141.470 ;
        RECT 105.275 141.070 105.565 141.115 ;
        RECT 103.880 140.930 105.565 141.070 ;
        RECT 98.450 140.730 98.590 140.885 ;
        RECT 103.880 140.870 104.200 140.930 ;
        RECT 104.800 140.870 105.120 140.930 ;
        RECT 105.275 140.885 105.565 140.930 ;
        RECT 105.735 140.885 106.025 141.115 ;
        RECT 106.195 140.885 106.485 141.115 ;
        RECT 107.115 141.070 107.405 141.115 ;
        RECT 108.480 141.070 108.800 141.130 ;
        RECT 115.470 141.115 115.610 141.950 ;
        RECT 117.235 141.950 119.840 142.090 ;
        RECT 117.235 141.905 117.525 141.950 ;
        RECT 119.520 141.890 119.840 141.950 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 107.115 140.930 108.800 141.070 ;
        RECT 107.115 140.885 107.405 140.930 ;
        RECT 99.740 140.730 100.060 140.790 ;
        RECT 98.450 140.590 100.060 140.730 ;
        RECT 106.270 140.730 106.410 140.885 ;
        RECT 108.480 140.870 108.800 140.930 ;
        RECT 115.395 140.885 115.685 141.115 ;
        RECT 117.680 140.870 118.000 141.130 ;
        RECT 119.535 140.885 119.825 141.115 ;
        RECT 108.020 140.730 108.340 140.790 ;
        RECT 110.795 140.730 111.085 140.775 ;
        RECT 106.270 140.590 111.085 140.730 ;
        RECT 99.740 140.530 100.060 140.590 ;
        RECT 108.020 140.530 108.340 140.590 ;
        RECT 110.795 140.545 111.085 140.590 ;
        RECT 112.160 140.730 112.480 140.790 ;
        RECT 119.610 140.730 119.750 140.885 ;
        RECT 112.160 140.590 119.750 140.730 ;
        RECT 112.160 140.530 112.480 140.590 ;
        RECT 100.200 140.390 100.520 140.450 ;
        RECT 97.070 140.250 100.520 140.390 ;
        RECT 95.140 140.190 95.460 140.250 ;
        RECT 95.615 140.205 95.905 140.250 ;
        RECT 100.200 140.190 100.520 140.250 ;
        RECT 103.880 140.190 104.200 140.450 ;
        RECT 111.240 140.190 111.560 140.450 ;
        RECT 113.080 140.190 113.400 140.450 ;
        RECT 118.140 140.190 118.460 140.450 ;
        RECT 120.455 140.390 120.745 140.435 ;
        RECT 121.820 140.390 122.140 140.450 ;
        RECT 120.455 140.250 122.140 140.390 ;
        RECT 120.455 140.205 120.745 140.250 ;
        RECT 121.820 140.190 122.140 140.250 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 11.010 139.570 125.890 140.050 ;
        RECT 14.640 139.170 14.960 139.430 ;
        RECT 17.400 139.170 17.720 139.430 ;
        RECT 19.240 139.170 19.560 139.430 ;
        RECT 29.375 139.185 29.665 139.415 ;
        RECT 34.880 139.370 35.200 139.430 ;
        RECT 34.880 139.230 37.410 139.370 ;
        RECT 19.700 139.075 20.020 139.090 ;
        RECT 16.955 139.030 17.245 139.075 ;
        RECT 19.700 139.030 20.235 139.075 ;
        RECT 16.955 138.890 20.235 139.030 ;
        RECT 16.955 138.845 17.245 138.890 ;
        RECT 19.700 138.845 20.235 138.890 ;
        RECT 21.950 139.030 22.240 139.075 ;
        RECT 23.380 139.030 23.700 139.090 ;
        RECT 25.210 139.030 25.500 139.075 ;
        RECT 21.950 138.890 25.500 139.030 ;
        RECT 21.950 138.845 22.240 138.890 ;
        RECT 19.700 138.830 20.020 138.845 ;
        RECT 23.380 138.830 23.700 138.890 ;
        RECT 25.210 138.845 25.500 138.890 ;
        RECT 26.130 139.030 26.420 139.075 ;
        RECT 27.990 139.030 28.280 139.075 ;
        RECT 26.130 138.890 28.280 139.030 ;
        RECT 26.130 138.845 26.420 138.890 ;
        RECT 27.990 138.845 28.280 138.890 ;
        RECT 15.100 138.490 15.420 138.750 ;
        RECT 23.810 138.690 24.100 138.735 ;
        RECT 26.130 138.690 26.345 138.845 ;
        RECT 23.810 138.550 26.345 138.690 ;
        RECT 27.075 138.690 27.365 138.735 ;
        RECT 29.450 138.690 29.590 139.185 ;
        RECT 34.880 139.170 35.200 139.230 ;
        RECT 33.500 139.030 33.820 139.090 ;
        RECT 37.270 139.030 37.410 139.230 ;
        RECT 37.640 139.170 37.960 139.430 ;
        RECT 38.115 139.185 38.405 139.415 ;
        RECT 51.915 139.370 52.205 139.415 ;
        RECT 52.360 139.370 52.680 139.430 ;
        RECT 51.915 139.230 52.680 139.370 ;
        RECT 51.915 139.185 52.205 139.230 ;
        RECT 38.190 139.030 38.330 139.185 ;
        RECT 52.360 139.170 52.680 139.230 ;
        RECT 55.135 139.370 55.425 139.415 ;
        RECT 55.580 139.370 55.900 139.430 ;
        RECT 62.940 139.370 63.260 139.430 ;
        RECT 55.135 139.230 63.260 139.370 ;
        RECT 55.135 139.185 55.425 139.230 ;
        RECT 55.580 139.170 55.900 139.230 ;
        RECT 62.940 139.170 63.260 139.230 ;
        RECT 67.540 139.170 67.860 139.430 ;
        RECT 71.220 139.170 71.540 139.430 ;
        RECT 72.615 139.370 72.905 139.415 ;
        RECT 79.960 139.370 80.280 139.430 ;
        RECT 72.615 139.230 80.280 139.370 ;
        RECT 72.615 139.185 72.905 139.230 ;
        RECT 33.500 138.890 36.950 139.030 ;
        RECT 37.270 138.890 38.330 139.030 ;
        RECT 44.095 139.030 44.385 139.075 ;
        RECT 47.315 139.030 47.605 139.075 ;
        RECT 44.095 138.890 47.605 139.030 ;
        RECT 33.500 138.830 33.820 138.890 ;
        RECT 27.075 138.550 29.590 138.690 ;
        RECT 29.820 138.690 30.140 138.750 ;
        RECT 36.810 138.735 36.950 138.890 ;
        RECT 44.095 138.845 44.385 138.890 ;
        RECT 47.315 138.845 47.605 138.890 ;
        RECT 30.295 138.690 30.585 138.735 ;
        RECT 33.055 138.690 33.345 138.735 ;
        RECT 35.815 138.690 36.105 138.735 ;
        RECT 29.820 138.550 30.585 138.690 ;
        RECT 23.810 138.505 24.100 138.550 ;
        RECT 27.075 138.505 27.365 138.550 ;
        RECT 29.820 138.490 30.140 138.550 ;
        RECT 30.295 138.505 30.585 138.550 ;
        RECT 32.210 138.550 36.105 138.690 ;
        RECT 16.480 138.150 16.800 138.410 ;
        RECT 27.980 138.350 28.300 138.410 ;
        RECT 28.915 138.350 29.205 138.395 ;
        RECT 27.980 138.210 29.205 138.350 ;
        RECT 27.980 138.150 28.300 138.210 ;
        RECT 28.915 138.165 29.205 138.210 ;
        RECT 30.740 138.350 31.060 138.410 ;
        RECT 31.675 138.350 31.965 138.395 ;
        RECT 30.740 138.210 31.965 138.350 ;
        RECT 30.740 138.150 31.060 138.210 ;
        RECT 31.675 138.165 31.965 138.210 ;
        RECT 23.810 138.010 24.100 138.055 ;
        RECT 26.590 138.010 26.880 138.055 ;
        RECT 28.450 138.010 28.740 138.055 ;
        RECT 23.810 137.870 28.740 138.010 ;
        RECT 23.810 137.825 24.100 137.870 ;
        RECT 26.590 137.825 26.880 137.870 ;
        RECT 28.450 137.825 28.740 137.870 ;
        RECT 27.520 137.670 27.840 137.730 ;
        RECT 32.210 137.670 32.350 138.550 ;
        RECT 33.055 138.505 33.345 138.550 ;
        RECT 35.815 138.505 36.105 138.550 ;
        RECT 36.735 138.690 37.025 138.735 ;
        RECT 39.035 138.690 39.325 138.735 ;
        RECT 41.780 138.690 42.100 138.750 ;
        RECT 36.735 138.550 42.100 138.690 ;
        RECT 36.735 138.505 37.025 138.550 ;
        RECT 39.035 138.505 39.325 138.550 ;
        RECT 41.780 138.490 42.100 138.550 ;
        RECT 45.000 138.490 45.320 138.750 ;
        RECT 45.475 138.505 45.765 138.735 ;
        RECT 48.220 138.690 48.540 138.750 ;
        RECT 48.695 138.690 48.985 138.735 ;
        RECT 48.220 138.550 48.985 138.690 ;
        RECT 32.580 138.350 32.900 138.410 ;
        RECT 39.955 138.350 40.245 138.395 ;
        RECT 32.580 138.210 40.245 138.350 ;
        RECT 32.580 138.150 32.900 138.210 ;
        RECT 39.955 138.165 40.245 138.210 ;
        RECT 44.540 138.350 44.860 138.410 ;
        RECT 45.550 138.350 45.690 138.505 ;
        RECT 48.220 138.490 48.540 138.550 ;
        RECT 48.695 138.505 48.985 138.550 ;
        RECT 49.155 138.505 49.445 138.735 ;
        RECT 44.540 138.210 45.690 138.350 ;
        RECT 44.540 138.150 44.860 138.210 ;
        RECT 49.230 138.010 49.370 138.505 ;
        RECT 49.600 138.490 49.920 138.750 ;
        RECT 50.520 138.490 50.840 138.750 ;
        RECT 50.980 138.690 51.300 138.750 ;
        RECT 52.360 138.690 52.680 138.750 ;
        RECT 50.980 138.550 52.680 138.690 ;
        RECT 50.980 138.490 51.300 138.550 ;
        RECT 52.360 138.490 52.680 138.550 ;
        RECT 61.560 138.490 61.880 138.750 ;
        RECT 63.030 138.735 63.170 139.170 ;
        RECT 66.175 139.030 66.465 139.075 ;
        RECT 69.855 139.030 70.145 139.075 ;
        RECT 72.140 139.030 72.460 139.090 ;
        RECT 66.175 138.890 68.690 139.030 ;
        RECT 66.175 138.845 66.465 138.890 ;
        RECT 62.955 138.505 63.245 138.735 ;
        RECT 64.320 138.690 64.640 138.750 ;
        RECT 68.550 138.735 68.690 138.890 ;
        RECT 69.855 138.890 72.460 139.030 ;
        RECT 69.855 138.845 70.145 138.890 ;
        RECT 72.140 138.830 72.460 138.890 ;
        RECT 67.095 138.690 67.385 138.735 ;
        RECT 64.320 138.550 67.385 138.690 ;
        RECT 64.320 138.490 64.640 138.550 ;
        RECT 67.095 138.505 67.385 138.550 ;
        RECT 68.475 138.505 68.765 138.735 ;
        RECT 69.380 138.490 69.700 138.750 ;
        RECT 70.315 138.505 70.605 138.735 ;
        RECT 49.690 138.350 49.830 138.490 ;
        RECT 55.580 138.350 55.900 138.410 ;
        RECT 49.690 138.210 55.900 138.350 ;
        RECT 55.580 138.150 55.900 138.210 ;
        RECT 56.500 138.150 56.820 138.410 ;
        RECT 57.880 138.350 58.200 138.410 ;
        RECT 70.390 138.350 70.530 138.505 ;
        RECT 71.680 138.490 72.000 138.750 ;
        RECT 57.880 138.210 70.530 138.350 ;
        RECT 57.880 138.150 58.200 138.210 ;
        RECT 51.900 138.010 52.220 138.070 ;
        RECT 53.295 138.010 53.585 138.055 ;
        RECT 72.690 138.010 72.830 139.185 ;
        RECT 79.960 139.170 80.280 139.230 ;
        RECT 85.955 139.370 86.245 139.415 ;
        RECT 86.400 139.370 86.720 139.430 ;
        RECT 85.955 139.230 86.720 139.370 ;
        RECT 85.955 139.185 86.245 139.230 ;
        RECT 86.400 139.170 86.720 139.230 ;
        RECT 88.255 139.370 88.545 139.415 ;
        RECT 89.160 139.370 89.480 139.430 ;
        RECT 104.815 139.370 105.105 139.415 ;
        RECT 88.255 139.230 89.480 139.370 ;
        RECT 88.255 139.185 88.545 139.230 ;
        RECT 89.160 139.170 89.480 139.230 ;
        RECT 103.050 139.230 105.105 139.370 ;
        RECT 80.050 139.030 80.190 139.170 ;
        RECT 87.780 139.030 88.100 139.090 ;
        RECT 79.590 138.890 80.190 139.030 ;
        RECT 86.490 138.890 88.100 139.030 ;
        RECT 79.040 138.490 79.360 138.750 ;
        RECT 79.590 138.735 79.730 138.890 ;
        RECT 79.515 138.505 79.805 138.735 ;
        RECT 79.975 138.690 80.265 138.735 ;
        RECT 80.420 138.690 80.740 138.750 ;
        RECT 79.975 138.550 80.740 138.690 ;
        RECT 79.975 138.505 80.265 138.550 ;
        RECT 80.420 138.490 80.740 138.550 ;
        RECT 80.895 138.690 81.185 138.735 ;
        RECT 81.340 138.690 81.660 138.750 ;
        RECT 86.490 138.735 86.630 138.890 ;
        RECT 87.780 138.830 88.100 138.890 ;
        RECT 101.595 139.030 101.885 139.075 ;
        RECT 103.050 139.030 103.190 139.230 ;
        RECT 104.815 139.185 105.105 139.230 ;
        RECT 109.400 139.370 109.720 139.430 ;
        RECT 110.335 139.370 110.625 139.415 ;
        RECT 109.400 139.230 110.625 139.370 ;
        RECT 109.400 139.170 109.720 139.230 ;
        RECT 110.335 139.185 110.625 139.230 ;
        RECT 112.160 139.170 112.480 139.430 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 101.595 138.890 103.190 139.030 ;
        RECT 103.880 139.030 104.200 139.090 ;
        RECT 104.355 139.030 104.645 139.075 ;
        RECT 109.875 139.030 110.165 139.075 ;
        RECT 111.240 139.030 111.560 139.090 ;
        RECT 114.705 139.030 114.995 139.075 ;
        RECT 103.880 138.890 104.645 139.030 ;
        RECT 101.595 138.845 101.885 138.890 ;
        RECT 103.880 138.830 104.200 138.890 ;
        RECT 104.355 138.845 104.645 138.890 ;
        RECT 107.190 138.890 114.995 139.030 ;
        RECT 80.895 138.550 81.660 138.690 ;
        RECT 80.895 138.505 81.185 138.550 ;
        RECT 80.970 138.350 81.110 138.505 ;
        RECT 81.340 138.490 81.660 138.550 ;
        RECT 86.415 138.505 86.705 138.735 ;
        RECT 86.860 138.690 87.180 138.750 ;
        RECT 87.335 138.690 87.625 138.735 ;
        RECT 86.860 138.550 87.625 138.690 ;
        RECT 86.860 138.490 87.180 138.550 ;
        RECT 87.335 138.505 87.625 138.550 ;
        RECT 96.060 138.690 96.380 138.750 ;
        RECT 100.215 138.690 100.505 138.735 ;
        RECT 96.060 138.550 100.505 138.690 ;
        RECT 96.060 138.490 96.380 138.550 ;
        RECT 100.215 138.505 100.505 138.550 ;
        RECT 102.960 138.490 103.280 138.750 ;
        RECT 103.420 138.490 103.740 138.750 ;
        RECT 104.800 138.690 105.120 138.750 ;
        RECT 106.195 138.690 106.485 138.735 ;
        RECT 104.800 138.550 106.485 138.690 ;
        RECT 104.800 138.490 105.120 138.550 ;
        RECT 106.195 138.505 106.485 138.550 ;
        RECT 106.640 138.490 106.960 138.750 ;
        RECT 107.190 138.735 107.330 138.890 ;
        RECT 109.875 138.845 110.165 138.890 ;
        RECT 111.240 138.830 111.560 138.890 ;
        RECT 114.705 138.845 114.995 138.890 ;
        RECT 116.710 139.030 117.000 139.075 ;
        RECT 118.140 139.030 118.460 139.090 ;
        RECT 119.970 139.030 120.260 139.075 ;
        RECT 116.710 138.890 120.260 139.030 ;
        RECT 116.710 138.845 117.000 138.890 ;
        RECT 118.140 138.830 118.460 138.890 ;
        RECT 119.970 138.845 120.260 138.890 ;
        RECT 120.890 139.030 121.180 139.075 ;
        RECT 122.750 139.030 123.040 139.075 ;
        RECT 120.890 138.890 123.040 139.030 ;
        RECT 120.890 138.845 121.180 138.890 ;
        RECT 122.750 138.845 123.040 138.890 ;
        RECT 107.115 138.505 107.405 138.735 ;
        RECT 108.035 138.690 108.325 138.735 ;
        RECT 108.480 138.690 108.800 138.750 ;
        RECT 108.035 138.550 108.800 138.690 ;
        RECT 108.035 138.505 108.325 138.550 ;
        RECT 108.480 138.490 108.800 138.550 ;
        RECT 113.095 138.690 113.385 138.735 ;
        RECT 117.680 138.690 118.000 138.750 ;
        RECT 113.095 138.550 118.000 138.690 ;
        RECT 113.095 138.505 113.385 138.550 ;
        RECT 117.680 138.490 118.000 138.550 ;
        RECT 118.570 138.690 118.860 138.735 ;
        RECT 120.890 138.690 121.105 138.845 ;
        RECT 118.570 138.550 121.105 138.690 ;
        RECT 118.570 138.505 118.860 138.550 ;
        RECT 121.820 138.490 122.140 138.750 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 80.510 138.210 81.110 138.350 ;
        RECT 99.280 138.350 99.600 138.410 ;
        RECT 100.675 138.350 100.965 138.395 ;
        RECT 99.280 138.210 100.965 138.350 ;
        RECT 80.510 138.070 80.650 138.210 ;
        RECT 99.280 138.150 99.600 138.210 ;
        RECT 100.675 138.165 100.965 138.210 ;
        RECT 108.940 138.150 109.260 138.410 ;
        RECT 122.280 138.350 122.600 138.410 ;
        RECT 123.675 138.350 123.965 138.395 ;
        RECT 122.280 138.210 123.965 138.350 ;
        RECT 122.280 138.150 122.600 138.210 ;
        RECT 123.675 138.165 123.965 138.210 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 49.230 137.870 50.290 138.010 ;
        RECT 50.150 137.730 50.290 137.870 ;
        RECT 51.900 137.870 53.585 138.010 ;
        RECT 51.900 137.810 52.220 137.870 ;
        RECT 53.295 137.825 53.585 137.870 ;
        RECT 53.830 137.870 72.830 138.010 ;
        RECT 73.060 138.010 73.380 138.070 ;
        RECT 78.580 138.010 78.900 138.070 ;
        RECT 80.420 138.010 80.740 138.070 ;
        RECT 73.060 137.870 80.740 138.010 ;
        RECT 27.520 137.530 32.350 137.670 ;
        RECT 34.895 137.670 35.185 137.715 ;
        RECT 38.100 137.670 38.420 137.730 ;
        RECT 34.895 137.530 38.420 137.670 ;
        RECT 27.520 137.470 27.840 137.530 ;
        RECT 34.895 137.485 35.185 137.530 ;
        RECT 38.100 137.470 38.420 137.530 ;
        RECT 43.160 137.670 43.480 137.730 ;
        RECT 44.095 137.670 44.385 137.715 ;
        RECT 43.160 137.530 44.385 137.670 ;
        RECT 43.160 137.470 43.480 137.530 ;
        RECT 44.095 137.485 44.385 137.530 ;
        RECT 46.395 137.670 46.685 137.715 ;
        RECT 48.680 137.670 49.000 137.730 ;
        RECT 46.395 137.530 49.000 137.670 ;
        RECT 46.395 137.485 46.685 137.530 ;
        RECT 48.680 137.470 49.000 137.530 ;
        RECT 50.060 137.670 50.380 137.730 ;
        RECT 53.830 137.670 53.970 137.870 ;
        RECT 73.060 137.810 73.380 137.870 ;
        RECT 78.580 137.810 78.900 137.870 ;
        RECT 80.420 137.810 80.740 137.870 ;
        RECT 118.570 138.010 118.860 138.055 ;
        RECT 121.350 138.010 121.640 138.055 ;
        RECT 123.210 138.010 123.500 138.055 ;
        RECT 118.570 137.870 123.500 138.010 ;
        RECT 118.570 137.825 118.860 137.870 ;
        RECT 121.350 137.825 121.640 137.870 ;
        RECT 123.210 137.825 123.500 137.870 ;
        RECT 50.060 137.530 53.970 137.670 ;
        RECT 62.495 137.670 62.785 137.715 ;
        RECT 65.240 137.670 65.560 137.730 ;
        RECT 62.495 137.530 65.560 137.670 ;
        RECT 50.060 137.470 50.380 137.530 ;
        RECT 62.495 137.485 62.785 137.530 ;
        RECT 65.240 137.470 65.560 137.530 ;
        RECT 77.675 137.670 77.965 137.715 ;
        RECT 78.120 137.670 78.440 137.730 ;
        RECT 77.675 137.530 78.440 137.670 ;
        RECT 77.675 137.485 77.965 137.530 ;
        RECT 78.120 137.470 78.440 137.530 ;
        RECT 99.295 137.670 99.585 137.715 ;
        RECT 100.200 137.670 100.520 137.730 ;
        RECT 99.295 137.530 100.520 137.670 ;
        RECT 99.295 137.485 99.585 137.530 ;
        RECT 100.200 137.470 100.520 137.530 ;
        RECT 101.580 137.470 101.900 137.730 ;
        RECT 102.055 137.670 102.345 137.715 ;
        RECT 103.880 137.670 104.200 137.730 ;
        RECT 102.055 137.530 104.200 137.670 ;
        RECT 102.055 137.485 102.345 137.530 ;
        RECT 103.880 137.470 104.200 137.530 ;
        RECT 104.340 137.470 104.660 137.730 ;
        RECT 113.555 137.670 113.845 137.715 ;
        RECT 114.000 137.670 114.320 137.730 ;
        RECT 113.555 137.530 114.320 137.670 ;
        RECT 113.555 137.485 113.845 137.530 ;
        RECT 114.000 137.470 114.320 137.530 ;
        RECT 11.810 136.850 125.890 137.330 ;
        RECT 27.520 136.695 27.840 136.710 ;
        RECT 27.520 136.465 28.055 136.695 ;
        RECT 50.520 136.650 50.840 136.710 ;
        RECT 51.440 136.650 51.760 136.710 ;
        RECT 73.060 136.650 73.380 136.710 ;
        RECT 50.520 136.510 73.380 136.650 ;
        RECT 27.520 136.450 27.840 136.465 ;
        RECT 50.520 136.450 50.840 136.510 ;
        RECT 51.440 136.450 51.760 136.510 ;
        RECT 73.060 136.450 73.380 136.510 ;
        RECT 73.520 136.650 73.840 136.710 ;
        RECT 76.755 136.650 77.045 136.695 ;
        RECT 73.520 136.510 77.045 136.650 ;
        RECT 73.520 136.450 73.840 136.510 ;
        RECT 76.755 136.465 77.045 136.510 ;
        RECT 86.415 136.650 86.705 136.695 ;
        RECT 86.860 136.650 87.180 136.710 ;
        RECT 86.415 136.510 87.180 136.650 ;
        RECT 86.415 136.465 86.705 136.510 ;
        RECT 86.860 136.450 87.180 136.510 ;
        RECT 31.630 136.310 31.920 136.355 ;
        RECT 34.410 136.310 34.700 136.355 ;
        RECT 36.270 136.310 36.560 136.355 ;
        RECT 31.630 136.170 36.560 136.310 ;
        RECT 31.630 136.125 31.920 136.170 ;
        RECT 34.410 136.125 34.700 136.170 ;
        RECT 36.270 136.125 36.560 136.170 ;
        RECT 37.195 136.125 37.485 136.355 ;
        RECT 108.940 136.310 109.260 136.370 ;
        RECT 83.270 136.170 93.530 136.310 ;
        RECT 16.480 135.970 16.800 136.030 ;
        RECT 18.795 135.970 19.085 136.015 ;
        RECT 30.740 135.970 31.060 136.030 ;
        RECT 37.270 135.970 37.410 136.125 ;
        RECT 83.270 136.030 83.410 136.170 ;
        RECT 16.480 135.830 31.060 135.970 ;
        RECT 16.480 135.770 16.800 135.830 ;
        RECT 18.795 135.785 19.085 135.830 ;
        RECT 30.740 135.770 31.060 135.830 ;
        RECT 36.350 135.830 37.410 135.970 ;
        RECT 56.040 135.970 56.360 136.030 ;
        RECT 61.575 135.970 61.865 136.015 ;
        RECT 69.380 135.970 69.700 136.030 ;
        RECT 56.040 135.830 69.700 135.970 ;
        RECT 17.400 135.630 17.720 135.690 ;
        RECT 19.255 135.630 19.545 135.675 ;
        RECT 17.400 135.490 19.545 135.630 ;
        RECT 17.400 135.430 17.720 135.490 ;
        RECT 19.255 135.445 19.545 135.490 ;
        RECT 31.630 135.630 31.920 135.675 ;
        RECT 34.895 135.630 35.185 135.675 ;
        RECT 36.350 135.630 36.490 135.830 ;
        RECT 56.040 135.770 56.360 135.830 ;
        RECT 61.575 135.785 61.865 135.830 ;
        RECT 69.380 135.770 69.700 135.830 ;
        RECT 81.800 135.970 82.120 136.030 ;
        RECT 83.180 135.970 83.500 136.030 ;
        RECT 81.800 135.830 83.500 135.970 ;
        RECT 81.800 135.770 82.120 135.830 ;
        RECT 83.180 135.770 83.500 135.830 ;
        RECT 84.115 135.970 84.405 136.015 ;
        RECT 84.560 135.970 84.880 136.030 ;
        RECT 93.390 136.015 93.530 136.170 ;
        RECT 102.590 136.170 109.260 136.310 ;
        RECT 102.590 136.015 102.730 136.170 ;
        RECT 108.940 136.110 109.260 136.170 ;
        RECT 115.810 136.310 116.100 136.355 ;
        RECT 118.590 136.310 118.880 136.355 ;
        RECT 120.450 136.310 120.740 136.355 ;
        RECT 115.810 136.170 120.740 136.310 ;
        RECT 115.810 136.125 116.100 136.170 ;
        RECT 118.590 136.125 118.880 136.170 ;
        RECT 120.450 136.125 120.740 136.170 ;
        RECT 84.115 135.830 84.880 135.970 ;
        RECT 84.115 135.785 84.405 135.830 ;
        RECT 84.560 135.770 84.880 135.830 ;
        RECT 93.315 135.970 93.605 136.015 ;
        RECT 102.515 135.970 102.805 136.015 ;
        RECT 108.020 135.970 108.340 136.030 ;
        RECT 111.945 135.970 112.235 136.015 ;
        RECT 93.315 135.830 102.805 135.970 ;
        RECT 93.315 135.785 93.605 135.830 ;
        RECT 102.515 135.785 102.805 135.830 ;
        RECT 103.970 135.830 112.235 135.970 ;
        RECT 31.630 135.490 34.165 135.630 ;
        RECT 31.630 135.445 31.920 135.490 ;
        RECT 29.770 135.290 30.060 135.335 ;
        RECT 31.200 135.290 31.520 135.350 ;
        RECT 33.950 135.335 34.165 135.490 ;
        RECT 34.895 135.490 36.490 135.630 ;
        RECT 34.895 135.445 35.185 135.490 ;
        RECT 36.735 135.445 37.025 135.675 ;
        RECT 33.030 135.290 33.320 135.335 ;
        RECT 29.770 135.150 33.320 135.290 ;
        RECT 29.770 135.105 30.060 135.150 ;
        RECT 31.200 135.090 31.520 135.150 ;
        RECT 33.030 135.105 33.320 135.150 ;
        RECT 33.950 135.290 34.240 135.335 ;
        RECT 35.810 135.290 36.100 135.335 ;
        RECT 33.950 135.150 36.100 135.290 ;
        RECT 33.950 135.105 34.240 135.150 ;
        RECT 35.810 135.105 36.100 135.150 ;
        RECT 19.700 134.750 20.020 135.010 ;
        RECT 21.555 134.950 21.845 134.995 ;
        RECT 24.300 134.950 24.620 135.010 ;
        RECT 21.555 134.810 24.620 134.950 ;
        RECT 21.555 134.765 21.845 134.810 ;
        RECT 24.300 134.750 24.620 134.810 ;
        RECT 27.980 134.950 28.300 135.010 ;
        RECT 36.810 134.950 36.950 135.445 ;
        RECT 38.100 135.430 38.420 135.690 ;
        RECT 60.180 135.630 60.500 135.690 ;
        RECT 62.940 135.630 63.260 135.690 ;
        RECT 65.715 135.630 66.005 135.675 ;
        RECT 60.180 135.490 63.260 135.630 ;
        RECT 60.180 135.430 60.500 135.490 ;
        RECT 62.940 135.430 63.260 135.490 ;
        RECT 64.870 135.490 66.005 135.630 ;
        RECT 27.980 134.810 36.950 134.950 ;
        RECT 58.800 134.950 59.120 135.010 ;
        RECT 62.480 134.950 62.800 135.010 ;
        RECT 64.870 134.995 65.010 135.490 ;
        RECT 65.715 135.445 66.005 135.490 ;
        RECT 76.740 135.430 77.060 135.690 ;
        RECT 77.215 135.630 77.505 135.675 ;
        RECT 77.660 135.630 77.980 135.690 ;
        RECT 77.215 135.490 77.980 135.630 ;
        RECT 77.215 135.445 77.505 135.490 ;
        RECT 77.660 135.430 77.980 135.490 ;
        RECT 78.120 135.430 78.440 135.690 ;
        RECT 87.780 135.630 88.100 135.690 ;
        RECT 92.840 135.630 93.160 135.690 ;
        RECT 103.970 135.675 104.110 135.830 ;
        RECT 108.020 135.770 108.340 135.830 ;
        RECT 111.945 135.785 112.235 135.830 ;
        RECT 100.675 135.630 100.965 135.675 ;
        RECT 87.780 135.490 100.965 135.630 ;
        RECT 87.780 135.430 88.100 135.490 ;
        RECT 92.840 135.430 93.160 135.490 ;
        RECT 100.675 135.445 100.965 135.490 ;
        RECT 103.895 135.445 104.185 135.675 ;
        RECT 107.115 135.630 107.405 135.675 ;
        RECT 105.810 135.490 107.405 135.630 ;
        RECT 94.695 135.290 94.985 135.335 ;
        RECT 99.280 135.290 99.600 135.350 ;
        RECT 103.435 135.290 103.725 135.335 ;
        RECT 94.695 135.150 103.725 135.290 ;
        RECT 94.695 135.105 94.985 135.150 ;
        RECT 99.280 135.090 99.600 135.150 ;
        RECT 103.435 135.105 103.725 135.150 ;
        RECT 58.800 134.810 62.800 134.950 ;
        RECT 27.980 134.750 28.300 134.810 ;
        RECT 58.800 134.750 59.120 134.810 ;
        RECT 62.480 134.750 62.800 134.810 ;
        RECT 64.795 134.765 65.085 134.995 ;
        RECT 66.635 134.950 66.925 134.995 ;
        RECT 70.300 134.950 70.620 135.010 ;
        RECT 66.635 134.810 70.620 134.950 ;
        RECT 66.635 134.765 66.925 134.810 ;
        RECT 70.300 134.750 70.620 134.810 ;
        RECT 74.440 134.950 74.760 135.010 ;
        RECT 75.835 134.950 76.125 134.995 ;
        RECT 74.440 134.810 76.125 134.950 ;
        RECT 74.440 134.750 74.760 134.810 ;
        RECT 75.835 134.765 76.125 134.810 ;
        RECT 84.100 134.950 84.420 135.010 ;
        RECT 84.575 134.950 84.865 134.995 ;
        RECT 84.100 134.810 84.865 134.950 ;
        RECT 84.100 134.750 84.420 134.810 ;
        RECT 84.575 134.765 84.865 134.810 ;
        RECT 94.220 134.750 94.540 135.010 ;
        RECT 96.060 134.950 96.380 135.010 ;
        RECT 96.535 134.950 96.825 134.995 ;
        RECT 96.060 134.810 96.825 134.950 ;
        RECT 96.060 134.750 96.380 134.810 ;
        RECT 96.535 134.765 96.825 134.810 ;
        RECT 101.120 134.750 101.440 135.010 ;
        RECT 105.810 134.995 105.950 135.490 ;
        RECT 107.115 135.445 107.405 135.490 ;
        RECT 115.810 135.630 116.100 135.675 ;
        RECT 115.810 135.490 118.345 135.630 ;
        RECT 115.810 135.445 116.100 135.490 ;
        RECT 114.000 135.335 114.320 135.350 ;
        RECT 118.130 135.335 118.345 135.490 ;
        RECT 119.060 135.430 119.380 135.690 ;
        RECT 120.915 135.445 121.205 135.675 ;
        RECT 113.950 135.290 114.320 135.335 ;
        RECT 117.210 135.290 117.500 135.335 ;
        RECT 113.950 135.150 117.500 135.290 ;
        RECT 113.950 135.105 114.320 135.150 ;
        RECT 117.210 135.105 117.500 135.150 ;
        RECT 118.130 135.290 118.420 135.335 ;
        RECT 119.990 135.290 120.280 135.335 ;
        RECT 118.130 135.150 120.280 135.290 ;
        RECT 118.130 135.105 118.420 135.150 ;
        RECT 119.990 135.105 120.280 135.150 ;
        RECT 114.000 135.090 114.320 135.105 ;
        RECT 105.735 134.765 106.025 134.995 ;
        RECT 106.180 134.750 106.500 135.010 ;
        RECT 108.020 134.950 108.340 135.010 ;
        RECT 120.990 134.950 121.130 135.445 ;
        RECT 121.820 134.950 122.140 135.010 ;
        RECT 108.020 134.810 122.140 134.950 ;
        RECT 108.020 134.750 108.340 134.810 ;
        RECT 121.820 134.750 122.140 134.810 ;
        RECT 11.010 134.130 125.890 134.610 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 23.395 133.745 23.685 133.975 ;
        RECT 15.970 133.590 16.260 133.635 ;
        RECT 17.400 133.590 17.720 133.650 ;
        RECT 19.230 133.590 19.520 133.635 ;
        RECT 15.970 133.450 19.520 133.590 ;
        RECT 15.970 133.405 16.260 133.450 ;
        RECT 17.400 133.390 17.720 133.450 ;
        RECT 19.230 133.405 19.520 133.450 ;
        RECT 20.150 133.590 20.440 133.635 ;
        RECT 22.010 133.590 22.300 133.635 ;
        RECT 20.150 133.450 22.300 133.590 ;
        RECT 20.150 133.405 20.440 133.450 ;
        RECT 22.010 133.405 22.300 133.450 ;
        RECT 17.830 133.250 18.120 133.295 ;
        RECT 20.150 133.250 20.365 133.405 ;
        RECT 17.830 133.110 20.365 133.250 ;
        RECT 21.095 133.250 21.385 133.295 ;
        RECT 23.470 133.250 23.610 133.745 ;
        RECT 31.200 133.730 31.520 133.990 ;
        RECT 43.160 133.730 43.480 133.990 ;
        RECT 43.635 133.930 43.925 133.975 ;
        RECT 55.135 133.930 55.425 133.975 ;
        RECT 55.580 133.930 55.900 133.990 ;
        RECT 59.720 133.930 60.040 133.990 ;
        RECT 43.635 133.790 54.890 133.930 ;
        RECT 43.635 133.745 43.925 133.790 ;
        RECT 45.935 133.590 46.225 133.635 ;
        RECT 48.235 133.590 48.525 133.635 ;
        RECT 54.750 133.590 54.890 133.790 ;
        RECT 55.135 133.790 55.900 133.930 ;
        RECT 55.135 133.745 55.425 133.790 ;
        RECT 55.580 133.730 55.900 133.790 ;
        RECT 56.130 133.790 60.040 133.930 ;
        RECT 56.130 133.590 56.270 133.790 ;
        RECT 59.720 133.730 60.040 133.790 ;
        RECT 61.805 133.930 62.095 133.975 ;
        RECT 62.480 133.930 62.800 133.990 ;
        RECT 71.220 133.930 71.540 133.990 ;
        RECT 79.960 133.930 80.280 133.990 ;
        RECT 61.805 133.790 62.800 133.930 ;
        RECT 61.805 133.745 62.095 133.790 ;
        RECT 62.480 133.730 62.800 133.790 ;
        RECT 63.030 133.790 71.540 133.930 ;
        RECT 63.030 133.590 63.170 133.790 ;
        RECT 71.220 133.730 71.540 133.790 ;
        RECT 79.590 133.790 80.280 133.930 ;
        RECT 45.935 133.450 48.525 133.590 ;
        RECT 45.935 133.405 46.225 133.450 ;
        RECT 48.235 133.405 48.525 133.450 ;
        RECT 50.610 133.450 52.130 133.590 ;
        RECT 54.750 133.450 56.270 133.590 ;
        RECT 56.590 133.450 63.170 133.590 ;
        RECT 63.810 133.590 64.100 133.635 ;
        RECT 64.780 133.590 65.100 133.650 ;
        RECT 67.070 133.590 67.360 133.635 ;
        RECT 63.810 133.450 67.360 133.590 ;
        RECT 21.095 133.110 23.610 133.250 ;
        RECT 17.830 133.065 18.120 133.110 ;
        RECT 21.095 133.065 21.385 133.110 ;
        RECT 24.300 133.050 24.620 133.310 ;
        RECT 29.375 133.250 29.665 133.295 ;
        RECT 29.820 133.250 30.140 133.310 ;
        RECT 30.755 133.250 31.045 133.295 ;
        RECT 29.375 133.110 31.045 133.250 ;
        RECT 29.375 133.065 29.665 133.110 ;
        RECT 29.820 133.050 30.140 133.110 ;
        RECT 30.755 133.065 31.045 133.110 ;
        RECT 42.255 133.065 42.545 133.295 ;
        RECT 42.700 133.250 43.020 133.310 ;
        RECT 44.555 133.250 44.845 133.295 ;
        RECT 42.700 133.110 44.845 133.250 ;
        RECT 22.935 132.910 23.225 132.955 ;
        RECT 27.980 132.910 28.300 132.970 ;
        RECT 22.935 132.770 28.300 132.910 ;
        RECT 22.935 132.725 23.225 132.770 ;
        RECT 27.980 132.710 28.300 132.770 ;
        RECT 41.335 132.725 41.625 132.955 ;
        RECT 42.330 132.910 42.470 133.065 ;
        RECT 42.700 133.050 43.020 133.110 ;
        RECT 44.555 133.065 44.845 133.110 ;
        RECT 49.615 133.065 49.905 133.295 ;
        RECT 43.160 132.910 43.480 132.970 ;
        RECT 42.330 132.770 43.480 132.910 ;
        RECT 17.830 132.570 18.120 132.615 ;
        RECT 20.610 132.570 20.900 132.615 ;
        RECT 22.470 132.570 22.760 132.615 ;
        RECT 41.410 132.570 41.550 132.725 ;
        RECT 43.160 132.710 43.480 132.770 ;
        RECT 45.460 132.710 45.780 132.970 ;
        RECT 45.920 132.910 46.240 132.970 ;
        RECT 48.220 132.910 48.540 132.970 ;
        RECT 49.690 132.910 49.830 133.065 ;
        RECT 50.060 133.050 50.380 133.310 ;
        RECT 50.610 133.295 50.750 133.450 ;
        RECT 50.535 133.065 50.825 133.295 ;
        RECT 51.440 133.050 51.760 133.310 ;
        RECT 51.990 133.250 52.130 133.450 ;
        RECT 51.990 133.110 54.890 133.250 ;
        RECT 45.920 132.770 49.830 132.910 ;
        RECT 45.920 132.710 46.240 132.770 ;
        RECT 48.220 132.710 48.540 132.770 ;
        RECT 54.200 132.710 54.520 132.970 ;
        RECT 54.750 132.955 54.890 133.110 ;
        RECT 54.675 132.910 54.965 132.955 ;
        RECT 55.580 132.910 55.900 132.970 ;
        RECT 54.675 132.770 55.900 132.910 ;
        RECT 54.675 132.725 54.965 132.770 ;
        RECT 55.580 132.710 55.900 132.770 ;
        RECT 17.830 132.430 22.760 132.570 ;
        RECT 17.830 132.385 18.120 132.430 ;
        RECT 20.610 132.385 20.900 132.430 ;
        RECT 22.470 132.385 22.760 132.430 ;
        RECT 23.010 132.430 41.550 132.570 ;
        RECT 41.780 132.570 42.100 132.630 ;
        RECT 56.590 132.570 56.730 133.450 ;
        RECT 63.810 133.405 64.100 133.450 ;
        RECT 64.780 133.390 65.100 133.450 ;
        RECT 67.070 133.405 67.360 133.450 ;
        RECT 67.990 133.590 68.280 133.635 ;
        RECT 69.850 133.590 70.140 133.635 ;
        RECT 67.990 133.450 70.140 133.590 ;
        RECT 67.990 133.405 68.280 133.450 ;
        RECT 69.850 133.405 70.140 133.450 ;
        RECT 57.895 133.250 58.185 133.295 ;
        RECT 57.050 133.110 58.185 133.250 ;
        RECT 57.050 132.615 57.190 133.110 ;
        RECT 57.895 133.065 58.185 133.110 ;
        RECT 65.670 133.250 65.960 133.295 ;
        RECT 67.990 133.250 68.205 133.405 ;
        RECT 65.670 133.110 68.205 133.250 ;
        RECT 68.935 133.250 69.225 133.295 ;
        RECT 70.300 133.250 70.620 133.310 ;
        RECT 68.935 133.110 70.620 133.250 ;
        RECT 65.670 133.065 65.960 133.110 ;
        RECT 68.935 133.065 69.225 133.110 ;
        RECT 70.300 133.050 70.620 133.110 ;
        RECT 70.760 133.050 71.080 133.310 ;
        RECT 79.040 133.050 79.360 133.310 ;
        RECT 79.590 133.295 79.730 133.790 ;
        RECT 79.960 133.730 80.280 133.790 ;
        RECT 86.415 133.745 86.705 133.975 ;
        RECT 98.605 133.930 98.895 133.975 ;
        RECT 99.280 133.930 99.600 133.990 ;
        RECT 98.605 133.790 99.600 133.930 ;
        RECT 98.605 133.745 98.895 133.790 ;
        RECT 84.100 133.590 84.420 133.650 ;
        RECT 80.050 133.450 84.420 133.590 ;
        RECT 80.050 133.295 80.190 133.450 ;
        RECT 84.100 133.390 84.420 133.450 ;
        RECT 79.515 133.065 79.805 133.295 ;
        RECT 79.975 133.065 80.265 133.295 ;
        RECT 80.420 133.250 80.740 133.310 ;
        RECT 80.895 133.250 81.185 133.295 ;
        RECT 80.420 133.110 81.185 133.250 ;
        RECT 80.420 133.050 80.740 133.110 ;
        RECT 80.895 133.065 81.185 133.110 ;
        RECT 81.340 133.250 81.660 133.310 ;
        RECT 84.575 133.250 84.865 133.295 ;
        RECT 81.340 133.110 84.865 133.250 ;
        RECT 86.490 133.250 86.630 133.745 ;
        RECT 99.280 133.730 99.600 133.790 ;
        RECT 105.260 133.930 105.580 133.990 ;
        RECT 108.035 133.930 108.325 133.975 ;
        RECT 105.260 133.790 108.325 133.930 ;
        RECT 105.260 133.730 105.580 133.790 ;
        RECT 108.035 133.745 108.325 133.790 ;
        RECT 118.155 133.930 118.445 133.975 ;
        RECT 119.060 133.930 119.380 133.990 ;
        RECT 118.155 133.790 119.380 133.930 ;
        RECT 118.155 133.745 118.445 133.790 ;
        RECT 119.060 133.730 119.380 133.790 ;
        RECT 90.950 133.590 91.240 133.635 ;
        RECT 93.300 133.590 93.620 133.650 ;
        RECT 94.210 133.590 94.500 133.635 ;
        RECT 90.950 133.450 94.500 133.590 ;
        RECT 90.950 133.405 91.240 133.450 ;
        RECT 93.300 133.390 93.620 133.450 ;
        RECT 94.210 133.405 94.500 133.450 ;
        RECT 95.130 133.590 95.420 133.635 ;
        RECT 96.990 133.590 97.280 133.635 ;
        RECT 95.130 133.450 97.280 133.590 ;
        RECT 95.130 133.405 95.420 133.450 ;
        RECT 96.990 133.405 97.280 133.450 ;
        RECT 100.610 133.590 100.900 133.635 ;
        RECT 101.120 133.590 101.440 133.650 ;
        RECT 103.870 133.590 104.160 133.635 ;
        RECT 100.610 133.450 104.160 133.590 ;
        RECT 100.610 133.405 100.900 133.450 ;
        RECT 87.335 133.250 87.625 133.295 ;
        RECT 86.490 133.110 87.625 133.250 ;
        RECT 61.100 132.910 61.420 132.970 ;
        RECT 70.850 132.910 70.990 133.050 ;
        RECT 61.100 132.770 70.990 132.910 ;
        RECT 80.970 132.910 81.110 133.065 ;
        RECT 81.340 133.050 81.660 133.110 ;
        RECT 84.575 133.065 84.865 133.110 ;
        RECT 87.335 133.065 87.625 133.110 ;
        RECT 92.810 133.250 93.100 133.295 ;
        RECT 95.130 133.250 95.345 133.405 ;
        RECT 101.120 133.390 101.440 133.450 ;
        RECT 103.870 133.405 104.160 133.450 ;
        RECT 104.790 133.590 105.080 133.635 ;
        RECT 106.650 133.590 106.940 133.635 ;
        RECT 104.790 133.450 106.940 133.590 ;
        RECT 104.790 133.405 105.080 133.450 ;
        RECT 106.650 133.405 106.940 133.450 ;
        RECT 92.810 133.110 95.345 133.250 ;
        RECT 95.600 133.250 95.920 133.310 ;
        RECT 96.075 133.250 96.365 133.295 ;
        RECT 95.600 133.110 96.365 133.250 ;
        RECT 92.810 133.065 93.100 133.110 ;
        RECT 81.800 132.910 82.120 132.970 ;
        RECT 80.970 132.770 82.120 132.910 ;
        RECT 61.100 132.710 61.420 132.770 ;
        RECT 81.800 132.710 82.120 132.770 ;
        RECT 83.180 132.710 83.500 132.970 ;
        RECT 84.100 132.710 84.420 132.970 ;
        RECT 84.650 132.910 84.790 133.065 ;
        RECT 95.600 133.050 95.920 133.110 ;
        RECT 96.075 133.065 96.365 133.110 ;
        RECT 97.915 133.250 98.205 133.295 ;
        RECT 98.360 133.250 98.680 133.310 ;
        RECT 97.915 133.110 98.680 133.250 ;
        RECT 97.915 133.065 98.205 133.110 ;
        RECT 98.360 133.050 98.680 133.110 ;
        RECT 102.470 133.250 102.760 133.295 ;
        RECT 104.790 133.250 105.005 133.405 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 102.470 133.110 105.005 133.250 ;
        RECT 105.735 133.250 106.025 133.295 ;
        RECT 106.180 133.250 106.500 133.310 ;
        RECT 105.735 133.110 106.500 133.250 ;
        RECT 102.470 133.065 102.760 133.110 ;
        RECT 105.735 133.065 106.025 133.110 ;
        RECT 106.180 133.050 106.500 133.110 ;
        RECT 107.100 133.250 107.420 133.310 ;
        RECT 108.955 133.250 109.245 133.295 ;
        RECT 107.100 133.110 109.245 133.250 ;
        RECT 107.100 133.050 107.420 133.110 ;
        RECT 108.955 133.065 109.245 133.110 ;
        RECT 113.080 133.250 113.400 133.310 ;
        RECT 117.235 133.250 117.525 133.295 ;
        RECT 113.080 133.110 117.525 133.250 ;
        RECT 113.080 133.050 113.400 133.110 ;
        RECT 117.235 133.065 117.525 133.110 ;
        RECT 88.945 132.910 89.235 132.955 ;
        RECT 94.220 132.910 94.540 132.970 ;
        RECT 84.650 132.770 94.540 132.910 ;
        RECT 98.450 132.910 98.590 133.050 ;
        RECT 107.575 132.910 107.865 132.955 ;
        RECT 108.020 132.910 108.340 132.970 ;
        RECT 98.450 132.770 108.340 132.910 ;
        RECT 88.945 132.725 89.235 132.770 ;
        RECT 94.220 132.710 94.540 132.770 ;
        RECT 107.575 132.725 107.865 132.770 ;
        RECT 108.020 132.710 108.340 132.770 ;
        RECT 109.875 132.910 110.165 132.955 ;
        RECT 110.320 132.910 110.640 132.970 ;
        RECT 109.875 132.770 110.640 132.910 ;
        RECT 109.875 132.725 110.165 132.770 ;
        RECT 110.320 132.710 110.640 132.770 ;
        RECT 41.780 132.430 56.730 132.570 ;
        RECT 13.965 132.230 14.255 132.275 ;
        RECT 19.700 132.230 20.020 132.290 ;
        RECT 23.010 132.230 23.150 132.430 ;
        RECT 41.780 132.370 42.100 132.430 ;
        RECT 56.975 132.385 57.265 132.615 ;
        RECT 65.670 132.570 65.960 132.615 ;
        RECT 68.450 132.570 68.740 132.615 ;
        RECT 70.310 132.570 70.600 132.615 ;
        RECT 65.670 132.430 70.600 132.570 ;
        RECT 65.670 132.385 65.960 132.430 ;
        RECT 68.450 132.385 68.740 132.430 ;
        RECT 70.310 132.385 70.600 132.430 ;
        RECT 92.810 132.570 93.100 132.615 ;
        RECT 95.590 132.570 95.880 132.615 ;
        RECT 97.450 132.570 97.740 132.615 ;
        RECT 92.810 132.430 97.740 132.570 ;
        RECT 92.810 132.385 93.100 132.430 ;
        RECT 95.590 132.385 95.880 132.430 ;
        RECT 97.450 132.385 97.740 132.430 ;
        RECT 102.470 132.570 102.760 132.615 ;
        RECT 105.250 132.570 105.540 132.615 ;
        RECT 107.110 132.570 107.400 132.615 ;
        RECT 102.470 132.430 107.400 132.570 ;
        RECT 102.470 132.385 102.760 132.430 ;
        RECT 105.250 132.385 105.540 132.430 ;
        RECT 107.110 132.385 107.400 132.430 ;
        RECT 13.965 132.090 23.150 132.230 ;
        RECT 29.835 132.230 30.125 132.275 ;
        RECT 30.280 132.230 30.600 132.290 ;
        RECT 29.835 132.090 30.600 132.230 ;
        RECT 13.965 132.045 14.255 132.090 ;
        RECT 19.700 132.030 20.020 132.090 ;
        RECT 29.835 132.045 30.125 132.090 ;
        RECT 30.280 132.030 30.600 132.090 ;
        RECT 41.320 132.230 41.640 132.290 ;
        RECT 44.555 132.230 44.845 132.275 ;
        RECT 41.320 132.090 44.845 132.230 ;
        RECT 41.320 132.030 41.640 132.090 ;
        RECT 44.555 132.045 44.845 132.090 ;
        RECT 54.200 132.230 54.520 132.290 ;
        RECT 56.040 132.230 56.360 132.290 ;
        RECT 54.200 132.090 56.360 132.230 ;
        RECT 54.200 132.030 54.520 132.090 ;
        RECT 56.040 132.030 56.360 132.090 ;
        RECT 58.815 132.230 59.105 132.275 ;
        RECT 59.260 132.230 59.580 132.290 ;
        RECT 58.815 132.090 59.580 132.230 ;
        RECT 58.815 132.045 59.105 132.090 ;
        RECT 59.260 132.030 59.580 132.090 ;
        RECT 75.820 132.230 76.140 132.290 ;
        RECT 77.675 132.230 77.965 132.275 ;
        RECT 75.820 132.090 77.965 132.230 ;
        RECT 75.820 132.030 76.140 132.090 ;
        RECT 77.675 132.045 77.965 132.090 ;
        RECT 88.240 132.030 88.560 132.290 ;
        RECT 11.810 131.410 125.890 131.890 ;
        RECT 17.400 131.010 17.720 131.270 ;
        RECT 31.200 131.210 31.520 131.270 ;
        RECT 32.580 131.210 32.900 131.270 ;
        RECT 35.585 131.210 35.875 131.255 ;
        RECT 19.330 131.070 32.350 131.210 ;
        RECT 19.330 130.575 19.470 131.070 ;
        RECT 31.200 131.010 31.520 131.070 ;
        RECT 27.080 130.870 27.370 130.915 ;
        RECT 28.940 130.870 29.230 130.915 ;
        RECT 31.720 130.870 32.010 130.915 ;
        RECT 27.080 130.730 32.010 130.870 ;
        RECT 32.210 130.870 32.350 131.070 ;
        RECT 32.580 131.070 35.875 131.210 ;
        RECT 32.580 131.010 32.900 131.070 ;
        RECT 35.585 131.025 35.875 131.070 ;
        RECT 41.320 131.010 41.640 131.270 ;
        RECT 41.795 131.025 42.085 131.255 ;
        RECT 43.160 131.210 43.480 131.270 ;
        RECT 43.160 131.070 61.330 131.210 ;
        RECT 37.195 130.870 37.485 130.915 ;
        RECT 41.870 130.870 42.010 131.025 ;
        RECT 43.160 131.010 43.480 131.070 ;
        RECT 43.250 130.870 43.390 131.010 ;
        RECT 32.210 130.730 37.485 130.870 ;
        RECT 27.080 130.685 27.370 130.730 ;
        RECT 28.940 130.685 29.230 130.730 ;
        RECT 31.720 130.685 32.010 130.730 ;
        RECT 37.195 130.685 37.485 130.730 ;
        RECT 38.650 130.730 42.010 130.870 ;
        RECT 42.790 130.730 43.390 130.870 ;
        RECT 56.010 130.870 56.300 130.915 ;
        RECT 58.790 130.870 59.080 130.915 ;
        RECT 60.650 130.870 60.940 130.915 ;
        RECT 56.010 130.730 60.940 130.870 ;
        RECT 61.190 130.870 61.330 131.070 ;
        RECT 64.780 131.010 65.100 131.270 ;
        RECT 70.775 131.210 71.065 131.255 ;
        RECT 71.220 131.210 71.540 131.270 ;
        RECT 66.480 131.070 70.530 131.210 ;
        RECT 66.480 130.870 66.620 131.070 ;
        RECT 61.190 130.730 66.620 130.870 ;
        RECT 19.255 130.345 19.545 130.575 ;
        RECT 19.700 130.330 20.020 130.590 ;
        RECT 30.740 130.530 31.060 130.590 ;
        RECT 38.650 130.530 38.790 130.730 ;
        RECT 42.255 130.530 42.545 130.575 ;
        RECT 30.740 130.390 38.790 130.530 ;
        RECT 39.110 130.390 42.545 130.530 ;
        RECT 30.740 130.330 31.060 130.390 ;
        RECT 15.100 130.190 15.420 130.250 ;
        RECT 16.940 130.190 17.260 130.250 ;
        RECT 15.100 130.050 17.260 130.190 ;
        RECT 15.100 129.990 15.420 130.050 ;
        RECT 16.940 129.990 17.260 130.050 ;
        RECT 26.615 130.190 26.905 130.235 ;
        RECT 27.980 130.190 28.300 130.250 ;
        RECT 26.615 130.050 28.300 130.190 ;
        RECT 26.615 130.005 26.905 130.050 ;
        RECT 27.980 129.990 28.300 130.050 ;
        RECT 28.440 129.990 28.760 130.250 ;
        RECT 31.720 130.190 32.010 130.235 ;
        RECT 29.475 130.050 32.010 130.190 ;
        RECT 20.160 129.850 20.480 129.910 ;
        RECT 29.475 129.895 29.690 130.050 ;
        RECT 31.720 130.005 32.010 130.050 ;
        RECT 34.420 130.190 34.740 130.250 ;
        RECT 39.110 130.190 39.250 130.390 ;
        RECT 42.255 130.345 42.545 130.390 ;
        RECT 34.420 130.050 39.250 130.190 ;
        RECT 34.420 129.990 34.740 130.050 ;
        RECT 39.495 130.005 39.785 130.235 ;
        RECT 40.415 130.190 40.705 130.235 ;
        RECT 42.790 130.190 42.930 130.730 ;
        RECT 56.010 130.685 56.300 130.730 ;
        RECT 58.790 130.685 59.080 130.730 ;
        RECT 60.650 130.685 60.940 130.730 ;
        RECT 47.300 130.530 47.620 130.590 ;
        RECT 43.250 130.390 47.620 130.530 ;
        RECT 43.250 130.235 43.390 130.390 ;
        RECT 47.300 130.330 47.620 130.390 ;
        RECT 59.260 130.330 59.580 130.590 ;
        RECT 66.480 130.530 66.620 130.730 ;
        RECT 67.555 130.870 67.845 130.915 ;
        RECT 70.390 130.870 70.530 131.070 ;
        RECT 70.775 131.070 71.540 131.210 ;
        RECT 70.775 131.025 71.065 131.070 ;
        RECT 71.220 131.010 71.540 131.070 ;
        RECT 73.520 131.010 73.840 131.270 ;
        RECT 76.280 131.010 76.600 131.270 ;
        RECT 83.425 131.210 83.715 131.255 ;
        RECT 84.100 131.210 84.420 131.270 ;
        RECT 83.425 131.070 84.420 131.210 ;
        RECT 83.425 131.025 83.715 131.070 ;
        RECT 84.100 131.010 84.420 131.070 ;
        RECT 93.300 131.010 93.620 131.270 ;
        RECT 95.600 131.010 95.920 131.270 ;
        RECT 98.820 131.210 99.140 131.270 ;
        RECT 100.675 131.210 100.965 131.255 ;
        RECT 98.820 131.070 100.965 131.210 ;
        RECT 98.820 131.010 99.140 131.070 ;
        RECT 100.675 131.025 100.965 131.070 ;
        RECT 101.580 131.210 101.900 131.270 ;
        RECT 106.655 131.210 106.945 131.255 ;
        RECT 101.580 131.070 106.945 131.210 ;
        RECT 101.580 131.010 101.900 131.070 ;
        RECT 106.655 131.025 106.945 131.070 ;
        RECT 107.560 131.210 107.880 131.270 ;
        RECT 108.955 131.210 109.245 131.255 ;
        RECT 107.560 131.070 109.245 131.210 ;
        RECT 107.560 131.010 107.880 131.070 ;
        RECT 108.955 131.025 109.245 131.070 ;
        RECT 78.135 130.870 78.425 130.915 ;
        RECT 85.020 130.870 85.340 130.930 ;
        RECT 67.555 130.730 69.150 130.870 ;
        RECT 70.390 130.730 72.830 130.870 ;
        RECT 67.555 130.685 67.845 130.730 ;
        RECT 68.015 130.530 68.305 130.575 ;
        RECT 66.480 130.390 68.305 130.530 ;
        RECT 68.015 130.345 68.305 130.390 ;
        RECT 40.415 130.050 42.930 130.190 ;
        RECT 40.415 130.005 40.705 130.050 ;
        RECT 43.175 130.005 43.465 130.235 ;
        RECT 27.540 129.850 27.830 129.895 ;
        RECT 29.400 129.850 29.690 129.895 ;
        RECT 20.160 129.710 25.450 129.850 ;
        RECT 20.160 129.650 20.480 129.710 ;
        RECT 22.015 129.510 22.305 129.555 ;
        RECT 24.760 129.510 25.080 129.570 ;
        RECT 22.015 129.370 25.080 129.510 ;
        RECT 25.310 129.510 25.450 129.710 ;
        RECT 27.540 129.710 29.690 129.850 ;
        RECT 27.540 129.665 27.830 129.710 ;
        RECT 29.400 129.665 29.690 129.710 ;
        RECT 30.280 129.895 30.600 129.910 ;
        RECT 30.280 129.850 30.610 129.895 ;
        RECT 33.580 129.850 33.870 129.895 ;
        RECT 30.280 129.710 33.870 129.850 ;
        RECT 30.280 129.665 30.610 129.710 ;
        RECT 33.580 129.665 33.870 129.710 ;
        RECT 38.100 129.850 38.420 129.910 ;
        RECT 38.575 129.850 38.865 129.895 ;
        RECT 38.100 129.710 38.865 129.850 ;
        RECT 30.280 129.650 30.600 129.665 ;
        RECT 38.100 129.650 38.420 129.710 ;
        RECT 38.575 129.665 38.865 129.710 ;
        RECT 39.570 129.510 39.710 130.005 ;
        RECT 45.920 129.990 46.240 130.250 ;
        RECT 46.395 130.005 46.685 130.235 ;
        RECT 41.780 129.650 42.100 129.910 ;
        RECT 46.470 129.850 46.610 130.005 ;
        RECT 46.840 129.990 47.160 130.250 ;
        RECT 47.760 130.190 48.080 130.250 ;
        RECT 51.440 130.190 51.760 130.250 ;
        RECT 52.360 130.190 52.680 130.250 ;
        RECT 47.760 130.050 52.680 130.190 ;
        RECT 47.760 129.990 48.080 130.050 ;
        RECT 51.440 129.990 51.760 130.050 ;
        RECT 52.360 129.990 52.680 130.050 ;
        RECT 56.010 130.190 56.300 130.235 ;
        RECT 56.010 130.050 58.545 130.190 ;
        RECT 56.010 130.005 56.300 130.050 ;
        RECT 50.060 129.850 50.380 129.910 ;
        RECT 46.470 129.710 50.380 129.850 ;
        RECT 50.060 129.650 50.380 129.710 ;
        RECT 54.150 129.850 54.440 129.895 ;
        RECT 55.120 129.850 55.440 129.910 ;
        RECT 58.330 129.895 58.545 130.050 ;
        RECT 61.100 129.990 61.420 130.250 ;
        RECT 64.320 129.990 64.640 130.250 ;
        RECT 65.240 130.190 65.560 130.250 ;
        RECT 69.010 130.235 69.150 130.730 ;
        RECT 66.635 130.190 66.925 130.235 ;
        RECT 65.240 130.050 66.925 130.190 ;
        RECT 65.240 129.990 65.560 130.050 ;
        RECT 66.635 130.005 66.925 130.050 ;
        RECT 68.935 130.190 69.225 130.235 ;
        RECT 71.220 130.190 71.540 130.250 ;
        RECT 72.690 130.235 72.830 130.730 ;
        RECT 78.135 130.730 85.340 130.870 ;
        RECT 78.135 130.685 78.425 130.730 ;
        RECT 85.020 130.670 85.340 130.730 ;
        RECT 87.290 130.870 87.580 130.915 ;
        RECT 90.070 130.870 90.360 130.915 ;
        RECT 91.930 130.870 92.220 130.915 ;
        RECT 87.290 130.730 92.220 130.870 ;
        RECT 87.290 130.685 87.580 130.730 ;
        RECT 90.070 130.685 90.360 130.730 ;
        RECT 91.930 130.685 92.220 130.730 ;
        RECT 76.740 130.330 77.060 130.590 ;
        RECT 88.240 130.530 88.560 130.590 ;
        RECT 90.555 130.530 90.845 130.575 ;
        RECT 88.240 130.390 90.845 130.530 ;
        RECT 88.240 130.330 88.560 130.390 ;
        RECT 90.555 130.345 90.845 130.390 ;
        RECT 107.650 130.390 110.090 130.530 ;
        RECT 68.935 130.050 71.540 130.190 ;
        RECT 68.935 130.005 69.225 130.050 ;
        RECT 57.410 129.850 57.700 129.895 ;
        RECT 54.150 129.710 57.700 129.850 ;
        RECT 54.150 129.665 54.440 129.710 ;
        RECT 55.120 129.650 55.440 129.710 ;
        RECT 57.410 129.665 57.700 129.710 ;
        RECT 58.330 129.850 58.620 129.895 ;
        RECT 60.190 129.850 60.480 129.895 ;
        RECT 58.330 129.710 60.480 129.850 ;
        RECT 66.710 129.850 66.850 130.005 ;
        RECT 71.220 129.990 71.540 130.050 ;
        RECT 72.155 130.005 72.445 130.235 ;
        RECT 72.615 130.190 72.905 130.235 ;
        RECT 75.360 130.190 75.680 130.250 ;
        RECT 72.615 130.050 75.680 130.190 ;
        RECT 72.615 130.005 72.905 130.050 ;
        RECT 70.315 129.850 70.605 129.895 ;
        RECT 66.710 129.710 70.605 129.850 ;
        RECT 72.230 129.850 72.370 130.005 ;
        RECT 75.360 129.990 75.680 130.050 ;
        RECT 75.820 129.990 76.140 130.250 ;
        RECT 77.200 129.990 77.520 130.250 ;
        RECT 79.040 130.190 79.360 130.250 ;
        RECT 79.975 130.190 80.265 130.235 ;
        RECT 79.040 130.050 80.265 130.190 ;
        RECT 79.040 129.990 79.360 130.050 ;
        RECT 79.975 130.005 80.265 130.050 ;
        RECT 80.420 129.990 80.740 130.250 ;
        RECT 80.895 130.190 81.185 130.235 ;
        RECT 81.340 130.190 81.660 130.250 ;
        RECT 80.895 130.050 81.660 130.190 ;
        RECT 80.895 130.005 81.185 130.050 ;
        RECT 81.340 129.990 81.660 130.050 ;
        RECT 81.800 129.990 82.120 130.250 ;
        RECT 87.290 130.190 87.580 130.235 ;
        RECT 91.920 130.190 92.240 130.250 ;
        RECT 92.395 130.190 92.685 130.235 ;
        RECT 87.290 130.050 89.825 130.190 ;
        RECT 87.290 130.005 87.580 130.050 ;
        RECT 73.520 129.850 73.840 129.910 ;
        RECT 72.230 129.710 73.840 129.850 ;
        RECT 58.330 129.665 58.620 129.710 ;
        RECT 60.190 129.665 60.480 129.710 ;
        RECT 70.315 129.665 70.605 129.710 ;
        RECT 73.520 129.650 73.840 129.710 ;
        RECT 85.430 129.850 85.720 129.895 ;
        RECT 86.860 129.850 87.180 129.910 ;
        RECT 89.610 129.895 89.825 130.050 ;
        RECT 91.920 130.050 92.685 130.190 ;
        RECT 91.920 129.990 92.240 130.050 ;
        RECT 92.395 130.005 92.685 130.050 ;
        RECT 92.840 130.190 93.160 130.250 ;
        RECT 93.775 130.190 94.065 130.235 ;
        RECT 94.680 130.190 95.000 130.250 ;
        RECT 92.840 130.050 95.000 130.190 ;
        RECT 92.840 129.990 93.160 130.050 ;
        RECT 93.775 130.005 94.065 130.050 ;
        RECT 94.680 129.990 95.000 130.050 ;
        RECT 96.060 130.190 96.380 130.250 ;
        RECT 96.535 130.190 96.825 130.235 ;
        RECT 96.060 130.050 96.825 130.190 ;
        RECT 96.060 129.990 96.380 130.050 ;
        RECT 96.535 130.005 96.825 130.050 ;
        RECT 101.580 129.990 101.900 130.250 ;
        RECT 102.040 129.990 102.360 130.250 ;
        RECT 106.640 130.190 106.960 130.250 ;
        RECT 107.650 130.235 107.790 130.390 ;
        RECT 107.575 130.190 107.865 130.235 ;
        RECT 106.640 130.050 107.865 130.190 ;
        RECT 106.640 129.990 106.960 130.050 ;
        RECT 107.575 130.005 107.865 130.050 ;
        RECT 108.480 129.990 108.800 130.250 ;
        RECT 109.950 130.235 110.090 130.390 ;
        RECT 109.875 130.005 110.165 130.235 ;
        RECT 110.320 129.990 110.640 130.250 ;
        RECT 88.690 129.850 88.980 129.895 ;
        RECT 85.430 129.710 88.980 129.850 ;
        RECT 85.430 129.665 85.720 129.710 ;
        RECT 86.860 129.650 87.180 129.710 ;
        RECT 88.690 129.665 88.980 129.710 ;
        RECT 89.610 129.850 89.900 129.895 ;
        RECT 91.470 129.850 91.760 129.895 ;
        RECT 89.610 129.710 91.760 129.850 ;
        RECT 89.610 129.665 89.900 129.710 ;
        RECT 91.470 129.665 91.760 129.710 ;
        RECT 104.815 129.850 105.105 129.895 ;
        RECT 108.020 129.850 108.340 129.910 ;
        RECT 104.815 129.710 108.340 129.850 ;
        RECT 104.815 129.665 105.105 129.710 ;
        RECT 108.020 129.650 108.340 129.710 ;
        RECT 25.310 129.370 39.710 129.510 ;
        RECT 42.240 129.510 42.560 129.570 ;
        RECT 44.095 129.510 44.385 129.555 ;
        RECT 42.240 129.370 44.385 129.510 ;
        RECT 22.015 129.325 22.305 129.370 ;
        RECT 24.760 129.310 25.080 129.370 ;
        RECT 42.240 129.310 42.560 129.370 ;
        RECT 44.095 129.325 44.385 129.370 ;
        RECT 44.540 129.310 44.860 129.570 ;
        RECT 52.145 129.510 52.435 129.555 ;
        RECT 55.580 129.510 55.900 129.570 ;
        RECT 57.880 129.510 58.200 129.570 ;
        RECT 52.145 129.370 58.200 129.510 ;
        RECT 52.145 129.325 52.435 129.370 ;
        RECT 55.580 129.310 55.900 129.370 ;
        RECT 57.880 129.310 58.200 129.370 ;
        RECT 78.595 129.510 78.885 129.555 ;
        RECT 79.040 129.510 79.360 129.570 ;
        RECT 78.595 129.370 79.360 129.510 ;
        RECT 78.595 129.325 78.885 129.370 ;
        RECT 79.040 129.310 79.360 129.370 ;
        RECT 11.010 128.690 125.890 129.170 ;
        RECT 14.425 128.490 14.715 128.535 ;
        RECT 20.160 128.490 20.480 128.550 ;
        RECT 14.425 128.350 20.480 128.490 ;
        RECT 14.425 128.305 14.715 128.350 ;
        RECT 20.160 128.290 20.480 128.350 ;
        RECT 23.855 128.305 24.145 128.535 ;
        RECT 27.075 128.490 27.365 128.535 ;
        RECT 28.440 128.490 28.760 128.550 ;
        RECT 27.075 128.350 28.760 128.490 ;
        RECT 27.075 128.305 27.365 128.350 ;
        RECT 16.430 128.150 16.720 128.195 ;
        RECT 17.400 128.150 17.720 128.210 ;
        RECT 19.690 128.150 19.980 128.195 ;
        RECT 16.430 128.010 19.980 128.150 ;
        RECT 16.430 127.965 16.720 128.010 ;
        RECT 17.400 127.950 17.720 128.010 ;
        RECT 19.690 127.965 19.980 128.010 ;
        RECT 20.610 128.150 20.900 128.195 ;
        RECT 22.470 128.150 22.760 128.195 ;
        RECT 20.610 128.010 22.760 128.150 ;
        RECT 20.610 127.965 20.900 128.010 ;
        RECT 22.470 127.965 22.760 128.010 ;
        RECT 18.290 127.810 18.580 127.855 ;
        RECT 20.610 127.810 20.825 127.965 ;
        RECT 18.290 127.670 20.825 127.810 ;
        RECT 21.555 127.810 21.845 127.855 ;
        RECT 23.930 127.810 24.070 128.305 ;
        RECT 28.440 128.290 28.760 128.350 ;
        RECT 29.835 128.305 30.125 128.535 ;
        RECT 31.675 128.490 31.965 128.535 ;
        RECT 32.580 128.490 32.900 128.550 ;
        RECT 31.675 128.350 32.900 128.490 ;
        RECT 31.675 128.305 31.965 128.350 ;
        RECT 29.910 128.150 30.050 128.305 ;
        RECT 32.580 128.290 32.900 128.350 ;
        RECT 39.955 128.490 40.245 128.535 ;
        RECT 41.780 128.490 42.100 128.550 ;
        RECT 39.955 128.350 42.100 128.490 ;
        RECT 39.955 128.305 40.245 128.350 ;
        RECT 41.780 128.290 42.100 128.350 ;
        RECT 55.120 128.290 55.440 128.550 ;
        RECT 57.880 128.290 58.200 128.550 ;
        RECT 63.415 128.490 63.705 128.535 ;
        RECT 65.240 128.490 65.560 128.550 ;
        RECT 63.415 128.350 65.560 128.490 ;
        RECT 63.415 128.305 63.705 128.350 ;
        RECT 65.240 128.290 65.560 128.350 ;
        RECT 71.680 128.490 72.000 128.550 ;
        RECT 86.860 128.490 87.180 128.550 ;
        RECT 88.255 128.490 88.545 128.535 ;
        RECT 71.680 128.350 79.730 128.490 ;
        RECT 71.680 128.290 72.000 128.350 ;
        RECT 61.100 128.150 61.420 128.210 ;
        RECT 26.230 128.010 30.050 128.150 ;
        RECT 53.370 128.010 61.420 128.150 ;
        RECT 21.555 127.670 24.070 127.810 ;
        RECT 18.290 127.625 18.580 127.670 ;
        RECT 21.555 127.625 21.845 127.670 ;
        RECT 24.760 127.610 25.080 127.870 ;
        RECT 26.230 127.855 26.370 128.010 ;
        RECT 26.155 127.625 26.445 127.855 ;
        RECT 27.060 127.810 27.380 127.870 ;
        RECT 27.535 127.810 27.825 127.855 ;
        RECT 27.060 127.670 27.825 127.810 ;
        RECT 27.060 127.610 27.380 127.670 ;
        RECT 27.535 127.625 27.825 127.670 ;
        RECT 28.440 127.610 28.760 127.870 ;
        RECT 35.800 127.810 36.120 127.870 ;
        RECT 38.115 127.810 38.405 127.855 ;
        RECT 35.800 127.670 38.405 127.810 ;
        RECT 35.800 127.610 36.120 127.670 ;
        RECT 38.115 127.625 38.405 127.670 ;
        RECT 38.560 127.610 38.880 127.870 ;
        RECT 39.495 127.810 39.785 127.855 ;
        RECT 39.940 127.810 40.260 127.870 ;
        RECT 41.335 127.810 41.625 127.855 ;
        RECT 39.495 127.670 40.260 127.810 ;
        RECT 39.495 127.625 39.785 127.670 ;
        RECT 39.940 127.610 40.260 127.670 ;
        RECT 40.950 127.670 41.625 127.810 ;
        RECT 23.395 127.470 23.685 127.515 ;
        RECT 27.980 127.470 28.300 127.530 ;
        RECT 23.395 127.330 28.300 127.470 ;
        RECT 23.395 127.285 23.685 127.330 ;
        RECT 27.980 127.270 28.300 127.330 ;
        RECT 28.900 127.470 29.220 127.530 ;
        RECT 32.135 127.470 32.425 127.515 ;
        RECT 28.900 127.330 32.425 127.470 ;
        RECT 28.900 127.270 29.220 127.330 ;
        RECT 32.135 127.285 32.425 127.330 ;
        RECT 32.595 127.285 32.885 127.515 ;
        RECT 18.290 127.130 18.580 127.175 ;
        RECT 21.070 127.130 21.360 127.175 ;
        RECT 22.930 127.130 23.220 127.175 ;
        RECT 18.290 126.990 23.220 127.130 ;
        RECT 18.290 126.945 18.580 126.990 ;
        RECT 21.070 126.945 21.360 126.990 ;
        RECT 22.930 126.945 23.220 126.990 ;
        RECT 30.280 127.130 30.600 127.190 ;
        RECT 31.200 127.130 31.520 127.190 ;
        RECT 32.670 127.130 32.810 127.285 ;
        RECT 30.280 126.990 32.810 127.130 ;
        RECT 38.100 127.130 38.420 127.190 ;
        RECT 40.950 127.130 41.090 127.670 ;
        RECT 41.335 127.625 41.625 127.670 ;
        RECT 41.780 127.610 42.100 127.870 ;
        RECT 42.255 127.625 42.545 127.855 ;
        RECT 43.175 127.810 43.465 127.855 ;
        RECT 47.760 127.810 48.080 127.870 ;
        RECT 43.175 127.670 48.080 127.810 ;
        RECT 43.175 127.625 43.465 127.670 ;
        RECT 42.330 127.470 42.470 127.625 ;
        RECT 47.760 127.610 48.080 127.670 ;
        RECT 52.820 127.810 53.140 127.870 ;
        RECT 53.370 127.855 53.510 128.010 ;
        RECT 61.100 127.950 61.420 128.010 ;
        RECT 74.900 128.150 75.220 128.210 ;
        RECT 74.900 128.010 77.890 128.150 ;
        RECT 74.900 127.950 75.220 128.010 ;
        RECT 53.295 127.810 53.585 127.855 ;
        RECT 52.820 127.670 53.585 127.810 ;
        RECT 52.820 127.610 53.140 127.670 ;
        RECT 53.295 127.625 53.585 127.670 ;
        RECT 54.675 127.625 54.965 127.855 ;
        RECT 62.495 127.810 62.785 127.855 ;
        RECT 59.810 127.670 62.785 127.810 ;
        RECT 51.900 127.470 52.220 127.530 ;
        RECT 54.750 127.470 54.890 127.625 ;
        RECT 42.330 127.330 51.670 127.470 ;
        RECT 45.920 127.130 46.240 127.190 ;
        RECT 38.100 126.990 39.710 127.130 ;
        RECT 40.950 126.990 46.240 127.130 ;
        RECT 51.530 127.130 51.670 127.330 ;
        RECT 51.900 127.330 54.890 127.470 ;
        RECT 56.040 127.470 56.360 127.530 ;
        RECT 56.515 127.470 56.805 127.515 ;
        RECT 56.040 127.330 56.805 127.470 ;
        RECT 51.900 127.270 52.220 127.330 ;
        RECT 56.040 127.270 56.360 127.330 ;
        RECT 56.515 127.285 56.805 127.330 ;
        RECT 57.435 127.470 57.725 127.515 ;
        RECT 58.340 127.470 58.660 127.530 ;
        RECT 57.435 127.330 58.660 127.470 ;
        RECT 57.435 127.285 57.725 127.330 ;
        RECT 58.340 127.270 58.660 127.330 ;
        RECT 53.280 127.130 53.600 127.190 ;
        RECT 59.810 127.175 59.950 127.670 ;
        RECT 62.495 127.625 62.785 127.670 ;
        RECT 63.875 127.625 64.165 127.855 ;
        RECT 61.100 127.470 61.420 127.530 ;
        RECT 63.950 127.470 64.090 127.625 ;
        RECT 71.220 127.610 71.540 127.870 ;
        RECT 75.360 127.610 75.680 127.870 ;
        RECT 76.280 127.610 76.600 127.870 ;
        RECT 77.750 127.855 77.890 128.010 ;
        RECT 79.040 127.950 79.360 128.210 ;
        RECT 79.590 128.150 79.730 128.350 ;
        RECT 86.860 128.350 88.545 128.490 ;
        RECT 86.860 128.290 87.180 128.350 ;
        RECT 88.255 128.305 88.545 128.350 ;
        RECT 93.760 128.490 94.080 128.550 ;
        RECT 94.235 128.490 94.525 128.535 ;
        RECT 93.760 128.350 94.525 128.490 ;
        RECT 93.760 128.290 94.080 128.350 ;
        RECT 94.235 128.305 94.525 128.350 ;
        RECT 104.340 128.490 104.660 128.550 ;
        RECT 105.735 128.490 106.025 128.535 ;
        RECT 104.340 128.350 106.025 128.490 ;
        RECT 104.340 128.290 104.660 128.350 ;
        RECT 105.735 128.305 106.025 128.350 ;
        RECT 92.840 128.150 93.160 128.210 ;
        RECT 96.535 128.150 96.825 128.195 ;
        RECT 79.590 128.010 92.610 128.150 ;
        RECT 77.675 127.625 77.965 127.855 ;
        RECT 80.435 127.810 80.725 127.855 ;
        RECT 78.210 127.670 80.725 127.810 ;
        RECT 61.100 127.330 64.090 127.470 ;
        RECT 61.100 127.270 61.420 127.330 ;
        RECT 72.140 127.270 72.460 127.530 ;
        RECT 72.600 127.470 72.920 127.530 ;
        RECT 74.455 127.470 74.745 127.515 ;
        RECT 72.600 127.330 74.745 127.470 ;
        RECT 75.450 127.470 75.590 127.610 ;
        RECT 78.210 127.530 78.350 127.670 ;
        RECT 80.435 127.625 80.725 127.670 ;
        RECT 87.780 127.810 88.100 127.870 ;
        RECT 88.715 127.810 89.005 127.855 ;
        RECT 87.780 127.670 89.005 127.810 ;
        RECT 87.780 127.610 88.100 127.670 ;
        RECT 88.715 127.625 89.005 127.670 ;
        RECT 91.920 127.610 92.240 127.870 ;
        RECT 92.470 127.810 92.610 128.010 ;
        RECT 92.840 128.010 96.825 128.150 ;
        RECT 92.840 127.950 93.160 128.010 ;
        RECT 96.535 127.965 96.825 128.010 ;
        RECT 105.275 128.150 105.565 128.195 ;
        RECT 108.020 128.150 108.340 128.210 ;
        RECT 119.520 128.195 119.840 128.210 ;
        RECT 105.275 128.010 108.340 128.150 ;
        RECT 105.275 127.965 105.565 128.010 ;
        RECT 108.020 127.950 108.340 128.010 ;
        RECT 116.250 128.150 116.540 128.195 ;
        RECT 119.510 128.150 119.840 128.195 ;
        RECT 116.250 128.010 119.840 128.150 ;
        RECT 116.250 127.965 116.540 128.010 ;
        RECT 119.510 127.965 119.840 128.010 ;
        RECT 119.520 127.950 119.840 127.965 ;
        RECT 120.430 128.150 120.720 128.195 ;
        RECT 122.290 128.150 122.580 128.195 ;
        RECT 120.430 128.010 122.580 128.150 ;
        RECT 120.430 127.965 120.720 128.010 ;
        RECT 122.290 127.965 122.580 128.010 ;
        RECT 95.155 127.810 95.445 127.855 ;
        RECT 101.580 127.810 101.900 127.870 ;
        RECT 106.640 127.810 106.960 127.870 ;
        RECT 92.470 127.670 106.960 127.810 ;
        RECT 95.155 127.625 95.445 127.670 ;
        RECT 101.580 127.610 101.900 127.670 ;
        RECT 106.640 127.610 106.960 127.670 ;
        RECT 110.335 127.810 110.625 127.855 ;
        RECT 110.780 127.810 111.100 127.870 ;
        RECT 114.460 127.855 114.780 127.870 ;
        RECT 114.245 127.810 114.780 127.855 ;
        RECT 110.335 127.670 114.780 127.810 ;
        RECT 110.335 127.625 110.625 127.670 ;
        RECT 110.780 127.610 111.100 127.670 ;
        RECT 114.245 127.625 114.780 127.670 ;
        RECT 118.110 127.810 118.400 127.855 ;
        RECT 120.430 127.810 120.645 127.965 ;
        RECT 122.740 127.810 123.060 127.870 ;
        RECT 118.110 127.670 120.645 127.810 ;
        RECT 121.450 127.670 123.060 127.810 ;
        RECT 118.110 127.625 118.400 127.670 ;
        RECT 114.460 127.610 114.780 127.625 ;
        RECT 78.120 127.470 78.440 127.530 ;
        RECT 75.450 127.330 78.440 127.470 ;
        RECT 72.600 127.270 72.920 127.330 ;
        RECT 74.455 127.285 74.745 127.330 ;
        RECT 78.120 127.270 78.440 127.330 ;
        RECT 78.595 127.470 78.885 127.515 ;
        RECT 80.880 127.470 81.200 127.530 ;
        RECT 78.595 127.330 81.200 127.470 ;
        RECT 78.595 127.285 78.885 127.330 ;
        RECT 80.880 127.270 81.200 127.330 ;
        RECT 81.340 127.270 81.660 127.530 ;
        RECT 96.060 127.270 96.380 127.530 ;
        RECT 107.560 127.270 107.880 127.530 ;
        RECT 108.955 127.285 109.245 127.515 ;
        RECT 51.530 126.990 53.600 127.130 ;
        RECT 30.280 126.930 30.600 126.990 ;
        RECT 31.200 126.930 31.520 126.990 ;
        RECT 38.100 126.930 38.420 126.990 ;
        RECT 29.360 126.590 29.680 126.850 ;
        RECT 37.195 126.790 37.485 126.835 ;
        RECT 37.640 126.790 37.960 126.850 ;
        RECT 37.195 126.650 37.960 126.790 ;
        RECT 37.195 126.605 37.485 126.650 ;
        RECT 37.640 126.590 37.960 126.650 ;
        RECT 39.020 126.590 39.340 126.850 ;
        RECT 39.570 126.790 39.710 126.990 ;
        RECT 45.920 126.930 46.240 126.990 ;
        RECT 53.280 126.930 53.600 126.990 ;
        RECT 59.735 126.945 60.025 127.175 ;
        RECT 76.755 127.130 77.045 127.175 ;
        RECT 87.780 127.130 88.100 127.190 ;
        RECT 60.270 126.990 66.620 127.130 ;
        RECT 60.270 126.790 60.410 126.990 ;
        RECT 39.570 126.650 60.410 126.790 ;
        RECT 63.400 126.790 63.720 126.850 ;
        RECT 64.335 126.790 64.625 126.835 ;
        RECT 63.400 126.650 64.625 126.790 ;
        RECT 66.480 126.790 66.620 126.990 ;
        RECT 76.755 126.990 88.100 127.130 ;
        RECT 76.755 126.945 77.045 126.990 ;
        RECT 87.780 126.930 88.100 126.990 ;
        RECT 106.180 127.130 106.500 127.190 ;
        RECT 109.030 127.130 109.170 127.285 ;
        RECT 109.860 127.270 110.180 127.530 ;
        RECT 121.450 127.515 121.590 127.670 ;
        RECT 122.740 127.610 123.060 127.670 ;
        RECT 121.375 127.285 121.665 127.515 ;
        RECT 121.820 127.470 122.140 127.530 ;
        RECT 123.215 127.470 123.505 127.515 ;
        RECT 121.820 127.330 123.505 127.470 ;
        RECT 121.820 127.270 122.140 127.330 ;
        RECT 123.215 127.285 123.505 127.330 ;
        RECT 106.180 126.990 109.170 127.130 ;
        RECT 118.110 127.130 118.400 127.175 ;
        RECT 120.890 127.130 121.180 127.175 ;
        RECT 122.750 127.130 123.040 127.175 ;
        RECT 118.110 126.990 123.040 127.130 ;
        RECT 106.180 126.930 106.500 126.990 ;
        RECT 118.110 126.945 118.400 126.990 ;
        RECT 120.890 126.945 121.180 126.990 ;
        RECT 122.750 126.945 123.040 126.990 ;
        RECT 70.300 126.790 70.620 126.850 ;
        RECT 66.480 126.650 70.620 126.790 ;
        RECT 63.400 126.590 63.720 126.650 ;
        RECT 64.335 126.605 64.625 126.650 ;
        RECT 70.300 126.590 70.620 126.650 ;
        RECT 77.660 126.590 77.980 126.850 ;
        RECT 79.500 126.590 79.820 126.850 ;
        RECT 112.175 126.790 112.465 126.835 ;
        RECT 124.120 126.790 124.440 126.850 ;
        RECT 112.175 126.650 124.440 126.790 ;
        RECT 112.175 126.605 112.465 126.650 ;
        RECT 124.120 126.590 124.440 126.650 ;
        RECT 11.810 125.970 125.890 126.450 ;
        RECT 17.400 125.570 17.720 125.830 ;
        RECT 29.360 125.770 29.680 125.830 ;
        RECT 39.035 125.770 39.325 125.815 ;
        RECT 43.160 125.770 43.480 125.830 ;
        RECT 29.360 125.630 39.325 125.770 ;
        RECT 29.360 125.570 29.680 125.630 ;
        RECT 39.035 125.585 39.325 125.630 ;
        RECT 39.570 125.630 43.480 125.770 ;
        RECT 20.160 125.430 20.480 125.490 ;
        RECT 19.790 125.290 20.480 125.430 ;
        RECT 19.790 125.135 19.930 125.290 ;
        RECT 20.160 125.230 20.480 125.290 ;
        RECT 28.440 125.430 28.760 125.490 ;
        RECT 39.570 125.430 39.710 125.630 ;
        RECT 43.160 125.570 43.480 125.630 ;
        RECT 44.080 125.570 44.400 125.830 ;
        RECT 49.600 125.570 49.920 125.830 ;
        RECT 77.660 125.570 77.980 125.830 ;
        RECT 86.415 125.770 86.705 125.815 ;
        RECT 91.920 125.770 92.240 125.830 ;
        RECT 122.740 125.770 123.060 125.830 ;
        RECT 123.215 125.770 123.505 125.815 ;
        RECT 86.415 125.630 92.240 125.770 ;
        RECT 86.415 125.585 86.705 125.630 ;
        RECT 91.920 125.570 92.240 125.630 ;
        RECT 114.780 125.630 121.590 125.770 ;
        RECT 28.440 125.290 39.710 125.430 ;
        RECT 41.795 125.430 42.085 125.475 ;
        RECT 46.380 125.430 46.700 125.490 ;
        RECT 41.795 125.290 46.700 125.430 ;
        RECT 28.440 125.230 28.760 125.290 ;
        RECT 19.255 124.905 19.545 125.135 ;
        RECT 19.715 124.905 20.005 125.135 ;
        RECT 27.075 125.090 27.365 125.135 ;
        RECT 28.900 125.090 29.220 125.150 ;
        RECT 20.250 124.950 26.370 125.090 ;
        RECT 16.940 124.550 17.260 124.810 ;
        RECT 19.330 124.750 19.470 124.905 ;
        RECT 20.250 124.750 20.390 124.950 ;
        RECT 22.935 124.750 23.225 124.795 ;
        RECT 19.330 124.610 20.390 124.750 ;
        RECT 22.090 124.610 23.225 124.750 ;
        RECT 20.160 123.870 20.480 124.130 ;
        RECT 22.090 124.115 22.230 124.610 ;
        RECT 22.935 124.565 23.225 124.610 ;
        RECT 26.230 124.410 26.370 124.950 ;
        RECT 27.075 124.950 29.220 125.090 ;
        RECT 27.075 124.905 27.365 124.950 ;
        RECT 28.900 124.890 29.220 124.950 ;
        RECT 27.995 124.750 28.285 124.795 ;
        RECT 29.450 124.750 29.590 125.290 ;
        RECT 41.795 125.245 42.085 125.290 ;
        RECT 46.380 125.230 46.700 125.290 ;
        RECT 50.060 125.430 50.380 125.490 ;
        RECT 61.990 125.430 62.280 125.475 ;
        RECT 64.770 125.430 65.060 125.475 ;
        RECT 66.630 125.430 66.920 125.475 ;
        RECT 50.060 125.290 51.670 125.430 ;
        RECT 50.060 125.230 50.380 125.290 ;
        RECT 39.480 124.890 39.800 125.150 ;
        RECT 43.620 124.890 43.940 125.150 ;
        RECT 44.540 125.090 44.860 125.150 ;
        RECT 44.170 124.950 44.860 125.090 ;
        RECT 27.995 124.610 29.590 124.750 ;
        RECT 27.995 124.565 28.285 124.610 ;
        RECT 38.100 124.550 38.420 124.810 ;
        RECT 40.415 124.750 40.705 124.795 ;
        RECT 41.320 124.750 41.640 124.810 ;
        RECT 40.415 124.610 41.640 124.750 ;
        RECT 40.415 124.565 40.705 124.610 ;
        RECT 41.320 124.550 41.640 124.610 ;
        RECT 42.700 124.550 43.020 124.810 ;
        RECT 44.170 124.750 44.310 124.950 ;
        RECT 44.540 124.890 44.860 124.950 ;
        RECT 46.010 124.950 51.210 125.090 ;
        RECT 46.010 124.810 46.150 124.950 ;
        RECT 43.710 124.610 44.310 124.750 ;
        RECT 28.915 124.410 29.205 124.455 ;
        RECT 30.740 124.410 31.060 124.470 ;
        RECT 26.230 124.270 28.670 124.410 ;
        RECT 28.530 124.130 28.670 124.270 ;
        RECT 28.915 124.270 31.060 124.410 ;
        RECT 28.915 124.225 29.205 124.270 ;
        RECT 30.740 124.210 31.060 124.270 ;
        RECT 39.035 124.410 39.325 124.455 ;
        RECT 43.710 124.410 43.850 124.610 ;
        RECT 45.920 124.550 46.240 124.810 ;
        RECT 46.395 124.565 46.685 124.795 ;
        RECT 46.855 124.565 47.145 124.795 ;
        RECT 39.035 124.270 43.850 124.410 ;
        RECT 44.095 124.410 44.385 124.455 ;
        RECT 44.555 124.410 44.845 124.455 ;
        RECT 44.095 124.270 44.845 124.410 ;
        RECT 39.035 124.225 39.325 124.270 ;
        RECT 44.095 124.225 44.385 124.270 ;
        RECT 44.555 124.225 44.845 124.270 ;
        RECT 22.015 123.885 22.305 124.115 ;
        RECT 23.380 124.070 23.700 124.130 ;
        RECT 23.855 124.070 24.145 124.115 ;
        RECT 23.380 123.930 24.145 124.070 ;
        RECT 23.380 123.870 23.700 123.930 ;
        RECT 23.855 123.885 24.145 123.930 ;
        RECT 28.440 124.070 28.760 124.130 ;
        RECT 30.280 124.070 30.600 124.130 ;
        RECT 28.440 123.930 30.600 124.070 ;
        RECT 28.440 123.870 28.760 123.930 ;
        RECT 30.280 123.870 30.600 123.930 ;
        RECT 31.200 124.070 31.520 124.130 ;
        RECT 31.675 124.070 31.965 124.115 ;
        RECT 31.200 123.930 31.965 124.070 ;
        RECT 31.200 123.870 31.520 123.930 ;
        RECT 31.675 123.885 31.965 123.930 ;
        RECT 41.335 124.070 41.625 124.115 ;
        RECT 42.700 124.070 43.020 124.130 ;
        RECT 41.335 123.930 43.020 124.070 ;
        RECT 46.470 124.070 46.610 124.565 ;
        RECT 46.930 124.410 47.070 124.565 ;
        RECT 47.760 124.550 48.080 124.810 ;
        RECT 51.070 124.795 51.210 124.950 ;
        RECT 51.530 124.795 51.670 125.290 ;
        RECT 61.990 125.290 66.920 125.430 ;
        RECT 61.990 125.245 62.280 125.290 ;
        RECT 64.770 125.245 65.060 125.290 ;
        RECT 66.630 125.245 66.920 125.290 ;
        RECT 103.895 125.245 104.185 125.475 ;
        RECT 111.715 125.430 112.005 125.475 ;
        RECT 114.780 125.430 114.920 125.630 ;
        RECT 111.715 125.290 114.920 125.430 ;
        RECT 116.270 125.430 116.560 125.475 ;
        RECT 119.050 125.430 119.340 125.475 ;
        RECT 120.910 125.430 121.200 125.475 ;
        RECT 116.270 125.290 121.200 125.430 ;
        RECT 121.450 125.430 121.590 125.630 ;
        RECT 122.740 125.630 123.505 125.770 ;
        RECT 122.740 125.570 123.060 125.630 ;
        RECT 123.215 125.585 123.505 125.630 ;
        RECT 121.450 125.290 122.970 125.430 ;
        RECT 111.715 125.245 112.005 125.290 ;
        RECT 116.270 125.245 116.560 125.290 ;
        RECT 119.050 125.245 119.340 125.290 ;
        RECT 120.910 125.245 121.200 125.290 ;
        RECT 58.340 125.135 58.660 125.150 ;
        RECT 58.125 125.090 58.660 125.135 ;
        RECT 51.990 124.950 58.660 125.090 ;
        RECT 51.990 124.795 52.130 124.950 ;
        RECT 58.125 124.905 58.660 124.950 ;
        RECT 58.340 124.890 58.660 124.905 ;
        RECT 65.240 124.890 65.560 125.150 ;
        RECT 65.700 125.090 66.020 125.150 ;
        RECT 67.095 125.090 67.385 125.135 ;
        RECT 65.700 124.950 67.385 125.090 ;
        RECT 65.700 124.890 66.020 124.950 ;
        RECT 67.095 124.905 67.385 124.950 ;
        RECT 101.120 124.890 101.440 125.150 ;
        RECT 50.995 124.565 51.285 124.795 ;
        RECT 51.455 124.565 51.745 124.795 ;
        RECT 51.915 124.565 52.205 124.795 ;
        RECT 52.360 124.750 52.680 124.810 ;
        RECT 52.835 124.750 53.125 124.795 ;
        RECT 52.360 124.610 53.125 124.750 ;
        RECT 52.360 124.550 52.680 124.610 ;
        RECT 52.835 124.565 53.125 124.610 ;
        RECT 61.990 124.750 62.280 124.795 ;
        RECT 70.300 124.750 70.620 124.810 ;
        RECT 71.235 124.750 71.525 124.795 ;
        RECT 61.990 124.610 64.525 124.750 ;
        RECT 61.990 124.565 62.280 124.610 ;
        RECT 53.280 124.410 53.600 124.470 ;
        RECT 63.400 124.455 63.720 124.470 ;
        RECT 46.930 124.270 53.600 124.410 ;
        RECT 53.280 124.210 53.600 124.270 ;
        RECT 60.130 124.410 60.420 124.455 ;
        RECT 63.390 124.410 63.720 124.455 ;
        RECT 60.130 124.270 63.720 124.410 ;
        RECT 60.130 124.225 60.420 124.270 ;
        RECT 63.390 124.225 63.720 124.270 ;
        RECT 64.310 124.455 64.525 124.610 ;
        RECT 70.300 124.610 71.525 124.750 ;
        RECT 70.300 124.550 70.620 124.610 ;
        RECT 71.235 124.565 71.525 124.610 ;
        RECT 78.120 124.750 78.440 124.810 ;
        RECT 78.595 124.750 78.885 124.795 ;
        RECT 78.120 124.610 78.885 124.750 ;
        RECT 78.120 124.550 78.440 124.610 ;
        RECT 78.595 124.565 78.885 124.610 ;
        RECT 79.055 124.565 79.345 124.795 ;
        RECT 64.310 124.410 64.600 124.455 ;
        RECT 66.170 124.410 66.460 124.455 ;
        RECT 64.310 124.270 66.460 124.410 ;
        RECT 64.310 124.225 64.600 124.270 ;
        RECT 66.170 124.225 66.460 124.270 ;
        RECT 75.360 124.410 75.680 124.470 ;
        RECT 79.130 124.410 79.270 124.565 ;
        RECT 92.840 124.550 93.160 124.810 ;
        RECT 103.970 124.750 104.110 125.245 ;
        RECT 106.180 125.090 106.500 125.150 ;
        RECT 108.495 125.090 108.785 125.135 ;
        RECT 106.180 124.950 108.785 125.090 ;
        RECT 106.180 124.890 106.500 124.950 ;
        RECT 108.495 124.905 108.785 124.950 ;
        RECT 121.375 125.090 121.665 125.135 ;
        RECT 121.820 125.090 122.140 125.150 ;
        RECT 121.375 124.950 122.140 125.090 ;
        RECT 121.375 124.905 121.665 124.950 ;
        RECT 121.820 124.890 122.140 124.950 ;
        RECT 104.815 124.750 105.105 124.795 ;
        RECT 103.970 124.610 105.105 124.750 ;
        RECT 104.815 124.565 105.105 124.610 ;
        RECT 109.860 124.750 110.180 124.810 ;
        RECT 122.830 124.795 122.970 125.290 ;
        RECT 112.405 124.750 112.695 124.795 ;
        RECT 109.860 124.610 112.695 124.750 ;
        RECT 109.860 124.550 110.180 124.610 ;
        RECT 112.405 124.565 112.695 124.610 ;
        RECT 116.270 124.750 116.560 124.795 ;
        RECT 119.535 124.750 119.825 124.795 ;
        RECT 116.270 124.610 118.805 124.750 ;
        RECT 116.270 124.565 116.560 124.610 ;
        RECT 87.320 124.410 87.640 124.470 ;
        RECT 93.760 124.410 94.080 124.470 ;
        RECT 117.680 124.455 118.000 124.470 ;
        RECT 109.415 124.410 109.705 124.455 ;
        RECT 75.360 124.270 94.080 124.410 ;
        RECT 63.400 124.210 63.720 124.225 ;
        RECT 75.360 124.210 75.680 124.270 ;
        RECT 87.320 124.210 87.640 124.270 ;
        RECT 93.760 124.210 94.080 124.270 ;
        RECT 102.130 124.270 109.705 124.410 ;
        RECT 102.130 124.130 102.270 124.270 ;
        RECT 109.415 124.225 109.705 124.270 ;
        RECT 114.410 124.410 114.700 124.455 ;
        RECT 117.670 124.410 118.000 124.455 ;
        RECT 114.410 124.270 118.000 124.410 ;
        RECT 114.410 124.225 114.700 124.270 ;
        RECT 117.670 124.225 118.000 124.270 ;
        RECT 118.590 124.455 118.805 124.610 ;
        RECT 119.535 124.610 121.130 124.750 ;
        RECT 119.535 124.565 119.825 124.610 ;
        RECT 118.590 124.410 118.880 124.455 ;
        RECT 120.450 124.410 120.740 124.455 ;
        RECT 118.590 124.270 120.740 124.410 ;
        RECT 118.590 124.225 118.880 124.270 ;
        RECT 120.450 124.225 120.740 124.270 ;
        RECT 117.680 124.210 118.000 124.225 ;
        RECT 50.060 124.070 50.380 124.130 ;
        RECT 46.470 123.930 50.380 124.070 ;
        RECT 41.335 123.885 41.625 123.930 ;
        RECT 42.700 123.870 43.020 123.930 ;
        RECT 50.060 123.870 50.380 123.930 ;
        RECT 71.680 123.870 72.000 124.130 ;
        RECT 81.340 124.070 81.660 124.130 ;
        RECT 83.180 124.070 83.500 124.130 ;
        RECT 101.595 124.070 101.885 124.115 ;
        RECT 81.340 123.930 101.885 124.070 ;
        RECT 81.340 123.870 81.660 123.930 ;
        RECT 83.180 123.870 83.500 123.930 ;
        RECT 101.595 123.885 101.885 123.930 ;
        RECT 102.040 123.870 102.360 124.130 ;
        RECT 105.735 124.070 106.025 124.115 ;
        RECT 106.640 124.070 106.960 124.130 ;
        RECT 105.735 123.930 106.960 124.070 ;
        RECT 120.990 124.070 121.130 124.610 ;
        RECT 122.755 124.565 123.045 124.795 ;
        RECT 124.120 124.550 124.440 124.810 ;
        RECT 121.835 124.070 122.125 124.115 ;
        RECT 120.990 123.930 122.125 124.070 ;
        RECT 105.735 123.885 106.025 123.930 ;
        RECT 106.640 123.870 106.960 123.930 ;
        RECT 121.835 123.885 122.125 123.930 ;
        RECT 11.010 123.250 125.890 123.730 ;
        RECT 27.980 123.050 28.300 123.110 ;
        RECT 31.200 123.050 31.520 123.110 ;
        RECT 27.150 122.910 34.650 123.050 ;
        RECT 16.020 122.710 16.340 122.770 ;
        RECT 16.890 122.710 17.180 122.755 ;
        RECT 20.150 122.710 20.440 122.755 ;
        RECT 16.020 122.570 20.440 122.710 ;
        RECT 16.020 122.510 16.340 122.570 ;
        RECT 16.890 122.525 17.180 122.570 ;
        RECT 20.150 122.525 20.440 122.570 ;
        RECT 21.070 122.710 21.360 122.755 ;
        RECT 22.930 122.710 23.220 122.755 ;
        RECT 21.070 122.570 23.220 122.710 ;
        RECT 21.070 122.525 21.360 122.570 ;
        RECT 22.930 122.525 23.220 122.570 ;
        RECT 14.885 122.370 15.175 122.415 ;
        RECT 17.860 122.370 18.180 122.430 ;
        RECT 14.885 122.230 18.180 122.370 ;
        RECT 14.885 122.185 15.175 122.230 ;
        RECT 17.860 122.170 18.180 122.230 ;
        RECT 18.750 122.370 19.040 122.415 ;
        RECT 21.070 122.370 21.285 122.525 ;
        RECT 18.750 122.230 21.285 122.370 ;
        RECT 23.855 122.370 24.145 122.415 ;
        RECT 27.150 122.370 27.290 122.910 ;
        RECT 27.980 122.850 28.300 122.910 ;
        RECT 31.200 122.850 31.520 122.910 ;
        RECT 27.520 122.755 27.840 122.770 ;
        RECT 27.470 122.710 27.840 122.755 ;
        RECT 30.730 122.710 31.020 122.755 ;
        RECT 27.470 122.570 31.020 122.710 ;
        RECT 27.470 122.525 27.840 122.570 ;
        RECT 30.730 122.525 31.020 122.570 ;
        RECT 31.650 122.710 31.940 122.755 ;
        RECT 33.510 122.710 33.800 122.755 ;
        RECT 31.650 122.570 33.800 122.710 ;
        RECT 31.650 122.525 31.940 122.570 ;
        RECT 33.510 122.525 33.800 122.570 ;
        RECT 27.520 122.510 27.840 122.525 ;
        RECT 23.855 122.230 27.290 122.370 ;
        RECT 29.330 122.370 29.620 122.415 ;
        RECT 31.650 122.370 31.865 122.525 ;
        RECT 34.510 122.415 34.650 122.910 ;
        RECT 38.100 122.850 38.420 123.110 ;
        RECT 39.020 123.050 39.340 123.110 ;
        RECT 40.415 123.050 40.705 123.095 ;
        RECT 39.020 122.910 40.705 123.050 ;
        RECT 39.020 122.850 39.340 122.910 ;
        RECT 40.415 122.865 40.705 122.910 ;
        RECT 41.320 123.050 41.640 123.110 ;
        RECT 43.160 123.050 43.480 123.110 ;
        RECT 41.320 122.910 43.480 123.050 ;
        RECT 41.320 122.850 41.640 122.910 ;
        RECT 43.160 122.850 43.480 122.910 ;
        RECT 44.080 123.050 44.400 123.110 ;
        RECT 44.555 123.050 44.845 123.095 ;
        RECT 44.080 122.910 44.845 123.050 ;
        RECT 44.080 122.850 44.400 122.910 ;
        RECT 44.555 122.865 44.845 122.910 ;
        RECT 58.340 122.850 58.660 123.110 ;
        RECT 60.195 122.865 60.485 123.095 ;
        RECT 71.925 123.050 72.215 123.095 ;
        RECT 72.600 123.050 72.920 123.110 ;
        RECT 71.925 122.910 72.920 123.050 ;
        RECT 71.925 122.865 72.215 122.910 ;
        RECT 34.880 122.710 35.200 122.770 ;
        RECT 36.735 122.710 37.025 122.755 ;
        RECT 34.880 122.570 37.025 122.710 ;
        RECT 38.190 122.710 38.330 122.850 ;
        RECT 45.475 122.710 45.765 122.755 ;
        RECT 38.190 122.570 45.765 122.710 ;
        RECT 34.880 122.510 35.200 122.570 ;
        RECT 36.735 122.525 37.025 122.570 ;
        RECT 45.475 122.525 45.765 122.570 ;
        RECT 32.595 122.370 32.885 122.415 ;
        RECT 29.330 122.230 31.865 122.370 ;
        RECT 32.210 122.230 32.885 122.370 ;
        RECT 18.750 122.185 19.040 122.230 ;
        RECT 23.855 122.185 24.145 122.230 ;
        RECT 29.330 122.185 29.620 122.230 ;
        RECT 22.015 122.030 22.305 122.075 ;
        RECT 22.920 122.030 23.240 122.090 ;
        RECT 22.015 121.890 23.240 122.030 ;
        RECT 22.015 121.845 22.305 121.890 ;
        RECT 22.920 121.830 23.240 121.890 ;
        RECT 25.465 122.030 25.755 122.075 ;
        RECT 28.900 122.030 29.220 122.090 ;
        RECT 25.465 121.890 29.220 122.030 ;
        RECT 25.465 121.845 25.755 121.890 ;
        RECT 28.900 121.830 29.220 121.890 ;
        RECT 30.740 122.030 31.060 122.090 ;
        RECT 32.210 122.030 32.350 122.230 ;
        RECT 32.595 122.185 32.885 122.230 ;
        RECT 34.435 122.370 34.725 122.415 ;
        RECT 34.435 122.230 37.870 122.370 ;
        RECT 34.435 122.185 34.725 122.230 ;
        RECT 30.740 121.890 32.350 122.030 ;
        RECT 37.730 122.030 37.870 122.230 ;
        RECT 38.100 122.170 38.420 122.430 ;
        RECT 38.560 122.170 38.880 122.430 ;
        RECT 41.320 122.170 41.640 122.430 ;
        RECT 42.255 122.370 42.545 122.415 ;
        RECT 42.255 122.230 43.390 122.370 ;
        RECT 42.255 122.185 42.545 122.230 ;
        RECT 41.780 122.030 42.100 122.090 ;
        RECT 42.715 122.030 43.005 122.075 ;
        RECT 37.730 121.890 41.550 122.030 ;
        RECT 30.740 121.830 31.060 121.890 ;
        RECT 41.410 121.750 41.550 121.890 ;
        RECT 41.780 121.890 43.005 122.030 ;
        RECT 41.780 121.830 42.100 121.890 ;
        RECT 42.715 121.845 43.005 121.890 ;
        RECT 18.750 121.690 19.040 121.735 ;
        RECT 21.530 121.690 21.820 121.735 ;
        RECT 23.390 121.690 23.680 121.735 ;
        RECT 18.750 121.550 23.680 121.690 ;
        RECT 18.750 121.505 19.040 121.550 ;
        RECT 21.530 121.505 21.820 121.550 ;
        RECT 23.390 121.505 23.680 121.550 ;
        RECT 29.330 121.690 29.620 121.735 ;
        RECT 32.110 121.690 32.400 121.735 ;
        RECT 33.970 121.690 34.260 121.735 ;
        RECT 29.330 121.550 34.260 121.690 ;
        RECT 29.330 121.505 29.620 121.550 ;
        RECT 32.110 121.505 32.400 121.550 ;
        RECT 33.970 121.505 34.260 121.550 ;
        RECT 34.510 121.550 40.170 121.690 ;
        RECT 20.160 121.350 20.480 121.410 ;
        RECT 34.510 121.350 34.650 121.550 ;
        RECT 20.160 121.210 34.650 121.350 ;
        RECT 39.020 121.350 39.340 121.410 ;
        RECT 39.495 121.350 39.785 121.395 ;
        RECT 39.020 121.210 39.785 121.350 ;
        RECT 40.030 121.350 40.170 121.550 ;
        RECT 41.320 121.490 41.640 121.750 ;
        RECT 43.250 121.350 43.390 122.230 ;
        RECT 43.620 122.170 43.940 122.430 ;
        RECT 53.280 122.370 53.600 122.430 ;
        RECT 57.895 122.370 58.185 122.415 ;
        RECT 53.280 122.230 58.185 122.370 ;
        RECT 60.270 122.370 60.410 122.865 ;
        RECT 72.600 122.850 72.920 122.910 ;
        RECT 83.180 122.850 83.500 123.110 ;
        RECT 87.320 123.095 87.640 123.110 ;
        RECT 87.320 122.865 87.855 123.095 ;
        RECT 94.680 123.050 95.000 123.110 ;
        RECT 99.525 123.050 99.815 123.095 ;
        RECT 102.040 123.050 102.360 123.110 ;
        RECT 94.680 122.910 97.670 123.050 ;
        RECT 87.320 122.850 87.640 122.865 ;
        RECT 94.680 122.850 95.000 122.910 ;
        RECT 77.200 122.755 77.520 122.770 ;
        RECT 73.930 122.710 74.220 122.755 ;
        RECT 77.190 122.710 77.520 122.755 ;
        RECT 73.930 122.570 77.520 122.710 ;
        RECT 73.930 122.525 74.220 122.570 ;
        RECT 77.190 122.525 77.520 122.570 ;
        RECT 77.200 122.510 77.520 122.525 ;
        RECT 78.110 122.710 78.400 122.755 ;
        RECT 79.970 122.710 80.260 122.755 ;
        RECT 82.735 122.710 83.025 122.755 ;
        RECT 78.110 122.570 80.260 122.710 ;
        RECT 78.110 122.525 78.400 122.570 ;
        RECT 79.970 122.525 80.260 122.570 ;
        RECT 80.510 122.570 83.025 122.710 ;
        RECT 61.575 122.370 61.865 122.415 ;
        RECT 60.270 122.230 61.865 122.370 ;
        RECT 53.280 122.170 53.600 122.230 ;
        RECT 57.895 122.185 58.185 122.230 ;
        RECT 61.575 122.185 61.865 122.230 ;
        RECT 75.790 122.370 76.080 122.415 ;
        RECT 78.110 122.370 78.325 122.525 ;
        RECT 75.790 122.230 78.325 122.370 ;
        RECT 75.790 122.185 76.080 122.230 ;
        RECT 79.040 122.170 79.360 122.430 ;
        RECT 80.510 122.370 80.650 122.570 ;
        RECT 82.735 122.525 83.025 122.570 ;
        RECT 84.560 122.710 84.880 122.770 ;
        RECT 89.620 122.755 89.940 122.770 ;
        RECT 89.570 122.710 89.940 122.755 ;
        RECT 92.830 122.710 93.120 122.755 ;
        RECT 84.560 122.570 85.710 122.710 ;
        RECT 84.560 122.510 84.880 122.570 ;
        RECT 85.570 122.415 85.710 122.570 ;
        RECT 89.570 122.570 93.120 122.710 ;
        RECT 89.570 122.525 89.940 122.570 ;
        RECT 92.830 122.525 93.120 122.570 ;
        RECT 93.750 122.710 94.040 122.755 ;
        RECT 95.610 122.710 95.900 122.755 ;
        RECT 93.750 122.570 95.900 122.710 ;
        RECT 93.750 122.525 94.040 122.570 ;
        RECT 95.610 122.525 95.900 122.570 ;
        RECT 89.620 122.510 89.940 122.525 ;
        RECT 79.590 122.230 80.650 122.370 ;
        RECT 80.895 122.370 81.185 122.415 ;
        RECT 80.895 122.230 85.250 122.370 ;
        RECT 56.040 122.030 56.360 122.090 ;
        RECT 56.975 122.030 57.265 122.075 ;
        RECT 56.040 121.890 57.265 122.030 ;
        RECT 56.040 121.830 56.360 121.890 ;
        RECT 56.975 121.845 57.265 121.890 ;
        RECT 73.520 122.030 73.840 122.090 ;
        RECT 76.740 122.030 77.060 122.090 ;
        RECT 79.590 122.030 79.730 122.230 ;
        RECT 80.895 122.185 81.185 122.230 ;
        RECT 81.815 122.030 82.105 122.075 ;
        RECT 73.520 121.890 79.730 122.030 ;
        RECT 81.430 121.890 82.105 122.030 ;
        RECT 85.110 122.030 85.250 122.230 ;
        RECT 85.495 122.185 85.785 122.415 ;
        RECT 85.940 122.170 86.260 122.430 ;
        RECT 91.430 122.370 91.720 122.415 ;
        RECT 93.750 122.370 93.965 122.525 ;
        RECT 91.430 122.230 93.965 122.370 ;
        RECT 91.430 122.185 91.720 122.230 ;
        RECT 94.680 122.170 95.000 122.430 ;
        RECT 97.530 122.370 97.670 122.910 ;
        RECT 99.525 122.910 102.360 123.050 ;
        RECT 99.525 122.865 99.815 122.910 ;
        RECT 102.040 122.850 102.360 122.910 ;
        RECT 114.460 122.850 114.780 123.110 ;
        RECT 117.680 122.850 118.000 123.110 ;
        RECT 119.075 123.050 119.365 123.095 ;
        RECT 119.520 123.050 119.840 123.110 ;
        RECT 119.075 122.910 119.840 123.050 ;
        RECT 119.075 122.865 119.365 122.910 ;
        RECT 119.520 122.850 119.840 122.910 ;
        RECT 98.375 122.710 98.665 122.755 ;
        RECT 101.530 122.710 101.820 122.755 ;
        RECT 104.790 122.710 105.080 122.755 ;
        RECT 98.375 122.570 105.080 122.710 ;
        RECT 98.375 122.525 98.665 122.570 ;
        RECT 101.530 122.525 101.820 122.570 ;
        RECT 104.790 122.525 105.080 122.570 ;
        RECT 105.710 122.710 106.000 122.755 ;
        RECT 107.570 122.710 107.860 122.755 ;
        RECT 105.710 122.570 107.860 122.710 ;
        RECT 105.710 122.525 106.000 122.570 ;
        RECT 107.570 122.525 107.860 122.570 ;
        RECT 97.915 122.370 98.205 122.415 ;
        RECT 97.530 122.230 98.205 122.370 ;
        RECT 97.915 122.185 98.205 122.230 ;
        RECT 103.390 122.370 103.680 122.415 ;
        RECT 105.710 122.370 105.925 122.525 ;
        RECT 103.390 122.230 105.925 122.370 ;
        RECT 103.390 122.185 103.680 122.230 ;
        RECT 91.920 122.030 92.240 122.090 ;
        RECT 96.535 122.030 96.825 122.075 ;
        RECT 85.110 121.890 96.825 122.030 ;
        RECT 97.990 122.030 98.130 122.185 ;
        RECT 106.180 122.170 106.500 122.430 ;
        RECT 106.640 122.170 106.960 122.430 ;
        RECT 108.020 122.370 108.340 122.430 ;
        RECT 108.495 122.370 108.785 122.415 ;
        RECT 108.020 122.230 108.785 122.370 ;
        RECT 108.020 122.170 108.340 122.230 ;
        RECT 108.495 122.185 108.785 122.230 ;
        RECT 113.540 122.370 113.860 122.430 ;
        RECT 114.935 122.370 115.225 122.415 ;
        RECT 113.540 122.230 115.225 122.370 ;
        RECT 113.540 122.170 113.860 122.230 ;
        RECT 114.935 122.185 115.225 122.230 ;
        RECT 116.300 122.370 116.620 122.430 ;
        RECT 118.155 122.370 118.445 122.415 ;
        RECT 118.615 122.370 118.905 122.415 ;
        RECT 116.300 122.230 118.905 122.370 ;
        RECT 116.300 122.170 116.620 122.230 ;
        RECT 118.155 122.185 118.445 122.230 ;
        RECT 118.615 122.185 118.905 122.230 ;
        RECT 104.340 122.030 104.660 122.090 ;
        RECT 97.990 121.890 104.660 122.030 ;
        RECT 106.270 122.030 106.410 122.170 ;
        RECT 114.015 122.030 114.305 122.075 ;
        RECT 106.270 121.890 114.305 122.030 ;
        RECT 73.520 121.830 73.840 121.890 ;
        RECT 76.740 121.830 77.060 121.890 ;
        RECT 75.790 121.690 76.080 121.735 ;
        RECT 78.570 121.690 78.860 121.735 ;
        RECT 80.430 121.690 80.720 121.735 ;
        RECT 75.790 121.550 80.720 121.690 ;
        RECT 75.790 121.505 76.080 121.550 ;
        RECT 78.570 121.505 78.860 121.550 ;
        RECT 80.430 121.505 80.720 121.550 ;
        RECT 40.030 121.210 43.390 121.350 ;
        RECT 20.160 121.150 20.480 121.210 ;
        RECT 39.020 121.150 39.340 121.210 ;
        RECT 39.495 121.165 39.785 121.210 ;
        RECT 51.900 121.150 52.220 121.410 ;
        RECT 52.820 121.350 53.140 121.410 ;
        RECT 53.740 121.350 54.060 121.410 ;
        RECT 52.820 121.210 54.060 121.350 ;
        RECT 52.820 121.150 53.140 121.210 ;
        RECT 53.740 121.150 54.060 121.210 ;
        RECT 62.495 121.350 62.785 121.395 ;
        RECT 63.860 121.350 64.180 121.410 ;
        RECT 62.495 121.210 64.180 121.350 ;
        RECT 62.495 121.165 62.785 121.210 ;
        RECT 63.860 121.150 64.180 121.210 ;
        RECT 71.680 121.350 72.000 121.410 ;
        RECT 81.430 121.350 81.570 121.890 ;
        RECT 81.815 121.845 82.105 121.890 ;
        RECT 91.920 121.830 92.240 121.890 ;
        RECT 96.535 121.845 96.825 121.890 ;
        RECT 104.340 121.830 104.660 121.890 ;
        RECT 114.015 121.845 114.305 121.890 ;
        RECT 91.430 121.690 91.720 121.735 ;
        RECT 94.210 121.690 94.500 121.735 ;
        RECT 96.070 121.690 96.360 121.735 ;
        RECT 91.430 121.550 96.360 121.690 ;
        RECT 91.430 121.505 91.720 121.550 ;
        RECT 94.210 121.505 94.500 121.550 ;
        RECT 96.070 121.505 96.360 121.550 ;
        RECT 103.390 121.690 103.680 121.735 ;
        RECT 106.170 121.690 106.460 121.735 ;
        RECT 108.030 121.690 108.320 121.735 ;
        RECT 103.390 121.550 108.320 121.690 ;
        RECT 103.390 121.505 103.680 121.550 ;
        RECT 106.170 121.505 106.460 121.550 ;
        RECT 108.030 121.505 108.320 121.550 ;
        RECT 71.680 121.210 81.570 121.350 ;
        RECT 85.035 121.350 85.325 121.395 ;
        RECT 85.480 121.350 85.800 121.410 ;
        RECT 85.035 121.210 85.800 121.350 ;
        RECT 71.680 121.150 72.000 121.210 ;
        RECT 85.035 121.165 85.325 121.210 ;
        RECT 85.480 121.150 85.800 121.210 ;
        RECT 116.775 121.350 117.065 121.395 ;
        RECT 118.140 121.350 118.460 121.410 ;
        RECT 116.775 121.210 118.460 121.350 ;
        RECT 116.775 121.165 117.065 121.210 ;
        RECT 118.140 121.150 118.460 121.210 ;
        RECT 11.810 120.530 125.890 121.010 ;
        RECT 16.020 120.130 16.340 120.390 ;
        RECT 19.790 120.190 22.690 120.330 ;
        RECT 19.790 119.990 19.930 120.190 ;
        RECT 19.330 119.850 19.930 119.990 ;
        RECT 19.330 119.695 19.470 119.850 ;
        RECT 22.015 119.805 22.305 120.035 ;
        RECT 22.550 119.990 22.690 120.190 ;
        RECT 22.920 120.130 23.240 120.390 ;
        RECT 28.440 120.330 28.760 120.390 ;
        RECT 71.680 120.330 72.000 120.390 ;
        RECT 77.200 120.330 77.520 120.390 ;
        RECT 79.515 120.330 79.805 120.375 ;
        RECT 23.470 120.190 28.760 120.330 ;
        RECT 23.470 119.990 23.610 120.190 ;
        RECT 28.440 120.130 28.760 120.190 ;
        RECT 70.850 120.190 76.050 120.330 ;
        RECT 22.550 119.850 23.610 119.990 ;
        RECT 25.235 119.990 25.525 120.035 ;
        RECT 27.520 119.990 27.840 120.050 ;
        RECT 29.820 119.990 30.140 120.050 ;
        RECT 34.880 119.990 35.200 120.050 ;
        RECT 25.235 119.850 27.840 119.990 ;
        RECT 25.235 119.805 25.525 119.850 ;
        RECT 19.255 119.465 19.545 119.695 ;
        RECT 19.715 119.650 20.005 119.695 ;
        RECT 20.160 119.650 20.480 119.710 ;
        RECT 19.715 119.510 20.480 119.650 ;
        RECT 19.715 119.465 20.005 119.510 ;
        RECT 20.160 119.450 20.480 119.510 ;
        RECT 15.575 119.310 15.865 119.355 ;
        RECT 16.940 119.310 17.260 119.370 ;
        RECT 22.090 119.310 22.230 119.805 ;
        RECT 27.520 119.790 27.840 119.850 ;
        RECT 28.070 119.850 35.200 119.990 ;
        RECT 28.070 119.650 28.210 119.850 ;
        RECT 29.820 119.790 30.140 119.850 ;
        RECT 34.880 119.790 35.200 119.850 ;
        RECT 35.770 119.990 36.060 120.035 ;
        RECT 38.550 119.990 38.840 120.035 ;
        RECT 40.410 119.990 40.700 120.035 ;
        RECT 51.440 119.990 51.760 120.050 ;
        RECT 60.610 119.990 60.900 120.035 ;
        RECT 63.390 119.990 63.680 120.035 ;
        RECT 65.250 119.990 65.540 120.035 ;
        RECT 35.770 119.850 40.700 119.990 ;
        RECT 35.770 119.805 36.060 119.850 ;
        RECT 38.550 119.805 38.840 119.850 ;
        RECT 40.410 119.805 40.700 119.850 ;
        RECT 50.610 119.850 60.410 119.990 ;
        RECT 26.230 119.510 28.210 119.650 ;
        RECT 26.230 119.355 26.370 119.510 ;
        RECT 28.440 119.450 28.760 119.710 ;
        RECT 31.660 119.695 31.980 119.710 ;
        RECT 31.660 119.650 32.195 119.695 ;
        RECT 28.990 119.510 32.195 119.650 ;
        RECT 23.855 119.310 24.145 119.355 ;
        RECT 15.575 119.170 18.320 119.310 ;
        RECT 22.090 119.170 24.145 119.310 ;
        RECT 15.575 119.125 15.865 119.170 ;
        RECT 16.940 119.110 17.260 119.170 ;
        RECT 18.180 118.970 18.320 119.170 ;
        RECT 23.855 119.125 24.145 119.170 ;
        RECT 24.775 119.310 25.065 119.355 ;
        RECT 26.155 119.310 26.445 119.355 ;
        RECT 24.775 119.170 26.445 119.310 ;
        RECT 24.775 119.125 25.065 119.170 ;
        RECT 26.155 119.125 26.445 119.170 ;
        RECT 27.060 119.310 27.380 119.370 ;
        RECT 28.990 119.355 29.130 119.510 ;
        RECT 31.660 119.465 32.195 119.510 ;
        RECT 31.660 119.450 31.980 119.465 ;
        RECT 39.020 119.450 39.340 119.710 ;
        RECT 28.915 119.310 29.205 119.355 ;
        RECT 27.060 119.170 29.205 119.310 ;
        RECT 24.850 118.970 24.990 119.125 ;
        RECT 27.060 119.110 27.380 119.170 ;
        RECT 28.915 119.125 29.205 119.170 ;
        RECT 35.770 119.310 36.060 119.355 ;
        RECT 40.875 119.310 41.165 119.355 ;
        RECT 41.320 119.310 41.640 119.370 ;
        RECT 50.610 119.355 50.750 119.850 ;
        RECT 51.440 119.790 51.760 119.850 ;
        RECT 51.915 119.650 52.205 119.695 ;
        RECT 53.740 119.650 54.060 119.710 ;
        RECT 56.040 119.650 56.360 119.710 ;
        RECT 51.915 119.510 56.360 119.650 ;
        RECT 60.270 119.650 60.410 119.850 ;
        RECT 60.610 119.850 65.540 119.990 ;
        RECT 60.610 119.805 60.900 119.850 ;
        RECT 63.390 119.805 63.680 119.850 ;
        RECT 65.250 119.805 65.540 119.850 ;
        RECT 61.100 119.650 61.420 119.710 ;
        RECT 60.270 119.510 61.420 119.650 ;
        RECT 51.915 119.465 52.205 119.510 ;
        RECT 53.740 119.450 54.060 119.510 ;
        RECT 56.040 119.450 56.360 119.510 ;
        RECT 61.100 119.450 61.420 119.510 ;
        RECT 63.860 119.450 64.180 119.710 ;
        RECT 70.850 119.695 70.990 120.190 ;
        RECT 71.680 120.130 72.000 120.190 ;
        RECT 73.535 119.990 73.825 120.035 ;
        RECT 74.900 119.990 75.220 120.050 ;
        RECT 73.535 119.850 75.220 119.990 ;
        RECT 73.535 119.805 73.825 119.850 ;
        RECT 74.900 119.790 75.220 119.850 ;
        RECT 70.775 119.465 71.065 119.695 ;
        RECT 71.235 119.650 71.525 119.695 ;
        RECT 75.360 119.650 75.680 119.710 ;
        RECT 75.910 119.695 76.050 120.190 ;
        RECT 77.200 120.190 79.805 120.330 ;
        RECT 77.200 120.130 77.520 120.190 ;
        RECT 79.515 120.145 79.805 120.190 ;
        RECT 82.505 120.330 82.795 120.375 ;
        RECT 84.100 120.330 84.420 120.390 ;
        RECT 94.680 120.330 95.000 120.390 ;
        RECT 96.075 120.330 96.365 120.375 ;
        RECT 101.120 120.330 101.440 120.390 ;
        RECT 82.505 120.190 84.420 120.330 ;
        RECT 82.505 120.145 82.795 120.190 ;
        RECT 84.100 120.130 84.420 120.190 ;
        RECT 86.030 120.190 92.150 120.330 ;
        RECT 80.420 119.990 80.740 120.050 ;
        RECT 84.560 119.990 84.880 120.050 ;
        RECT 80.420 119.850 84.880 119.990 ;
        RECT 80.420 119.790 80.740 119.850 ;
        RECT 84.560 119.790 84.880 119.850 ;
        RECT 71.235 119.510 75.680 119.650 ;
        RECT 71.235 119.465 71.525 119.510 ;
        RECT 75.360 119.450 75.680 119.510 ;
        RECT 75.835 119.650 76.125 119.695 ;
        RECT 86.030 119.650 86.170 120.190 ;
        RECT 86.370 119.990 86.660 120.035 ;
        RECT 89.150 119.990 89.440 120.035 ;
        RECT 91.010 119.990 91.300 120.035 ;
        RECT 86.370 119.850 91.300 119.990 ;
        RECT 92.010 119.990 92.150 120.190 ;
        RECT 94.680 120.190 96.365 120.330 ;
        RECT 94.680 120.130 95.000 120.190 ;
        RECT 96.075 120.145 96.365 120.190 ;
        RECT 99.830 120.190 101.440 120.330 ;
        RECT 99.830 119.990 99.970 120.190 ;
        RECT 101.120 120.130 101.440 120.190 ;
        RECT 92.010 119.850 99.970 119.990 ;
        RECT 86.370 119.805 86.660 119.850 ;
        RECT 89.150 119.805 89.440 119.850 ;
        RECT 91.010 119.805 91.300 119.850 ;
        RECT 75.835 119.510 86.170 119.650 ;
        RECT 88.700 119.650 89.020 119.710 ;
        RECT 89.635 119.650 89.925 119.695 ;
        RECT 88.700 119.510 89.925 119.650 ;
        RECT 75.835 119.465 76.125 119.510 ;
        RECT 88.700 119.450 89.020 119.510 ;
        RECT 89.635 119.465 89.925 119.510 ;
        RECT 91.475 119.650 91.765 119.695 ;
        RECT 91.920 119.650 92.240 119.710 ;
        RECT 92.470 119.695 92.610 119.850 ;
        RECT 100.215 119.805 100.505 120.035 ;
        RECT 91.475 119.510 92.240 119.650 ;
        RECT 91.475 119.465 91.765 119.510 ;
        RECT 91.920 119.450 92.240 119.510 ;
        RECT 92.395 119.465 92.685 119.695 ;
        RECT 94.220 119.650 94.540 119.710 ;
        RECT 96.060 119.650 96.380 119.710 ;
        RECT 94.220 119.510 97.670 119.650 ;
        RECT 94.220 119.450 94.540 119.510 ;
        RECT 96.060 119.450 96.380 119.510 ;
        RECT 35.770 119.170 38.305 119.310 ;
        RECT 35.770 119.125 36.060 119.170 ;
        RECT 38.090 119.015 38.305 119.170 ;
        RECT 40.875 119.170 41.640 119.310 ;
        RECT 40.875 119.125 41.165 119.170 ;
        RECT 41.320 119.110 41.640 119.170 ;
        RECT 50.535 119.125 50.825 119.355 ;
        RECT 52.835 119.310 53.125 119.355 ;
        RECT 53.280 119.310 53.600 119.370 ;
        RECT 56.745 119.310 57.035 119.355 ;
        RECT 52.835 119.170 57.035 119.310 ;
        RECT 52.835 119.125 53.125 119.170 ;
        RECT 53.280 119.110 53.600 119.170 ;
        RECT 56.745 119.125 57.035 119.170 ;
        RECT 60.610 119.310 60.900 119.355 ;
        RECT 65.240 119.310 65.560 119.370 ;
        RECT 65.715 119.310 66.005 119.355 ;
        RECT 60.610 119.170 63.145 119.310 ;
        RECT 60.610 119.125 60.900 119.170 ;
        RECT 18.180 118.830 24.990 118.970 ;
        RECT 26.615 118.970 26.905 119.015 ;
        RECT 33.910 118.970 34.200 119.015 ;
        RECT 37.170 118.970 37.460 119.015 ;
        RECT 26.615 118.830 37.460 118.970 ;
        RECT 26.615 118.785 26.905 118.830 ;
        RECT 33.910 118.785 34.200 118.830 ;
        RECT 37.170 118.785 37.460 118.830 ;
        RECT 38.090 118.970 38.380 119.015 ;
        RECT 39.950 118.970 40.240 119.015 ;
        RECT 38.090 118.830 40.240 118.970 ;
        RECT 38.090 118.785 38.380 118.830 ;
        RECT 39.950 118.785 40.240 118.830 ;
        RECT 46.840 118.970 47.160 119.030 ;
        RECT 51.440 118.970 51.760 119.030 ;
        RECT 52.375 118.970 52.665 119.015 ;
        RECT 46.840 118.830 52.665 118.970 ;
        RECT 46.840 118.770 47.160 118.830 ;
        RECT 51.440 118.770 51.760 118.830 ;
        RECT 52.375 118.785 52.665 118.830 ;
        RECT 58.750 118.970 59.040 119.015 ;
        RECT 60.180 118.970 60.500 119.030 ;
        RECT 62.930 119.015 63.145 119.170 ;
        RECT 65.240 119.170 66.005 119.310 ;
        RECT 65.240 119.110 65.560 119.170 ;
        RECT 65.715 119.125 66.005 119.170 ;
        RECT 67.080 119.310 67.400 119.370 ;
        RECT 68.475 119.310 68.765 119.355 ;
        RECT 67.080 119.170 68.765 119.310 ;
        RECT 67.080 119.110 67.400 119.170 ;
        RECT 68.475 119.125 68.765 119.170 ;
        RECT 71.695 119.310 71.985 119.355 ;
        RECT 72.600 119.310 72.920 119.370 ;
        RECT 76.295 119.310 76.585 119.355 ;
        RECT 79.975 119.310 80.265 119.355 ;
        RECT 80.420 119.310 80.740 119.370 ;
        RECT 71.695 119.170 76.585 119.310 ;
        RECT 71.695 119.125 71.985 119.170 ;
        RECT 62.010 118.970 62.300 119.015 ;
        RECT 58.750 118.830 62.300 118.970 ;
        RECT 58.750 118.785 59.040 118.830 ;
        RECT 60.180 118.770 60.500 118.830 ;
        RECT 62.010 118.785 62.300 118.830 ;
        RECT 62.930 118.970 63.220 119.015 ;
        RECT 64.790 118.970 65.080 119.015 ;
        RECT 62.930 118.830 65.080 118.970 ;
        RECT 68.550 118.970 68.690 119.125 ;
        RECT 72.600 119.110 72.920 119.170 ;
        RECT 76.295 119.125 76.585 119.170 ;
        RECT 77.290 119.170 80.740 119.310 ;
        RECT 68.550 118.830 74.670 118.970 ;
        RECT 62.930 118.785 63.220 118.830 ;
        RECT 64.790 118.785 65.080 118.830 ;
        RECT 17.400 118.430 17.720 118.690 ;
        RECT 17.860 118.630 18.180 118.690 ;
        RECT 20.175 118.630 20.465 118.675 ;
        RECT 27.520 118.630 27.840 118.690 ;
        RECT 17.860 118.490 27.840 118.630 ;
        RECT 17.860 118.430 18.180 118.490 ;
        RECT 20.175 118.445 20.465 118.490 ;
        RECT 27.520 118.430 27.840 118.490 ;
        RECT 28.900 118.630 29.220 118.690 ;
        RECT 29.375 118.630 29.665 118.675 ;
        RECT 28.900 118.490 29.665 118.630 ;
        RECT 28.900 118.430 29.220 118.490 ;
        RECT 29.375 118.445 29.665 118.490 ;
        RECT 31.200 118.430 31.520 118.690 ;
        RECT 50.060 118.430 50.380 118.690 ;
        RECT 54.675 118.630 54.965 118.675 ;
        RECT 56.040 118.630 56.360 118.690 ;
        RECT 54.675 118.490 56.360 118.630 ;
        RECT 54.675 118.445 54.965 118.490 ;
        RECT 56.040 118.430 56.360 118.490 ;
        RECT 68.935 118.630 69.225 118.675 ;
        RECT 73.980 118.630 74.300 118.690 ;
        RECT 68.935 118.490 74.300 118.630 ;
        RECT 74.530 118.630 74.670 118.830 ;
        RECT 76.740 118.770 77.060 119.030 ;
        RECT 77.290 118.630 77.430 119.170 ;
        RECT 79.975 119.125 80.265 119.170 ;
        RECT 80.420 119.110 80.740 119.170 ;
        RECT 81.340 119.110 81.660 119.370 ;
        RECT 86.370 119.310 86.660 119.355 ;
        RECT 86.370 119.170 88.905 119.310 ;
        RECT 86.370 119.125 86.660 119.170 ;
        RECT 77.660 118.970 77.980 119.030 ;
        RECT 80.895 118.970 81.185 119.015 ;
        RECT 77.660 118.830 81.185 118.970 ;
        RECT 77.660 118.770 77.980 118.830 ;
        RECT 80.895 118.785 81.185 118.830 ;
        RECT 84.510 118.970 84.800 119.015 ;
        RECT 85.940 118.970 86.260 119.030 ;
        RECT 88.690 119.015 88.905 119.170 ;
        RECT 93.760 119.110 94.080 119.370 ;
        RECT 96.995 119.310 97.285 119.355 ;
        RECT 95.690 119.170 97.285 119.310 ;
        RECT 87.770 118.970 88.060 119.015 ;
        RECT 84.510 118.830 88.060 118.970 ;
        RECT 84.510 118.785 84.800 118.830 ;
        RECT 85.940 118.770 86.260 118.830 ;
        RECT 87.770 118.785 88.060 118.830 ;
        RECT 88.690 118.970 88.980 119.015 ;
        RECT 90.550 118.970 90.840 119.015 ;
        RECT 88.690 118.830 90.840 118.970 ;
        RECT 88.690 118.785 88.980 118.830 ;
        RECT 90.550 118.785 90.840 118.830 ;
        RECT 74.530 118.490 77.430 118.630 ;
        RECT 78.120 118.630 78.440 118.690 ;
        RECT 78.595 118.630 78.885 118.675 ;
        RECT 78.120 118.490 78.885 118.630 ;
        RECT 68.935 118.445 69.225 118.490 ;
        RECT 73.980 118.430 74.300 118.490 ;
        RECT 78.120 118.430 78.440 118.490 ;
        RECT 78.595 118.445 78.885 118.490 ;
        RECT 93.315 118.630 93.605 118.675 ;
        RECT 94.220 118.630 94.540 118.690 ;
        RECT 95.690 118.675 95.830 119.170 ;
        RECT 96.995 119.125 97.285 119.170 ;
        RECT 97.530 118.970 97.670 119.510 ;
        RECT 99.295 119.310 99.585 119.355 ;
        RECT 100.290 119.310 100.430 119.805 ;
        RECT 101.210 119.650 101.350 120.130 ;
        RECT 104.340 119.990 104.660 120.050 ;
        RECT 116.300 119.990 116.620 120.050 ;
        RECT 104.340 119.850 116.620 119.990 ;
        RECT 104.340 119.790 104.660 119.850 ;
        RECT 116.300 119.790 116.620 119.850 ;
        RECT 117.190 119.990 117.480 120.035 ;
        RECT 119.970 119.990 120.260 120.035 ;
        RECT 121.830 119.990 122.120 120.035 ;
        RECT 117.190 119.850 122.120 119.990 ;
        RECT 117.190 119.805 117.480 119.850 ;
        RECT 119.970 119.805 120.260 119.850 ;
        RECT 121.830 119.805 122.120 119.850 ;
        RECT 102.975 119.650 103.265 119.695 ;
        RECT 106.180 119.650 106.500 119.710 ;
        RECT 101.210 119.510 106.500 119.650 ;
        RECT 102.975 119.465 103.265 119.510 ;
        RECT 106.180 119.450 106.500 119.510 ;
        RECT 107.115 119.650 107.405 119.695 ;
        RECT 108.480 119.650 108.800 119.710 ;
        RECT 113.540 119.695 113.860 119.710 ;
        RECT 113.325 119.650 113.860 119.695 ;
        RECT 107.115 119.510 113.860 119.650 ;
        RECT 107.115 119.465 107.405 119.510 ;
        RECT 108.480 119.450 108.800 119.510 ;
        RECT 113.325 119.465 113.860 119.510 ;
        RECT 113.540 119.450 113.860 119.465 ;
        RECT 99.295 119.170 100.430 119.310 ;
        RECT 99.295 119.125 99.585 119.170 ;
        RECT 104.340 119.110 104.660 119.370 ;
        RECT 107.560 119.110 107.880 119.370 ;
        RECT 117.190 119.310 117.480 119.355 ;
        RECT 117.190 119.170 119.725 119.310 ;
        RECT 117.190 119.125 117.480 119.170 ;
        RECT 102.055 118.970 102.345 119.015 ;
        RECT 97.530 118.830 102.345 118.970 ;
        RECT 102.055 118.785 102.345 118.830 ;
        RECT 102.500 118.970 102.820 119.030 ;
        RECT 107.650 118.970 107.790 119.110 ;
        RECT 102.500 118.830 107.790 118.970 ;
        RECT 115.330 118.970 115.620 119.015 ;
        RECT 116.760 118.970 117.080 119.030 ;
        RECT 119.510 119.015 119.725 119.170 ;
        RECT 120.440 119.110 120.760 119.370 ;
        RECT 121.820 119.310 122.140 119.370 ;
        RECT 122.295 119.310 122.585 119.355 ;
        RECT 123.660 119.310 123.980 119.370 ;
        RECT 121.820 119.170 123.980 119.310 ;
        RECT 121.820 119.110 122.140 119.170 ;
        RECT 122.295 119.125 122.585 119.170 ;
        RECT 123.660 119.110 123.980 119.170 ;
        RECT 118.590 118.970 118.880 119.015 ;
        RECT 115.330 118.830 118.880 118.970 ;
        RECT 102.500 118.770 102.820 118.830 ;
        RECT 115.330 118.785 115.620 118.830 ;
        RECT 116.760 118.770 117.080 118.830 ;
        RECT 118.590 118.785 118.880 118.830 ;
        RECT 119.510 118.970 119.800 119.015 ;
        RECT 121.370 118.970 121.660 119.015 ;
        RECT 119.510 118.830 121.660 118.970 ;
        RECT 119.510 118.785 119.800 118.830 ;
        RECT 121.370 118.785 121.660 118.830 ;
        RECT 93.315 118.490 94.540 118.630 ;
        RECT 93.315 118.445 93.605 118.490 ;
        RECT 94.220 118.430 94.540 118.490 ;
        RECT 95.615 118.445 95.905 118.675 ;
        RECT 98.360 118.430 98.680 118.690 ;
        RECT 104.800 118.430 105.120 118.690 ;
        RECT 109.415 118.630 109.705 118.675 ;
        RECT 111.700 118.630 112.020 118.690 ;
        RECT 109.415 118.490 112.020 118.630 ;
        RECT 109.415 118.445 109.705 118.490 ;
        RECT 111.700 118.430 112.020 118.490 ;
        RECT 11.010 117.810 125.890 118.290 ;
        RECT 16.265 117.610 16.555 117.655 ;
        RECT 20.160 117.610 20.480 117.670 ;
        RECT 16.265 117.470 20.480 117.610 ;
        RECT 16.265 117.425 16.555 117.470 ;
        RECT 20.160 117.410 20.480 117.470 ;
        RECT 30.740 117.410 31.060 117.670 ;
        RECT 34.895 117.610 35.185 117.655 ;
        RECT 38.560 117.610 38.880 117.670 ;
        RECT 34.895 117.470 38.880 117.610 ;
        RECT 34.895 117.425 35.185 117.470 ;
        RECT 38.560 117.410 38.880 117.470 ;
        RECT 46.840 117.610 47.160 117.670 ;
        RECT 48.005 117.610 48.295 117.655 ;
        RECT 46.840 117.470 48.295 117.610 ;
        RECT 46.840 117.410 47.160 117.470 ;
        RECT 48.005 117.425 48.295 117.470 ;
        RECT 52.820 117.610 53.140 117.670 ;
        RECT 52.820 117.470 56.730 117.610 ;
        RECT 52.820 117.410 53.140 117.470 ;
        RECT 17.400 117.270 17.720 117.330 ;
        RECT 18.270 117.270 18.560 117.315 ;
        RECT 21.530 117.270 21.820 117.315 ;
        RECT 17.400 117.130 21.820 117.270 ;
        RECT 17.400 117.070 17.720 117.130 ;
        RECT 18.270 117.085 18.560 117.130 ;
        RECT 21.530 117.085 21.820 117.130 ;
        RECT 22.450 117.270 22.740 117.315 ;
        RECT 24.310 117.270 24.600 117.315 ;
        RECT 22.450 117.130 24.600 117.270 ;
        RECT 22.450 117.085 22.740 117.130 ;
        RECT 24.310 117.085 24.600 117.130 ;
        RECT 31.660 117.270 31.980 117.330 ;
        RECT 50.060 117.315 50.380 117.330 ;
        RECT 33.055 117.270 33.345 117.315 ;
        RECT 31.660 117.130 33.345 117.270 ;
        RECT 20.130 116.930 20.420 116.975 ;
        RECT 22.450 116.930 22.665 117.085 ;
        RECT 31.660 117.070 31.980 117.130 ;
        RECT 33.055 117.085 33.345 117.130 ;
        RECT 50.010 117.270 50.380 117.315 ;
        RECT 53.270 117.270 53.560 117.315 ;
        RECT 50.010 117.130 53.560 117.270 ;
        RECT 50.010 117.085 50.380 117.130 ;
        RECT 53.270 117.085 53.560 117.130 ;
        RECT 54.190 117.270 54.480 117.315 ;
        RECT 56.050 117.270 56.340 117.315 ;
        RECT 54.190 117.130 56.340 117.270 ;
        RECT 56.590 117.270 56.730 117.470 ;
        RECT 60.180 117.410 60.500 117.670 ;
        RECT 62.940 117.410 63.260 117.670 ;
        RECT 72.140 117.610 72.460 117.670 ;
        RECT 77.660 117.610 77.980 117.670 ;
        RECT 72.140 117.470 77.980 117.610 ;
        RECT 72.140 117.410 72.460 117.470 ;
        RECT 77.660 117.410 77.980 117.470 ;
        RECT 79.040 117.610 79.360 117.670 ;
        RECT 81.355 117.610 81.645 117.655 ;
        RECT 79.040 117.470 81.645 117.610 ;
        RECT 79.040 117.410 79.360 117.470 ;
        RECT 81.355 117.425 81.645 117.470 ;
        RECT 86.415 117.610 86.705 117.655 ;
        RECT 88.700 117.610 89.020 117.670 ;
        RECT 86.415 117.470 89.020 117.610 ;
        RECT 86.415 117.425 86.705 117.470 ;
        RECT 88.700 117.410 89.020 117.470 ;
        RECT 89.175 117.610 89.465 117.655 ;
        RECT 89.620 117.610 89.940 117.670 ;
        RECT 89.175 117.470 89.940 117.610 ;
        RECT 89.175 117.425 89.465 117.470 ;
        RECT 89.620 117.410 89.940 117.470 ;
        RECT 90.785 117.610 91.075 117.655 ;
        RECT 94.220 117.610 94.540 117.670 ;
        RECT 90.785 117.470 94.540 117.610 ;
        RECT 90.785 117.425 91.075 117.470 ;
        RECT 94.220 117.410 94.540 117.470 ;
        RECT 101.365 117.610 101.655 117.655 ;
        RECT 102.500 117.610 102.820 117.670 ;
        RECT 101.365 117.470 102.820 117.610 ;
        RECT 101.365 117.425 101.655 117.470 ;
        RECT 102.500 117.410 102.820 117.470 ;
        RECT 110.795 117.425 111.085 117.655 ;
        RECT 73.980 117.315 74.300 117.330 ;
        RECT 63.415 117.270 63.705 117.315 ;
        RECT 56.590 117.130 63.705 117.270 ;
        RECT 54.190 117.085 54.480 117.130 ;
        RECT 56.050 117.085 56.340 117.130 ;
        RECT 63.415 117.085 63.705 117.130 ;
        RECT 73.930 117.270 74.300 117.315 ;
        RECT 77.190 117.270 77.480 117.315 ;
        RECT 73.930 117.130 77.480 117.270 ;
        RECT 73.930 117.085 74.300 117.130 ;
        RECT 77.190 117.085 77.480 117.130 ;
        RECT 78.110 117.270 78.400 117.315 ;
        RECT 79.970 117.270 80.260 117.315 ;
        RECT 78.110 117.130 80.260 117.270 ;
        RECT 78.110 117.085 78.400 117.130 ;
        RECT 79.970 117.085 80.260 117.130 ;
        RECT 84.560 117.270 84.880 117.330 ;
        RECT 87.795 117.270 88.085 117.315 ;
        RECT 92.790 117.270 93.080 117.315 ;
        RECT 96.050 117.270 96.340 117.315 ;
        RECT 84.560 117.130 87.550 117.270 ;
        RECT 50.060 117.070 50.380 117.085 ;
        RECT 20.130 116.790 22.665 116.930 ;
        RECT 20.130 116.745 20.420 116.790 ;
        RECT 23.380 116.730 23.700 116.990 ;
        RECT 29.835 116.930 30.125 116.975 ;
        RECT 31.200 116.930 31.520 116.990 ;
        RECT 32.595 116.930 32.885 116.975 ;
        RECT 41.780 116.930 42.100 116.990 ;
        RECT 29.835 116.790 31.520 116.930 ;
        RECT 29.835 116.745 30.125 116.790 ;
        RECT 31.200 116.730 31.520 116.790 ;
        RECT 31.750 116.790 42.100 116.930 ;
        RECT 25.235 116.590 25.525 116.635 ;
        RECT 27.060 116.590 27.380 116.650 ;
        RECT 25.235 116.450 27.380 116.590 ;
        RECT 25.235 116.405 25.525 116.450 ;
        RECT 27.060 116.390 27.380 116.450 ;
        RECT 27.520 116.590 27.840 116.650 ;
        RECT 31.750 116.590 31.890 116.790 ;
        RECT 32.595 116.745 32.885 116.790 ;
        RECT 41.780 116.730 42.100 116.790 ;
        RECT 47.315 116.930 47.605 116.975 ;
        RECT 47.760 116.930 48.080 116.990 ;
        RECT 47.315 116.790 48.080 116.930 ;
        RECT 47.315 116.745 47.605 116.790 ;
        RECT 47.760 116.730 48.080 116.790 ;
        RECT 51.870 116.930 52.160 116.975 ;
        RECT 54.190 116.930 54.405 117.085 ;
        RECT 73.980 117.070 74.300 117.085 ;
        RECT 51.870 116.790 54.405 116.930 ;
        RECT 55.135 116.930 55.425 116.975 ;
        RECT 55.580 116.930 55.900 116.990 ;
        RECT 55.135 116.790 55.900 116.930 ;
        RECT 51.870 116.745 52.160 116.790 ;
        RECT 55.135 116.745 55.425 116.790 ;
        RECT 55.580 116.730 55.900 116.790 ;
        RECT 59.735 116.930 60.025 116.975 ;
        RECT 61.100 116.930 61.420 116.990 ;
        RECT 65.240 116.930 65.560 116.990 ;
        RECT 59.735 116.790 61.420 116.930 ;
        RECT 59.735 116.745 60.025 116.790 ;
        RECT 61.100 116.730 61.420 116.790 ;
        RECT 62.110 116.790 65.560 116.930 ;
        RECT 27.520 116.450 31.890 116.590 ;
        RECT 27.520 116.390 27.840 116.450 ;
        RECT 32.135 116.405 32.425 116.635 ;
        RECT 52.360 116.590 52.680 116.650 ;
        RECT 56.975 116.590 57.265 116.635 ;
        RECT 62.110 116.590 62.250 116.790 ;
        RECT 65.240 116.730 65.560 116.790 ;
        RECT 65.715 116.745 66.005 116.975 ;
        RECT 75.790 116.930 76.080 116.975 ;
        RECT 78.110 116.930 78.325 117.085 ;
        RECT 84.560 117.070 84.880 117.130 ;
        RECT 82.275 116.930 82.565 116.975 ;
        RECT 75.790 116.790 78.325 116.930 ;
        RECT 78.670 116.790 82.565 116.930 ;
        RECT 75.790 116.745 76.080 116.790 ;
        RECT 52.360 116.450 62.250 116.590 ;
        RECT 20.130 116.250 20.420 116.295 ;
        RECT 22.910 116.250 23.200 116.295 ;
        RECT 24.770 116.250 25.060 116.295 ;
        RECT 20.130 116.110 25.060 116.250 ;
        RECT 20.130 116.065 20.420 116.110 ;
        RECT 22.910 116.065 23.200 116.110 ;
        RECT 24.770 116.065 25.060 116.110 ;
        RECT 28.440 116.250 28.760 116.310 ;
        RECT 32.210 116.250 32.350 116.405 ;
        RECT 52.360 116.390 52.680 116.450 ;
        RECT 56.975 116.405 57.265 116.450 ;
        RECT 62.495 116.405 62.785 116.635 ;
        RECT 65.790 116.590 65.930 116.745 ;
        RECT 65.330 116.450 65.930 116.590 ;
        RECT 71.925 116.590 72.215 116.635 ;
        RECT 73.520 116.590 73.840 116.650 ;
        RECT 71.925 116.450 73.840 116.590 ;
        RECT 28.440 116.110 32.350 116.250 ;
        RECT 51.870 116.250 52.160 116.295 ;
        RECT 54.650 116.250 54.940 116.295 ;
        RECT 56.510 116.250 56.800 116.295 ;
        RECT 51.870 116.110 56.800 116.250 ;
        RECT 28.440 116.050 28.760 116.110 ;
        RECT 51.870 116.065 52.160 116.110 ;
        RECT 54.650 116.065 54.940 116.110 ;
        RECT 56.510 116.065 56.800 116.110 ;
        RECT 46.380 115.710 46.700 115.970 ;
        RECT 53.280 115.910 53.600 115.970 ;
        RECT 62.570 115.910 62.710 116.405 ;
        RECT 65.330 116.295 65.470 116.450 ;
        RECT 71.925 116.405 72.215 116.450 ;
        RECT 73.520 116.390 73.840 116.450 ;
        RECT 74.900 116.590 75.220 116.650 ;
        RECT 78.670 116.590 78.810 116.790 ;
        RECT 82.275 116.745 82.565 116.790 ;
        RECT 85.480 116.730 85.800 116.990 ;
        RECT 87.410 116.975 87.550 117.130 ;
        RECT 87.795 117.130 96.340 117.270 ;
        RECT 87.795 117.085 88.085 117.130 ;
        RECT 92.790 117.085 93.080 117.130 ;
        RECT 96.050 117.085 96.340 117.130 ;
        RECT 96.970 117.270 97.260 117.315 ;
        RECT 98.830 117.270 99.120 117.315 ;
        RECT 96.970 117.130 99.120 117.270 ;
        RECT 96.970 117.085 97.260 117.130 ;
        RECT 98.830 117.085 99.120 117.130 ;
        RECT 103.370 117.270 103.660 117.315 ;
        RECT 104.800 117.270 105.120 117.330 ;
        RECT 106.630 117.270 106.920 117.315 ;
        RECT 103.370 117.130 106.920 117.270 ;
        RECT 103.370 117.085 103.660 117.130 ;
        RECT 87.335 116.930 87.625 116.975 ;
        RECT 88.715 116.930 89.005 116.975 ;
        RECT 87.335 116.790 89.005 116.930 ;
        RECT 87.335 116.745 87.625 116.790 ;
        RECT 88.715 116.745 89.005 116.790 ;
        RECT 94.650 116.930 94.940 116.975 ;
        RECT 96.970 116.930 97.185 117.085 ;
        RECT 104.800 117.070 105.120 117.130 ;
        RECT 106.630 117.085 106.920 117.130 ;
        RECT 107.550 117.270 107.840 117.315 ;
        RECT 109.410 117.270 109.700 117.315 ;
        RECT 107.550 117.130 109.700 117.270 ;
        RECT 107.550 117.085 107.840 117.130 ;
        RECT 109.410 117.085 109.700 117.130 ;
        RECT 94.650 116.790 97.185 116.930 ;
        RECT 97.915 116.930 98.205 116.975 ;
        RECT 98.360 116.930 98.680 116.990 ;
        RECT 97.915 116.790 98.680 116.930 ;
        RECT 94.650 116.745 94.940 116.790 ;
        RECT 97.915 116.745 98.205 116.790 ;
        RECT 98.360 116.730 98.680 116.790 ;
        RECT 105.230 116.930 105.520 116.975 ;
        RECT 107.550 116.930 107.765 117.085 ;
        RECT 105.230 116.790 107.765 116.930 ;
        RECT 105.230 116.745 105.520 116.790 ;
        RECT 108.020 116.730 108.340 116.990 ;
        RECT 108.495 116.930 108.785 116.975 ;
        RECT 110.870 116.930 111.010 117.425 ;
        RECT 116.760 117.410 117.080 117.670 ;
        RECT 119.075 117.610 119.365 117.655 ;
        RECT 120.440 117.610 120.760 117.670 ;
        RECT 119.075 117.470 120.760 117.610 ;
        RECT 119.075 117.425 119.365 117.470 ;
        RECT 120.440 117.410 120.760 117.470 ;
        RECT 108.495 116.790 111.010 116.930 ;
        RECT 108.495 116.745 108.785 116.790 ;
        RECT 111.700 116.730 112.020 116.990 ;
        RECT 116.300 116.730 116.620 116.990 ;
        RECT 118.140 116.730 118.460 116.990 ;
        RECT 74.900 116.450 78.810 116.590 ;
        RECT 74.900 116.390 75.220 116.450 ;
        RECT 79.040 116.390 79.360 116.650 ;
        RECT 80.895 116.590 81.185 116.635 ;
        RECT 91.920 116.590 92.240 116.650 ;
        RECT 99.755 116.590 100.045 116.635 ;
        RECT 80.895 116.450 100.045 116.590 ;
        RECT 108.110 116.590 108.250 116.730 ;
        RECT 110.320 116.590 110.640 116.650 ;
        RECT 108.110 116.450 110.640 116.590 ;
        RECT 80.895 116.405 81.185 116.450 ;
        RECT 91.920 116.390 92.240 116.450 ;
        RECT 99.755 116.405 100.045 116.450 ;
        RECT 110.320 116.390 110.640 116.450 ;
        RECT 65.255 116.065 65.545 116.295 ;
        RECT 75.790 116.250 76.080 116.295 ;
        RECT 78.570 116.250 78.860 116.295 ;
        RECT 80.430 116.250 80.720 116.295 ;
        RECT 75.790 116.110 80.720 116.250 ;
        RECT 75.790 116.065 76.080 116.110 ;
        RECT 78.570 116.065 78.860 116.110 ;
        RECT 80.430 116.065 80.720 116.110 ;
        RECT 94.650 116.250 94.940 116.295 ;
        RECT 97.430 116.250 97.720 116.295 ;
        RECT 99.290 116.250 99.580 116.295 ;
        RECT 94.650 116.110 99.580 116.250 ;
        RECT 94.650 116.065 94.940 116.110 ;
        RECT 97.430 116.065 97.720 116.110 ;
        RECT 99.290 116.065 99.580 116.110 ;
        RECT 105.230 116.250 105.520 116.295 ;
        RECT 108.010 116.250 108.300 116.295 ;
        RECT 109.870 116.250 110.160 116.295 ;
        RECT 105.230 116.110 110.160 116.250 ;
        RECT 105.230 116.065 105.520 116.110 ;
        RECT 108.010 116.065 108.300 116.110 ;
        RECT 109.870 116.065 110.160 116.110 ;
        RECT 53.280 115.770 62.710 115.910 ;
        RECT 66.635 115.910 66.925 115.955 ;
        RECT 68.000 115.910 68.320 115.970 ;
        RECT 66.635 115.770 68.320 115.910 ;
        RECT 53.280 115.710 53.600 115.770 ;
        RECT 66.635 115.725 66.925 115.770 ;
        RECT 68.000 115.710 68.320 115.770 ;
        RECT 11.810 115.090 125.890 115.570 ;
        RECT 47.760 114.890 48.080 114.950 ;
        RECT 49.615 114.890 49.905 114.935 ;
        RECT 47.760 114.750 49.905 114.890 ;
        RECT 47.760 114.690 48.080 114.750 ;
        RECT 49.615 114.705 49.905 114.750 ;
        RECT 55.135 114.890 55.425 114.935 ;
        RECT 55.580 114.890 55.900 114.950 ;
        RECT 55.135 114.750 55.900 114.890 ;
        RECT 55.135 114.705 55.425 114.750 ;
        RECT 55.580 114.690 55.900 114.750 ;
        RECT 60.885 114.890 61.175 114.935 ;
        RECT 62.940 114.890 63.260 114.950 ;
        RECT 60.885 114.750 63.260 114.890 ;
        RECT 60.885 114.705 61.175 114.750 ;
        RECT 62.940 114.690 63.260 114.750 ;
        RECT 79.040 114.690 79.360 114.950 ;
        RECT 64.750 114.550 65.040 114.595 ;
        RECT 67.530 114.550 67.820 114.595 ;
        RECT 69.390 114.550 69.680 114.595 ;
        RECT 64.750 114.410 69.680 114.550 ;
        RECT 64.750 114.365 65.040 114.410 ;
        RECT 67.530 114.365 67.820 114.410 ;
        RECT 69.390 114.365 69.680 114.410 ;
        RECT 81.340 114.550 81.660 114.610 ;
        RECT 123.215 114.550 123.505 114.595 ;
        RECT 81.340 114.410 123.505 114.550 ;
        RECT 81.340 114.350 81.660 114.410 ;
        RECT 123.215 114.365 123.505 114.410 ;
        RECT 52.835 114.210 53.125 114.255 ;
        RECT 53.280 114.210 53.600 114.270 ;
        RECT 52.835 114.070 53.600 114.210 ;
        RECT 52.835 114.025 53.125 114.070 ;
        RECT 53.280 114.010 53.600 114.070 ;
        RECT 65.240 114.210 65.560 114.270 ;
        RECT 65.240 114.070 67.770 114.210 ;
        RECT 65.240 114.010 65.560 114.070 ;
        RECT 24.300 113.870 24.620 113.930 ;
        RECT 24.775 113.870 25.065 113.915 ;
        RECT 24.300 113.730 25.065 113.870 ;
        RECT 24.300 113.670 24.620 113.730 ;
        RECT 24.775 113.685 25.065 113.730 ;
        RECT 46.855 113.685 47.145 113.915 ;
        RECT 38.560 113.530 38.880 113.590 ;
        RECT 46.930 113.530 47.070 113.685 ;
        RECT 51.440 113.670 51.760 113.930 ;
        RECT 54.215 113.870 54.505 113.915 ;
        RECT 56.040 113.870 56.360 113.930 ;
        RECT 54.215 113.730 56.360 113.870 ;
        RECT 54.215 113.685 54.505 113.730 ;
        RECT 56.040 113.670 56.360 113.730 ;
        RECT 64.750 113.870 65.040 113.915 ;
        RECT 67.630 113.870 67.770 114.070 ;
        RECT 68.000 114.010 68.320 114.270 ;
        RECT 69.855 113.870 70.145 113.915 ;
        RECT 64.750 113.730 67.285 113.870 ;
        RECT 67.630 113.730 70.145 113.870 ;
        RECT 64.750 113.685 65.040 113.730 ;
        RECT 51.915 113.530 52.205 113.575 ;
        RECT 52.820 113.530 53.140 113.590 ;
        RECT 38.560 113.390 48.910 113.530 ;
        RECT 38.560 113.330 38.880 113.390 ;
        RECT 25.695 113.190 25.985 113.235 ;
        RECT 31.660 113.190 31.980 113.250 ;
        RECT 25.695 113.050 31.980 113.190 ;
        RECT 25.695 113.005 25.985 113.050 ;
        RECT 31.660 112.990 31.980 113.050 ;
        RECT 47.315 113.190 47.605 113.235 ;
        RECT 48.220 113.190 48.540 113.250 ;
        RECT 47.315 113.050 48.540 113.190 ;
        RECT 48.770 113.190 48.910 113.390 ;
        RECT 51.915 113.390 53.140 113.530 ;
        RECT 51.915 113.345 52.205 113.390 ;
        RECT 52.820 113.330 53.140 113.390 ;
        RECT 62.890 113.530 63.180 113.575 ;
        RECT 64.320 113.530 64.640 113.590 ;
        RECT 67.070 113.575 67.285 113.730 ;
        RECT 69.855 113.685 70.145 113.730 ;
        RECT 78.120 113.670 78.440 113.930 ;
        RECT 114.920 113.870 115.240 113.930 ;
        RECT 116.315 113.870 116.605 113.915 ;
        RECT 114.920 113.730 116.605 113.870 ;
        RECT 114.920 113.670 115.240 113.730 ;
        RECT 116.315 113.685 116.605 113.730 ;
        RECT 117.220 113.870 117.540 113.930 ;
        RECT 118.615 113.870 118.905 113.915 ;
        RECT 117.220 113.730 118.905 113.870 ;
        RECT 117.220 113.670 117.540 113.730 ;
        RECT 118.615 113.685 118.905 113.730 ;
        RECT 119.060 113.670 119.380 113.930 ;
        RECT 124.120 113.670 124.440 113.930 ;
        RECT 66.150 113.530 66.440 113.575 ;
        RECT 62.890 113.390 66.440 113.530 ;
        RECT 62.890 113.345 63.180 113.390 ;
        RECT 64.320 113.330 64.640 113.390 ;
        RECT 66.150 113.345 66.440 113.390 ;
        RECT 67.070 113.530 67.360 113.575 ;
        RECT 68.930 113.530 69.220 113.575 ;
        RECT 67.070 113.390 69.220 113.530 ;
        RECT 67.070 113.345 67.360 113.390 ;
        RECT 68.930 113.345 69.220 113.390 ;
        RECT 116.760 113.330 117.080 113.590 ;
        RECT 64.780 113.190 65.100 113.250 ;
        RECT 48.770 113.050 65.100 113.190 ;
        RECT 47.315 113.005 47.605 113.050 ;
        RECT 48.220 112.990 48.540 113.050 ;
        RECT 64.780 112.990 65.100 113.050 ;
        RECT 115.380 113.190 115.700 113.250 ;
        RECT 117.695 113.190 117.985 113.235 ;
        RECT 115.380 113.050 117.985 113.190 ;
        RECT 115.380 112.990 115.700 113.050 ;
        RECT 117.695 113.005 117.985 113.050 ;
        RECT 119.980 112.990 120.300 113.250 ;
        RECT 11.010 112.370 125.890 112.850 ;
        RECT 28.915 111.985 29.205 112.215 ;
        RECT 37.640 112.170 37.960 112.230 ;
        RECT 50.520 112.170 50.840 112.230 ;
        RECT 31.290 112.030 37.410 112.170 ;
        RECT 19.815 111.830 20.105 111.875 ;
        RECT 22.000 111.830 22.320 111.890 ;
        RECT 23.055 111.830 23.705 111.875 ;
        RECT 19.815 111.690 23.705 111.830 ;
        RECT 19.815 111.645 20.405 111.690 ;
        RECT 20.115 111.330 20.405 111.645 ;
        RECT 22.000 111.630 22.320 111.690 ;
        RECT 23.055 111.645 23.705 111.690 ;
        RECT 25.695 111.830 25.985 111.875 ;
        RECT 28.990 111.830 29.130 111.985 ;
        RECT 25.695 111.690 29.130 111.830 ;
        RECT 29.360 111.830 29.680 111.890 ;
        RECT 31.290 111.830 31.430 112.030 ;
        RECT 37.270 111.890 37.410 112.030 ;
        RECT 37.640 112.030 50.840 112.170 ;
        RECT 37.640 111.970 37.960 112.030 ;
        RECT 50.520 111.970 50.840 112.030 ;
        RECT 52.820 112.170 53.140 112.230 ;
        RECT 53.525 112.170 53.815 112.215 ;
        RECT 52.820 112.030 53.815 112.170 ;
        RECT 52.820 111.970 53.140 112.030 ;
        RECT 53.525 111.985 53.815 112.030 ;
        RECT 64.320 112.170 64.640 112.230 ;
        RECT 64.795 112.170 65.085 112.215 ;
        RECT 64.320 112.030 65.085 112.170 ;
        RECT 64.320 111.970 64.640 112.030 ;
        RECT 64.795 111.985 65.085 112.030 ;
        RECT 29.360 111.690 31.430 111.830 ;
        RECT 25.695 111.645 25.985 111.690 ;
        RECT 29.360 111.630 29.680 111.690 ;
        RECT 21.195 111.490 21.485 111.535 ;
        RECT 24.775 111.490 25.065 111.535 ;
        RECT 26.610 111.490 26.900 111.535 ;
        RECT 21.195 111.350 26.900 111.490 ;
        RECT 21.195 111.305 21.485 111.350 ;
        RECT 24.775 111.305 25.065 111.350 ;
        RECT 26.610 111.305 26.900 111.350 ;
        RECT 29.835 111.490 30.125 111.535 ;
        RECT 30.280 111.490 30.600 111.550 ;
        RECT 31.290 111.535 31.430 111.690 ;
        RECT 37.180 111.830 37.500 111.890 ;
        RECT 48.220 111.875 48.540 111.890 ;
        RECT 45.480 111.830 45.770 111.875 ;
        RECT 47.340 111.830 47.630 111.875 ;
        RECT 37.180 111.690 39.710 111.830 ;
        RECT 37.180 111.630 37.500 111.690 ;
        RECT 29.835 111.350 30.600 111.490 ;
        RECT 29.835 111.305 30.125 111.350 ;
        RECT 30.280 111.290 30.600 111.350 ;
        RECT 31.215 111.305 31.505 111.535 ;
        RECT 33.040 111.490 33.360 111.550 ;
        RECT 33.515 111.490 33.805 111.535 ;
        RECT 33.040 111.350 33.805 111.490 ;
        RECT 33.040 111.290 33.360 111.350 ;
        RECT 33.515 111.305 33.805 111.350 ;
        RECT 33.960 111.290 34.280 111.550 ;
        RECT 38.560 111.290 38.880 111.550 ;
        RECT 39.570 111.535 39.710 111.690 ;
        RECT 45.480 111.690 47.630 111.830 ;
        RECT 45.480 111.645 45.770 111.690 ;
        RECT 47.340 111.645 47.630 111.690 ;
        RECT 39.495 111.305 39.785 111.535 ;
        RECT 41.795 111.490 42.085 111.535 ;
        RECT 42.240 111.490 42.560 111.550 ;
        RECT 41.795 111.350 42.560 111.490 ;
        RECT 41.795 111.305 42.085 111.350 ;
        RECT 42.240 111.290 42.560 111.350 ;
        RECT 42.700 111.290 43.020 111.550 ;
        RECT 46.380 111.290 46.700 111.550 ;
        RECT 47.415 111.490 47.630 111.645 ;
        RECT 48.220 111.830 48.550 111.875 ;
        RECT 51.520 111.830 51.810 111.875 ;
        RECT 100.200 111.830 100.520 111.890 ;
        RECT 114.920 111.830 115.240 111.890 ;
        RECT 48.220 111.690 51.810 111.830 ;
        RECT 48.220 111.645 48.550 111.690 ;
        RECT 51.520 111.645 51.810 111.690 ;
        RECT 66.480 111.690 76.050 111.830 ;
        RECT 48.220 111.630 48.540 111.645 ;
        RECT 49.660 111.490 49.950 111.535 ;
        RECT 47.415 111.350 49.950 111.490 ;
        RECT 49.660 111.305 49.950 111.350 ;
        RECT 59.720 111.490 60.040 111.550 ;
        RECT 61.575 111.490 61.865 111.535 ;
        RECT 59.720 111.350 61.865 111.490 ;
        RECT 59.720 111.290 60.040 111.350 ;
        RECT 61.575 111.305 61.865 111.350 ;
        RECT 64.780 111.490 65.100 111.550 ;
        RECT 65.255 111.490 65.545 111.535 ;
        RECT 66.480 111.490 66.620 111.690 ;
        RECT 64.780 111.350 66.620 111.490 ;
        RECT 64.780 111.290 65.100 111.350 ;
        RECT 65.255 111.305 65.545 111.350 ;
        RECT 74.440 111.290 74.760 111.550 ;
        RECT 75.910 111.535 76.050 111.690 ;
        RECT 100.200 111.690 106.870 111.830 ;
        RECT 100.200 111.630 100.520 111.690 ;
        RECT 75.835 111.305 76.125 111.535 ;
        RECT 95.140 111.490 95.460 111.550 ;
        RECT 97.455 111.490 97.745 111.535 ;
        RECT 95.140 111.350 97.745 111.490 ;
        RECT 95.140 111.290 95.460 111.350 ;
        RECT 97.455 111.305 97.745 111.350 ;
        RECT 101.120 111.490 101.440 111.550 ;
        RECT 101.595 111.490 101.885 111.535 ;
        RECT 101.120 111.350 101.885 111.490 ;
        RECT 101.120 111.290 101.440 111.350 ;
        RECT 101.595 111.305 101.885 111.350 ;
        RECT 16.940 110.950 17.260 111.210 ;
        RECT 27.060 111.150 27.380 111.210 ;
        RECT 39.020 111.150 39.340 111.210 ;
        RECT 41.320 111.150 41.640 111.210 ;
        RECT 44.555 111.150 44.845 111.195 ;
        RECT 27.060 111.010 44.845 111.150 ;
        RECT 27.060 110.950 27.380 111.010 ;
        RECT 39.020 110.950 39.340 111.010 ;
        RECT 41.320 110.950 41.640 111.010 ;
        RECT 44.555 110.965 44.845 111.010 ;
        RECT 77.200 110.950 77.520 111.210 ;
        RECT 101.670 111.150 101.810 111.305 ;
        RECT 103.880 111.290 104.200 111.550 ;
        RECT 106.730 111.535 106.870 111.690 ;
        RECT 111.330 111.690 115.240 111.830 ;
        RECT 111.330 111.535 111.470 111.690 ;
        RECT 114.920 111.630 115.240 111.690 ;
        RECT 115.380 111.630 115.700 111.890 ;
        RECT 116.760 111.830 117.080 111.890 ;
        RECT 117.675 111.830 118.325 111.875 ;
        RECT 121.275 111.830 121.565 111.875 ;
        RECT 116.760 111.690 121.565 111.830 ;
        RECT 116.760 111.630 117.080 111.690 ;
        RECT 117.675 111.645 118.325 111.690 ;
        RECT 120.975 111.645 121.565 111.690 ;
        RECT 106.195 111.305 106.485 111.535 ;
        RECT 106.655 111.305 106.945 111.535 ;
        RECT 111.255 111.305 111.545 111.535 ;
        RECT 114.480 111.490 114.770 111.535 ;
        RECT 116.315 111.490 116.605 111.535 ;
        RECT 119.895 111.490 120.185 111.535 ;
        RECT 114.480 111.350 120.185 111.490 ;
        RECT 114.480 111.305 114.770 111.350 ;
        RECT 116.315 111.305 116.605 111.350 ;
        RECT 119.895 111.305 120.185 111.350 ;
        RECT 120.975 111.330 121.265 111.645 ;
        RECT 106.270 111.150 106.410 111.305 ;
        RECT 111.330 111.150 111.470 111.305 ;
        RECT 101.670 111.010 111.470 111.150 ;
        RECT 114.015 110.965 114.305 111.195 ;
        RECT 21.195 110.810 21.485 110.855 ;
        RECT 24.315 110.810 24.605 110.855 ;
        RECT 26.205 110.810 26.495 110.855 ;
        RECT 21.195 110.670 26.495 110.810 ;
        RECT 21.195 110.625 21.485 110.670 ;
        RECT 24.315 110.625 24.605 110.670 ;
        RECT 26.205 110.625 26.495 110.670 ;
        RECT 38.560 110.810 38.880 110.870 ;
        RECT 40.875 110.810 41.165 110.855 ;
        RECT 38.560 110.670 41.165 110.810 ;
        RECT 38.560 110.610 38.880 110.670 ;
        RECT 40.875 110.625 41.165 110.670 ;
        RECT 45.020 110.810 45.310 110.855 ;
        RECT 46.880 110.810 47.170 110.855 ;
        RECT 49.660 110.810 49.950 110.855 ;
        RECT 45.020 110.670 49.950 110.810 ;
        RECT 45.020 110.625 45.310 110.670 ;
        RECT 46.880 110.625 47.170 110.670 ;
        RECT 49.660 110.625 49.950 110.670 ;
        RECT 110.320 110.810 110.640 110.870 ;
        RECT 114.090 110.810 114.230 110.965 ;
        RECT 124.120 110.950 124.440 111.210 ;
        RECT 110.320 110.670 114.230 110.810 ;
        RECT 114.885 110.810 115.175 110.855 ;
        RECT 116.775 110.810 117.065 110.855 ;
        RECT 119.895 110.810 120.185 110.855 ;
        RECT 114.885 110.670 120.185 110.810 ;
        RECT 110.320 110.610 110.640 110.670 ;
        RECT 114.885 110.625 115.175 110.670 ;
        RECT 116.775 110.625 117.065 110.670 ;
        RECT 119.895 110.625 120.185 110.670 ;
        RECT 30.740 110.270 31.060 110.530 ;
        RECT 31.200 110.470 31.520 110.530 ;
        RECT 32.595 110.470 32.885 110.515 ;
        RECT 31.200 110.330 32.885 110.470 ;
        RECT 31.200 110.270 31.520 110.330 ;
        RECT 32.595 110.285 32.885 110.330 ;
        RECT 34.420 110.470 34.740 110.530 ;
        RECT 34.895 110.470 35.185 110.515 ;
        RECT 34.420 110.330 35.185 110.470 ;
        RECT 34.420 110.270 34.740 110.330 ;
        RECT 34.895 110.285 35.185 110.330 ;
        RECT 39.940 110.270 40.260 110.530 ;
        RECT 43.635 110.470 43.925 110.515 ;
        RECT 44.540 110.470 44.860 110.530 ;
        RECT 43.635 110.330 44.860 110.470 ;
        RECT 43.635 110.285 43.925 110.330 ;
        RECT 44.540 110.270 44.860 110.330 ;
        RECT 62.480 110.270 62.800 110.530 ;
        RECT 75.360 110.270 75.680 110.530 ;
        RECT 97.900 110.470 98.220 110.530 ;
        RECT 98.375 110.470 98.665 110.515 ;
        RECT 97.900 110.330 98.665 110.470 ;
        RECT 97.900 110.270 98.220 110.330 ;
        RECT 98.375 110.285 98.665 110.330 ;
        RECT 101.580 110.470 101.900 110.530 ;
        RECT 102.055 110.470 102.345 110.515 ;
        RECT 101.580 110.330 102.345 110.470 ;
        RECT 101.580 110.270 101.900 110.330 ;
        RECT 102.055 110.285 102.345 110.330 ;
        RECT 104.815 110.470 105.105 110.515 ;
        RECT 105.260 110.470 105.580 110.530 ;
        RECT 104.815 110.330 105.580 110.470 ;
        RECT 104.815 110.285 105.105 110.330 ;
        RECT 105.260 110.270 105.580 110.330 ;
        RECT 105.720 110.270 106.040 110.530 ;
        RECT 107.560 110.270 107.880 110.530 ;
        RECT 111.715 110.470 112.005 110.515 ;
        RECT 115.380 110.470 115.700 110.530 ;
        RECT 111.715 110.330 115.700 110.470 ;
        RECT 111.715 110.285 112.005 110.330 ;
        RECT 115.380 110.270 115.700 110.330 ;
        RECT 11.810 109.650 125.890 110.130 ;
        RECT 21.555 109.450 21.845 109.495 ;
        RECT 22.000 109.450 22.320 109.510 ;
        RECT 29.360 109.450 29.680 109.510 ;
        RECT 21.555 109.310 22.320 109.450 ;
        RECT 21.555 109.265 21.845 109.310 ;
        RECT 22.000 109.250 22.320 109.310 ;
        RECT 25.310 109.310 29.680 109.450 ;
        RECT 25.310 108.770 25.450 109.310 ;
        RECT 29.360 109.250 29.680 109.310 ;
        RECT 42.700 109.450 43.020 109.510 ;
        RECT 47.775 109.450 48.065 109.495 ;
        RECT 42.700 109.310 48.065 109.450 ;
        RECT 42.700 109.250 43.020 109.310 ;
        RECT 47.775 109.265 48.065 109.310 ;
        RECT 48.680 109.450 49.000 109.510 ;
        RECT 91.920 109.450 92.240 109.510 ;
        RECT 112.175 109.450 112.465 109.495 ;
        RECT 122.280 109.450 122.600 109.510 ;
        RECT 48.680 109.310 67.310 109.450 ;
        RECT 48.680 109.250 49.000 109.310 ;
        RECT 29.935 109.110 30.225 109.155 ;
        RECT 33.055 109.110 33.345 109.155 ;
        RECT 34.945 109.110 35.235 109.155 ;
        RECT 39.020 109.110 39.340 109.170 ;
        RECT 29.935 108.970 35.235 109.110 ;
        RECT 29.935 108.925 30.225 108.970 ;
        RECT 33.055 108.925 33.345 108.970 ;
        RECT 34.945 108.925 35.235 108.970 ;
        RECT 35.890 108.970 39.340 109.110 ;
        RECT 22.090 108.630 25.450 108.770 ;
        RECT 19.240 108.230 19.560 108.490 ;
        RECT 22.090 108.475 22.230 108.630 ;
        RECT 19.715 108.430 20.005 108.475 ;
        RECT 22.015 108.430 22.305 108.475 ;
        RECT 19.715 108.290 22.305 108.430 ;
        RECT 19.715 108.245 20.005 108.290 ;
        RECT 22.015 108.245 22.305 108.290 ;
        RECT 22.460 108.430 22.780 108.490 ;
        RECT 25.310 108.475 25.450 108.630 ;
        RECT 25.695 108.770 25.985 108.815 ;
        RECT 29.360 108.770 29.680 108.830 ;
        RECT 25.695 108.630 29.680 108.770 ;
        RECT 25.695 108.585 25.985 108.630 ;
        RECT 29.360 108.570 29.680 108.630 ;
        RECT 34.420 108.570 34.740 108.830 ;
        RECT 35.890 108.815 36.030 108.970 ;
        RECT 39.020 108.910 39.340 108.970 ;
        RECT 40.515 109.110 40.805 109.155 ;
        RECT 43.635 109.110 43.925 109.155 ;
        RECT 45.525 109.110 45.815 109.155 ;
        RECT 40.515 108.970 45.815 109.110 ;
        RECT 40.515 108.925 40.805 108.970 ;
        RECT 43.635 108.925 43.925 108.970 ;
        RECT 45.525 108.925 45.815 108.970 ;
        RECT 60.755 109.110 61.045 109.155 ;
        RECT 63.875 109.110 64.165 109.155 ;
        RECT 65.765 109.110 66.055 109.155 ;
        RECT 60.755 108.970 66.055 109.110 ;
        RECT 60.755 108.925 61.045 108.970 ;
        RECT 63.875 108.925 64.165 108.970 ;
        RECT 65.765 108.925 66.055 108.970 ;
        RECT 35.815 108.585 36.105 108.815 ;
        RECT 36.275 108.770 36.565 108.815 ;
        RECT 41.780 108.770 42.100 108.830 ;
        RECT 36.275 108.630 42.100 108.770 ;
        RECT 36.275 108.585 36.565 108.630 ;
        RECT 41.780 108.570 42.100 108.630 ;
        RECT 44.540 108.770 44.860 108.830 ;
        RECT 45.015 108.770 45.305 108.815 ;
        RECT 44.540 108.630 45.305 108.770 ;
        RECT 44.540 108.570 44.860 108.630 ;
        RECT 45.015 108.585 45.305 108.630 ;
        RECT 46.395 108.770 46.685 108.815 ;
        RECT 51.900 108.770 52.220 108.830 ;
        RECT 46.395 108.630 52.220 108.770 ;
        RECT 46.395 108.585 46.685 108.630 ;
        RECT 51.900 108.570 52.220 108.630 ;
        RECT 56.515 108.770 56.805 108.815 ;
        RECT 59.260 108.770 59.580 108.830 ;
        RECT 56.515 108.630 59.580 108.770 ;
        RECT 56.515 108.585 56.805 108.630 ;
        RECT 59.260 108.570 59.580 108.630 ;
        RECT 62.480 108.770 62.800 108.830 ;
        RECT 65.255 108.770 65.545 108.815 ;
        RECT 62.480 108.630 65.545 108.770 ;
        RECT 62.480 108.570 62.800 108.630 ;
        RECT 65.255 108.585 65.545 108.630 ;
        RECT 66.620 108.570 66.940 108.830 ;
        RECT 24.775 108.430 25.065 108.475 ;
        RECT 22.460 108.290 25.065 108.430 ;
        RECT 22.460 108.230 22.780 108.290 ;
        RECT 24.775 108.245 25.065 108.290 ;
        RECT 25.235 108.245 25.525 108.475 ;
        RECT 28.855 108.135 29.145 108.450 ;
        RECT 29.935 108.430 30.225 108.475 ;
        RECT 33.515 108.430 33.805 108.475 ;
        RECT 35.350 108.430 35.640 108.475 ;
        RECT 29.935 108.290 35.640 108.430 ;
        RECT 29.935 108.245 30.225 108.290 ;
        RECT 33.515 108.245 33.805 108.290 ;
        RECT 35.350 108.245 35.640 108.290 ;
        RECT 28.555 108.090 29.145 108.135 ;
        RECT 30.740 108.090 31.060 108.150 ;
        RECT 39.435 108.135 39.725 108.450 ;
        RECT 40.515 108.430 40.805 108.475 ;
        RECT 44.095 108.430 44.385 108.475 ;
        RECT 45.930 108.430 46.220 108.475 ;
        RECT 40.515 108.290 46.220 108.430 ;
        RECT 40.515 108.245 40.805 108.290 ;
        RECT 44.095 108.245 44.385 108.290 ;
        RECT 45.930 108.245 46.220 108.290 ;
        RECT 46.840 108.230 47.160 108.490 ;
        RECT 50.520 108.230 50.840 108.490 ;
        RECT 55.135 108.360 55.425 108.475 ;
        RECT 55.025 108.245 55.425 108.360 ;
        RECT 55.025 108.220 55.350 108.245 ;
        RECT 55.580 108.230 55.900 108.490 ;
        RECT 67.170 108.475 67.310 109.310 ;
        RECT 91.920 109.310 99.050 109.450 ;
        RECT 91.920 109.250 92.240 109.310 ;
        RECT 77.660 109.110 77.980 109.170 ;
        RECT 74.530 108.970 77.980 109.110 ;
        RECT 74.530 108.815 74.670 108.970 ;
        RECT 77.660 108.910 77.980 108.970 ;
        RECT 78.695 109.110 78.985 109.155 ;
        RECT 81.815 109.110 82.105 109.155 ;
        RECT 83.705 109.110 83.995 109.155 ;
        RECT 87.320 109.110 87.640 109.170 ;
        RECT 92.010 109.110 92.150 109.250 ;
        RECT 78.695 108.970 83.995 109.110 ;
        RECT 78.695 108.925 78.985 108.970 ;
        RECT 81.815 108.925 82.105 108.970 ;
        RECT 83.705 108.925 83.995 108.970 ;
        RECT 84.650 108.970 92.150 109.110 ;
        RECT 93.415 109.110 93.705 109.155 ;
        RECT 96.535 109.110 96.825 109.155 ;
        RECT 98.425 109.110 98.715 109.155 ;
        RECT 93.415 108.970 98.715 109.110 ;
        RECT 74.455 108.585 74.745 108.815 ;
        RECT 75.360 108.770 75.680 108.830 ;
        RECT 84.650 108.815 84.790 108.970 ;
        RECT 87.320 108.910 87.640 108.970 ;
        RECT 93.415 108.925 93.705 108.970 ;
        RECT 96.535 108.925 96.825 108.970 ;
        RECT 98.425 108.925 98.715 108.970 ;
        RECT 83.195 108.770 83.485 108.815 ;
        RECT 75.360 108.630 83.485 108.770 ;
        RECT 75.360 108.570 75.680 108.630 ;
        RECT 83.195 108.585 83.485 108.630 ;
        RECT 84.575 108.585 84.865 108.815 ;
        RECT 89.175 108.770 89.465 108.815 ;
        RECT 95.600 108.770 95.920 108.830 ;
        RECT 89.175 108.630 95.920 108.770 ;
        RECT 89.175 108.585 89.465 108.630 ;
        RECT 95.600 108.570 95.920 108.630 ;
        RECT 97.900 108.570 98.220 108.830 ;
        RECT 98.910 108.770 99.050 109.310 ;
        RECT 112.175 109.310 122.600 109.450 ;
        RECT 112.175 109.265 112.465 109.310 ;
        RECT 122.280 109.250 122.600 109.310 ;
        RECT 104.915 109.110 105.205 109.155 ;
        RECT 108.035 109.110 108.325 109.155 ;
        RECT 109.925 109.110 110.215 109.155 ;
        RECT 104.915 108.970 110.215 109.110 ;
        RECT 104.915 108.925 105.205 108.970 ;
        RECT 108.035 108.925 108.325 108.970 ;
        RECT 109.925 108.925 110.215 108.970 ;
        RECT 117.795 109.110 118.085 109.155 ;
        RECT 120.915 109.110 121.205 109.155 ;
        RECT 122.805 109.110 123.095 109.155 ;
        RECT 117.795 108.970 123.095 109.110 ;
        RECT 117.795 108.925 118.085 108.970 ;
        RECT 120.915 108.925 121.205 108.970 ;
        RECT 122.805 108.925 123.095 108.970 ;
        RECT 99.295 108.770 99.585 108.815 ;
        RECT 98.910 108.630 99.585 108.770 ;
        RECT 99.295 108.585 99.585 108.630 ;
        RECT 100.675 108.770 100.965 108.815 ;
        RECT 107.100 108.770 107.420 108.830 ;
        RECT 100.675 108.630 107.420 108.770 ;
        RECT 100.675 108.585 100.965 108.630 ;
        RECT 107.100 108.570 107.420 108.630 ;
        RECT 107.560 108.770 107.880 108.830 ;
        RECT 109.415 108.770 109.705 108.815 ;
        RECT 107.560 108.630 109.705 108.770 ;
        RECT 107.560 108.570 107.880 108.630 ;
        RECT 109.415 108.585 109.705 108.630 ;
        RECT 113.555 108.770 113.845 108.815 ;
        RECT 118.600 108.770 118.920 108.830 ;
        RECT 113.555 108.630 118.920 108.770 ;
        RECT 113.555 108.585 113.845 108.630 ;
        RECT 118.600 108.570 118.920 108.630 ;
        RECT 119.980 108.770 120.300 108.830 ;
        RECT 122.295 108.770 122.585 108.815 ;
        RECT 119.980 108.630 122.585 108.770 ;
        RECT 119.980 108.570 120.300 108.630 ;
        RECT 122.295 108.585 122.585 108.630 ;
        RECT 123.660 108.570 123.980 108.830 ;
        RECT 31.795 108.090 32.445 108.135 ;
        RECT 28.555 107.950 32.445 108.090 ;
        RECT 28.555 107.905 28.845 107.950 ;
        RECT 30.740 107.890 31.060 107.950 ;
        RECT 31.795 107.905 32.445 107.950 ;
        RECT 39.135 108.090 39.725 108.135 ;
        RECT 39.940 108.090 40.260 108.150 ;
        RECT 42.375 108.090 43.025 108.135 ;
        RECT 39.135 107.950 43.025 108.090 ;
        RECT 55.210 108.090 55.350 108.220 ;
        RECT 56.040 108.090 56.360 108.150 ;
        RECT 59.675 108.135 59.965 108.450 ;
        RECT 60.755 108.430 61.045 108.475 ;
        RECT 64.335 108.430 64.625 108.475 ;
        RECT 66.170 108.430 66.460 108.475 ;
        RECT 60.755 108.290 66.460 108.430 ;
        RECT 60.755 108.245 61.045 108.290 ;
        RECT 64.335 108.245 64.625 108.290 ;
        RECT 66.170 108.245 66.460 108.290 ;
        RECT 67.095 108.245 67.385 108.475 ;
        RECT 72.600 108.230 72.920 108.490 ;
        RECT 55.210 107.950 56.360 108.090 ;
        RECT 39.135 107.905 39.425 107.950 ;
        RECT 39.940 107.890 40.260 107.950 ;
        RECT 42.375 107.905 43.025 107.950 ;
        RECT 56.040 107.890 56.360 107.950 ;
        RECT 59.375 108.090 59.965 108.135 ;
        RECT 60.180 108.090 60.500 108.150 ;
        RECT 62.615 108.090 63.265 108.135 ;
        RECT 59.375 107.950 63.265 108.090 ;
        RECT 59.375 107.905 59.665 107.950 ;
        RECT 60.180 107.890 60.500 107.950 ;
        RECT 62.615 107.905 63.265 107.950 ;
        RECT 73.060 108.090 73.380 108.150 ;
        RECT 77.615 108.135 77.905 108.450 ;
        RECT 78.695 108.430 78.985 108.475 ;
        RECT 82.275 108.430 82.565 108.475 ;
        RECT 84.110 108.430 84.400 108.475 ;
        RECT 78.695 108.290 84.400 108.430 ;
        RECT 78.695 108.245 78.985 108.290 ;
        RECT 82.275 108.245 82.565 108.290 ;
        RECT 84.110 108.245 84.400 108.290 ;
        RECT 85.020 108.430 85.340 108.490 ;
        RECT 85.955 108.430 86.245 108.475 ;
        RECT 85.020 108.290 86.245 108.430 ;
        RECT 85.020 108.230 85.340 108.290 ;
        RECT 85.955 108.245 86.245 108.290 ;
        RECT 87.780 108.230 88.100 108.490 ;
        RECT 92.335 108.135 92.625 108.450 ;
        RECT 93.415 108.430 93.705 108.475 ;
        RECT 96.995 108.430 97.285 108.475 ;
        RECT 98.830 108.430 99.120 108.475 ;
        RECT 93.415 108.290 99.120 108.430 ;
        RECT 93.415 108.245 93.705 108.290 ;
        RECT 96.995 108.245 97.285 108.290 ;
        RECT 98.830 108.245 99.120 108.290 ;
        RECT 77.315 108.090 77.905 108.135 ;
        RECT 80.555 108.090 81.205 108.135 ;
        RECT 73.060 107.950 81.205 108.090 ;
        RECT 73.060 107.890 73.380 107.950 ;
        RECT 77.315 107.905 77.605 107.950 ;
        RECT 80.555 107.905 81.205 107.950 ;
        RECT 92.035 108.090 92.625 108.135 ;
        RECT 95.140 108.135 95.460 108.150 ;
        RECT 103.835 108.135 104.125 108.450 ;
        RECT 104.915 108.430 105.205 108.475 ;
        RECT 108.495 108.430 108.785 108.475 ;
        RECT 110.330 108.430 110.620 108.475 ;
        RECT 104.915 108.290 110.620 108.430 ;
        RECT 104.915 108.245 105.205 108.290 ;
        RECT 108.495 108.245 108.785 108.290 ;
        RECT 110.330 108.245 110.620 108.290 ;
        RECT 110.780 108.230 111.100 108.490 ;
        RECT 111.255 108.245 111.545 108.475 ;
        RECT 95.140 108.090 95.925 108.135 ;
        RECT 92.035 107.950 95.925 108.090 ;
        RECT 92.035 107.905 92.325 107.950 ;
        RECT 95.140 107.905 95.925 107.950 ;
        RECT 103.535 108.090 104.125 108.135 ;
        RECT 105.720 108.090 106.040 108.150 ;
        RECT 106.775 108.090 107.425 108.135 ;
        RECT 103.535 107.950 107.425 108.090 ;
        RECT 103.535 107.905 103.825 107.950 ;
        RECT 95.140 107.890 95.460 107.905 ;
        RECT 105.720 107.890 106.040 107.950 ;
        RECT 106.775 107.905 107.425 107.950 ;
        RECT 51.440 107.550 51.760 107.810 ;
        RECT 68.015 107.750 68.305 107.795 ;
        RECT 70.300 107.750 70.620 107.810 ;
        RECT 68.015 107.610 70.620 107.750 ;
        RECT 68.015 107.565 68.305 107.610 ;
        RECT 70.300 107.550 70.620 107.610 ;
        RECT 73.535 107.750 73.825 107.795 ;
        RECT 79.500 107.750 79.820 107.810 ;
        RECT 73.535 107.610 79.820 107.750 ;
        RECT 73.535 107.565 73.825 107.610 ;
        RECT 79.500 107.550 79.820 107.610 ;
        RECT 85.020 107.550 85.340 107.810 ;
        RECT 88.700 107.550 89.020 107.810 ;
        RECT 100.660 107.750 100.980 107.810 ;
        RECT 111.330 107.750 111.470 108.245 ;
        RECT 116.715 108.135 117.005 108.450 ;
        RECT 117.795 108.430 118.085 108.475 ;
        RECT 121.375 108.430 121.665 108.475 ;
        RECT 123.210 108.430 123.500 108.475 ;
        RECT 117.795 108.290 123.500 108.430 ;
        RECT 117.795 108.245 118.085 108.290 ;
        RECT 121.375 108.245 121.665 108.290 ;
        RECT 123.210 108.245 123.500 108.290 ;
        RECT 116.415 108.090 117.005 108.135 ;
        RECT 117.220 108.090 117.540 108.150 ;
        RECT 119.655 108.090 120.305 108.135 ;
        RECT 116.415 107.950 120.305 108.090 ;
        RECT 116.415 107.905 116.705 107.950 ;
        RECT 117.220 107.890 117.540 107.950 ;
        RECT 119.655 107.905 120.305 107.950 ;
        RECT 100.660 107.610 111.470 107.750 ;
        RECT 100.660 107.550 100.980 107.610 ;
        RECT 11.010 106.930 125.890 107.410 ;
        RECT 31.200 106.730 31.520 106.790 ;
        RECT 23.010 106.590 31.520 106.730 ;
        RECT 17.055 106.390 17.345 106.435 ;
        RECT 20.295 106.390 20.945 106.435 ;
        RECT 22.460 106.390 22.780 106.450 ;
        RECT 23.010 106.435 23.150 106.590 ;
        RECT 31.200 106.530 31.520 106.590 ;
        RECT 66.160 106.730 66.480 106.790 ;
        RECT 77.200 106.730 77.520 106.790 ;
        RECT 85.955 106.730 86.245 106.775 ;
        RECT 66.160 106.590 71.910 106.730 ;
        RECT 66.160 106.530 66.480 106.590 ;
        RECT 17.055 106.250 22.780 106.390 ;
        RECT 17.055 106.205 17.645 106.250 ;
        RECT 20.295 106.205 20.945 106.250 ;
        RECT 17.355 105.890 17.645 106.205 ;
        RECT 22.460 106.190 22.780 106.250 ;
        RECT 22.935 106.205 23.225 106.435 ;
        RECT 28.435 106.390 29.085 106.435 ;
        RECT 32.035 106.390 32.325 106.435 ;
        RECT 36.735 106.390 37.025 106.435 ;
        RECT 28.435 106.250 37.025 106.390 ;
        RECT 28.435 106.205 29.085 106.250 ;
        RECT 31.735 106.205 32.325 106.250 ;
        RECT 36.735 106.205 37.025 106.250 ;
        RECT 41.335 106.390 41.625 106.435 ;
        RECT 42.700 106.390 43.020 106.450 ;
        RECT 41.335 106.250 43.020 106.390 ;
        RECT 41.335 106.205 41.625 106.250 ;
        RECT 18.435 106.050 18.725 106.095 ;
        RECT 22.015 106.050 22.305 106.095 ;
        RECT 23.850 106.050 24.140 106.095 ;
        RECT 18.435 105.910 24.140 106.050 ;
        RECT 18.435 105.865 18.725 105.910 ;
        RECT 22.015 105.865 22.305 105.910 ;
        RECT 23.850 105.865 24.140 105.910 ;
        RECT 25.240 106.050 25.530 106.095 ;
        RECT 27.075 106.050 27.365 106.095 ;
        RECT 30.655 106.050 30.945 106.095 ;
        RECT 25.240 105.910 30.945 106.050 ;
        RECT 25.240 105.865 25.530 105.910 ;
        RECT 27.075 105.865 27.365 105.910 ;
        RECT 30.655 105.865 30.945 105.910 ;
        RECT 31.735 105.890 32.025 106.205 ;
        RECT 42.700 106.190 43.020 106.250 ;
        RECT 43.615 106.390 44.265 106.435 ;
        RECT 47.215 106.390 47.505 106.435 ;
        RECT 43.615 106.250 47.505 106.390 ;
        RECT 43.615 106.205 44.265 106.250 ;
        RECT 46.915 106.205 47.505 106.250 ;
        RECT 51.440 106.390 51.760 106.450 ;
        RECT 51.915 106.390 52.205 106.435 ;
        RECT 51.440 106.250 52.205 106.390 ;
        RECT 46.915 106.110 47.205 106.205 ;
        RECT 51.440 106.190 51.760 106.250 ;
        RECT 51.915 106.205 52.205 106.250 ;
        RECT 54.195 106.390 54.845 106.435 ;
        RECT 55.580 106.390 55.900 106.450 ;
        RECT 57.795 106.390 58.085 106.435 ;
        RECT 54.195 106.250 58.085 106.390 ;
        RECT 54.195 106.205 54.845 106.250 ;
        RECT 55.580 106.190 55.900 106.250 ;
        RECT 57.495 106.205 58.085 106.250 ;
        RECT 62.480 106.390 62.800 106.450 ;
        RECT 64.435 106.390 64.725 106.435 ;
        RECT 67.675 106.390 68.325 106.435 ;
        RECT 62.480 106.250 68.325 106.390 ;
        RECT 37.180 105.850 37.500 106.110 ;
        RECT 39.020 106.050 39.340 106.110 ;
        RECT 39.955 106.050 40.245 106.095 ;
        RECT 39.020 105.910 40.245 106.050 ;
        RECT 39.020 105.850 39.340 105.910 ;
        RECT 39.955 105.865 40.245 105.910 ;
        RECT 40.420 106.050 40.710 106.095 ;
        RECT 42.255 106.050 42.545 106.095 ;
        RECT 45.835 106.050 46.125 106.095 ;
        RECT 40.420 105.910 46.125 106.050 ;
        RECT 40.420 105.865 40.710 105.910 ;
        RECT 42.255 105.865 42.545 105.910 ;
        RECT 45.835 105.865 46.125 105.910 ;
        RECT 46.840 105.890 47.205 106.110 ;
        RECT 51.000 106.050 51.290 106.095 ;
        RECT 52.835 106.050 53.125 106.095 ;
        RECT 56.415 106.050 56.705 106.095 ;
        RECT 51.000 105.910 56.705 106.050 ;
        RECT 46.840 105.850 47.160 105.890 ;
        RECT 51.000 105.865 51.290 105.910 ;
        RECT 52.835 105.865 53.125 105.910 ;
        RECT 56.415 105.865 56.705 105.910 ;
        RECT 57.495 105.890 57.785 106.205 ;
        RECT 62.480 106.190 62.800 106.250 ;
        RECT 64.435 106.205 65.025 106.250 ;
        RECT 67.675 106.205 68.325 106.250 ;
        RECT 64.735 105.890 65.025 106.205 ;
        RECT 70.300 106.190 70.620 106.450 ;
        RECT 71.770 106.095 71.910 106.590 ;
        RECT 77.200 106.590 85.250 106.730 ;
        RECT 77.200 106.530 77.520 106.590 ;
        RECT 75.015 106.390 75.305 106.435 ;
        RECT 78.255 106.390 78.905 106.435 ;
        RECT 75.015 106.250 78.905 106.390 ;
        RECT 75.015 106.205 75.605 106.250 ;
        RECT 78.255 106.205 78.905 106.250 ;
        RECT 79.500 106.390 79.820 106.450 ;
        RECT 80.895 106.390 81.185 106.435 ;
        RECT 79.500 106.250 81.185 106.390 ;
        RECT 75.315 106.110 75.605 106.205 ;
        RECT 79.500 106.190 79.820 106.250 ;
        RECT 80.895 106.205 81.185 106.250 ;
        RECT 65.815 106.050 66.105 106.095 ;
        RECT 69.395 106.050 69.685 106.095 ;
        RECT 71.230 106.050 71.520 106.095 ;
        RECT 65.815 105.910 71.520 106.050 ;
        RECT 65.815 105.865 66.105 105.910 ;
        RECT 69.395 105.865 69.685 105.910 ;
        RECT 71.230 105.865 71.520 105.910 ;
        RECT 71.695 105.865 71.985 106.095 ;
        RECT 75.315 105.890 75.680 106.110 ;
        RECT 85.110 106.095 85.250 106.590 ;
        RECT 85.955 106.590 90.770 106.730 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 85.955 106.545 86.245 106.590 ;
        RECT 88.700 106.190 89.020 106.450 ;
        RECT 90.630 106.390 90.770 106.590 ;
        RECT 90.995 106.390 91.645 106.435 ;
        RECT 94.595 106.390 94.885 106.435 ;
        RECT 90.630 106.250 94.885 106.390 ;
        RECT 90.995 106.205 91.645 106.250 ;
        RECT 94.295 106.205 94.885 106.250 ;
        RECT 100.775 106.390 101.065 106.435 ;
        RECT 101.580 106.390 101.900 106.450 ;
        RECT 104.015 106.390 104.665 106.435 ;
        RECT 100.775 106.250 104.665 106.390 ;
        RECT 100.775 106.205 101.365 106.250 ;
        RECT 75.360 105.850 75.680 105.890 ;
        RECT 76.395 106.050 76.685 106.095 ;
        RECT 79.975 106.050 80.265 106.095 ;
        RECT 81.810 106.050 82.100 106.095 ;
        RECT 76.395 105.910 82.100 106.050 ;
        RECT 76.395 105.865 76.685 105.910 ;
        RECT 79.975 105.865 80.265 105.910 ;
        RECT 81.810 105.865 82.100 105.910 ;
        RECT 85.035 106.050 85.325 106.095 ;
        RECT 85.495 106.050 85.785 106.095 ;
        RECT 86.860 106.050 87.180 106.110 ;
        RECT 85.035 105.910 87.180 106.050 ;
        RECT 85.035 105.865 85.325 105.910 ;
        RECT 85.495 105.865 85.785 105.910 ;
        RECT 86.860 105.850 87.180 105.910 ;
        RECT 87.320 105.850 87.640 106.110 ;
        RECT 87.800 106.050 88.090 106.095 ;
        RECT 89.635 106.050 89.925 106.095 ;
        RECT 93.215 106.050 93.505 106.095 ;
        RECT 87.800 105.910 93.505 106.050 ;
        RECT 87.800 105.865 88.090 105.910 ;
        RECT 89.635 105.865 89.925 105.910 ;
        RECT 93.215 105.865 93.505 105.910 ;
        RECT 94.295 105.890 94.585 106.205 ;
        RECT 101.075 105.890 101.365 106.205 ;
        RECT 101.580 106.190 101.900 106.250 ;
        RECT 104.015 106.205 104.665 106.250 ;
        RECT 105.260 106.390 105.580 106.450 ;
        RECT 106.655 106.390 106.945 106.435 ;
        RECT 105.260 106.250 106.945 106.390 ;
        RECT 105.260 106.190 105.580 106.250 ;
        RECT 106.655 106.205 106.945 106.250 ;
        RECT 115.380 106.390 115.700 106.450 ;
        RECT 115.955 106.390 116.245 106.435 ;
        RECT 119.195 106.390 119.845 106.435 ;
        RECT 115.380 106.250 119.845 106.390 ;
        RECT 115.380 106.190 115.700 106.250 ;
        RECT 115.955 106.205 116.545 106.250 ;
        RECT 119.195 106.205 119.845 106.250 ;
        RECT 121.835 106.390 122.125 106.435 ;
        RECT 122.280 106.390 122.600 106.450 ;
        RECT 121.835 106.250 122.600 106.390 ;
        RECT 121.835 106.205 122.125 106.250 ;
        RECT 102.155 106.050 102.445 106.095 ;
        RECT 105.735 106.050 106.025 106.095 ;
        RECT 107.570 106.050 107.860 106.095 ;
        RECT 102.155 105.910 107.860 106.050 ;
        RECT 102.155 105.865 102.445 105.910 ;
        RECT 105.735 105.865 106.025 105.910 ;
        RECT 107.570 105.865 107.860 105.910 ;
        RECT 108.035 106.050 108.325 106.095 ;
        RECT 110.320 106.050 110.640 106.110 ;
        RECT 108.035 105.910 110.640 106.050 ;
        RECT 108.035 105.865 108.325 105.910 ;
        RECT 110.320 105.850 110.640 105.910 ;
        RECT 116.255 105.890 116.545 106.205 ;
        RECT 122.280 106.190 122.600 106.250 ;
        RECT 117.335 106.050 117.625 106.095 ;
        RECT 120.915 106.050 121.205 106.095 ;
        RECT 122.750 106.050 123.040 106.095 ;
        RECT 117.335 105.910 123.040 106.050 ;
        RECT 117.335 105.865 117.625 105.910 ;
        RECT 120.915 105.865 121.205 105.910 ;
        RECT 122.750 105.865 123.040 105.910 ;
        RECT 123.215 106.050 123.505 106.095 ;
        RECT 123.660 106.050 123.980 106.110 ;
        RECT 123.215 105.910 123.980 106.050 ;
        RECT 123.215 105.865 123.505 105.910 ;
        RECT 123.660 105.850 123.980 105.910 ;
        RECT 14.195 105.525 14.485 105.755 ;
        RECT 24.315 105.710 24.605 105.755 ;
        RECT 24.775 105.710 25.065 105.755 ;
        RECT 26.600 105.710 26.920 105.770 ;
        RECT 24.315 105.570 26.920 105.710 ;
        RECT 24.315 105.525 24.605 105.570 ;
        RECT 24.775 105.525 25.065 105.570 ;
        RECT 14.270 105.030 14.410 105.525 ;
        RECT 26.600 105.510 26.920 105.570 ;
        RECT 34.895 105.710 35.185 105.755 ;
        RECT 35.800 105.710 36.120 105.770 ;
        RECT 34.895 105.570 36.120 105.710 ;
        RECT 37.270 105.710 37.410 105.850 ;
        RECT 39.480 105.710 39.800 105.770 ;
        RECT 37.270 105.570 39.800 105.710 ;
        RECT 34.895 105.525 35.185 105.570 ;
        RECT 35.800 105.510 36.120 105.570 ;
        RECT 39.480 105.510 39.800 105.570 ;
        RECT 47.760 105.710 48.080 105.770 ;
        RECT 50.075 105.710 50.365 105.755 ;
        RECT 47.760 105.570 50.365 105.710 ;
        RECT 47.760 105.510 48.080 105.570 ;
        RECT 50.075 105.525 50.365 105.570 ;
        RECT 50.535 105.710 50.825 105.755 ;
        RECT 51.900 105.710 52.220 105.770 ;
        RECT 50.535 105.570 52.220 105.710 ;
        RECT 50.535 105.525 50.825 105.570 ;
        RECT 51.900 105.510 52.220 105.570 ;
        RECT 55.580 105.710 55.900 105.770 ;
        RECT 60.655 105.710 60.945 105.755 ;
        RECT 55.580 105.570 60.945 105.710 ;
        RECT 55.580 105.510 55.900 105.570 ;
        RECT 60.655 105.525 60.945 105.570 ;
        RECT 61.575 105.710 61.865 105.755 ;
        RECT 65.240 105.710 65.560 105.770 ;
        RECT 72.155 105.710 72.445 105.755 ;
        RECT 61.575 105.570 65.560 105.710 ;
        RECT 61.575 105.525 61.865 105.570 ;
        RECT 65.240 105.510 65.560 105.570 ;
        RECT 71.770 105.570 72.445 105.710 ;
        RECT 71.770 105.430 71.910 105.570 ;
        RECT 72.155 105.525 72.445 105.570 ;
        RECT 82.275 105.710 82.565 105.755 ;
        RECT 87.410 105.710 87.550 105.850 ;
        RECT 82.275 105.570 87.550 105.710 ;
        RECT 91.460 105.710 91.780 105.770 ;
        RECT 97.455 105.710 97.745 105.755 ;
        RECT 91.460 105.570 97.745 105.710 ;
        RECT 82.275 105.525 82.565 105.570 ;
        RECT 91.460 105.510 91.780 105.570 ;
        RECT 97.455 105.525 97.745 105.570 ;
        RECT 97.915 105.710 98.205 105.755 ;
        RECT 101.580 105.710 101.900 105.770 ;
        RECT 97.915 105.570 101.900 105.710 ;
        RECT 97.915 105.525 98.205 105.570 ;
        RECT 101.580 105.510 101.900 105.570 ;
        RECT 113.080 105.510 113.400 105.770 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 18.435 105.370 18.725 105.415 ;
        RECT 21.555 105.370 21.845 105.415 ;
        RECT 23.445 105.370 23.735 105.415 ;
        RECT 18.435 105.230 23.735 105.370 ;
        RECT 18.435 105.185 18.725 105.230 ;
        RECT 21.555 105.185 21.845 105.230 ;
        RECT 23.445 105.185 23.735 105.230 ;
        RECT 25.645 105.370 25.935 105.415 ;
        RECT 27.535 105.370 27.825 105.415 ;
        RECT 30.655 105.370 30.945 105.415 ;
        RECT 25.645 105.230 30.945 105.370 ;
        RECT 25.645 105.185 25.935 105.230 ;
        RECT 27.535 105.185 27.825 105.230 ;
        RECT 30.655 105.185 30.945 105.230 ;
        RECT 40.825 105.370 41.115 105.415 ;
        RECT 42.715 105.370 43.005 105.415 ;
        RECT 45.835 105.370 46.125 105.415 ;
        RECT 40.825 105.230 46.125 105.370 ;
        RECT 40.825 105.185 41.115 105.230 ;
        RECT 42.715 105.185 43.005 105.230 ;
        RECT 45.835 105.185 46.125 105.230 ;
        RECT 51.405 105.370 51.695 105.415 ;
        RECT 53.295 105.370 53.585 105.415 ;
        RECT 56.415 105.370 56.705 105.415 ;
        RECT 51.405 105.230 56.705 105.370 ;
        RECT 51.405 105.185 51.695 105.230 ;
        RECT 53.295 105.185 53.585 105.230 ;
        RECT 56.415 105.185 56.705 105.230 ;
        RECT 65.815 105.370 66.105 105.415 ;
        RECT 68.935 105.370 69.225 105.415 ;
        RECT 70.825 105.370 71.115 105.415 ;
        RECT 65.815 105.230 71.115 105.370 ;
        RECT 65.815 105.185 66.105 105.230 ;
        RECT 68.935 105.185 69.225 105.230 ;
        RECT 70.825 105.185 71.115 105.230 ;
        RECT 71.680 105.170 72.000 105.430 ;
        RECT 76.395 105.370 76.685 105.415 ;
        RECT 79.515 105.370 79.805 105.415 ;
        RECT 81.405 105.370 81.695 105.415 ;
        RECT 76.395 105.230 81.695 105.370 ;
        RECT 76.395 105.185 76.685 105.230 ;
        RECT 79.515 105.185 79.805 105.230 ;
        RECT 81.405 105.185 81.695 105.230 ;
        RECT 88.205 105.370 88.495 105.415 ;
        RECT 90.095 105.370 90.385 105.415 ;
        RECT 93.215 105.370 93.505 105.415 ;
        RECT 88.205 105.230 93.505 105.370 ;
        RECT 88.205 105.185 88.495 105.230 ;
        RECT 90.095 105.185 90.385 105.230 ;
        RECT 93.215 105.185 93.505 105.230 ;
        RECT 102.155 105.370 102.445 105.415 ;
        RECT 105.275 105.370 105.565 105.415 ;
        RECT 107.165 105.370 107.455 105.415 ;
        RECT 102.155 105.230 107.455 105.370 ;
        RECT 102.155 105.185 102.445 105.230 ;
        RECT 105.275 105.185 105.565 105.230 ;
        RECT 107.165 105.185 107.455 105.230 ;
        RECT 117.335 105.370 117.625 105.415 ;
        RECT 120.455 105.370 120.745 105.415 ;
        RECT 122.345 105.370 122.635 105.415 ;
        RECT 117.335 105.230 122.635 105.370 ;
        RECT 117.335 105.185 117.625 105.230 ;
        RECT 120.455 105.185 120.745 105.230 ;
        RECT 122.345 105.185 122.635 105.230 ;
        RECT 23.840 105.030 24.160 105.090 ;
        RECT 14.270 104.890 24.160 105.030 ;
        RECT 23.840 104.830 24.160 104.890 ;
        RECT 26.095 105.030 26.385 105.075 ;
        RECT 38.560 105.030 38.880 105.090 ;
        RECT 26.095 104.890 38.880 105.030 ;
        RECT 26.095 104.845 26.385 104.890 ;
        RECT 38.560 104.830 38.880 104.890 ;
        RECT 84.560 104.830 84.880 105.090 ;
        RECT 11.810 104.210 125.890 104.690 ;
        RECT 46.840 104.010 47.160 104.070 ;
        RECT 47.315 104.010 47.605 104.055 ;
        RECT 46.840 103.870 47.605 104.010 ;
        RECT 46.840 103.810 47.160 103.870 ;
        RECT 47.315 103.825 47.605 103.870 ;
        RECT 60.180 103.810 60.500 104.070 ;
        RECT 62.480 103.810 62.800 104.070 ;
        RECT 73.060 103.810 73.380 104.070 ;
        RECT 75.360 103.810 75.680 104.070 ;
        RECT 95.140 103.810 95.460 104.070 ;
        RECT 117.220 103.810 117.540 104.070 ;
        RECT 27.175 103.670 27.465 103.715 ;
        RECT 30.295 103.670 30.585 103.715 ;
        RECT 32.185 103.670 32.475 103.715 ;
        RECT 27.175 103.530 32.475 103.670 ;
        RECT 27.175 103.485 27.465 103.530 ;
        RECT 30.295 103.485 30.585 103.530 ;
        RECT 32.185 103.485 32.475 103.530 ;
        RECT 80.535 103.670 80.825 103.715 ;
        RECT 83.655 103.670 83.945 103.715 ;
        RECT 85.545 103.670 85.835 103.715 ;
        RECT 80.535 103.530 85.835 103.670 ;
        RECT 80.535 103.485 80.825 103.530 ;
        RECT 83.655 103.485 83.945 103.530 ;
        RECT 85.545 103.485 85.835 103.530 ;
        RECT 31.660 103.130 31.980 103.390 ;
        RECT 85.020 103.130 85.340 103.390 ;
        RECT 86.415 103.330 86.705 103.375 ;
        RECT 87.320 103.330 87.640 103.390 ;
        RECT 86.415 103.190 87.640 103.330 ;
        RECT 86.415 103.145 86.705 103.190 ;
        RECT 87.320 103.130 87.640 103.190 ;
        RECT 19.240 102.990 19.560 103.050 ;
        RECT 26.095 102.990 26.385 103.010 ;
        RECT 19.240 102.850 26.385 102.990 ;
        RECT 19.240 102.790 19.560 102.850 ;
        RECT 13.260 102.650 13.580 102.710 ;
        RECT 26.095 102.695 26.385 102.850 ;
        RECT 27.175 102.990 27.465 103.035 ;
        RECT 30.755 102.990 31.045 103.035 ;
        RECT 32.590 102.990 32.880 103.035 ;
        RECT 27.175 102.850 32.880 102.990 ;
        RECT 27.175 102.805 27.465 102.850 ;
        RECT 30.755 102.805 31.045 102.850 ;
        RECT 32.590 102.805 32.880 102.850 ;
        RECT 33.055 102.805 33.345 103.035 ;
        RECT 39.480 102.990 39.800 103.050 ;
        RECT 47.775 102.990 48.065 103.035 ;
        RECT 56.040 102.990 56.360 103.050 ;
        RECT 59.735 102.990 60.025 103.035 ;
        RECT 62.035 102.990 62.325 103.035 ;
        RECT 39.480 102.850 62.325 102.990 ;
        RECT 22.935 102.650 23.225 102.695 ;
        RECT 13.260 102.510 23.225 102.650 ;
        RECT 13.260 102.450 13.580 102.510 ;
        RECT 22.935 102.465 23.225 102.510 ;
        RECT 25.795 102.650 26.385 102.695 ;
        RECT 29.035 102.650 29.685 102.695 ;
        RECT 25.795 102.510 29.685 102.650 ;
        RECT 25.795 102.465 26.085 102.510 ;
        RECT 29.035 102.465 29.685 102.510 ;
        RECT 27.060 102.310 27.380 102.370 ;
        RECT 33.130 102.310 33.270 102.805 ;
        RECT 39.480 102.790 39.800 102.850 ;
        RECT 47.775 102.805 48.065 102.850 ;
        RECT 56.040 102.790 56.360 102.850 ;
        RECT 59.735 102.805 60.025 102.850 ;
        RECT 62.035 102.805 62.325 102.850 ;
        RECT 73.535 102.990 73.825 103.035 ;
        RECT 74.915 102.990 75.205 103.035 ;
        RECT 77.200 102.990 77.520 103.050 ;
        RECT 73.535 102.850 77.520 102.990 ;
        RECT 73.535 102.805 73.825 102.850 ;
        RECT 74.915 102.805 75.205 102.850 ;
        RECT 77.200 102.790 77.520 102.850 ;
        RECT 79.455 102.695 79.745 103.010 ;
        RECT 80.535 102.990 80.825 103.035 ;
        RECT 84.115 102.990 84.405 103.035 ;
        RECT 85.950 102.990 86.240 103.035 ;
        RECT 80.535 102.850 86.240 102.990 ;
        RECT 80.535 102.805 80.825 102.850 ;
        RECT 84.115 102.805 84.405 102.850 ;
        RECT 85.950 102.805 86.240 102.850 ;
        RECT 86.860 102.990 87.180 103.050 ;
        RECT 95.615 102.990 95.905 103.035 ;
        RECT 101.120 102.990 101.440 103.050 ;
        RECT 116.775 102.990 117.065 103.035 ;
        RECT 86.860 102.850 117.065 102.990 ;
        RECT 86.860 102.790 87.180 102.850 ;
        RECT 95.615 102.805 95.905 102.850 ;
        RECT 101.120 102.790 101.440 102.850 ;
        RECT 116.775 102.805 117.065 102.850 ;
        RECT 76.295 102.465 76.585 102.695 ;
        RECT 79.155 102.650 79.745 102.695 ;
        RECT 82.395 102.650 83.045 102.695 ;
        RECT 84.560 102.650 84.880 102.710 ;
        RECT 79.155 102.510 84.880 102.650 ;
        RECT 79.155 102.465 79.445 102.510 ;
        RECT 82.395 102.465 83.045 102.510 ;
        RECT 27.060 102.170 33.270 102.310 ;
        RECT 76.370 102.310 76.510 102.465 ;
        RECT 84.560 102.450 84.880 102.510 ;
        RECT 83.640 102.310 83.960 102.370 ;
        RECT 76.370 102.170 83.960 102.310 ;
        RECT 27.060 102.110 27.380 102.170 ;
        RECT 83.640 102.110 83.960 102.170 ;
        RECT 11.010 101.490 125.890 101.970 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 11.040 215.785 12.580 216.155 ;
        RECT 39.560 215.785 41.100 216.155 ;
        RECT 68.080 215.785 69.620 216.155 ;
        RECT 96.600 215.785 98.140 216.155 ;
        RECT 25.300 213.065 26.840 213.435 ;
        RECT 53.820 213.065 55.360 213.435 ;
        RECT 82.340 213.065 83.880 213.435 ;
        RECT 110.860 213.065 112.400 213.435 ;
        RECT 11.040 210.345 12.580 210.715 ;
        RECT 39.560 210.345 41.100 210.715 ;
        RECT 68.080 210.345 69.620 210.715 ;
        RECT 96.600 210.345 98.140 210.715 ;
        RECT 25.300 207.625 26.840 207.995 ;
        RECT 53.820 207.625 55.360 207.995 ;
        RECT 82.340 207.625 83.880 207.995 ;
        RECT 110.860 207.625 112.400 207.995 ;
        RECT 11.040 204.905 12.580 205.275 ;
        RECT 39.560 204.905 41.100 205.275 ;
        RECT 68.080 204.905 69.620 205.275 ;
        RECT 96.600 204.905 98.140 205.275 ;
        RECT 25.300 202.185 26.840 202.555 ;
        RECT 53.820 202.185 55.360 202.555 ;
        RECT 82.340 202.185 83.880 202.555 ;
        RECT 110.860 202.185 112.400 202.555 ;
        RECT 11.040 199.465 12.580 199.835 ;
        RECT 39.560 199.465 41.100 199.835 ;
        RECT 68.080 199.465 69.620 199.835 ;
        RECT 96.600 199.465 98.140 199.835 ;
        RECT 65.270 198.640 65.530 198.960 ;
        RECT 64.810 197.280 65.070 197.600 ;
        RECT 25.300 196.745 26.840 197.115 ;
        RECT 53.820 196.745 55.360 197.115 ;
        RECT 62.970 195.580 63.230 195.900 ;
        RECT 57.450 195.240 57.710 195.560 ;
        RECT 11.040 194.025 12.580 194.395 ;
        RECT 39.560 194.025 41.100 194.395 ;
        RECT 25.300 191.305 26.840 191.675 ;
        RECT 53.820 191.305 55.360 191.675 ;
        RECT 11.040 188.585 12.580 188.955 ;
        RECT 39.560 188.585 41.100 188.955 ;
        RECT 32.150 187.420 32.410 187.740 ;
        RECT 51.010 187.650 51.270 187.740 ;
        RECT 50.610 187.510 51.270 187.650 ;
        RECT 25.300 185.865 26.840 186.235 ;
        RECT 32.210 184.680 32.350 187.420 ;
        RECT 47.330 187.080 47.590 187.400 ;
        RECT 43.650 186.400 43.910 186.720 ;
        RECT 43.710 185.020 43.850 186.400 ;
        RECT 35.370 184.700 35.630 185.020 ;
        RECT 43.650 184.700 43.910 185.020 ;
        RECT 32.150 184.360 32.410 184.680 ;
        RECT 33.990 184.360 34.250 184.680 ;
        RECT 11.040 183.145 12.580 183.515 ;
        RECT 25.300 180.425 26.840 180.795 ;
        RECT 11.040 177.705 12.580 178.075 ;
        RECT 32.210 176.860 32.350 184.360 ;
        RECT 32.150 176.540 32.410 176.860 ;
        RECT 30.310 175.520 30.570 175.840 ;
        RECT 25.300 174.985 26.840 175.355 ;
        RECT 23.410 173.480 23.670 173.800 ;
        RECT 22.030 173.140 22.290 173.460 ;
        RECT 11.040 172.265 12.580 172.635 ;
        RECT 17.430 171.100 17.690 171.420 ;
        RECT 17.490 169.380 17.630 171.100 ;
        RECT 21.110 170.760 21.370 171.080 ;
        RECT 17.430 169.060 17.690 169.380 ;
        RECT 11.040 166.825 12.580 167.195 ;
        RECT 21.170 166.660 21.310 170.760 ;
        RECT 22.090 169.380 22.230 173.140 ;
        RECT 22.030 169.060 22.290 169.380 ;
        RECT 23.470 168.360 23.610 173.480 ;
        RECT 30.370 173.460 30.510 175.520 ;
        RECT 32.210 174.140 32.350 176.540 ;
        RECT 32.150 173.820 32.410 174.140 ;
        RECT 34.050 173.460 34.190 184.360 ;
        RECT 35.430 182.980 35.570 184.700 ;
        RECT 38.590 183.740 38.850 184.000 ;
        RECT 38.190 183.680 38.850 183.740 ;
        RECT 42.730 183.680 42.990 184.000 ;
        RECT 38.190 183.600 38.790 183.680 ;
        RECT 35.370 182.660 35.630 182.980 ;
        RECT 36.750 176.540 37.010 176.860 ;
        RECT 30.310 173.140 30.570 173.460 ;
        RECT 33.990 173.140 34.250 173.460 ;
        RECT 24.790 172.800 25.050 173.120 ;
        RECT 27.090 172.800 27.350 173.120 ;
        RECT 27.550 172.800 27.810 173.120 ;
        RECT 33.530 172.800 33.790 173.120 ;
        RECT 23.870 170.080 24.130 170.400 ;
        RECT 23.410 168.040 23.670 168.360 ;
        RECT 22.950 167.360 23.210 167.680 ;
        RECT 21.110 166.340 21.370 166.660 ;
        RECT 23.010 165.980 23.150 167.360 ;
        RECT 23.930 166.660 24.070 170.080 ;
        RECT 24.330 168.380 24.590 168.700 ;
        RECT 24.390 167.420 24.530 168.380 ;
        RECT 24.850 168.360 24.990 172.800 ;
        RECT 25.300 169.545 26.840 169.915 ;
        RECT 24.790 168.040 25.050 168.360 ;
        RECT 27.150 168.100 27.290 172.800 ;
        RECT 27.610 168.700 27.750 172.800 ;
        RECT 33.590 171.080 33.730 172.800 ;
        RECT 32.150 170.760 32.410 171.080 ;
        RECT 33.530 170.760 33.790 171.080 ;
        RECT 32.210 170.400 32.350 170.760 ;
        RECT 34.050 170.740 34.190 173.140 ;
        RECT 34.910 172.800 35.170 173.120 ;
        RECT 34.970 172.100 35.110 172.800 ;
        RECT 34.910 171.780 35.170 172.100 ;
        RECT 36.290 171.440 36.550 171.760 ;
        RECT 34.910 170.760 35.170 171.080 ;
        RECT 33.990 170.420 34.250 170.740 ;
        RECT 32.150 170.080 32.410 170.400 ;
        RECT 33.530 170.080 33.790 170.400 ;
        RECT 27.550 168.380 27.810 168.700 ;
        RECT 32.150 168.380 32.410 168.700 ;
        RECT 27.150 167.960 27.750 168.100 ;
        RECT 24.390 167.280 24.990 167.420 ;
        RECT 23.870 166.340 24.130 166.660 ;
        RECT 22.950 165.660 23.210 165.980 ;
        RECT 11.040 161.385 12.580 161.755 ;
        RECT 23.930 161.220 24.070 166.340 ;
        RECT 24.330 165.660 24.590 165.980 ;
        RECT 23.870 160.900 24.130 161.220 ;
        RECT 22.490 160.220 22.750 160.540 ;
        RECT 22.030 157.160 22.290 157.480 ;
        RECT 13.750 156.820 14.010 157.140 ;
        RECT 11.040 155.945 12.580 156.315 ;
        RECT 13.810 155.780 13.950 156.820 ;
        RECT 13.750 155.460 14.010 155.780 ;
        RECT 21.570 155.120 21.830 155.440 ;
        RECT 14.210 154.780 14.470 155.100 ;
        RECT 16.510 154.780 16.770 155.100 ;
        RECT 11.040 150.505 12.580 150.875 ;
        RECT 14.270 149.660 14.410 154.780 ;
        RECT 16.570 150.340 16.710 154.780 ;
        RECT 19.270 154.440 19.530 154.760 ;
        RECT 17.430 151.380 17.690 151.700 ;
        RECT 17.490 150.340 17.630 151.380 ;
        RECT 19.330 150.340 19.470 154.440 ;
        RECT 21.630 153.820 21.770 155.120 ;
        RECT 22.090 154.670 22.230 157.160 ;
        RECT 22.550 155.440 22.690 160.220 ;
        RECT 22.950 159.880 23.210 160.200 ;
        RECT 23.010 156.660 23.150 159.880 ;
        RECT 23.410 159.200 23.670 159.520 ;
        RECT 23.470 157.480 23.610 159.200 ;
        RECT 23.410 157.160 23.670 157.480 ;
        RECT 23.010 156.520 23.610 156.660 ;
        RECT 22.490 155.120 22.750 155.440 ;
        RECT 23.470 155.180 23.610 156.520 ;
        RECT 23.470 155.040 24.070 155.180 ;
        RECT 23.410 154.670 23.670 154.760 ;
        RECT 22.090 154.530 23.670 154.670 ;
        RECT 21.630 153.680 22.230 153.820 ;
        RECT 21.570 151.040 21.830 151.360 ;
        RECT 21.630 150.340 21.770 151.040 ;
        RECT 16.510 150.020 16.770 150.340 ;
        RECT 17.430 150.020 17.690 150.340 ;
        RECT 19.270 150.020 19.530 150.340 ;
        RECT 21.570 150.020 21.830 150.340 ;
        RECT 14.210 149.340 14.470 149.660 ;
        RECT 22.090 149.320 22.230 153.680 ;
        RECT 23.010 152.040 23.150 154.530 ;
        RECT 23.410 154.440 23.670 154.530 ;
        RECT 23.400 153.565 23.680 153.935 ;
        RECT 22.950 151.720 23.210 152.040 ;
        RECT 22.030 149.000 22.290 149.320 ;
        RECT 22.090 147.280 22.230 149.000 ;
        RECT 22.030 146.960 22.290 147.280 ;
        RECT 11.040 145.065 12.580 145.435 ;
        RECT 14.670 144.240 14.930 144.560 ;
        RECT 11.040 139.625 12.580 139.995 ;
        RECT 14.730 139.460 14.870 144.240 ;
        RECT 23.010 144.220 23.150 151.720 ;
        RECT 23.470 144.560 23.610 153.565 ;
        RECT 23.930 152.720 24.070 155.040 ;
        RECT 24.390 154.615 24.530 165.660 ;
        RECT 24.850 165.640 24.990 167.280 ;
        RECT 27.610 165.980 27.750 167.960 ;
        RECT 27.550 165.660 27.810 165.980 ;
        RECT 24.790 165.320 25.050 165.640 ;
        RECT 24.850 160.200 24.990 165.320 ;
        RECT 28.010 164.640 28.270 164.960 ;
        RECT 25.300 164.105 26.840 164.475 ;
        RECT 28.070 163.260 28.210 164.640 ;
        RECT 32.210 164.020 32.350 168.380 ;
        RECT 32.610 167.360 32.870 167.680 ;
        RECT 31.750 163.880 32.350 164.020 ;
        RECT 32.670 163.940 32.810 167.360 ;
        RECT 33.070 165.320 33.330 165.640 ;
        RECT 33.130 163.940 33.270 165.320 ;
        RECT 28.010 162.940 28.270 163.260 ;
        RECT 28.070 161.220 28.210 162.940 ;
        RECT 28.010 160.900 28.270 161.220 ;
        RECT 24.790 159.880 25.050 160.200 ;
        RECT 25.300 158.665 26.840 159.035 ;
        RECT 31.750 158.500 31.890 163.880 ;
        RECT 32.610 163.620 32.870 163.940 ;
        RECT 33.070 163.620 33.330 163.940 ;
        RECT 33.590 160.200 33.730 170.080 ;
        RECT 34.050 168.700 34.190 170.420 ;
        RECT 33.990 168.380 34.250 168.700 ;
        RECT 34.050 168.100 34.190 168.380 ;
        RECT 34.050 167.960 34.650 168.100 ;
        RECT 34.970 168.020 35.110 170.760 ;
        RECT 35.830 170.420 36.090 170.740 ;
        RECT 35.890 169.040 36.030 170.420 ;
        RECT 36.350 169.380 36.490 171.440 ;
        RECT 36.290 169.060 36.550 169.380 ;
        RECT 35.830 168.720 36.090 169.040 ;
        RECT 36.810 168.360 36.950 176.540 ;
        RECT 37.670 170.080 37.930 170.400 ;
        RECT 37.730 168.700 37.870 170.080 ;
        RECT 37.670 168.380 37.930 168.700 ;
        RECT 36.750 168.040 37.010 168.360 ;
        RECT 34.510 165.980 34.650 167.960 ;
        RECT 34.910 167.700 35.170 168.020 ;
        RECT 34.450 165.660 34.710 165.980 ;
        RECT 34.970 165.300 35.110 167.700 ;
        RECT 36.750 166.000 37.010 166.320 ;
        RECT 34.910 164.980 35.170 165.300 ;
        RECT 36.280 164.445 36.560 164.815 ;
        RECT 34.910 162.600 35.170 162.920 ;
        RECT 34.450 161.920 34.710 162.240 ;
        RECT 33.530 159.880 33.790 160.200 ;
        RECT 33.070 159.540 33.330 159.860 ;
        RECT 31.690 158.180 31.950 158.500 ;
        RECT 30.310 157.160 30.570 157.480 ;
        RECT 27.090 156.480 27.350 156.800 ;
        RECT 24.790 154.780 25.050 155.100 ;
        RECT 24.320 154.245 24.600 154.615 ;
        RECT 24.330 153.760 24.590 154.080 ;
        RECT 23.870 152.400 24.130 152.720 ;
        RECT 23.930 149.320 24.070 152.400 ;
        RECT 24.390 152.380 24.530 153.760 ;
        RECT 24.850 153.060 24.990 154.780 ;
        RECT 25.300 153.225 26.840 153.595 ;
        RECT 24.790 152.740 25.050 153.060 ;
        RECT 24.330 152.060 24.590 152.380 ;
        RECT 27.150 151.700 27.290 156.480 ;
        RECT 28.010 154.780 28.270 155.100 ;
        RECT 27.550 153.760 27.810 154.080 ;
        RECT 24.790 151.610 25.050 151.700 ;
        RECT 24.790 151.470 25.450 151.610 ;
        RECT 24.790 151.380 25.050 151.470 ;
        RECT 25.310 150.000 25.450 151.470 ;
        RECT 27.090 151.380 27.350 151.700 ;
        RECT 27.610 150.000 27.750 153.760 ;
        RECT 28.070 150.340 28.210 154.780 ;
        RECT 30.370 153.060 30.510 157.160 ;
        RECT 30.310 152.740 30.570 153.060 ;
        RECT 28.930 151.040 29.190 151.360 ;
        RECT 28.990 150.340 29.130 151.040 ;
        RECT 28.010 150.020 28.270 150.340 ;
        RECT 28.930 150.020 29.190 150.340 ;
        RECT 25.250 149.680 25.510 150.000 ;
        RECT 27.550 149.680 27.810 150.000 ;
        RECT 30.370 149.660 30.510 152.740 ;
        RECT 33.130 150.340 33.270 159.540 ;
        RECT 33.990 158.180 34.250 158.500 ;
        RECT 34.050 155.440 34.190 158.180 ;
        RECT 33.530 155.120 33.790 155.440 ;
        RECT 33.990 155.120 34.250 155.440 ;
        RECT 33.590 150.340 33.730 155.120 ;
        RECT 31.690 150.020 31.950 150.340 ;
        RECT 33.070 150.020 33.330 150.340 ;
        RECT 33.530 150.020 33.790 150.340 ;
        RECT 30.310 149.340 30.570 149.660 ;
        RECT 23.870 149.000 24.130 149.320 ;
        RECT 31.750 148.640 31.890 150.020 ;
        RECT 31.690 148.320 31.950 148.640 ;
        RECT 25.300 147.785 26.840 148.155 ;
        RECT 33.130 147.620 33.270 150.020 ;
        RECT 33.070 147.300 33.330 147.620 ;
        RECT 31.690 144.580 31.950 144.900 ;
        RECT 23.410 144.240 23.670 144.560 ;
        RECT 22.950 143.900 23.210 144.220 ;
        RECT 22.030 143.560 22.290 143.880 ;
        RECT 17.430 142.880 17.690 143.200 ;
        RECT 17.490 141.500 17.630 142.880 ;
        RECT 22.090 142.180 22.230 143.560 ;
        RECT 24.790 143.220 25.050 143.540 ;
        RECT 22.030 141.860 22.290 142.180 ;
        RECT 17.430 141.180 17.690 141.500 ;
        RECT 19.730 141.180 19.990 141.500 ;
        RECT 15.130 140.500 15.390 140.820 ;
        RECT 14.670 139.140 14.930 139.460 ;
        RECT 15.190 138.780 15.330 140.500 ;
        RECT 17.490 139.460 17.630 141.180 ;
        RECT 19.270 140.840 19.530 141.160 ;
        RECT 19.330 139.460 19.470 140.840 ;
        RECT 17.430 139.140 17.690 139.460 ;
        RECT 19.270 139.140 19.530 139.460 ;
        RECT 15.130 138.460 15.390 138.780 ;
        RECT 11.040 134.185 12.580 134.555 ;
        RECT 15.190 130.280 15.330 138.460 ;
        RECT 16.510 138.120 16.770 138.440 ;
        RECT 16.570 136.060 16.710 138.120 ;
        RECT 16.510 135.740 16.770 136.060 ;
        RECT 17.490 135.720 17.630 139.140 ;
        RECT 19.790 139.120 19.930 141.180 ;
        RECT 23.410 140.160 23.670 140.480 ;
        RECT 23.470 139.120 23.610 140.160 ;
        RECT 19.730 138.800 19.990 139.120 ;
        RECT 23.410 138.800 23.670 139.120 ;
        RECT 17.430 135.400 17.690 135.720 ;
        RECT 19.730 134.720 19.990 135.040 ;
        RECT 24.330 134.720 24.590 135.040 ;
        RECT 17.430 133.360 17.690 133.680 ;
        RECT 17.490 131.300 17.630 133.360 ;
        RECT 19.790 132.320 19.930 134.720 ;
        RECT 24.390 133.340 24.530 134.720 ;
        RECT 24.330 133.020 24.590 133.340 ;
        RECT 24.850 132.740 24.990 143.220 ;
        RECT 25.300 142.345 26.840 142.715 ;
        RECT 30.770 141.180 31.030 141.500 ;
        RECT 27.550 140.160 27.810 140.480 ;
        RECT 29.850 140.160 30.110 140.480 ;
        RECT 27.610 137.760 27.750 140.160 ;
        RECT 29.910 138.780 30.050 140.160 ;
        RECT 29.850 138.460 30.110 138.780 ;
        RECT 30.830 138.440 30.970 141.180 ;
        RECT 28.010 138.120 28.270 138.440 ;
        RECT 30.770 138.120 31.030 138.440 ;
        RECT 27.550 137.440 27.810 137.760 ;
        RECT 25.300 136.905 26.840 137.275 ;
        RECT 27.610 136.740 27.750 137.440 ;
        RECT 27.550 136.420 27.810 136.740 ;
        RECT 28.070 135.040 28.210 138.120 ;
        RECT 30.830 136.060 30.970 138.120 ;
        RECT 30.770 135.740 31.030 136.060 ;
        RECT 28.010 134.720 28.270 135.040 ;
        RECT 28.070 133.000 28.210 134.720 ;
        RECT 29.850 133.020 30.110 133.340 ;
        RECT 24.390 132.600 24.990 132.740 ;
        RECT 28.010 132.680 28.270 133.000 ;
        RECT 19.730 132.000 19.990 132.320 ;
        RECT 17.430 130.980 17.690 131.300 ;
        RECT 19.790 130.620 19.930 132.000 ;
        RECT 19.730 130.300 19.990 130.620 ;
        RECT 15.130 129.960 15.390 130.280 ;
        RECT 16.970 129.960 17.230 130.280 ;
        RECT 11.040 128.745 12.580 129.115 ;
        RECT 17.030 124.840 17.170 129.960 ;
        RECT 20.190 129.620 20.450 129.940 ;
        RECT 20.250 128.580 20.390 129.620 ;
        RECT 20.190 128.260 20.450 128.580 ;
        RECT 17.430 127.920 17.690 128.240 ;
        RECT 17.490 125.860 17.630 127.920 ;
        RECT 17.430 125.540 17.690 125.860 ;
        RECT 20.250 125.520 20.390 128.260 ;
        RECT 20.190 125.200 20.450 125.520 ;
        RECT 16.970 124.520 17.230 124.840 ;
        RECT 11.040 123.305 12.580 123.675 ;
        RECT 16.050 122.480 16.310 122.800 ;
        RECT 16.110 120.420 16.250 122.480 ;
        RECT 16.050 120.100 16.310 120.420 ;
        RECT 17.030 119.400 17.170 124.520 ;
        RECT 20.190 123.840 20.450 124.160 ;
        RECT 23.410 123.840 23.670 124.160 ;
        RECT 17.890 122.140 18.150 122.460 ;
        RECT 16.970 119.080 17.230 119.400 ;
        RECT 17.950 118.720 18.090 122.140 ;
        RECT 20.250 121.440 20.390 123.840 ;
        RECT 22.950 121.800 23.210 122.120 ;
        RECT 20.190 121.120 20.450 121.440 ;
        RECT 20.250 119.740 20.390 121.120 ;
        RECT 23.010 120.420 23.150 121.800 ;
        RECT 22.950 120.100 23.210 120.420 ;
        RECT 20.190 119.420 20.450 119.740 ;
        RECT 17.430 118.400 17.690 118.720 ;
        RECT 17.890 118.400 18.150 118.720 ;
        RECT 11.040 117.865 12.580 118.235 ;
        RECT 17.490 117.360 17.630 118.400 ;
        RECT 20.250 117.700 20.390 119.420 ;
        RECT 20.190 117.380 20.450 117.700 ;
        RECT 17.430 117.040 17.690 117.360 ;
        RECT 23.470 117.020 23.610 123.840 ;
        RECT 23.410 116.700 23.670 117.020 ;
        RECT 24.390 113.960 24.530 132.600 ;
        RECT 25.300 131.465 26.840 131.835 ;
        RECT 28.070 130.280 28.210 132.680 ;
        RECT 28.010 129.960 28.270 130.280 ;
        RECT 28.470 129.960 28.730 130.280 ;
        RECT 24.790 129.280 25.050 129.600 ;
        RECT 24.850 127.900 24.990 129.280 ;
        RECT 24.790 127.580 25.050 127.900 ;
        RECT 27.090 127.580 27.350 127.900 ;
        RECT 25.300 126.025 26.840 126.395 ;
        RECT 25.300 120.585 26.840 120.955 ;
        RECT 27.150 119.400 27.290 127.580 ;
        RECT 28.070 127.560 28.210 129.960 ;
        RECT 28.530 128.580 28.670 129.960 ;
        RECT 28.470 128.260 28.730 128.580 ;
        RECT 28.470 127.580 28.730 127.900 ;
        RECT 28.010 127.240 28.270 127.560 ;
        RECT 28.070 123.140 28.210 127.240 ;
        RECT 28.530 125.520 28.670 127.580 ;
        RECT 28.930 127.240 29.190 127.560 ;
        RECT 28.470 125.200 28.730 125.520 ;
        RECT 28.990 125.180 29.130 127.240 ;
        RECT 29.390 126.560 29.650 126.880 ;
        RECT 29.450 125.860 29.590 126.560 ;
        RECT 29.390 125.540 29.650 125.860 ;
        RECT 28.930 124.860 29.190 125.180 ;
        RECT 28.470 123.840 28.730 124.160 ;
        RECT 28.010 122.820 28.270 123.140 ;
        RECT 27.550 122.480 27.810 122.800 ;
        RECT 27.610 120.080 27.750 122.480 ;
        RECT 28.530 120.420 28.670 123.840 ;
        RECT 28.990 122.120 29.130 124.860 ;
        RECT 28.930 121.800 29.190 122.120 ;
        RECT 28.470 120.100 28.730 120.420 ;
        RECT 27.550 119.760 27.810 120.080 ;
        RECT 28.530 119.740 28.670 120.100 ;
        RECT 28.470 119.420 28.730 119.740 ;
        RECT 27.090 119.080 27.350 119.400 ;
        RECT 27.550 118.400 27.810 118.720 ;
        RECT 27.610 116.680 27.750 118.400 ;
        RECT 27.090 116.360 27.350 116.680 ;
        RECT 27.550 116.360 27.810 116.680 ;
        RECT 25.300 115.145 26.840 115.515 ;
        RECT 24.330 113.640 24.590 113.960 ;
        RECT 11.040 112.425 12.580 112.795 ;
        RECT 22.030 111.600 22.290 111.920 ;
        RECT 16.970 110.920 17.230 111.240 ;
        RECT 11.040 106.985 12.580 107.355 ;
        RECT 13.290 102.420 13.550 102.740 ;
        RECT 11.040 101.545 12.580 101.915 ;
        RECT 11.900 100.100 12.180 100.690 ;
        RECT 13.350 100.100 13.490 102.420 ;
        RECT 11.900 99.960 13.490 100.100 ;
        RECT 17.030 100.100 17.170 110.920 ;
        RECT 22.090 109.540 22.230 111.600 ;
        RECT 27.150 111.240 27.290 116.360 ;
        RECT 28.530 116.340 28.670 119.420 ;
        RECT 28.990 118.720 29.130 121.800 ;
        RECT 29.910 120.080 30.050 133.020 ;
        RECT 30.310 132.000 30.570 132.320 ;
        RECT 30.370 129.940 30.510 132.000 ;
        RECT 30.830 131.210 30.970 135.740 ;
        RECT 31.230 135.060 31.490 135.380 ;
        RECT 31.290 134.020 31.430 135.060 ;
        RECT 31.230 133.700 31.490 134.020 ;
        RECT 31.230 131.210 31.490 131.300 ;
        RECT 30.830 131.070 31.490 131.210 ;
        RECT 31.230 130.980 31.490 131.070 ;
        RECT 30.770 130.300 31.030 130.620 ;
        RECT 30.310 129.620 30.570 129.940 ;
        RECT 30.310 126.900 30.570 127.220 ;
        RECT 30.370 124.160 30.510 126.900 ;
        RECT 30.830 124.500 30.970 130.300 ;
        RECT 31.290 127.220 31.430 130.980 ;
        RECT 31.230 126.900 31.490 127.220 ;
        RECT 30.770 124.180 31.030 124.500 ;
        RECT 30.310 123.840 30.570 124.160 ;
        RECT 31.230 123.840 31.490 124.160 ;
        RECT 31.290 123.140 31.430 123.840 ;
        RECT 31.230 122.820 31.490 123.140 ;
        RECT 31.750 122.540 31.890 144.580 ;
        RECT 33.990 142.880 34.250 143.200 ;
        RECT 34.050 142.180 34.190 142.880 ;
        RECT 33.990 141.860 34.250 142.180 ;
        RECT 33.070 141.520 33.330 141.840 ;
        RECT 32.610 138.120 32.870 138.440 ;
        RECT 32.670 131.300 32.810 138.120 ;
        RECT 32.610 130.980 32.870 131.300 ;
        RECT 32.670 128.580 32.810 130.980 ;
        RECT 32.610 128.260 32.870 128.580 ;
        RECT 30.370 122.400 31.890 122.540 ;
        RECT 29.850 119.760 30.110 120.080 ;
        RECT 28.930 118.400 29.190 118.720 ;
        RECT 28.470 116.020 28.730 116.340 ;
        RECT 29.390 111.600 29.650 111.920 ;
        RECT 27.090 110.920 27.350 111.240 ;
        RECT 25.300 109.705 26.840 110.075 ;
        RECT 22.030 109.220 22.290 109.540 ;
        RECT 19.270 108.200 19.530 108.520 ;
        RECT 22.490 108.200 22.750 108.520 ;
        RECT 19.330 103.080 19.470 108.200 ;
        RECT 22.550 106.480 22.690 108.200 ;
        RECT 22.490 106.160 22.750 106.480 ;
        RECT 26.630 105.710 26.890 105.800 ;
        RECT 27.150 105.710 27.290 110.920 ;
        RECT 29.450 109.540 29.590 111.600 ;
        RECT 30.370 111.580 30.510 122.400 ;
        RECT 30.770 121.800 31.030 122.120 ;
        RECT 30.830 117.700 30.970 121.800 ;
        RECT 31.690 119.420 31.950 119.740 ;
        RECT 31.230 118.400 31.490 118.720 ;
        RECT 30.770 117.380 31.030 117.700 ;
        RECT 31.290 117.020 31.430 118.400 ;
        RECT 31.750 117.360 31.890 119.420 ;
        RECT 31.690 117.040 31.950 117.360 ;
        RECT 31.230 116.700 31.490 117.020 ;
        RECT 31.690 112.960 31.950 113.280 ;
        RECT 30.310 111.260 30.570 111.580 ;
        RECT 30.770 110.240 31.030 110.560 ;
        RECT 31.230 110.240 31.490 110.560 ;
        RECT 29.390 109.220 29.650 109.540 ;
        RECT 29.390 108.770 29.650 108.860 ;
        RECT 29.390 108.630 30.050 108.770 ;
        RECT 29.390 108.540 29.650 108.630 ;
        RECT 26.630 105.570 27.290 105.710 ;
        RECT 26.630 105.480 26.890 105.570 ;
        RECT 23.870 104.800 24.130 105.120 ;
        RECT 19.270 102.760 19.530 103.080 ;
        RECT 23.930 100.690 24.070 104.800 ;
        RECT 25.300 104.265 26.840 104.635 ;
        RECT 27.150 102.400 27.290 105.570 ;
        RECT 27.090 102.080 27.350 102.400 ;
        RECT 29.910 100.690 30.050 108.630 ;
        RECT 30.830 108.180 30.970 110.240 ;
        RECT 30.770 107.860 31.030 108.180 ;
        RECT 31.290 106.820 31.430 110.240 ;
        RECT 31.230 106.500 31.490 106.820 ;
        RECT 31.750 103.420 31.890 112.960 ;
        RECT 33.130 111.580 33.270 141.520 ;
        RECT 33.530 140.840 33.790 141.160 ;
        RECT 33.590 139.120 33.730 140.840 ;
        RECT 33.990 140.160 34.250 140.480 ;
        RECT 33.530 138.800 33.790 139.120 ;
        RECT 34.050 111.580 34.190 140.160 ;
        RECT 34.510 130.280 34.650 161.920 ;
        RECT 34.970 161.220 35.110 162.600 ;
        RECT 36.350 161.980 36.490 164.445 ;
        RECT 36.810 162.920 36.950 166.000 ;
        RECT 37.210 165.320 37.470 165.640 ;
        RECT 37.270 162.920 37.410 165.320 ;
        RECT 37.670 164.640 37.930 164.960 ;
        RECT 36.750 162.600 37.010 162.920 ;
        RECT 37.210 162.600 37.470 162.920 ;
        RECT 36.350 161.840 36.950 161.980 ;
        RECT 34.910 160.900 35.170 161.220 ;
        RECT 35.830 157.840 36.090 158.160 ;
        RECT 35.370 154.100 35.630 154.420 ;
        RECT 34.910 153.760 35.170 154.080 ;
        RECT 34.970 148.980 35.110 153.760 ;
        RECT 34.910 148.660 35.170 148.980 ;
        RECT 34.910 141.860 35.170 142.180 ;
        RECT 34.970 139.460 35.110 141.860 ;
        RECT 35.430 141.160 35.570 154.100 ;
        RECT 35.370 140.840 35.630 141.160 ;
        RECT 34.910 139.140 35.170 139.460 ;
        RECT 34.450 129.960 34.710 130.280 ;
        RECT 35.890 127.900 36.030 157.840 ;
        RECT 36.290 157.335 36.550 157.480 ;
        RECT 36.280 156.965 36.560 157.335 ;
        RECT 36.810 156.660 36.950 161.840 ;
        RECT 37.210 160.220 37.470 160.540 ;
        RECT 37.270 158.500 37.410 160.220 ;
        RECT 37.210 158.180 37.470 158.500 ;
        RECT 37.270 157.480 37.410 158.180 ;
        RECT 37.210 157.160 37.470 157.480 ;
        RECT 36.350 156.520 36.950 156.660 ;
        RECT 36.350 141.500 36.490 156.520 ;
        RECT 37.210 156.480 37.470 156.800 ;
        RECT 36.750 154.780 37.010 155.100 ;
        RECT 36.810 152.380 36.950 154.780 ;
        RECT 36.750 152.060 37.010 152.380 ;
        RECT 36.750 144.240 37.010 144.560 ;
        RECT 36.810 143.735 36.950 144.240 ;
        RECT 36.740 143.365 37.020 143.735 ;
        RECT 37.270 141.500 37.410 156.480 ;
        RECT 37.730 148.380 37.870 164.640 ;
        RECT 38.190 157.480 38.330 183.600 ;
        RECT 39.560 183.145 41.100 183.515 ;
        RECT 42.790 181.960 42.930 183.680 ;
        RECT 43.710 182.640 43.850 184.700 ;
        RECT 45.490 183.680 45.750 184.000 ;
        RECT 43.650 182.320 43.910 182.640 ;
        RECT 41.350 181.640 41.610 181.960 ;
        RECT 42.730 181.640 42.990 181.960 ;
        RECT 41.410 179.240 41.550 181.640 ;
        RECT 41.350 178.920 41.610 179.240 ;
        RECT 39.560 177.705 41.100 178.075 ;
        RECT 39.560 172.265 41.100 172.635 ;
        RECT 39.050 168.720 39.310 169.040 ;
        RECT 39.110 168.360 39.250 168.720 ;
        RECT 39.050 168.040 39.310 168.360 ;
        RECT 39.560 166.825 41.100 167.195 ;
        RECT 39.970 166.340 40.230 166.660 ;
        RECT 40.890 166.340 41.150 166.660 ;
        RECT 40.030 165.980 40.170 166.340 ;
        RECT 40.950 165.980 41.090 166.340 ;
        RECT 39.970 165.660 40.230 165.980 ;
        RECT 40.890 165.660 41.150 165.980 ;
        RECT 38.590 164.640 38.850 164.960 ;
        RECT 38.130 157.160 38.390 157.480 ;
        RECT 38.650 156.800 38.790 164.640 ;
        RECT 39.050 162.260 39.310 162.580 ;
        RECT 39.110 157.335 39.250 162.260 ;
        RECT 39.560 161.385 41.100 161.755 ;
        RECT 41.410 160.880 41.550 178.920 ;
        RECT 43.190 170.760 43.450 171.080 ;
        RECT 43.250 169.380 43.390 170.760 ;
        RECT 43.190 169.060 43.450 169.380 ;
        RECT 41.810 162.600 42.070 162.920 ;
        RECT 41.350 160.560 41.610 160.880 ;
        RECT 39.510 159.880 39.770 160.200 ;
        RECT 39.570 157.820 39.710 159.880 ;
        RECT 39.970 159.375 40.230 159.520 ;
        RECT 39.960 159.005 40.240 159.375 ;
        RECT 39.510 157.500 39.770 157.820 ;
        RECT 39.040 156.965 39.320 157.335 ;
        RECT 38.590 156.480 38.850 156.800 ;
        RECT 39.560 155.945 41.100 156.315 ;
        RECT 38.130 153.760 38.390 154.080 ;
        RECT 38.190 152.040 38.330 153.760 ;
        RECT 41.870 152.040 42.010 162.600 ;
        RECT 42.270 160.220 42.530 160.540 ;
        RECT 42.330 157.480 42.470 160.220 ;
        RECT 43.710 157.480 43.850 182.320 ;
        RECT 45.550 182.300 45.690 183.680 ;
        RECT 47.390 182.980 47.530 187.080 ;
        RECT 47.790 184.700 48.050 185.020 ;
        RECT 47.330 182.660 47.590 182.980 ;
        RECT 45.490 181.980 45.750 182.300 ;
        RECT 47.330 181.980 47.590 182.300 ;
        RECT 47.390 179.240 47.530 181.980 ;
        RECT 47.850 181.960 47.990 184.700 ;
        RECT 48.250 183.680 48.510 184.000 ;
        RECT 48.310 182.980 48.450 183.680 ;
        RECT 50.610 182.980 50.750 187.510 ;
        RECT 51.010 187.420 51.270 187.510 ;
        RECT 57.510 187.400 57.650 195.240 ;
        RECT 59.750 194.900 60.010 195.220 ;
        RECT 59.810 188.420 59.950 194.900 ;
        RECT 63.030 193.180 63.170 195.580 ;
        RECT 63.430 194.900 63.690 195.220 ;
        RECT 63.490 193.860 63.630 194.900 ;
        RECT 63.430 193.540 63.690 193.860 ;
        RECT 64.870 193.180 65.010 197.280 ;
        RECT 65.330 196.580 65.470 198.640 ;
        RECT 71.710 197.960 71.970 198.280 ;
        RECT 71.250 197.280 71.510 197.600 ;
        RECT 65.270 196.260 65.530 196.580 ;
        RECT 69.870 194.560 70.130 194.880 ;
        RECT 68.080 194.025 69.620 194.395 ;
        RECT 69.930 193.180 70.070 194.560 ;
        RECT 71.310 193.860 71.450 197.280 ;
        RECT 71.770 196.240 71.910 197.960 ;
        RECT 82.340 196.745 83.880 197.115 ;
        RECT 110.860 196.745 112.400 197.115 ;
        RECT 71.710 195.920 71.970 196.240 ;
        RECT 71.250 193.540 71.510 193.860 ;
        RECT 62.970 192.860 63.230 193.180 ;
        RECT 64.810 192.860 65.070 193.180 ;
        RECT 67.110 192.860 67.370 193.180 ;
        RECT 69.870 193.090 70.130 193.180 ;
        RECT 69.870 192.950 70.530 193.090 ;
        RECT 69.870 192.860 70.130 192.950 ;
        RECT 59.750 188.100 60.010 188.420 ;
        RECT 57.450 187.080 57.710 187.400 ;
        RECT 51.010 186.400 51.270 186.720 ;
        RECT 53.310 186.400 53.570 186.720 ;
        RECT 55.610 186.400 55.870 186.720 ;
        RECT 51.070 184.680 51.210 186.400 ;
        RECT 53.370 185.020 53.510 186.400 ;
        RECT 53.820 185.865 55.360 186.235 ;
        RECT 53.310 184.700 53.570 185.020 ;
        RECT 51.010 184.360 51.270 184.680 ;
        RECT 48.250 182.660 48.510 182.980 ;
        RECT 50.550 182.660 50.810 182.980 ;
        RECT 55.670 182.640 55.810 186.400 ;
        RECT 57.510 184.680 57.650 187.080 ;
        RECT 63.030 184.680 63.170 192.860 ;
        RECT 64.870 190.120 65.010 192.860 ;
        RECT 65.730 190.140 65.990 190.460 ;
        RECT 64.810 189.800 65.070 190.120 ;
        RECT 65.790 187.400 65.930 190.140 ;
        RECT 65.730 187.080 65.990 187.400 ;
        RECT 66.190 184.700 66.450 185.020 ;
        RECT 57.450 184.360 57.710 184.680 ;
        RECT 60.670 184.360 60.930 184.680 ;
        RECT 62.510 184.360 62.770 184.680 ;
        RECT 62.970 184.360 63.230 184.680 ;
        RECT 55.610 182.320 55.870 182.640 ;
        RECT 60.730 181.960 60.870 184.360 ;
        RECT 62.570 182.640 62.710 184.360 ;
        RECT 62.510 182.320 62.770 182.640 ;
        RECT 47.790 181.640 48.050 181.960 ;
        RECT 58.370 181.640 58.630 181.960 ;
        RECT 60.670 181.640 60.930 181.960 ;
        RECT 47.850 179.580 47.990 181.640 ;
        RECT 53.820 180.425 55.360 180.795 ;
        RECT 58.430 180.260 58.570 181.640 ;
        RECT 58.370 179.940 58.630 180.260 ;
        RECT 47.790 179.260 48.050 179.580 ;
        RECT 58.370 179.260 58.630 179.580 ;
        RECT 47.330 178.920 47.590 179.240 ;
        RECT 45.490 178.240 45.750 178.560 ;
        RECT 45.950 178.240 46.210 178.560 ;
        RECT 45.550 177.540 45.690 178.240 ;
        RECT 45.490 177.220 45.750 177.540 ;
        RECT 45.550 172.860 45.690 177.220 ;
        RECT 46.010 173.800 46.150 178.240 ;
        RECT 46.870 176.200 47.130 176.520 ;
        RECT 46.930 174.820 47.070 176.200 ;
        RECT 46.870 174.500 47.130 174.820 ;
        RECT 45.950 173.480 46.210 173.800 ;
        RECT 45.550 172.720 46.610 172.860 ;
        RECT 45.030 168.380 45.290 168.700 ;
        RECT 44.570 165.660 44.830 165.980 ;
        RECT 44.630 165.300 44.770 165.660 ;
        RECT 44.570 164.980 44.830 165.300 ;
        RECT 45.090 163.260 45.230 168.380 ;
        RECT 46.470 168.360 46.610 172.720 ;
        RECT 46.870 171.100 47.130 171.420 ;
        RECT 46.410 168.040 46.670 168.360 ;
        RECT 45.490 166.340 45.750 166.660 ;
        RECT 45.550 165.980 45.690 166.340 ;
        RECT 45.490 165.660 45.750 165.980 ;
        RECT 45.950 164.815 46.210 164.960 ;
        RECT 45.940 164.445 46.220 164.815 ;
        RECT 45.030 162.940 45.290 163.260 ;
        RECT 45.950 159.540 46.210 159.860 ;
        RECT 46.010 157.480 46.150 159.540 ;
        RECT 42.270 157.160 42.530 157.480 ;
        RECT 43.650 157.160 43.910 157.480 ;
        RECT 45.950 157.160 46.210 157.480 ;
        RECT 42.330 155.440 42.470 157.160 ;
        RECT 45.490 156.820 45.750 157.140 ;
        RECT 42.730 156.480 42.990 156.800 ;
        RECT 44.570 156.480 44.830 156.800 ;
        RECT 42.270 155.120 42.530 155.440 ;
        RECT 42.270 153.760 42.530 154.080 ;
        RECT 38.130 151.720 38.390 152.040 ;
        RECT 41.810 151.895 42.070 152.040 ;
        RECT 41.350 151.380 41.610 151.700 ;
        RECT 41.800 151.525 42.080 151.895 ;
        RECT 39.560 150.505 41.100 150.875 ;
        RECT 40.430 149.340 40.690 149.660 ;
        RECT 40.890 149.570 41.150 149.660 ;
        RECT 41.410 149.570 41.550 151.380 ;
        RECT 41.870 149.660 42.010 151.525 ;
        RECT 40.890 149.430 41.550 149.570 ;
        RECT 40.890 149.340 41.150 149.430 ;
        RECT 41.810 149.340 42.070 149.660 ;
        RECT 37.730 148.240 38.330 148.380 ;
        RECT 38.590 148.320 38.850 148.640 ;
        RECT 38.190 144.220 38.330 148.240 ;
        RECT 38.130 143.900 38.390 144.220 ;
        RECT 37.670 141.860 37.930 142.180 ;
        RECT 36.290 141.180 36.550 141.500 ;
        RECT 37.210 141.180 37.470 141.500 ;
        RECT 37.730 139.460 37.870 141.860 ;
        RECT 38.130 141.520 38.390 141.840 ;
        RECT 38.190 141.160 38.330 141.520 ;
        RECT 38.130 140.840 38.390 141.160 ;
        RECT 37.670 139.140 37.930 139.460 ;
        RECT 38.130 137.440 38.390 137.760 ;
        RECT 38.190 135.720 38.330 137.440 ;
        RECT 38.130 135.400 38.390 135.720 ;
        RECT 38.130 129.620 38.390 129.940 ;
        RECT 35.830 127.580 36.090 127.900 ;
        RECT 38.190 127.220 38.330 129.620 ;
        RECT 38.650 127.900 38.790 148.320 ;
        RECT 40.490 146.600 40.630 149.340 ;
        RECT 40.890 148.660 41.150 148.980 ;
        RECT 41.350 148.660 41.610 148.980 ;
        RECT 40.950 146.940 41.090 148.660 ;
        RECT 40.890 146.620 41.150 146.940 ;
        RECT 40.430 146.280 40.690 146.600 ;
        RECT 39.050 145.600 39.310 145.920 ;
        RECT 39.110 128.150 39.250 145.600 ;
        RECT 39.560 145.065 41.100 145.435 ;
        RECT 41.410 144.810 41.550 148.660 ;
        RECT 41.870 146.600 42.010 149.340 ;
        RECT 41.810 146.280 42.070 146.600 ;
        RECT 40.950 144.670 41.550 144.810 ;
        RECT 40.950 143.540 41.090 144.670 ;
        RECT 41.340 144.045 41.620 144.415 ;
        RECT 41.350 143.900 41.610 144.045 ;
        RECT 40.890 143.220 41.150 143.540 ;
        RECT 41.810 142.880 42.070 143.200 ;
        RECT 41.870 142.180 42.010 142.880 ;
        RECT 41.810 141.860 42.070 142.180 ;
        RECT 39.970 141.180 40.230 141.500 ;
        RECT 40.030 140.480 40.170 141.180 ;
        RECT 41.810 140.840 42.070 141.160 ;
        RECT 39.970 140.160 40.230 140.480 ;
        RECT 39.560 139.625 41.100 139.995 ;
        RECT 41.870 138.780 42.010 140.840 ;
        RECT 41.810 138.460 42.070 138.780 ;
        RECT 39.560 134.185 41.100 134.555 ;
        RECT 41.870 132.660 42.010 138.460 ;
        RECT 41.810 132.340 42.070 132.660 ;
        RECT 41.350 132.000 41.610 132.320 ;
        RECT 41.410 131.300 41.550 132.000 ;
        RECT 41.350 130.980 41.610 131.300 ;
        RECT 42.330 130.700 42.470 153.760 ;
        RECT 42.790 133.340 42.930 156.480 ;
        RECT 44.110 151.380 44.370 151.700 ;
        RECT 43.650 151.040 43.910 151.360 ;
        RECT 43.190 149.340 43.450 149.660 ;
        RECT 43.250 147.620 43.390 149.340 ;
        RECT 43.190 147.300 43.450 147.620 ;
        RECT 43.190 145.600 43.450 145.920 ;
        RECT 43.250 144.560 43.390 145.600 ;
        RECT 43.190 144.240 43.450 144.560 ;
        RECT 43.190 143.735 43.450 143.880 ;
        RECT 43.180 143.365 43.460 143.735 ;
        RECT 43.190 137.440 43.450 137.760 ;
        RECT 43.250 134.020 43.390 137.440 ;
        RECT 43.190 133.700 43.450 134.020 ;
        RECT 42.730 133.020 42.990 133.340 ;
        RECT 43.190 132.680 43.450 133.000 ;
        RECT 43.250 131.300 43.390 132.680 ;
        RECT 43.190 130.980 43.450 131.300 ;
        RECT 41.410 130.560 42.470 130.700 ;
        RECT 39.560 128.745 41.100 129.115 ;
        RECT 39.110 128.010 39.710 128.150 ;
        RECT 38.590 127.580 38.850 127.900 ;
        RECT 38.130 126.900 38.390 127.220 ;
        RECT 37.670 126.560 37.930 126.880 ;
        RECT 39.050 126.560 39.310 126.880 ;
        RECT 34.910 122.480 35.170 122.800 ;
        RECT 34.970 120.080 35.110 122.480 ;
        RECT 34.910 119.760 35.170 120.080 ;
        RECT 37.730 112.260 37.870 126.560 ;
        RECT 38.120 125.005 38.400 125.375 ;
        RECT 38.190 124.840 38.330 125.005 ;
        RECT 38.130 124.520 38.390 124.840 ;
        RECT 38.190 123.140 38.330 124.520 ;
        RECT 39.110 123.140 39.250 126.560 ;
        RECT 39.570 125.180 39.710 128.010 ;
        RECT 39.970 127.580 40.230 127.900 ;
        RECT 40.030 127.415 40.170 127.580 ;
        RECT 39.960 127.045 40.240 127.415 ;
        RECT 39.510 124.860 39.770 125.180 ;
        RECT 41.410 124.840 41.550 130.560 ;
        RECT 41.810 129.620 42.070 129.940 ;
        RECT 41.870 128.580 42.010 129.620 ;
        RECT 42.270 129.280 42.530 129.600 ;
        RECT 41.810 128.260 42.070 128.580 ;
        RECT 41.800 127.725 42.080 128.095 ;
        RECT 41.810 127.580 42.070 127.725 ;
        RECT 41.350 124.520 41.610 124.840 ;
        RECT 39.560 123.305 41.100 123.675 ;
        RECT 38.130 122.820 38.390 123.140 ;
        RECT 39.050 122.820 39.310 123.140 ;
        RECT 41.350 122.820 41.610 123.140 ;
        RECT 41.410 122.460 41.550 122.820 ;
        RECT 38.130 122.140 38.390 122.460 ;
        RECT 38.590 122.140 38.850 122.460 ;
        RECT 41.350 122.140 41.610 122.460 ;
        RECT 38.190 117.100 38.330 122.140 ;
        RECT 38.650 117.700 38.790 122.140 ;
        RECT 41.810 121.800 42.070 122.120 ;
        RECT 41.350 121.460 41.610 121.780 ;
        RECT 39.050 121.120 39.310 121.440 ;
        RECT 39.110 119.740 39.250 121.120 ;
        RECT 39.050 119.420 39.310 119.740 ;
        RECT 41.410 119.400 41.550 121.460 ;
        RECT 41.350 119.080 41.610 119.400 ;
        RECT 39.560 117.865 41.100 118.235 ;
        RECT 38.590 117.380 38.850 117.700 ;
        RECT 38.190 116.960 38.790 117.100 ;
        RECT 38.650 113.620 38.790 116.960 ;
        RECT 38.590 113.300 38.850 113.620 ;
        RECT 37.670 111.940 37.930 112.260 ;
        RECT 37.210 111.600 37.470 111.920 ;
        RECT 33.070 111.260 33.330 111.580 ;
        RECT 33.990 111.260 34.250 111.580 ;
        RECT 34.450 110.240 34.710 110.560 ;
        RECT 34.510 108.860 34.650 110.240 ;
        RECT 34.450 108.540 34.710 108.860 ;
        RECT 37.270 106.140 37.410 111.600 ;
        RECT 38.650 111.580 38.790 113.300 ;
        RECT 39.560 112.425 41.100 112.795 ;
        RECT 38.590 111.260 38.850 111.580 ;
        RECT 41.410 111.240 41.550 119.080 ;
        RECT 41.870 117.020 42.010 121.800 ;
        RECT 41.810 116.700 42.070 117.020 ;
        RECT 42.330 111.580 42.470 129.280 ;
        RECT 42.720 128.405 43.000 128.775 ;
        RECT 42.790 124.840 42.930 128.405 ;
        RECT 43.250 125.860 43.390 130.980 ;
        RECT 43.190 125.540 43.450 125.860 ;
        RECT 42.730 124.520 42.990 124.840 ;
        RECT 42.730 123.840 42.990 124.160 ;
        RECT 42.790 111.580 42.930 123.840 ;
        RECT 43.250 123.140 43.390 125.540 ;
        RECT 43.710 125.180 43.850 151.040 ;
        RECT 44.170 149.660 44.310 151.380 ;
        RECT 44.110 149.340 44.370 149.660 ;
        RECT 44.170 147.280 44.310 149.340 ;
        RECT 44.110 146.960 44.370 147.280 ;
        RECT 44.110 146.280 44.370 146.600 ;
        RECT 44.170 144.220 44.310 146.280 ;
        RECT 44.110 143.900 44.370 144.220 ;
        RECT 44.630 138.440 44.770 156.480 ;
        RECT 45.550 155.100 45.690 156.820 ;
        RECT 46.010 155.780 46.150 157.160 ;
        RECT 45.950 155.460 46.210 155.780 ;
        RECT 46.470 155.100 46.610 168.040 ;
        RECT 46.930 167.680 47.070 171.100 ;
        RECT 46.870 167.360 47.130 167.680 ;
        RECT 46.930 156.800 47.070 167.360 ;
        RECT 47.390 157.480 47.530 178.920 ;
        RECT 53.310 178.240 53.570 178.560 ;
        RECT 53.370 173.120 53.510 178.240 ;
        RECT 56.070 176.540 56.330 176.860 ;
        RECT 53.820 174.985 55.360 175.355 ;
        RECT 55.610 174.050 55.870 174.140 ;
        RECT 56.130 174.050 56.270 176.540 ;
        RECT 56.530 175.520 56.790 175.840 ;
        RECT 55.610 173.910 56.270 174.050 ;
        RECT 55.610 173.820 55.870 173.910 ;
        RECT 51.470 172.800 51.730 173.120 ;
        RECT 53.310 172.800 53.570 173.120 ;
        RECT 56.130 172.860 56.270 173.910 ;
        RECT 56.590 173.460 56.730 175.520 ;
        RECT 56.530 173.140 56.790 173.460 ;
        RECT 51.530 171.760 51.670 172.800 ;
        RECT 53.370 172.100 53.510 172.800 ;
        RECT 56.130 172.720 56.730 172.860 ;
        RECT 53.310 171.780 53.570 172.100 ;
        RECT 51.470 171.440 51.730 171.760 ;
        RECT 52.850 171.330 53.110 171.420 ;
        RECT 52.450 171.190 53.110 171.330 ;
        RECT 52.450 169.380 52.590 171.190 ;
        RECT 52.850 171.100 53.110 171.190 ;
        RECT 52.390 169.060 52.650 169.380 ;
        RECT 48.250 168.040 48.510 168.360 ;
        RECT 48.310 165.980 48.450 168.040 ;
        RECT 53.370 167.420 53.510 171.780 ;
        RECT 53.820 169.545 55.360 169.915 ;
        RECT 55.610 169.060 55.870 169.380 ;
        RECT 52.450 167.280 53.510 167.420 ;
        RECT 55.150 167.360 55.410 167.680 ;
        RECT 48.250 165.660 48.510 165.980 ;
        RECT 52.450 164.700 52.590 167.280 ;
        RECT 52.850 166.340 53.110 166.660 ;
        RECT 52.910 165.380 53.050 166.340 ;
        RECT 55.210 166.320 55.350 167.360 ;
        RECT 55.150 166.000 55.410 166.320 ;
        RECT 54.230 165.890 54.490 165.980 ;
        RECT 54.230 165.750 54.890 165.890 ;
        RECT 54.230 165.660 54.490 165.750 ;
        RECT 54.750 165.550 54.890 165.750 ;
        RECT 55.670 165.550 55.810 169.060 ;
        RECT 56.590 168.360 56.730 172.720 ;
        RECT 57.450 171.100 57.710 171.420 ;
        RECT 56.530 168.040 56.790 168.360 ;
        RECT 54.750 165.410 55.810 165.550 ;
        RECT 52.910 165.240 53.510 165.380 ;
        RECT 52.450 164.560 53.050 164.700 ;
        RECT 52.390 162.940 52.650 163.260 ;
        RECT 47.790 162.260 48.050 162.580 ;
        RECT 47.850 160.880 47.990 162.260 ;
        RECT 47.790 160.560 48.050 160.880 ;
        RECT 48.240 160.365 48.520 160.735 ;
        RECT 47.330 157.160 47.590 157.480 ;
        RECT 47.790 157.160 48.050 157.480 ;
        RECT 46.870 156.480 47.130 156.800 ;
        RECT 47.850 155.100 47.990 157.160 ;
        RECT 48.310 157.140 48.450 160.365 ;
        RECT 52.450 159.520 52.590 162.940 ;
        RECT 50.090 159.200 50.350 159.520 ;
        RECT 52.390 159.200 52.650 159.520 ;
        RECT 48.250 156.820 48.510 157.140 ;
        RECT 49.630 156.480 49.890 156.800 ;
        RECT 49.690 155.100 49.830 156.480 ;
        RECT 45.490 154.780 45.750 155.100 ;
        RECT 46.410 154.780 46.670 155.100 ;
        RECT 47.790 154.780 48.050 155.100 ;
        RECT 49.630 154.780 49.890 155.100 ;
        RECT 47.330 153.760 47.590 154.080 ;
        RECT 46.410 151.380 46.670 151.700 ;
        RECT 45.490 151.040 45.750 151.360 ;
        RECT 45.550 149.660 45.690 151.040 ;
        RECT 45.490 149.340 45.750 149.660 ;
        RECT 45.030 148.320 45.290 148.640 ;
        RECT 45.090 138.780 45.230 148.320 ;
        RECT 45.550 146.600 45.690 149.340 ;
        RECT 45.490 146.280 45.750 146.600 ;
        RECT 45.490 145.600 45.750 145.920 ;
        RECT 45.030 138.460 45.290 138.780 ;
        RECT 44.570 138.120 44.830 138.440 ;
        RECT 45.550 133.000 45.690 145.600 ;
        RECT 46.470 141.840 46.610 151.380 ;
        RECT 46.870 143.220 47.130 143.540 ;
        RECT 46.410 141.520 46.670 141.840 ;
        RECT 46.930 141.500 47.070 143.220 ;
        RECT 46.870 141.180 47.130 141.500 ;
        RECT 45.490 132.680 45.750 133.000 ;
        RECT 45.950 132.680 46.210 133.000 ;
        RECT 46.010 130.280 46.150 132.680 ;
        RECT 47.390 130.620 47.530 153.760 ;
        RECT 50.150 143.200 50.290 159.200 ;
        RECT 52.450 157.820 52.590 159.200 ;
        RECT 52.390 157.500 52.650 157.820 ;
        RECT 51.470 155.460 51.730 155.780 ;
        RECT 51.530 155.100 51.670 155.460 ;
        RECT 51.470 154.780 51.730 155.100 ;
        RECT 52.390 154.780 52.650 155.100 ;
        RECT 51.530 154.420 51.670 154.780 ;
        RECT 51.930 154.440 52.190 154.760 ;
        RECT 51.470 154.100 51.730 154.420 ;
        RECT 50.550 152.400 50.810 152.720 ;
        RECT 50.610 143.620 50.750 152.400 ;
        RECT 51.990 152.380 52.130 154.440 ;
        RECT 52.450 153.060 52.590 154.780 ;
        RECT 52.390 152.740 52.650 153.060 ;
        RECT 51.930 152.060 52.190 152.380 ;
        RECT 51.990 151.780 52.130 152.060 ;
        RECT 52.450 152.040 52.590 152.740 ;
        RECT 51.530 151.640 52.130 151.780 ;
        RECT 52.390 151.720 52.650 152.040 ;
        RECT 51.530 149.660 51.670 151.640 ;
        RECT 51.470 149.340 51.730 149.660 ;
        RECT 52.450 149.320 52.590 151.720 ;
        RECT 52.910 150.340 53.050 164.560 ;
        RECT 53.370 163.340 53.510 165.240 ;
        RECT 53.820 164.105 55.360 164.475 ;
        RECT 53.370 163.260 53.970 163.340 ;
        RECT 53.310 163.200 53.970 163.260 ;
        RECT 53.310 162.940 53.570 163.200 ;
        RECT 53.310 162.260 53.570 162.580 ;
        RECT 53.370 161.220 53.510 162.260 ;
        RECT 53.310 160.900 53.570 161.220 ;
        RECT 53.370 157.900 53.510 160.900 ;
        RECT 53.830 160.540 53.970 163.200 ;
        RECT 53.770 160.220 54.030 160.540 ;
        RECT 54.220 160.365 54.500 160.735 ;
        RECT 55.670 160.540 55.810 165.410 ;
        RECT 54.290 160.200 54.430 160.365 ;
        RECT 55.610 160.220 55.870 160.540 ;
        RECT 54.230 159.880 54.490 160.200 ;
        RECT 56.070 159.880 56.330 160.200 ;
        RECT 56.130 159.520 56.270 159.880 ;
        RECT 56.070 159.200 56.330 159.520 ;
        RECT 53.820 158.665 55.360 159.035 ;
        RECT 53.370 157.820 53.970 157.900 ;
        RECT 53.310 157.760 53.970 157.820 ;
        RECT 53.310 157.500 53.570 157.760 ;
        RECT 53.310 156.820 53.570 157.140 ;
        RECT 53.370 152.040 53.510 156.820 ;
        RECT 53.830 155.100 53.970 157.760 ;
        RECT 56.590 156.660 56.730 168.040 ;
        RECT 57.510 166.660 57.650 171.100 ;
        RECT 58.430 171.080 58.570 179.260 ;
        RECT 60.730 176.520 60.870 181.640 ;
        RECT 63.030 179.580 63.170 184.360 ;
        RECT 66.250 181.280 66.390 184.700 ;
        RECT 67.170 184.680 67.310 192.860 ;
        RECT 69.410 192.520 69.670 192.840 ;
        RECT 67.570 191.840 67.830 192.160 ;
        RECT 67.630 188.420 67.770 191.840 ;
        RECT 69.470 190.800 69.610 192.520 ;
        RECT 69.870 192.180 70.130 192.500 ;
        RECT 69.930 190.800 70.070 192.180 ;
        RECT 69.410 190.480 69.670 190.800 ;
        RECT 69.870 190.480 70.130 190.800 ;
        RECT 69.470 190.120 69.610 190.480 ;
        RECT 69.410 189.800 69.670 190.120 ;
        RECT 68.080 188.585 69.620 188.955 ;
        RECT 67.570 188.100 67.830 188.420 ;
        RECT 69.930 187.400 70.070 190.480 ;
        RECT 70.390 189.780 70.530 192.950 ;
        RECT 70.790 190.820 71.050 191.140 ;
        RECT 70.330 189.460 70.590 189.780 ;
        RECT 70.390 188.420 70.530 189.460 ;
        RECT 70.330 188.100 70.590 188.420 ;
        RECT 69.870 187.080 70.130 187.400 ;
        RECT 70.330 187.080 70.590 187.400 ;
        RECT 69.870 186.400 70.130 186.720 ;
        RECT 69.930 185.360 70.070 186.400 ;
        RECT 70.390 185.700 70.530 187.080 ;
        RECT 70.330 185.380 70.590 185.700 ;
        RECT 69.870 185.040 70.130 185.360 ;
        RECT 67.110 184.360 67.370 184.680 ;
        RECT 68.080 183.145 69.620 183.515 ;
        RECT 66.190 180.960 66.450 181.280 ;
        RECT 67.110 180.960 67.370 181.280 ;
        RECT 62.970 179.260 63.230 179.580 ;
        RECT 64.350 178.920 64.610 179.240 ;
        RECT 60.670 176.200 60.930 176.520 ;
        RECT 60.730 173.800 60.870 176.200 ;
        RECT 64.410 176.180 64.550 178.920 ;
        RECT 64.350 175.860 64.610 176.180 ;
        RECT 61.590 174.160 61.850 174.480 ;
        RECT 59.750 173.480 60.010 173.800 ;
        RECT 60.670 173.480 60.930 173.800 ;
        RECT 59.810 172.100 59.950 173.480 ;
        RECT 60.730 172.100 60.870 173.480 ;
        RECT 59.750 171.780 60.010 172.100 ;
        RECT 60.670 171.780 60.930 172.100 ;
        RECT 58.370 170.760 58.630 171.080 ;
        RECT 58.430 166.660 58.570 170.760 ;
        RECT 60.210 170.080 60.470 170.400 ;
        RECT 60.270 168.020 60.410 170.080 ;
        RECT 60.210 167.700 60.470 168.020 ;
        RECT 57.450 166.340 57.710 166.660 ;
        RECT 58.370 166.340 58.630 166.660 ;
        RECT 57.450 162.260 57.710 162.580 ;
        RECT 56.990 161.920 57.250 162.240 ;
        RECT 57.050 157.820 57.190 161.920 ;
        RECT 56.990 157.500 57.250 157.820 ;
        RECT 57.050 157.140 57.190 157.500 ;
        RECT 56.990 156.820 57.250 157.140 ;
        RECT 56.590 156.520 57.190 156.660 ;
        RECT 57.050 155.100 57.190 156.520 ;
        RECT 57.510 155.780 57.650 162.260 ;
        RECT 58.430 160.540 58.570 166.340 ;
        RECT 60.210 166.000 60.470 166.320 ;
        RECT 59.750 165.550 60.010 165.640 ;
        RECT 60.270 165.550 60.410 166.000 ;
        RECT 60.730 165.640 60.870 171.780 ;
        RECT 59.750 165.410 60.410 165.550 ;
        RECT 59.750 165.320 60.010 165.410 ;
        RECT 60.670 165.320 60.930 165.640 ;
        RECT 60.730 163.260 60.870 165.320 ;
        RECT 60.670 162.940 60.930 163.260 ;
        RECT 60.730 160.880 60.870 162.940 ;
        RECT 60.670 160.560 60.930 160.880 ;
        RECT 58.370 160.220 58.630 160.540 ;
        RECT 57.910 159.880 58.170 160.200 ;
        RECT 57.970 157.820 58.110 159.880 ;
        RECT 57.910 157.500 58.170 157.820 ;
        RECT 58.830 156.820 59.090 157.140 ;
        RECT 58.890 155.780 59.030 156.820 ;
        RECT 59.290 156.480 59.550 156.800 ;
        RECT 57.450 155.460 57.710 155.780 ;
        RECT 58.830 155.460 59.090 155.780 ;
        RECT 59.350 155.100 59.490 156.480 ;
        RECT 53.770 154.780 54.030 155.100 ;
        RECT 55.610 154.780 55.870 155.100 ;
        RECT 56.990 154.780 57.250 155.100 ;
        RECT 59.290 154.780 59.550 155.100 ;
        RECT 53.820 153.225 55.360 153.595 ;
        RECT 55.670 152.040 55.810 154.780 ;
        RECT 57.050 152.720 57.190 154.780 ;
        RECT 56.990 152.400 57.250 152.720 ;
        RECT 57.450 152.400 57.710 152.720 ;
        RECT 53.310 151.720 53.570 152.040 ;
        RECT 54.230 151.720 54.490 152.040 ;
        RECT 55.610 151.720 55.870 152.040 ;
        RECT 52.850 150.020 53.110 150.340 ;
        RECT 54.290 149.660 54.430 151.720 ;
        RECT 54.230 149.340 54.490 149.660 ;
        RECT 52.390 149.000 52.650 149.320 ;
        RECT 57.510 148.980 57.650 152.400 ;
        RECT 58.830 149.680 59.090 150.000 ;
        RECT 57.450 148.660 57.710 148.980 ;
        RECT 53.820 147.785 55.360 148.155 ;
        RECT 58.890 146.600 59.030 149.680 ;
        RECT 60.670 149.000 60.930 149.320 ;
        RECT 59.290 146.960 59.550 147.280 ;
        RECT 53.770 146.280 54.030 146.600 ;
        RECT 54.690 146.280 54.950 146.600 ;
        RECT 56.530 146.280 56.790 146.600 ;
        RECT 58.370 146.280 58.630 146.600 ;
        RECT 58.830 146.280 59.090 146.600 ;
        RECT 52.390 145.600 52.650 145.920 ;
        RECT 52.450 144.900 52.590 145.600 ;
        RECT 52.390 144.580 52.650 144.900 ;
        RECT 53.830 144.220 53.970 146.280 ;
        RECT 51.930 143.900 52.190 144.220 ;
        RECT 53.770 143.900 54.030 144.220 ;
        RECT 50.610 143.480 51.210 143.620 ;
        RECT 50.090 142.880 50.350 143.200 ;
        RECT 49.630 140.160 49.890 140.480 ;
        RECT 48.240 138.605 48.520 138.975 ;
        RECT 49.690 138.780 49.830 140.160 ;
        RECT 51.070 138.780 51.210 143.480 ;
        RECT 48.250 138.460 48.510 138.605 ;
        RECT 49.630 138.460 49.890 138.780 ;
        RECT 50.550 138.460 50.810 138.780 ;
        RECT 51.010 138.460 51.270 138.780 ;
        RECT 48.310 133.000 48.450 138.460 ;
        RECT 48.710 137.440 48.970 137.760 ;
        RECT 50.090 137.440 50.350 137.760 ;
        RECT 48.250 132.680 48.510 133.000 ;
        RECT 47.330 130.300 47.590 130.620 ;
        RECT 45.950 129.960 46.210 130.280 ;
        RECT 46.870 129.960 47.130 130.280 ;
        RECT 47.790 129.960 48.050 130.280 ;
        RECT 44.570 129.280 44.830 129.600 ;
        RECT 44.110 125.540 44.370 125.860 ;
        RECT 43.650 124.860 43.910 125.180 ;
        RECT 44.170 123.140 44.310 125.540 ;
        RECT 44.630 125.180 44.770 129.280 ;
        RECT 46.010 127.220 46.150 129.960 ;
        RECT 45.950 126.900 46.210 127.220 ;
        RECT 44.570 124.860 44.830 125.180 ;
        RECT 46.010 124.840 46.150 126.900 ;
        RECT 46.410 125.200 46.670 125.520 ;
        RECT 45.950 124.520 46.210 124.840 ;
        RECT 43.190 122.820 43.450 123.140 ;
        RECT 44.110 122.820 44.370 123.140 ;
        RECT 43.250 122.370 43.390 122.820 ;
        RECT 43.650 122.370 43.910 122.460 ;
        RECT 43.250 122.230 43.910 122.370 ;
        RECT 43.650 122.140 43.910 122.230 ;
        RECT 46.470 117.100 46.610 125.200 ;
        RECT 46.930 119.060 47.070 129.960 ;
        RECT 47.850 127.900 47.990 129.960 ;
        RECT 47.790 127.580 48.050 127.900 ;
        RECT 47.850 124.840 47.990 127.580 ;
        RECT 47.790 124.520 48.050 124.840 ;
        RECT 46.870 118.740 47.130 119.060 ;
        RECT 46.930 117.700 47.070 118.740 ;
        RECT 46.870 117.380 47.130 117.700 ;
        RECT 46.470 116.960 47.070 117.100 ;
        RECT 46.410 115.680 46.670 116.000 ;
        RECT 46.470 111.580 46.610 115.680 ;
        RECT 42.270 111.260 42.530 111.580 ;
        RECT 42.730 111.260 42.990 111.580 ;
        RECT 46.410 111.260 46.670 111.580 ;
        RECT 39.050 110.920 39.310 111.240 ;
        RECT 41.350 110.920 41.610 111.240 ;
        RECT 38.590 110.580 38.850 110.900 ;
        RECT 37.210 105.820 37.470 106.140 ;
        RECT 35.830 105.480 36.090 105.800 ;
        RECT 31.690 103.100 31.950 103.420 ;
        RECT 35.890 100.690 36.030 105.480 ;
        RECT 38.650 105.120 38.790 110.580 ;
        RECT 39.110 109.200 39.250 110.920 ;
        RECT 39.970 110.240 40.230 110.560 ;
        RECT 44.570 110.240 44.830 110.560 ;
        RECT 39.050 108.880 39.310 109.200 ;
        RECT 39.110 106.140 39.250 108.880 ;
        RECT 40.030 108.180 40.170 110.240 ;
        RECT 42.730 109.220 42.990 109.540 ;
        RECT 41.810 108.540 42.070 108.860 ;
        RECT 39.970 107.860 40.230 108.180 ;
        RECT 39.560 106.985 41.100 107.355 ;
        RECT 39.050 105.820 39.310 106.140 ;
        RECT 39.510 105.480 39.770 105.800 ;
        RECT 38.590 104.800 38.850 105.120 ;
        RECT 39.570 103.080 39.710 105.480 ;
        RECT 39.510 102.760 39.770 103.080 ;
        RECT 39.560 101.545 41.100 101.915 ;
        RECT 41.870 100.690 42.010 108.540 ;
        RECT 42.790 106.480 42.930 109.220 ;
        RECT 44.630 108.860 44.770 110.240 ;
        RECT 44.570 108.540 44.830 108.860 ;
        RECT 46.930 108.520 47.070 116.960 ;
        RECT 47.790 116.700 48.050 117.020 ;
        RECT 47.850 114.980 47.990 116.700 ;
        RECT 47.790 114.660 48.050 114.980 ;
        RECT 48.250 112.960 48.510 113.280 ;
        RECT 48.310 111.920 48.450 112.960 ;
        RECT 48.250 111.600 48.510 111.920 ;
        RECT 48.770 109.540 48.910 137.440 ;
        RECT 50.150 133.340 50.290 137.440 ;
        RECT 50.610 136.740 50.750 138.460 ;
        RECT 51.990 138.100 52.130 143.900 ;
        RECT 54.750 143.110 54.890 146.280 ;
        RECT 55.150 145.940 55.410 146.260 ;
        RECT 55.210 144.220 55.350 145.940 ;
        RECT 56.590 144.220 56.730 146.280 ;
        RECT 57.910 145.600 58.170 145.920 ;
        RECT 57.970 144.415 58.110 145.600 ;
        RECT 58.430 144.560 58.570 146.280 ;
        RECT 55.150 143.900 55.410 144.220 ;
        RECT 56.530 143.900 56.790 144.220 ;
        RECT 57.900 144.045 58.180 144.415 ;
        RECT 58.370 144.240 58.630 144.560 ;
        RECT 57.450 143.560 57.710 143.880 ;
        RECT 54.750 142.970 55.810 143.110 ;
        RECT 53.820 142.345 55.360 142.715 ;
        RECT 52.390 140.500 52.650 140.820 ;
        RECT 52.450 139.460 52.590 140.500 ;
        RECT 55.670 139.460 55.810 142.970 ;
        RECT 56.070 142.880 56.330 143.200 ;
        RECT 56.130 141.500 56.270 142.880 ;
        RECT 56.070 141.180 56.330 141.500 ;
        RECT 52.390 139.140 52.650 139.460 ;
        RECT 55.610 139.140 55.870 139.460 ;
        RECT 52.390 138.460 52.650 138.780 ;
        RECT 51.930 137.780 52.190 138.100 ;
        RECT 52.450 136.820 52.590 138.460 ;
        RECT 55.610 138.120 55.870 138.440 ;
        RECT 56.530 138.350 56.790 138.440 ;
        RECT 57.510 138.350 57.650 143.560 ;
        RECT 57.970 138.440 58.110 144.045 ;
        RECT 58.830 143.900 59.090 144.220 ;
        RECT 56.130 138.210 57.650 138.350 ;
        RECT 53.820 136.905 55.360 137.275 ;
        RECT 50.550 136.420 50.810 136.740 ;
        RECT 51.470 136.420 51.730 136.740 ;
        RECT 51.990 136.680 52.590 136.820 ;
        RECT 51.530 133.340 51.670 136.420 ;
        RECT 50.090 133.020 50.350 133.340 ;
        RECT 51.470 133.020 51.730 133.340 ;
        RECT 50.150 129.940 50.290 133.020 ;
        RECT 51.530 130.280 51.670 133.020 ;
        RECT 51.470 129.960 51.730 130.280 ;
        RECT 50.090 129.620 50.350 129.940 ;
        RECT 50.150 128.095 50.290 129.620 ;
        RECT 50.080 127.725 50.360 128.095 ;
        RECT 49.620 127.045 49.900 127.415 ;
        RECT 49.690 125.860 49.830 127.045 ;
        RECT 49.630 125.540 49.890 125.860 ;
        RECT 50.150 125.520 50.290 127.725 ;
        RECT 51.990 127.560 52.130 136.680 ;
        RECT 55.670 134.020 55.810 138.120 ;
        RECT 56.130 136.060 56.270 138.210 ;
        RECT 56.530 138.120 56.790 138.210 ;
        RECT 57.910 138.120 58.170 138.440 ;
        RECT 56.070 135.740 56.330 136.060 ;
        RECT 55.610 133.700 55.870 134.020 ;
        RECT 54.230 132.680 54.490 133.000 ;
        RECT 55.610 132.680 55.870 133.000 ;
        RECT 54.290 132.320 54.430 132.680 ;
        RECT 54.230 132.000 54.490 132.320 ;
        RECT 53.820 131.465 55.360 131.835 ;
        RECT 52.390 129.960 52.650 130.280 ;
        RECT 51.930 127.240 52.190 127.560 ;
        RECT 50.090 125.200 50.350 125.520 ;
        RECT 50.150 124.160 50.290 125.200 ;
        RECT 50.090 123.840 50.350 124.160 ;
        RECT 51.990 123.220 52.130 127.240 ;
        RECT 52.450 124.840 52.590 129.960 ;
        RECT 55.150 129.620 55.410 129.940 ;
        RECT 55.210 128.580 55.350 129.620 ;
        RECT 55.670 129.600 55.810 132.680 ;
        RECT 56.130 132.320 56.270 135.740 ;
        RECT 58.890 135.040 59.030 143.900 ;
        RECT 59.350 141.160 59.490 146.960 ;
        RECT 59.750 145.940 60.010 146.260 ;
        RECT 59.810 141.160 59.950 145.940 ;
        RECT 60.730 144.900 60.870 149.000 ;
        RECT 61.120 148.805 61.400 149.175 ;
        RECT 61.190 147.620 61.330 148.805 ;
        RECT 61.130 147.300 61.390 147.620 ;
        RECT 60.670 144.580 60.930 144.900 ;
        RECT 61.130 143.220 61.390 143.540 ;
        RECT 61.190 141.160 61.330 143.220 ;
        RECT 59.290 140.840 59.550 141.160 ;
        RECT 59.750 140.840 60.010 141.160 ;
        RECT 60.210 140.840 60.470 141.160 ;
        RECT 61.130 140.840 61.390 141.160 ;
        RECT 60.270 135.720 60.410 140.840 ;
        RECT 61.650 138.780 61.790 174.160 ;
        RECT 62.050 171.100 62.310 171.420 ;
        RECT 62.110 168.360 62.250 171.100 ;
        RECT 64.410 170.740 64.550 175.860 ;
        RECT 66.250 173.800 66.390 180.960 ;
        RECT 66.190 173.480 66.450 173.800 ;
        RECT 66.250 171.420 66.390 173.480 ;
        RECT 66.190 171.100 66.450 171.420 ;
        RECT 64.350 170.420 64.610 170.740 ;
        RECT 62.050 168.040 62.310 168.360 ;
        RECT 62.110 155.100 62.250 168.040 ;
        RECT 62.510 165.660 62.770 165.980 ;
        RECT 62.570 163.940 62.710 165.660 ;
        RECT 62.510 163.620 62.770 163.940 ;
        RECT 63.430 162.600 63.690 162.920 ;
        RECT 62.510 159.200 62.770 159.520 ;
        RECT 62.570 157.820 62.710 159.200 ;
        RECT 62.510 157.500 62.770 157.820 ;
        RECT 63.490 155.780 63.630 162.600 ;
        RECT 63.430 155.460 63.690 155.780 ;
        RECT 62.050 154.780 62.310 155.100 ;
        RECT 64.410 149.660 64.550 170.420 ;
        RECT 65.270 162.600 65.530 162.920 ;
        RECT 65.330 157.480 65.470 162.600 ;
        RECT 66.190 161.920 66.450 162.240 ;
        RECT 66.250 160.540 66.390 161.920 ;
        RECT 66.190 160.220 66.450 160.540 ;
        RECT 66.250 157.480 66.390 160.220 ;
        RECT 66.650 159.200 66.910 159.520 ;
        RECT 65.270 157.160 65.530 157.480 ;
        RECT 66.190 157.160 66.450 157.480 ;
        RECT 64.350 149.340 64.610 149.660 ;
        RECT 63.890 148.320 64.150 148.640 ;
        RECT 63.950 144.560 64.090 148.320 ;
        RECT 63.890 144.240 64.150 144.560 ;
        RECT 62.970 140.160 63.230 140.480 ;
        RECT 63.030 139.460 63.170 140.160 ;
        RECT 62.970 139.140 63.230 139.460 ;
        RECT 64.410 138.780 64.550 149.340 ;
        RECT 65.330 143.880 65.470 157.160 ;
        RECT 66.710 151.360 66.850 159.200 ;
        RECT 67.170 152.380 67.310 180.960 ;
        RECT 68.080 177.705 69.620 178.075 ;
        RECT 67.570 176.540 67.830 176.860 ;
        RECT 67.630 174.140 67.770 176.540 ;
        RECT 70.330 175.520 70.590 175.840 ;
        RECT 67.570 173.820 67.830 174.140 ;
        RECT 69.870 173.140 70.130 173.460 ;
        RECT 68.080 172.265 69.620 172.635 ;
        RECT 69.930 171.420 70.070 173.140 ;
        RECT 69.870 171.100 70.130 171.420 ;
        RECT 69.870 167.360 70.130 167.680 ;
        RECT 68.080 166.825 69.620 167.195 ;
        RECT 69.930 165.980 70.070 167.360 ;
        RECT 68.950 165.660 69.210 165.980 ;
        RECT 69.410 165.660 69.670 165.980 ;
        RECT 69.870 165.660 70.130 165.980 ;
        RECT 69.010 163.600 69.150 165.660 ;
        RECT 68.950 163.280 69.210 163.600 ;
        RECT 69.470 162.920 69.610 165.660 ;
        RECT 69.410 162.600 69.670 162.920 ;
        RECT 68.080 161.385 69.620 161.755 ;
        RECT 68.950 160.900 69.210 161.220 ;
        RECT 69.010 160.735 69.150 160.900 ;
        RECT 68.940 160.365 69.220 160.735 ;
        RECT 69.410 160.450 69.670 160.540 ;
        RECT 69.930 160.450 70.070 165.660 ;
        RECT 70.390 163.260 70.530 175.520 ;
        RECT 70.850 163.940 70.990 190.820 ;
        RECT 71.250 189.800 71.510 190.120 ;
        RECT 71.310 185.020 71.450 189.800 ;
        RECT 71.250 184.700 71.510 185.020 ;
        RECT 71.250 183.680 71.510 184.000 ;
        RECT 71.310 182.640 71.450 183.680 ;
        RECT 71.250 182.320 71.510 182.640 ;
        RECT 71.770 182.300 71.910 195.920 ;
        RECT 79.530 195.580 79.790 195.900 ;
        RECT 84.590 195.580 84.850 195.900 ;
        RECT 75.390 194.560 75.650 194.880 ;
        RECT 75.850 194.560 76.110 194.880 ;
        RECT 75.450 193.520 75.590 194.560 ;
        RECT 75.390 193.200 75.650 193.520 ;
        RECT 74.010 192.520 74.270 192.840 ;
        RECT 72.170 191.840 72.430 192.160 ;
        RECT 72.230 190.460 72.370 191.840 ;
        RECT 72.170 190.140 72.430 190.460 ;
        RECT 73.550 189.295 73.810 189.440 ;
        RECT 73.540 188.925 73.820 189.295 ;
        RECT 74.070 187.740 74.210 192.520 ;
        RECT 75.390 189.800 75.650 190.120 ;
        RECT 74.470 189.120 74.730 189.440 ;
        RECT 73.550 187.420 73.810 187.740 ;
        RECT 74.010 187.420 74.270 187.740 ;
        RECT 72.630 186.400 72.890 186.720 ;
        RECT 72.170 185.040 72.430 185.360 ;
        RECT 71.710 181.980 71.970 182.300 ;
        RECT 72.230 181.960 72.370 185.040 ;
        RECT 72.690 184.680 72.830 186.400 ;
        RECT 73.610 184.680 73.750 187.420 ;
        RECT 74.530 186.720 74.670 189.120 ;
        RECT 75.450 187.740 75.590 189.800 ;
        RECT 75.910 189.780 76.050 194.560 ;
        RECT 79.590 191.140 79.730 195.580 ;
        RECT 80.910 194.900 81.170 195.220 ;
        RECT 80.970 193.860 81.110 194.900 ;
        RECT 80.910 193.540 81.170 193.860 ;
        RECT 84.650 193.180 84.790 195.580 ;
        RECT 85.050 194.560 85.310 194.880 ;
        RECT 85.110 193.180 85.250 194.560 ;
        RECT 96.600 194.025 98.140 194.395 ;
        RECT 98.850 193.200 99.110 193.520 ;
        RECT 103.450 193.200 103.710 193.520 ;
        RECT 84.590 192.860 84.850 193.180 ;
        RECT 85.050 192.860 85.310 193.180 ;
        RECT 91.030 192.860 91.290 193.180 ;
        RECT 81.830 192.520 82.090 192.840 ;
        RECT 81.890 191.140 82.030 192.520 ;
        RECT 82.340 191.305 83.880 191.675 ;
        RECT 79.530 190.820 79.790 191.140 ;
        RECT 81.830 190.820 82.090 191.140 ;
        RECT 91.090 190.120 91.230 192.860 ;
        RECT 98.910 191.140 99.050 193.200 ;
        RECT 100.230 191.840 100.490 192.160 ;
        RECT 98.850 190.820 99.110 191.140 ;
        RECT 76.310 189.800 76.570 190.120 ;
        RECT 80.450 189.800 80.710 190.120 ;
        RECT 91.030 189.800 91.290 190.120 ;
        RECT 91.950 189.800 92.210 190.120 ;
        RECT 75.850 189.460 76.110 189.780 ;
        RECT 76.370 187.740 76.510 189.800 ;
        RECT 80.510 188.420 80.650 189.800 ;
        RECT 91.030 189.120 91.290 189.440 ;
        RECT 80.450 188.100 80.710 188.420 ;
        RECT 89.650 188.100 89.910 188.420 ;
        RECT 75.390 187.420 75.650 187.740 ;
        RECT 76.310 187.420 76.570 187.740 ;
        RECT 74.470 186.400 74.730 186.720 ;
        RECT 72.630 184.360 72.890 184.680 ;
        RECT 73.550 184.360 73.810 184.680 ;
        RECT 72.170 181.640 72.430 181.960 ;
        RECT 72.170 176.540 72.430 176.860 ;
        RECT 72.230 174.140 72.370 176.540 ;
        RECT 72.690 176.520 72.830 184.360 ;
        RECT 73.090 183.680 73.350 184.000 ;
        RECT 73.150 177.200 73.290 183.680 ;
        RECT 73.610 177.540 73.750 184.360 ;
        RECT 73.550 177.220 73.810 177.540 ;
        RECT 73.090 176.880 73.350 177.200 ;
        RECT 72.630 176.200 72.890 176.520 ;
        RECT 71.250 173.820 71.510 174.140 ;
        RECT 72.170 173.820 72.430 174.140 ;
        RECT 71.310 171.420 71.450 173.820 ;
        RECT 72.690 173.460 72.830 176.200 ;
        RECT 73.150 174.480 73.290 176.880 ;
        RECT 73.610 175.580 73.750 177.220 ;
        RECT 75.450 177.200 75.590 187.420 ;
        RECT 75.850 184.020 76.110 184.340 ;
        RECT 75.910 181.280 76.050 184.020 ;
        RECT 76.370 184.000 76.510 187.420 ;
        RECT 87.810 187.080 88.070 187.400 ;
        RECT 82.340 185.865 83.880 186.235 ;
        RECT 82.750 184.700 83.010 185.020 ;
        RECT 76.310 183.680 76.570 184.000 ;
        RECT 81.830 183.680 82.090 184.000 ;
        RECT 75.850 180.960 76.110 181.280 ;
        RECT 78.150 180.960 78.410 181.280 ;
        RECT 75.910 179.580 76.050 180.960 ;
        RECT 78.210 180.260 78.350 180.960 ;
        RECT 78.150 179.940 78.410 180.260 ;
        RECT 75.850 179.260 76.110 179.580 ;
        RECT 81.890 178.900 82.030 183.680 ;
        RECT 82.810 182.640 82.950 184.700 ;
        RECT 82.750 182.320 83.010 182.640 ;
        RECT 87.870 181.960 88.010 187.080 ;
        RECT 89.190 186.400 89.450 186.720 ;
        RECT 89.250 185.020 89.390 186.400 ;
        RECT 89.710 185.020 89.850 188.100 ;
        RECT 91.090 188.080 91.230 189.120 ;
        RECT 91.030 187.760 91.290 188.080 ;
        RECT 92.010 185.700 92.150 189.800 ;
        RECT 93.330 189.120 93.590 189.440 ;
        RECT 93.390 188.080 93.530 189.120 ;
        RECT 96.600 188.585 98.140 188.955 ;
        RECT 93.330 187.760 93.590 188.080 ;
        RECT 100.290 187.400 100.430 191.840 ;
        RECT 103.510 190.460 103.650 193.200 ;
        RECT 107.590 192.860 107.850 193.180 ;
        RECT 103.910 192.520 104.170 192.840 ;
        RECT 103.450 190.140 103.710 190.460 ;
        RECT 102.530 189.120 102.790 189.440 ;
        RECT 102.590 187.740 102.730 189.120 ;
        RECT 102.530 187.420 102.790 187.740 ;
        RECT 100.230 187.080 100.490 187.400 ;
        RECT 101.610 187.080 101.870 187.400 ;
        RECT 91.950 185.380 92.210 185.700 ;
        RECT 94.710 185.040 94.970 185.360 ;
        RECT 89.190 184.700 89.450 185.020 ;
        RECT 89.650 184.700 89.910 185.020 ;
        RECT 87.810 181.640 88.070 181.960 ;
        RECT 82.340 180.425 83.880 180.795 ;
        RECT 87.870 179.580 88.010 181.640 ;
        RECT 87.810 179.260 88.070 179.580 ;
        RECT 86.430 178.920 86.690 179.240 ;
        RECT 75.850 178.580 76.110 178.900 ;
        RECT 81.830 178.580 82.090 178.900 ;
        RECT 75.390 176.880 75.650 177.200 ;
        RECT 75.910 176.520 76.050 178.580 ;
        RECT 78.150 178.240 78.410 178.560 ;
        RECT 78.210 177.200 78.350 178.240 ;
        RECT 86.490 177.540 86.630 178.920 ;
        RECT 86.430 177.220 86.690 177.540 ;
        RECT 76.310 176.880 76.570 177.200 ;
        RECT 78.150 176.880 78.410 177.200 ;
        RECT 84.590 176.880 84.850 177.200 ;
        RECT 87.870 176.940 88.010 179.260 ;
        RECT 75.850 176.200 76.110 176.520 ;
        RECT 73.610 175.440 74.210 175.580 ;
        RECT 74.070 174.820 74.210 175.440 ;
        RECT 73.550 174.500 73.810 174.820 ;
        RECT 74.010 174.500 74.270 174.820 ;
        RECT 73.090 174.160 73.350 174.480 ;
        RECT 72.630 173.140 72.890 173.460 ;
        RECT 72.690 171.420 72.830 173.140 ;
        RECT 73.150 173.120 73.290 174.160 ;
        RECT 73.090 172.800 73.350 173.120 ;
        RECT 73.150 171.760 73.290 172.800 ;
        RECT 73.090 171.440 73.350 171.760 ;
        RECT 71.250 171.100 71.510 171.420 ;
        RECT 72.630 171.100 72.890 171.420 ;
        RECT 71.710 170.420 71.970 170.740 ;
        RECT 71.250 168.720 71.510 169.040 ;
        RECT 71.310 166.660 71.450 168.720 ;
        RECT 71.770 168.020 71.910 170.420 ;
        RECT 72.630 170.080 72.890 170.400 ;
        RECT 73.090 170.080 73.350 170.400 ;
        RECT 72.690 168.360 72.830 170.080 ;
        RECT 72.630 168.040 72.890 168.360 ;
        RECT 71.710 167.700 71.970 168.020 ;
        RECT 71.770 166.660 71.910 167.700 ;
        RECT 71.250 166.340 71.510 166.660 ;
        RECT 71.710 166.340 71.970 166.660 ;
        RECT 72.690 166.320 72.830 168.040 ;
        RECT 72.630 166.000 72.890 166.320 ;
        RECT 72.170 164.980 72.430 165.300 ;
        RECT 70.790 163.620 71.050 163.940 ;
        RECT 70.330 162.940 70.590 163.260 ;
        RECT 70.850 160.540 70.990 163.620 ;
        RECT 71.710 162.940 71.970 163.260 ;
        RECT 71.770 160.540 71.910 162.940 ;
        RECT 72.230 162.920 72.370 164.980 ;
        RECT 72.690 164.020 72.830 166.000 ;
        RECT 73.150 165.980 73.290 170.080 ;
        RECT 73.090 165.660 73.350 165.980 ;
        RECT 72.690 163.880 73.290 164.020 ;
        RECT 72.630 163.280 72.890 163.600 ;
        RECT 72.170 162.600 72.430 162.920 ;
        RECT 69.410 160.310 70.070 160.450 ;
        RECT 69.410 160.220 69.670 160.310 ;
        RECT 70.790 160.220 71.050 160.540 ;
        RECT 71.710 160.220 71.970 160.540 ;
        RECT 70.850 157.480 70.990 160.220 ;
        RECT 71.250 159.880 71.510 160.200 ;
        RECT 71.310 159.520 71.450 159.880 ;
        RECT 71.250 159.200 71.510 159.520 ;
        RECT 70.790 157.160 71.050 157.480 ;
        RECT 67.570 156.480 67.830 156.800 ;
        RECT 69.870 156.480 70.130 156.800 ;
        RECT 70.330 156.480 70.590 156.800 ;
        RECT 67.630 154.420 67.770 156.480 ;
        RECT 68.080 155.945 69.620 156.315 ;
        RECT 69.930 155.100 70.070 156.480 ;
        RECT 69.870 154.780 70.130 155.100 ;
        RECT 68.030 154.440 68.290 154.760 ;
        RECT 67.570 154.100 67.830 154.420 ;
        RECT 67.630 153.060 67.770 154.100 ;
        RECT 67.570 152.740 67.830 153.060 ;
        RECT 67.110 152.060 67.370 152.380 ;
        RECT 68.090 151.780 68.230 154.440 ;
        RECT 69.930 153.820 70.070 154.780 ;
        RECT 69.470 153.680 70.070 153.820 ;
        RECT 69.470 152.040 69.610 153.680 ;
        RECT 70.390 152.040 70.530 156.480 ;
        RECT 71.310 155.440 71.450 159.200 ;
        RECT 71.770 157.480 71.910 160.220 ;
        RECT 71.710 157.160 71.970 157.480 ;
        RECT 71.250 155.120 71.510 155.440 ;
        RECT 67.170 151.700 68.230 151.780 ;
        RECT 69.410 151.720 69.670 152.040 ;
        RECT 70.330 151.895 70.590 152.040 ;
        RECT 67.110 151.640 68.230 151.700 ;
        RECT 67.110 151.380 67.370 151.640 ;
        RECT 70.320 151.525 70.600 151.895 ;
        RECT 66.650 151.040 66.910 151.360 ;
        RECT 65.270 143.560 65.530 143.880 ;
        RECT 61.590 138.460 61.850 138.780 ;
        RECT 64.350 138.460 64.610 138.780 ;
        RECT 60.210 135.400 60.470 135.720 ;
        RECT 62.970 135.400 63.230 135.720 ;
        RECT 58.830 134.720 59.090 135.040 ;
        RECT 62.510 134.720 62.770 135.040 ;
        RECT 62.570 134.020 62.710 134.720 ;
        RECT 59.750 133.700 60.010 134.020 ;
        RECT 62.510 133.700 62.770 134.020 ;
        RECT 56.070 132.000 56.330 132.320 ;
        RECT 59.290 132.000 59.550 132.320 ;
        RECT 55.610 129.280 55.870 129.600 ;
        RECT 55.150 128.260 55.410 128.580 ;
        RECT 52.850 127.580 53.110 127.900 ;
        RECT 52.390 124.520 52.650 124.840 ;
        RECT 51.530 123.080 52.130 123.220 ;
        RECT 51.530 120.080 51.670 123.080 ;
        RECT 52.910 121.860 53.050 127.580 ;
        RECT 56.130 127.560 56.270 132.000 ;
        RECT 59.350 130.620 59.490 132.000 ;
        RECT 59.290 130.300 59.550 130.620 ;
        RECT 57.910 129.280 58.170 129.600 ;
        RECT 57.970 128.580 58.110 129.280 ;
        RECT 57.910 128.260 58.170 128.580 ;
        RECT 56.070 127.240 56.330 127.560 ;
        RECT 58.370 127.240 58.630 127.560 ;
        RECT 53.310 126.900 53.570 127.220 ;
        RECT 53.370 125.090 53.510 126.900 ;
        RECT 53.820 126.025 55.360 126.395 ;
        RECT 53.370 124.950 53.970 125.090 ;
        RECT 53.310 124.180 53.570 124.500 ;
        RECT 53.370 122.460 53.510 124.180 ;
        RECT 53.310 122.140 53.570 122.460 ;
        RECT 51.990 121.720 53.050 121.860 ;
        RECT 51.990 121.440 52.130 121.720 ;
        RECT 51.930 121.120 52.190 121.440 ;
        RECT 52.850 121.120 53.110 121.440 ;
        RECT 51.470 119.760 51.730 120.080 ;
        RECT 51.470 118.740 51.730 119.060 ;
        RECT 50.090 118.400 50.350 118.720 ;
        RECT 50.150 117.360 50.290 118.400 ;
        RECT 50.090 117.040 50.350 117.360 ;
        RECT 51.530 113.960 51.670 118.740 ;
        RECT 51.990 116.420 52.130 121.120 ;
        RECT 52.910 117.700 53.050 121.120 ;
        RECT 53.370 119.400 53.510 122.140 ;
        RECT 53.830 121.440 53.970 124.950 ;
        RECT 56.130 122.120 56.270 127.240 ;
        RECT 58.430 125.180 58.570 127.240 ;
        RECT 58.370 124.860 58.630 125.180 ;
        RECT 58.430 123.140 58.570 124.860 ;
        RECT 58.370 122.820 58.630 123.140 ;
        RECT 56.070 121.800 56.330 122.120 ;
        RECT 53.770 121.120 54.030 121.440 ;
        RECT 53.820 120.585 55.360 120.955 ;
        RECT 56.130 119.740 56.270 121.800 ;
        RECT 53.770 119.420 54.030 119.740 ;
        RECT 56.070 119.420 56.330 119.740 ;
        RECT 53.310 119.080 53.570 119.400 ;
        RECT 53.830 118.630 53.970 119.420 ;
        RECT 53.370 118.490 53.970 118.630 ;
        RECT 52.850 117.380 53.110 117.700 ;
        RECT 52.390 116.420 52.650 116.680 ;
        RECT 51.990 116.360 52.650 116.420 ;
        RECT 51.990 116.280 52.590 116.360 ;
        RECT 51.470 113.640 51.730 113.960 ;
        RECT 50.550 111.940 50.810 112.260 ;
        RECT 48.710 109.220 48.970 109.540 ;
        RECT 50.610 108.520 50.750 111.940 ;
        RECT 51.990 108.860 52.130 116.280 ;
        RECT 52.910 113.620 53.050 117.380 ;
        RECT 53.370 116.000 53.510 118.490 ;
        RECT 56.070 118.400 56.330 118.720 ;
        RECT 55.610 116.700 55.870 117.020 ;
        RECT 53.310 115.680 53.570 116.000 ;
        RECT 53.370 114.300 53.510 115.680 ;
        RECT 53.820 115.145 55.360 115.515 ;
        RECT 55.670 114.980 55.810 116.700 ;
        RECT 55.610 114.660 55.870 114.980 ;
        RECT 53.310 113.980 53.570 114.300 ;
        RECT 56.130 113.960 56.270 118.400 ;
        RECT 56.070 113.640 56.330 113.960 ;
        RECT 52.850 113.300 53.110 113.620 ;
        RECT 52.910 112.260 53.050 113.300 ;
        RECT 52.850 111.940 53.110 112.260 ;
        RECT 59.810 111.580 59.950 133.700 ;
        RECT 61.130 132.680 61.390 133.000 ;
        RECT 61.190 130.280 61.330 132.680 ;
        RECT 61.130 129.960 61.390 130.280 ;
        RECT 61.190 128.240 61.330 129.960 ;
        RECT 61.130 127.920 61.390 128.240 ;
        RECT 61.130 127.240 61.390 127.560 ;
        RECT 61.190 119.740 61.330 127.240 ;
        RECT 61.130 119.420 61.390 119.740 ;
        RECT 60.210 118.740 60.470 119.060 ;
        RECT 60.270 117.700 60.410 118.740 ;
        RECT 60.210 117.380 60.470 117.700 ;
        RECT 61.190 117.020 61.330 119.420 ;
        RECT 63.030 117.700 63.170 135.400 ;
        RECT 64.410 130.280 64.550 138.460 ;
        RECT 65.270 137.440 65.530 137.760 ;
        RECT 64.810 133.360 65.070 133.680 ;
        RECT 64.870 131.300 65.010 133.360 ;
        RECT 64.810 130.980 65.070 131.300 ;
        RECT 65.330 130.280 65.470 137.440 ;
        RECT 64.350 130.190 64.610 130.280 ;
        RECT 64.350 130.050 65.010 130.190 ;
        RECT 64.350 129.960 64.610 130.050 ;
        RECT 63.430 126.560 63.690 126.880 ;
        RECT 63.490 124.500 63.630 126.560 ;
        RECT 63.430 124.180 63.690 124.500 ;
        RECT 63.890 121.120 64.150 121.440 ;
        RECT 63.950 119.740 64.090 121.120 ;
        RECT 63.890 119.420 64.150 119.740 ;
        RECT 62.970 117.380 63.230 117.700 ;
        RECT 61.130 116.700 61.390 117.020 ;
        RECT 63.030 114.980 63.170 117.380 ;
        RECT 62.970 114.660 63.230 114.980 ;
        RECT 64.350 113.300 64.610 113.620 ;
        RECT 64.410 112.260 64.550 113.300 ;
        RECT 64.870 113.280 65.010 130.050 ;
        RECT 65.270 129.960 65.530 130.280 ;
        RECT 65.270 128.260 65.530 128.580 ;
        RECT 65.330 125.180 65.470 128.260 ;
        RECT 65.270 124.860 65.530 125.180 ;
        RECT 65.730 124.860 65.990 125.180 ;
        RECT 65.270 119.310 65.530 119.400 ;
        RECT 65.790 119.310 65.930 124.860 ;
        RECT 67.170 119.400 67.310 151.380 ;
        RECT 68.080 150.505 69.620 150.875 ;
        RECT 69.870 150.020 70.130 150.340 ;
        RECT 68.080 145.065 69.620 145.435 ;
        RECT 69.930 144.300 70.070 150.020 ;
        RECT 71.770 149.660 71.910 157.160 ;
        RECT 72.230 154.500 72.370 162.600 ;
        RECT 72.690 160.880 72.830 163.280 ;
        RECT 73.150 163.260 73.290 163.880 ;
        RECT 73.090 162.940 73.350 163.260 ;
        RECT 73.090 161.920 73.350 162.240 ;
        RECT 72.630 160.560 72.890 160.880 ;
        RECT 72.630 155.460 72.890 155.780 ;
        RECT 72.690 155.100 72.830 155.460 ;
        RECT 72.630 154.780 72.890 155.100 ;
        RECT 72.230 154.360 72.830 154.500 ;
        RECT 72.170 153.760 72.430 154.080 ;
        RECT 72.230 152.720 72.370 153.760 ;
        RECT 72.170 152.400 72.430 152.720 ;
        RECT 72.170 151.720 72.430 152.040 ;
        RECT 72.230 151.360 72.370 151.720 ;
        RECT 72.170 151.040 72.430 151.360 ;
        RECT 71.710 149.340 71.970 149.660 ;
        RECT 70.330 148.320 70.590 148.640 ;
        RECT 71.710 148.320 71.970 148.640 ;
        RECT 69.010 144.160 70.070 144.300 ;
        RECT 70.390 144.220 70.530 148.320 ;
        RECT 71.770 147.620 71.910 148.320 ;
        RECT 71.710 147.300 71.970 147.620 ;
        RECT 70.790 146.620 71.050 146.940 ;
        RECT 70.850 144.560 70.990 146.620 ;
        RECT 70.790 144.240 71.050 144.560 ;
        RECT 69.010 142.180 69.150 144.160 ;
        RECT 70.330 143.900 70.590 144.220 ;
        RECT 69.870 142.880 70.130 143.200 ;
        RECT 68.950 141.860 69.210 142.180 ;
        RECT 67.570 140.500 67.830 140.820 ;
        RECT 67.630 139.460 67.770 140.500 ;
        RECT 69.010 140.480 69.150 141.860 ;
        RECT 68.950 140.160 69.210 140.480 ;
        RECT 68.080 139.625 69.620 139.995 ;
        RECT 67.570 139.140 67.830 139.460 ;
        RECT 69.410 138.690 69.670 138.780 ;
        RECT 69.930 138.690 70.070 142.880 ;
        RECT 71.250 141.180 71.510 141.500 ;
        RECT 70.790 140.840 71.050 141.160 ;
        RECT 69.410 138.550 70.070 138.690 ;
        RECT 69.410 138.460 69.670 138.550 ;
        RECT 69.470 136.060 69.610 138.460 ;
        RECT 69.410 135.740 69.670 136.060 ;
        RECT 70.330 134.720 70.590 135.040 ;
        RECT 68.080 134.185 69.620 134.555 ;
        RECT 70.390 133.340 70.530 134.720 ;
        RECT 70.850 133.340 70.990 140.840 ;
        RECT 71.310 139.460 71.450 141.180 ;
        RECT 71.250 139.140 71.510 139.460 ;
        RECT 71.770 138.780 71.910 147.300 ;
        RECT 72.690 146.600 72.830 154.360 ;
        RECT 73.150 153.060 73.290 161.920 ;
        RECT 73.090 152.740 73.350 153.060 ;
        RECT 73.090 149.340 73.350 149.660 ;
        RECT 73.150 146.940 73.290 149.340 ;
        RECT 73.610 148.640 73.750 174.500 ;
        RECT 74.010 173.140 74.270 173.460 ;
        RECT 74.070 168.700 74.210 173.140 ;
        RECT 75.910 171.760 76.050 176.200 ;
        RECT 76.370 174.140 76.510 176.880 ;
        RECT 77.230 175.860 77.490 176.180 ;
        RECT 77.290 174.820 77.430 175.860 ;
        RECT 77.230 174.500 77.490 174.820 ;
        RECT 76.310 173.820 76.570 174.140 ;
        RECT 77.290 173.800 77.430 174.500 ;
        RECT 77.230 173.480 77.490 173.800 ;
        RECT 75.850 171.440 76.110 171.760 ;
        RECT 76.770 170.080 77.030 170.400 ;
        RECT 74.010 168.380 74.270 168.700 ;
        RECT 74.070 165.980 74.210 168.380 ;
        RECT 74.010 165.660 74.270 165.980 ;
        RECT 76.830 164.960 76.970 170.080 ;
        RECT 76.770 164.640 77.030 164.960 ;
        RECT 77.690 164.640 77.950 164.960 ;
        RECT 77.230 162.940 77.490 163.260 ;
        RECT 77.290 161.220 77.430 162.940 ;
        RECT 76.310 160.900 76.570 161.220 ;
        RECT 77.230 160.900 77.490 161.220 ;
        RECT 76.370 158.500 76.510 160.900 ;
        RECT 77.750 160.540 77.890 164.640 ;
        RECT 77.690 160.220 77.950 160.540 ;
        RECT 77.230 159.880 77.490 160.200 ;
        RECT 76.770 159.200 77.030 159.520 ;
        RECT 76.310 158.180 76.570 158.500 ;
        RECT 76.300 156.965 76.580 157.335 ;
        RECT 76.310 156.820 76.570 156.965 ;
        RECT 74.010 156.480 74.270 156.800 ;
        RECT 74.070 155.100 74.210 156.480 ;
        RECT 74.010 154.780 74.270 155.100 ;
        RECT 74.930 153.760 75.190 154.080 ;
        RECT 74.010 151.040 74.270 151.360 ;
        RECT 73.550 148.320 73.810 148.640 ;
        RECT 73.090 146.620 73.350 146.940 ;
        RECT 73.610 146.600 73.750 148.320 ;
        RECT 72.630 146.510 72.890 146.600 ;
        RECT 72.230 146.370 72.890 146.510 ;
        RECT 72.230 139.120 72.370 146.370 ;
        RECT 72.630 146.280 72.890 146.370 ;
        RECT 73.550 146.280 73.810 146.600 ;
        RECT 73.090 145.940 73.350 146.260 ;
        RECT 73.150 144.415 73.290 145.940 ;
        RECT 73.080 144.045 73.360 144.415 ;
        RECT 74.070 141.500 74.210 151.040 ;
        RECT 74.460 147.445 74.740 147.815 ;
        RECT 74.530 147.280 74.670 147.445 ;
        RECT 74.470 146.960 74.730 147.280 ;
        RECT 74.530 144.220 74.670 146.960 ;
        RECT 74.470 143.900 74.730 144.220 ;
        RECT 74.010 141.180 74.270 141.500 ;
        RECT 72.170 138.800 72.430 139.120 ;
        RECT 71.710 138.460 71.970 138.780 ;
        RECT 71.250 133.700 71.510 134.020 ;
        RECT 70.330 133.020 70.590 133.340 ;
        RECT 70.790 133.020 71.050 133.340 ;
        RECT 71.310 131.300 71.450 133.700 ;
        RECT 71.250 131.210 71.510 131.300 ;
        RECT 71.250 131.070 71.910 131.210 ;
        RECT 71.250 130.980 71.510 131.070 ;
        RECT 71.250 129.960 71.510 130.280 ;
        RECT 68.080 128.745 69.620 129.115 ;
        RECT 71.310 127.900 71.450 129.960 ;
        RECT 71.770 128.580 71.910 131.070 ;
        RECT 71.710 128.260 71.970 128.580 ;
        RECT 71.250 127.580 71.510 127.900 ;
        RECT 72.230 127.560 72.370 138.800 ;
        RECT 73.090 137.780 73.350 138.100 ;
        RECT 73.150 136.740 73.290 137.780 ;
        RECT 73.090 136.420 73.350 136.740 ;
        RECT 73.550 136.420 73.810 136.740 ;
        RECT 73.610 131.300 73.750 136.420 ;
        RECT 74.470 134.720 74.730 135.040 ;
        RECT 73.550 130.980 73.810 131.300 ;
        RECT 73.550 129.620 73.810 129.940 ;
        RECT 72.170 127.240 72.430 127.560 ;
        RECT 72.630 127.240 72.890 127.560 ;
        RECT 70.330 126.560 70.590 126.880 ;
        RECT 70.390 124.840 70.530 126.560 ;
        RECT 70.330 124.520 70.590 124.840 ;
        RECT 71.710 123.840 71.970 124.160 ;
        RECT 68.080 123.305 69.620 123.675 ;
        RECT 71.770 121.440 71.910 123.840 ;
        RECT 71.710 121.120 71.970 121.440 ;
        RECT 71.770 120.420 71.910 121.120 ;
        RECT 71.710 120.100 71.970 120.420 ;
        RECT 65.270 119.170 65.930 119.310 ;
        RECT 65.270 119.080 65.530 119.170 ;
        RECT 67.110 119.080 67.370 119.400 ;
        RECT 65.330 117.020 65.470 119.080 ;
        RECT 68.080 117.865 69.620 118.235 ;
        RECT 72.230 117.700 72.370 127.240 ;
        RECT 72.690 123.140 72.830 127.240 ;
        RECT 72.630 122.820 72.890 123.140 ;
        RECT 72.690 119.400 72.830 122.820 ;
        RECT 73.610 122.120 73.750 129.620 ;
        RECT 73.550 121.800 73.810 122.120 ;
        RECT 72.630 119.080 72.890 119.400 ;
        RECT 72.170 117.380 72.430 117.700 ;
        RECT 65.270 116.700 65.530 117.020 ;
        RECT 65.330 114.300 65.470 116.700 ;
        RECT 73.610 116.680 73.750 121.800 ;
        RECT 74.010 118.400 74.270 118.720 ;
        RECT 74.070 117.360 74.210 118.400 ;
        RECT 74.010 117.040 74.270 117.360 ;
        RECT 73.550 116.360 73.810 116.680 ;
        RECT 68.030 115.680 68.290 116.000 ;
        RECT 68.090 114.300 68.230 115.680 ;
        RECT 72.620 114.805 72.900 115.175 ;
        RECT 65.270 113.980 65.530 114.300 ;
        RECT 68.030 113.980 68.290 114.300 ;
        RECT 64.810 112.960 65.070 113.280 ;
        RECT 64.350 111.940 64.610 112.260 ;
        RECT 64.870 111.580 65.010 112.960 ;
        RECT 59.750 111.260 60.010 111.580 ;
        RECT 64.810 111.260 65.070 111.580 ;
        RECT 62.510 110.240 62.770 110.560 ;
        RECT 53.820 109.705 55.360 110.075 ;
        RECT 62.570 108.860 62.710 110.240 ;
        RECT 51.930 108.540 52.190 108.860 ;
        RECT 59.290 108.770 59.550 108.860 ;
        RECT 59.290 108.630 59.950 108.770 ;
        RECT 59.290 108.540 59.550 108.630 ;
        RECT 46.870 108.200 47.130 108.520 ;
        RECT 50.550 108.200 50.810 108.520 ;
        RECT 51.470 107.520 51.730 107.840 ;
        RECT 51.530 106.480 51.670 107.520 ;
        RECT 42.730 106.160 42.990 106.480 ;
        RECT 51.470 106.160 51.730 106.480 ;
        RECT 46.870 105.820 47.130 106.140 ;
        RECT 46.930 104.100 47.070 105.820 ;
        RECT 51.990 105.800 52.130 108.540 ;
        RECT 55.610 108.200 55.870 108.520 ;
        RECT 55.670 106.480 55.810 108.200 ;
        RECT 56.070 107.860 56.330 108.180 ;
        RECT 55.610 106.160 55.870 106.480 ;
        RECT 47.790 105.480 48.050 105.800 ;
        RECT 51.930 105.480 52.190 105.800 ;
        RECT 55.610 105.480 55.870 105.800 ;
        RECT 46.870 103.780 47.130 104.100 ;
        RECT 47.850 100.690 47.990 105.480 ;
        RECT 53.820 104.265 55.360 104.635 ;
        RECT 17.880 100.100 18.160 100.690 ;
        RECT 17.030 99.960 18.160 100.100 ;
        RECT 11.900 98.690 12.180 99.960 ;
        RECT 17.880 98.690 18.160 99.960 ;
        RECT 23.860 98.690 24.140 100.690 ;
        RECT 29.840 98.690 30.120 100.690 ;
        RECT 35.820 98.690 36.100 100.690 ;
        RECT 41.800 98.690 42.080 100.690 ;
        RECT 47.780 98.690 48.060 100.690 ;
        RECT 53.760 100.100 54.040 100.690 ;
        RECT 55.670 100.100 55.810 105.480 ;
        RECT 56.130 103.080 56.270 107.860 ;
        RECT 56.070 102.760 56.330 103.080 ;
        RECT 59.810 100.690 59.950 108.630 ;
        RECT 62.510 108.540 62.770 108.860 ;
        RECT 65.330 108.360 65.470 113.980 ;
        RECT 68.080 112.425 69.620 112.795 ;
        RECT 66.650 108.770 66.910 108.860 ;
        RECT 66.250 108.630 66.910 108.770 ;
        RECT 66.250 108.360 66.390 108.630 ;
        RECT 66.650 108.540 66.910 108.630 ;
        RECT 72.690 108.520 72.830 114.805 ;
        RECT 74.530 111.580 74.670 134.720 ;
        RECT 74.990 128.240 75.130 153.760 ;
        RECT 76.310 151.040 76.570 151.360 ;
        RECT 75.390 147.300 75.650 147.620 ;
        RECT 75.450 144.560 75.590 147.300 ;
        RECT 75.390 144.240 75.650 144.560 ;
        RECT 75.390 140.335 75.650 140.480 ;
        RECT 75.380 139.965 75.660 140.335 ;
        RECT 76.370 134.780 76.510 151.040 ;
        RECT 76.830 141.160 76.970 159.200 ;
        RECT 77.290 157.140 77.430 159.880 ;
        RECT 77.690 159.540 77.950 159.860 ;
        RECT 77.750 157.480 77.890 159.540 ;
        RECT 77.690 157.160 77.950 157.480 ;
        RECT 77.230 156.820 77.490 157.140 ;
        RECT 77.290 154.760 77.430 156.820 ;
        RECT 77.750 155.100 77.890 157.160 ;
        RECT 78.210 156.660 78.350 176.880 ;
        RECT 79.530 176.540 79.790 176.860 ;
        RECT 79.590 173.120 79.730 176.540 ;
        RECT 84.130 176.200 84.390 176.520 ;
        RECT 79.990 175.520 80.250 175.840 ;
        RECT 80.050 174.140 80.190 175.520 ;
        RECT 82.340 174.985 83.880 175.355 ;
        RECT 84.190 174.820 84.330 176.200 ;
        RECT 84.650 176.180 84.790 176.880 ;
        RECT 87.870 176.800 88.470 176.940 ;
        RECT 88.330 176.520 88.470 176.800 ;
        RECT 88.270 176.200 88.530 176.520 ;
        RECT 84.590 175.860 84.850 176.180 ;
        RECT 84.650 174.820 84.790 175.860 ;
        RECT 85.050 175.520 85.310 175.840 ;
        RECT 84.130 174.500 84.390 174.820 ;
        RECT 84.590 174.500 84.850 174.820 ;
        RECT 79.990 173.820 80.250 174.140 ;
        RECT 79.530 172.800 79.790 173.120 ;
        RECT 78.610 167.360 78.870 167.680 ;
        RECT 78.670 164.960 78.810 167.360 ;
        RECT 78.610 164.640 78.870 164.960 ;
        RECT 78.670 163.260 78.810 164.640 ;
        RECT 78.610 162.940 78.870 163.260 ;
        RECT 78.610 161.920 78.870 162.240 ;
        RECT 78.670 161.220 78.810 161.920 ;
        RECT 78.610 160.900 78.870 161.220 ;
        RECT 79.070 160.900 79.330 161.220 ;
        RECT 78.670 157.480 78.810 160.900 ;
        RECT 78.610 157.160 78.870 157.480 ;
        RECT 79.130 156.800 79.270 160.900 ;
        RECT 78.210 156.520 78.810 156.660 ;
        RECT 77.690 154.780 77.950 155.100 ;
        RECT 77.230 154.440 77.490 154.760 ;
        RECT 77.230 153.760 77.490 154.080 ;
        RECT 76.770 140.840 77.030 141.160 ;
        RECT 76.770 135.575 77.030 135.720 ;
        RECT 76.760 135.205 77.040 135.575 ;
        RECT 76.370 134.640 76.970 134.780 ;
        RECT 75.850 132.000 76.110 132.320 ;
        RECT 75.910 130.280 76.050 132.000 ;
        RECT 76.310 130.980 76.570 131.300 ;
        RECT 75.390 129.960 75.650 130.280 ;
        RECT 75.850 129.960 76.110 130.280 ;
        RECT 74.930 127.920 75.190 128.240 ;
        RECT 75.450 127.900 75.590 129.960 ;
        RECT 76.370 127.900 76.510 130.980 ;
        RECT 76.830 130.620 76.970 134.640 ;
        RECT 76.770 130.300 77.030 130.620 ;
        RECT 77.290 130.280 77.430 153.760 ;
        RECT 78.150 152.740 78.410 153.060 ;
        RECT 78.210 152.040 78.350 152.740 ;
        RECT 77.690 151.720 77.950 152.040 ;
        RECT 78.150 151.720 78.410 152.040 ;
        RECT 77.750 149.660 77.890 151.720 ;
        RECT 78.210 149.660 78.350 151.720 ;
        RECT 78.670 149.660 78.810 156.520 ;
        RECT 79.070 156.480 79.330 156.800 ;
        RECT 79.130 155.100 79.270 156.480 ;
        RECT 79.070 154.780 79.330 155.100 ;
        RECT 79.590 154.500 79.730 172.800 ;
        RECT 82.340 169.545 83.880 169.915 ;
        RECT 83.670 167.700 83.930 168.020 ;
        RECT 83.730 167.535 83.870 167.700 ;
        RECT 83.660 167.165 83.940 167.535 ;
        RECT 80.450 164.640 80.710 164.960 ;
        RECT 80.510 163.940 80.650 164.640 ;
        RECT 82.340 164.105 83.880 164.475 ;
        RECT 80.450 163.620 80.710 163.940 ;
        RECT 81.370 159.880 81.630 160.200 ;
        RECT 84.130 159.880 84.390 160.200 ;
        RECT 81.430 158.500 81.570 159.880 ;
        RECT 82.340 158.665 83.880 159.035 ;
        RECT 84.190 158.500 84.330 159.880 ;
        RECT 81.370 158.180 81.630 158.500 ;
        RECT 84.130 158.180 84.390 158.500 ;
        RECT 79.990 157.160 80.250 157.480 ;
        RECT 80.050 155.100 80.190 157.160 ;
        RECT 84.650 156.660 84.790 174.500 ;
        RECT 85.110 171.420 85.250 175.520 ;
        RECT 88.330 174.140 88.470 176.200 ;
        RECT 89.250 175.840 89.390 184.700 ;
        RECT 89.190 175.520 89.450 175.840 ;
        RECT 89.250 174.480 89.390 175.520 ;
        RECT 89.190 174.160 89.450 174.480 ;
        RECT 88.270 173.820 88.530 174.140 ;
        RECT 86.890 173.140 87.150 173.460 ;
        RECT 86.950 172.100 87.090 173.140 ;
        RECT 86.890 171.780 87.150 172.100 ;
        RECT 85.050 171.100 85.310 171.420 ;
        RECT 87.350 170.760 87.610 171.080 ;
        RECT 86.890 170.420 87.150 170.740 ;
        RECT 86.950 166.660 87.090 170.420 ;
        RECT 87.410 169.380 87.550 170.760 ;
        RECT 88.330 169.380 88.470 173.820 ;
        RECT 89.710 171.760 89.850 184.700 ;
        RECT 94.770 182.300 94.910 185.040 ;
        RECT 96.600 183.145 98.140 183.515 ;
        RECT 94.710 181.980 94.970 182.300 ;
        RECT 94.770 177.620 94.910 181.980 ;
        RECT 97.470 180.960 97.730 181.280 ;
        RECT 97.530 179.240 97.670 180.960 ;
        RECT 98.390 179.260 98.650 179.580 ;
        RECT 97.470 178.920 97.730 179.240 ;
        RECT 96.600 177.705 98.140 178.075 ;
        RECT 94.310 177.540 94.910 177.620 ;
        RECT 94.250 177.480 94.910 177.540 ;
        RECT 94.250 177.220 94.510 177.480 ;
        RECT 89.650 171.440 89.910 171.760 ;
        RECT 88.730 171.100 88.990 171.420 ;
        RECT 92.410 171.100 92.670 171.420 ;
        RECT 87.350 169.060 87.610 169.380 ;
        RECT 88.270 169.060 88.530 169.380 ;
        RECT 87.410 168.700 87.550 169.060 ;
        RECT 87.350 168.380 87.610 168.700 ;
        RECT 86.890 166.340 87.150 166.660 ;
        RECT 88.330 165.980 88.470 169.060 ;
        RECT 88.270 165.660 88.530 165.980 ;
        RECT 88.270 162.600 88.530 162.920 ;
        RECT 88.330 161.220 88.470 162.600 ;
        RECT 88.270 160.900 88.530 161.220 ;
        RECT 88.790 160.880 88.930 171.100 ;
        RECT 92.470 169.040 92.610 171.100 ;
        RECT 92.410 168.720 92.670 169.040 ;
        RECT 94.770 168.360 94.910 177.480 ;
        RECT 97.470 176.880 97.730 177.200 ;
        RECT 97.530 174.820 97.670 176.880 ;
        RECT 98.450 174.820 98.590 179.260 ;
        RECT 100.690 178.240 100.950 178.560 ;
        RECT 100.750 176.940 100.890 178.240 ;
        RECT 100.750 176.800 101.350 176.940 ;
        RECT 101.210 176.520 101.350 176.800 ;
        RECT 101.150 176.200 101.410 176.520 ;
        RECT 97.470 174.500 97.730 174.820 ;
        RECT 98.390 174.500 98.650 174.820 ;
        RECT 101.210 174.140 101.350 176.200 ;
        RECT 101.150 173.820 101.410 174.140 ;
        RECT 96.600 172.265 98.140 172.635 ;
        RECT 100.690 171.100 100.950 171.420 ;
        RECT 95.170 170.420 95.430 170.740 ;
        RECT 94.710 168.040 94.970 168.360 ;
        RECT 92.870 167.360 93.130 167.680 ;
        RECT 90.110 165.660 90.370 165.980 ;
        RECT 90.170 163.260 90.310 165.660 ;
        RECT 90.110 162.940 90.370 163.260 ;
        RECT 90.170 162.240 90.310 162.940 ;
        RECT 92.930 162.580 93.070 167.360 ;
        RECT 94.770 166.660 94.910 168.040 ;
        RECT 94.710 166.340 94.970 166.660 ;
        RECT 92.870 162.260 93.130 162.580 ;
        RECT 89.650 161.920 89.910 162.240 ;
        RECT 90.110 161.920 90.370 162.240 ;
        RECT 93.790 161.920 94.050 162.240 ;
        RECT 89.710 161.220 89.850 161.920 ;
        RECT 89.650 160.900 89.910 161.220 ;
        RECT 88.730 160.560 88.990 160.880 ;
        RECT 93.330 160.220 93.590 160.540 ;
        RECT 89.190 159.200 89.450 159.520 ;
        RECT 91.950 159.200 92.210 159.520 ;
        RECT 89.250 157.140 89.390 159.200 ;
        RECT 92.010 157.820 92.150 159.200 ;
        RECT 91.950 157.500 92.210 157.820 ;
        RECT 93.390 157.480 93.530 160.220 ;
        RECT 93.850 157.820 93.990 161.920 ;
        RECT 94.710 160.560 94.970 160.880 ;
        RECT 94.250 159.200 94.510 159.520 ;
        RECT 93.790 157.500 94.050 157.820 ;
        RECT 93.330 157.160 93.590 157.480 ;
        RECT 89.190 156.820 89.450 157.140 ;
        RECT 84.190 156.520 84.790 156.660 ;
        RECT 79.990 154.780 80.250 155.100 ;
        RECT 79.130 154.360 79.730 154.500 ;
        RECT 79.130 152.040 79.270 154.360 ;
        RECT 82.340 153.225 83.880 153.595 ;
        RECT 81.830 152.740 82.090 153.060 ;
        RECT 81.890 152.040 82.030 152.740 ;
        RECT 84.190 152.380 84.330 156.520 ;
        RECT 88.270 152.740 88.530 153.060 ;
        RECT 84.130 152.060 84.390 152.380 ;
        RECT 79.070 151.720 79.330 152.040 ;
        RECT 81.830 151.720 82.090 152.040 ;
        RECT 79.530 151.040 79.790 151.360 ;
        RECT 80.910 151.040 81.170 151.360 ;
        RECT 79.590 149.660 79.730 151.040 ;
        RECT 77.690 149.340 77.950 149.660 ;
        RECT 78.150 149.340 78.410 149.660 ;
        RECT 78.610 149.340 78.870 149.660 ;
        RECT 79.530 149.340 79.790 149.660 ;
        RECT 77.690 148.320 77.950 148.640 ;
        RECT 77.750 135.720 77.890 148.320 ;
        RECT 78.610 145.600 78.870 145.920 ;
        RECT 78.670 138.100 78.810 145.600 ;
        RECT 80.450 143.900 80.710 144.220 ;
        RECT 79.070 142.880 79.330 143.200 ;
        RECT 79.130 141.160 79.270 142.880 ;
        RECT 79.530 141.860 79.790 142.180 ;
        RECT 79.070 140.840 79.330 141.160 ;
        RECT 79.130 138.975 79.270 140.840 ;
        RECT 79.060 138.605 79.340 138.975 ;
        RECT 79.070 138.460 79.330 138.605 ;
        RECT 78.610 137.780 78.870 138.100 ;
        RECT 78.150 137.440 78.410 137.760 ;
        RECT 78.210 135.720 78.350 137.440 ;
        RECT 77.690 135.400 77.950 135.720 ;
        RECT 78.150 135.400 78.410 135.720 ;
        RECT 79.130 133.340 79.270 138.460 ;
        RECT 79.070 133.020 79.330 133.340 ;
        RECT 79.130 130.280 79.270 133.020 ;
        RECT 77.230 129.960 77.490 130.280 ;
        RECT 79.070 129.960 79.330 130.280 ;
        RECT 79.070 129.280 79.330 129.600 ;
        RECT 79.130 128.240 79.270 129.280 ;
        RECT 79.070 127.920 79.330 128.240 ;
        RECT 75.390 127.580 75.650 127.900 ;
        RECT 76.310 127.580 76.570 127.900 ;
        RECT 78.150 127.240 78.410 127.560 ;
        RECT 77.690 126.560 77.950 126.880 ;
        RECT 77.750 125.860 77.890 126.560 ;
        RECT 77.690 125.540 77.950 125.860 ;
        RECT 78.210 124.840 78.350 127.240 ;
        RECT 79.590 126.880 79.730 141.860 ;
        RECT 80.510 141.160 80.650 143.900 ;
        RECT 79.990 140.840 80.250 141.160 ;
        RECT 80.450 140.840 80.710 141.160 ;
        RECT 80.050 139.460 80.190 140.840 ;
        RECT 80.450 140.160 80.710 140.480 ;
        RECT 79.990 139.140 80.250 139.460 ;
        RECT 80.050 134.020 80.190 139.140 ;
        RECT 80.510 138.780 80.650 140.160 ;
        RECT 80.450 138.460 80.710 138.780 ;
        RECT 80.450 137.780 80.710 138.100 ;
        RECT 79.990 133.700 80.250 134.020 ;
        RECT 80.050 130.190 80.190 133.700 ;
        RECT 80.510 133.340 80.650 137.780 ;
        RECT 80.450 133.020 80.710 133.340 ;
        RECT 80.450 130.190 80.710 130.280 ;
        RECT 80.050 130.050 80.710 130.190 ;
        RECT 80.450 129.960 80.710 130.050 ;
        RECT 80.970 127.560 81.110 151.040 ;
        RECT 88.330 149.660 88.470 152.740 ;
        RECT 92.870 149.680 93.130 150.000 ;
        RECT 88.270 149.570 88.530 149.660 ;
        RECT 87.870 149.430 88.530 149.570 ;
        RECT 82.340 147.785 83.880 148.155 ;
        RECT 84.130 145.940 84.390 146.260 ;
        RECT 83.210 145.600 83.470 145.920 ;
        RECT 83.270 144.220 83.410 145.600 ;
        RECT 83.670 144.240 83.930 144.560 ;
        RECT 83.210 143.900 83.470 144.220 ;
        RECT 83.730 143.880 83.870 144.240 ;
        RECT 81.830 143.560 82.090 143.880 ;
        RECT 83.670 143.560 83.930 143.880 ;
        RECT 81.370 140.840 81.630 141.160 ;
        RECT 81.430 138.780 81.570 140.840 ;
        RECT 81.370 138.460 81.630 138.780 ;
        RECT 81.890 136.060 82.030 143.560 ;
        RECT 84.190 143.200 84.330 145.940 ;
        RECT 85.970 144.300 86.230 144.560 ;
        RECT 86.890 144.300 87.150 144.560 ;
        RECT 85.970 144.240 87.150 144.300 ;
        RECT 84.590 143.900 84.850 144.220 ;
        RECT 86.030 144.160 87.090 144.240 ;
        RECT 84.130 142.880 84.390 143.200 ;
        RECT 82.340 142.345 83.880 142.715 ;
        RECT 84.650 140.480 84.790 143.900 ;
        RECT 86.430 140.500 86.690 140.820 ;
        RECT 84.590 140.160 84.850 140.480 ;
        RECT 82.340 136.905 83.880 137.275 ;
        RECT 84.650 136.060 84.790 140.160 ;
        RECT 86.490 139.460 86.630 140.500 ;
        RECT 86.430 139.140 86.690 139.460 ;
        RECT 87.870 139.120 88.010 149.430 ;
        RECT 88.270 149.340 88.530 149.430 ;
        RECT 88.270 148.320 88.530 148.640 ;
        RECT 90.570 148.320 90.830 148.640 ;
        RECT 88.330 146.260 88.470 148.320 ;
        RECT 90.110 146.280 90.370 146.600 ;
        RECT 88.270 145.940 88.530 146.260 ;
        RECT 90.170 144.900 90.310 146.280 ;
        RECT 90.630 145.920 90.770 148.320 ;
        RECT 92.930 147.620 93.070 149.680 ;
        RECT 92.870 147.300 93.130 147.620 ;
        RECT 93.390 146.600 93.530 157.160 ;
        RECT 94.310 156.800 94.450 159.200 ;
        RECT 94.770 158.500 94.910 160.560 ;
        RECT 94.710 158.180 94.970 158.500 ;
        RECT 94.250 156.480 94.510 156.800 ;
        RECT 94.710 151.040 94.970 151.360 ;
        RECT 91.950 146.280 92.210 146.600 ;
        RECT 93.330 146.280 93.590 146.600 ;
        RECT 94.250 146.280 94.510 146.600 ;
        RECT 90.570 145.600 90.830 145.920 ;
        RECT 90.630 144.900 90.770 145.600 ;
        RECT 90.110 144.580 90.370 144.900 ;
        RECT 90.570 144.580 90.830 144.900 ;
        RECT 92.010 141.500 92.150 146.280 ;
        RECT 94.310 144.900 94.450 146.280 ;
        RECT 94.250 144.580 94.510 144.900 ;
        RECT 93.790 141.860 94.050 142.180 ;
        RECT 91.950 141.180 92.210 141.500 ;
        RECT 89.190 140.840 89.450 141.160 ;
        RECT 89.250 139.460 89.390 140.840 ;
        RECT 89.190 139.140 89.450 139.460 ;
        RECT 87.810 138.800 88.070 139.120 ;
        RECT 86.890 138.460 87.150 138.780 ;
        RECT 86.950 136.740 87.090 138.460 ;
        RECT 86.890 136.420 87.150 136.740 ;
        RECT 81.830 135.740 82.090 136.060 ;
        RECT 83.210 135.740 83.470 136.060 ;
        RECT 84.590 135.740 84.850 136.060 ;
        RECT 81.370 133.020 81.630 133.340 ;
        RECT 81.430 130.280 81.570 133.020 ;
        RECT 83.270 133.000 83.410 135.740 ;
        RECT 87.870 135.720 88.010 138.800 ;
        RECT 87.810 135.400 88.070 135.720 ;
        RECT 84.130 134.720 84.390 135.040 ;
        RECT 84.190 133.680 84.330 134.720 ;
        RECT 84.130 133.360 84.390 133.680 ;
        RECT 84.190 133.000 84.330 133.360 ;
        RECT 81.830 132.680 82.090 133.000 ;
        RECT 83.210 132.680 83.470 133.000 ;
        RECT 84.130 132.680 84.390 133.000 ;
        RECT 81.890 130.280 82.030 132.680 ;
        RECT 82.340 131.465 83.880 131.835 ;
        RECT 84.190 131.300 84.330 132.680 ;
        RECT 84.130 130.980 84.390 131.300 ;
        RECT 85.050 130.640 85.310 130.960 ;
        RECT 81.370 129.960 81.630 130.280 ;
        RECT 81.830 129.960 82.090 130.280 ;
        RECT 80.910 127.240 81.170 127.560 ;
        RECT 81.370 127.240 81.630 127.560 ;
        RECT 79.530 126.560 79.790 126.880 ;
        RECT 78.150 124.520 78.410 124.840 ;
        RECT 75.390 124.180 75.650 124.500 ;
        RECT 74.930 119.760 75.190 120.080 ;
        RECT 74.990 116.680 75.130 119.760 ;
        RECT 75.450 119.740 75.590 124.180 ;
        RECT 81.430 124.160 81.570 127.240 ;
        RECT 82.340 126.025 83.880 126.395 ;
        RECT 81.370 123.840 81.630 124.160 ;
        RECT 83.210 123.840 83.470 124.160 ;
        RECT 83.270 123.140 83.410 123.840 ;
        RECT 83.210 122.820 83.470 123.140 ;
        RECT 77.230 122.480 77.490 122.800 ;
        RECT 76.770 121.800 77.030 122.120 ;
        RECT 75.390 119.420 75.650 119.740 ;
        RECT 76.830 119.060 76.970 121.800 ;
        RECT 77.290 120.420 77.430 122.480 ;
        RECT 79.070 122.140 79.330 122.460 ;
        RECT 77.230 120.100 77.490 120.420 ;
        RECT 76.770 118.740 77.030 119.060 ;
        RECT 77.690 118.740 77.950 119.060 ;
        RECT 77.750 117.700 77.890 118.740 ;
        RECT 78.150 118.400 78.410 118.720 ;
        RECT 77.690 117.380 77.950 117.700 ;
        RECT 74.930 116.360 75.190 116.680 ;
        RECT 78.210 113.960 78.350 118.400 ;
        RECT 79.130 117.700 79.270 122.140 ;
        RECT 83.270 121.860 83.410 122.820 ;
        RECT 84.590 122.480 84.850 122.800 ;
        RECT 83.270 121.720 84.330 121.860 ;
        RECT 82.340 120.585 83.880 120.955 ;
        RECT 84.190 120.420 84.330 121.720 ;
        RECT 84.130 120.100 84.390 120.420 ;
        RECT 84.650 120.080 84.790 122.480 ;
        RECT 80.450 119.760 80.710 120.080 ;
        RECT 84.590 119.760 84.850 120.080 ;
        RECT 80.510 119.400 80.650 119.760 ;
        RECT 80.450 119.080 80.710 119.400 ;
        RECT 81.370 119.080 81.630 119.400 ;
        RECT 79.070 117.380 79.330 117.700 ;
        RECT 79.070 116.360 79.330 116.680 ;
        RECT 79.130 114.980 79.270 116.360 ;
        RECT 79.070 114.660 79.330 114.980 ;
        RECT 81.430 114.640 81.570 119.080 ;
        RECT 84.650 117.360 84.790 119.760 ;
        RECT 84.590 117.040 84.850 117.360 ;
        RECT 82.340 115.145 83.880 115.515 ;
        RECT 81.370 114.320 81.630 114.640 ;
        RECT 78.150 113.640 78.410 113.960 ;
        RECT 74.470 111.260 74.730 111.580 ;
        RECT 77.230 110.920 77.490 111.240 ;
        RECT 75.390 110.240 75.650 110.560 ;
        RECT 75.450 108.860 75.590 110.240 ;
        RECT 75.390 108.540 75.650 108.860 ;
        RECT 65.330 108.220 66.390 108.360 ;
        RECT 60.210 107.860 60.470 108.180 ;
        RECT 60.270 104.100 60.410 107.860 ;
        RECT 66.250 106.820 66.390 108.220 ;
        RECT 72.630 108.200 72.890 108.520 ;
        RECT 73.090 107.860 73.350 108.180 ;
        RECT 70.330 107.520 70.590 107.840 ;
        RECT 68.080 106.985 69.620 107.355 ;
        RECT 66.190 106.500 66.450 106.820 ;
        RECT 70.390 106.480 70.530 107.520 ;
        RECT 62.510 106.160 62.770 106.480 ;
        RECT 70.330 106.160 70.590 106.480 ;
        RECT 62.570 104.100 62.710 106.160 ;
        RECT 65.270 105.540 65.530 105.800 ;
        RECT 65.270 105.480 65.930 105.540 ;
        RECT 65.330 105.400 65.930 105.480 ;
        RECT 60.210 103.780 60.470 104.100 ;
        RECT 62.510 103.780 62.770 104.100 ;
        RECT 65.790 100.690 65.930 105.400 ;
        RECT 71.710 105.140 71.970 105.460 ;
        RECT 68.080 101.545 69.620 101.915 ;
        RECT 71.770 100.690 71.910 105.140 ;
        RECT 73.150 104.100 73.290 107.860 ;
        RECT 77.290 106.820 77.430 110.920 ;
        RECT 82.340 109.705 83.880 110.075 ;
        RECT 77.690 108.880 77.950 109.200 ;
        RECT 77.230 106.500 77.490 106.820 ;
        RECT 75.390 105.820 75.650 106.140 ;
        RECT 75.450 104.100 75.590 105.820 ;
        RECT 73.090 103.780 73.350 104.100 ;
        RECT 75.390 103.780 75.650 104.100 ;
        RECT 77.290 103.080 77.430 106.500 ;
        RECT 77.230 102.760 77.490 103.080 ;
        RECT 77.750 100.690 77.890 108.880 ;
        RECT 85.110 108.520 85.250 130.640 ;
        RECT 86.890 129.620 87.150 129.940 ;
        RECT 86.950 128.580 87.090 129.620 ;
        RECT 86.890 128.260 87.150 128.580 ;
        RECT 87.870 127.900 88.010 135.400 ;
        RECT 88.270 132.000 88.530 132.320 ;
        RECT 88.330 130.620 88.470 132.000 ;
        RECT 88.270 130.300 88.530 130.620 ;
        RECT 92.010 130.280 92.150 141.180 ;
        RECT 92.870 135.400 93.130 135.720 ;
        RECT 92.930 130.280 93.070 135.400 ;
        RECT 93.330 133.360 93.590 133.680 ;
        RECT 93.390 131.300 93.530 133.360 ;
        RECT 93.330 130.980 93.590 131.300 ;
        RECT 91.950 129.960 92.210 130.280 ;
        RECT 92.870 129.960 93.130 130.280 ;
        RECT 92.010 127.900 92.150 129.960 ;
        RECT 93.850 128.580 93.990 141.860 ;
        RECT 94.770 141.160 94.910 151.040 ;
        RECT 95.230 146.940 95.370 170.420 ;
        RECT 99.770 170.080 100.030 170.400 ;
        RECT 96.090 168.380 96.350 168.700 ;
        RECT 95.620 167.165 95.900 167.535 ;
        RECT 95.690 166.320 95.830 167.165 ;
        RECT 95.630 166.000 95.890 166.320 ;
        RECT 96.150 165.640 96.290 168.380 ;
        RECT 98.390 167.360 98.650 167.680 ;
        RECT 96.600 166.825 98.140 167.195 ;
        RECT 98.450 166.660 98.590 167.360 ;
        RECT 98.390 166.340 98.650 166.660 ;
        RECT 96.090 165.320 96.350 165.640 ;
        RECT 96.150 157.820 96.290 165.320 ;
        RECT 98.450 163.340 98.590 166.340 ;
        RECT 99.830 163.940 99.970 170.080 ;
        RECT 100.750 169.380 100.890 171.100 ;
        RECT 100.690 169.060 100.950 169.380 ;
        RECT 99.770 163.620 100.030 163.940 ;
        RECT 97.990 163.260 98.590 163.340 ;
        RECT 101.210 163.260 101.350 173.820 ;
        RECT 101.670 168.360 101.810 187.080 ;
        RECT 102.070 186.400 102.330 186.720 ;
        RECT 102.130 184.680 102.270 186.400 ;
        RECT 103.510 184.680 103.650 190.140 ;
        RECT 103.970 185.700 104.110 192.520 ;
        RECT 106.210 191.840 106.470 192.160 ;
        RECT 106.270 189.780 106.410 191.840 ;
        RECT 106.210 189.460 106.470 189.780 ;
        RECT 107.650 188.420 107.790 192.860 ;
        RECT 109.890 192.520 110.150 192.840 ;
        RECT 109.430 191.840 109.690 192.160 ;
        RECT 109.490 190.460 109.630 191.840 ;
        RECT 109.950 191.140 110.090 192.520 ;
        RECT 110.860 191.305 112.400 191.675 ;
        RECT 109.890 190.820 110.150 191.140 ;
        RECT 109.430 190.140 109.690 190.460 ;
        RECT 114.030 190.140 114.290 190.460 ;
        RECT 107.590 188.100 107.850 188.420 ;
        RECT 109.890 187.420 110.150 187.740 ;
        RECT 106.210 187.080 106.470 187.400 ;
        RECT 104.370 186.400 104.630 186.720 ;
        RECT 103.910 185.380 104.170 185.700 ;
        RECT 102.070 184.360 102.330 184.680 ;
        RECT 103.450 184.360 103.710 184.680 ;
        RECT 103.510 182.300 103.650 184.360 ;
        RECT 103.450 181.980 103.710 182.300 ;
        RECT 104.430 181.960 104.570 186.400 ;
        RECT 105.290 183.680 105.550 184.000 ;
        RECT 105.350 182.300 105.490 183.680 ;
        RECT 106.270 182.640 106.410 187.080 ;
        RECT 109.950 182.980 110.090 187.420 ;
        RECT 112.650 186.400 112.910 186.720 ;
        RECT 110.860 185.865 112.400 186.235 ;
        RECT 112.710 185.020 112.850 186.400 ;
        RECT 114.090 185.020 114.230 190.140 ;
        RECT 112.650 184.700 112.910 185.020 ;
        RECT 114.030 184.700 114.290 185.020 ;
        RECT 109.890 182.660 110.150 182.980 ;
        RECT 106.210 182.320 106.470 182.640 ;
        RECT 105.290 181.980 105.550 182.300 ;
        RECT 104.370 181.640 104.630 181.960 ;
        RECT 102.530 180.960 102.790 181.280 ;
        RECT 102.590 178.900 102.730 180.960 ;
        RECT 102.530 178.580 102.790 178.900 ;
        RECT 102.990 175.520 103.250 175.840 ;
        RECT 103.050 173.800 103.190 175.520 ;
        RECT 102.990 173.480 103.250 173.800 ;
        RECT 106.270 171.420 106.410 182.320 ;
        RECT 107.590 181.980 107.850 182.300 ;
        RECT 106.670 181.640 106.930 181.960 ;
        RECT 106.730 178.560 106.870 181.640 ;
        RECT 107.130 180.960 107.390 181.280 ;
        RECT 106.670 178.240 106.930 178.560 ;
        RECT 106.730 176.520 106.870 178.240 ;
        RECT 107.190 176.860 107.330 180.960 ;
        RECT 107.130 176.540 107.390 176.860 ;
        RECT 106.670 176.200 106.930 176.520 ;
        RECT 105.750 171.100 106.010 171.420 ;
        RECT 106.210 171.100 106.470 171.420 ;
        RECT 103.450 170.760 103.710 171.080 ;
        RECT 102.990 170.420 103.250 170.740 ;
        RECT 102.070 168.720 102.330 169.040 ;
        RECT 101.610 168.040 101.870 168.360 ;
        RECT 97.930 163.200 98.590 163.260 ;
        RECT 97.930 162.940 98.190 163.200 ;
        RECT 99.770 162.940 100.030 163.260 ;
        RECT 101.150 162.940 101.410 163.260 ;
        RECT 96.600 161.385 98.140 161.755 ;
        RECT 99.310 159.200 99.570 159.520 ;
        RECT 96.090 157.500 96.350 157.820 ;
        RECT 96.090 156.820 96.350 157.140 ;
        RECT 95.170 146.620 95.430 146.940 ;
        RECT 94.710 140.840 94.970 141.160 ;
        RECT 95.170 140.160 95.430 140.480 ;
        RECT 94.250 134.720 94.510 135.040 ;
        RECT 94.310 133.000 94.450 134.720 ;
        RECT 94.250 132.680 94.510 133.000 ;
        RECT 94.710 129.960 94.970 130.280 ;
        RECT 93.790 128.260 94.050 128.580 ;
        RECT 92.870 127.920 93.130 128.240 ;
        RECT 87.810 127.580 88.070 127.900 ;
        RECT 91.950 127.580 92.210 127.900 ;
        RECT 87.810 126.900 88.070 127.220 ;
        RECT 87.350 124.180 87.610 124.500 ;
        RECT 87.410 123.140 87.550 124.180 ;
        RECT 87.350 122.820 87.610 123.140 ;
        RECT 85.970 122.140 86.230 122.460 ;
        RECT 85.510 121.120 85.770 121.440 ;
        RECT 85.570 117.020 85.710 121.120 ;
        RECT 86.030 119.060 86.170 122.140 ;
        RECT 85.970 118.740 86.230 119.060 ;
        RECT 85.510 116.700 85.770 117.020 ;
        RECT 87.350 108.880 87.610 109.200 ;
        RECT 85.050 108.200 85.310 108.520 ;
        RECT 79.530 107.520 79.790 107.840 ;
        RECT 85.050 107.520 85.310 107.840 ;
        RECT 79.590 106.480 79.730 107.520 ;
        RECT 79.530 106.160 79.790 106.480 ;
        RECT 84.590 104.800 84.850 105.120 ;
        RECT 82.340 104.265 83.880 104.635 ;
        RECT 84.650 102.740 84.790 104.800 ;
        RECT 85.110 103.420 85.250 107.520 ;
        RECT 87.410 106.140 87.550 108.880 ;
        RECT 87.870 108.520 88.010 126.900 ;
        RECT 92.010 125.860 92.150 127.580 ;
        RECT 91.950 125.540 92.210 125.860 ;
        RECT 89.650 122.480 89.910 122.800 ;
        RECT 88.730 119.420 88.990 119.740 ;
        RECT 88.790 117.700 88.930 119.420 ;
        RECT 89.710 117.700 89.850 122.480 ;
        RECT 92.010 122.120 92.150 125.540 ;
        RECT 92.930 125.375 93.070 127.920 ;
        RECT 92.860 125.005 93.140 125.375 ;
        RECT 92.930 124.840 93.070 125.005 ;
        RECT 92.870 124.520 93.130 124.840 ;
        RECT 93.790 124.180 94.050 124.500 ;
        RECT 91.950 121.800 92.210 122.120 ;
        RECT 92.010 119.740 92.150 121.800 ;
        RECT 91.950 119.420 92.210 119.740 ;
        RECT 88.730 117.380 88.990 117.700 ;
        RECT 89.650 117.380 89.910 117.700 ;
        RECT 92.010 116.680 92.150 119.420 ;
        RECT 93.850 119.400 93.990 124.180 ;
        RECT 94.770 123.140 94.910 129.960 ;
        RECT 94.710 122.820 94.970 123.140 ;
        RECT 94.710 122.140 94.970 122.460 ;
        RECT 94.770 120.420 94.910 122.140 ;
        RECT 94.710 120.100 94.970 120.420 ;
        RECT 94.250 119.420 94.510 119.740 ;
        RECT 93.790 119.080 94.050 119.400 ;
        RECT 94.310 118.720 94.450 119.420 ;
        RECT 94.250 118.400 94.510 118.720 ;
        RECT 94.310 117.700 94.450 118.400 ;
        RECT 94.250 117.380 94.510 117.700 ;
        RECT 91.950 116.360 92.210 116.680 ;
        RECT 92.010 109.540 92.150 116.360 ;
        RECT 95.230 111.580 95.370 140.160 ;
        RECT 96.150 138.780 96.290 156.820 ;
        RECT 98.390 156.480 98.650 156.800 ;
        RECT 96.600 155.945 98.140 156.315 ;
        RECT 97.930 155.460 98.190 155.780 ;
        RECT 97.470 154.100 97.730 154.420 ;
        RECT 97.530 152.040 97.670 154.100 ;
        RECT 97.990 152.040 98.130 155.460 ;
        RECT 98.450 152.040 98.590 156.480 ;
        RECT 98.850 154.780 99.110 155.100 ;
        RECT 98.910 152.040 99.050 154.780 ;
        RECT 97.470 151.720 97.730 152.040 ;
        RECT 97.930 151.720 98.190 152.040 ;
        RECT 98.390 151.720 98.650 152.040 ;
        RECT 98.850 151.720 99.110 152.040 ;
        RECT 96.600 150.505 98.140 150.875 ;
        RECT 98.910 150.340 99.050 151.720 ;
        RECT 98.850 150.020 99.110 150.340 ;
        RECT 96.550 149.000 96.810 149.320 ;
        RECT 98.390 149.000 98.650 149.320 ;
        RECT 96.610 147.620 96.750 149.000 ;
        RECT 96.550 147.300 96.810 147.620 ;
        RECT 96.600 145.065 98.140 145.435 ;
        RECT 97.470 143.220 97.730 143.540 ;
        RECT 97.530 141.160 97.670 143.220 ;
        RECT 97.930 142.880 98.190 143.200 ;
        RECT 97.990 142.180 98.130 142.880 ;
        RECT 97.930 141.860 98.190 142.180 ;
        RECT 97.990 141.160 98.130 141.860 ;
        RECT 97.470 140.840 97.730 141.160 ;
        RECT 97.930 140.840 98.190 141.160 ;
        RECT 96.600 139.625 98.140 139.995 ;
        RECT 96.090 138.460 96.350 138.780 ;
        RECT 96.090 134.720 96.350 135.040 ;
        RECT 95.630 133.020 95.890 133.340 ;
        RECT 95.690 131.300 95.830 133.020 ;
        RECT 95.630 130.980 95.890 131.300 ;
        RECT 96.150 130.280 96.290 134.720 ;
        RECT 96.600 134.185 98.140 134.555 ;
        RECT 98.450 133.340 98.590 149.000 ;
        RECT 98.850 147.300 99.110 147.620 ;
        RECT 98.390 133.020 98.650 133.340 ;
        RECT 98.910 131.300 99.050 147.300 ;
        RECT 99.370 138.440 99.510 159.200 ;
        RECT 99.830 154.080 99.970 162.940 ;
        RECT 102.130 162.920 102.270 168.720 ;
        RECT 102.530 164.640 102.790 164.960 ;
        RECT 102.070 162.600 102.330 162.920 ;
        RECT 100.230 161.920 100.490 162.240 ;
        RECT 99.770 153.760 100.030 154.080 ;
        RECT 99.770 140.500 100.030 140.820 ;
        RECT 99.310 138.120 99.570 138.440 ;
        RECT 99.830 137.670 99.970 140.500 ;
        RECT 100.290 140.480 100.430 161.920 ;
        RECT 102.590 160.200 102.730 164.640 ;
        RECT 100.690 159.880 100.950 160.200 ;
        RECT 102.530 159.880 102.790 160.200 ;
        RECT 100.750 158.500 100.890 159.880 ;
        RECT 100.690 158.180 100.950 158.500 ;
        RECT 102.590 157.140 102.730 159.880 ;
        RECT 102.530 156.820 102.790 157.140 ;
        RECT 103.050 156.660 103.190 170.420 ;
        RECT 103.510 168.360 103.650 170.760 ;
        RECT 105.810 169.040 105.950 171.100 ;
        RECT 105.750 168.720 106.010 169.040 ;
        RECT 103.450 168.040 103.710 168.360 ;
        RECT 103.510 162.830 103.650 168.040 ;
        RECT 105.810 162.920 105.950 168.720 ;
        RECT 106.210 167.360 106.470 167.680 ;
        RECT 103.910 162.830 104.170 162.920 ;
        RECT 103.510 162.690 104.170 162.830 ;
        RECT 103.910 162.600 104.170 162.690 ;
        RECT 105.750 162.600 106.010 162.920 ;
        RECT 103.450 161.920 103.710 162.240 ;
        RECT 102.590 156.520 103.190 156.660 ;
        RECT 100.690 151.040 100.950 151.360 ;
        RECT 102.070 151.040 102.330 151.360 ;
        RECT 100.750 146.600 100.890 151.040 ;
        RECT 100.690 146.280 100.950 146.600 ;
        RECT 102.130 144.220 102.270 151.040 ;
        RECT 102.070 143.900 102.330 144.220 ;
        RECT 102.590 143.880 102.730 156.520 ;
        RECT 102.990 154.100 103.250 154.420 ;
        RECT 102.530 143.560 102.790 143.880 ;
        RECT 100.690 142.880 100.950 143.200 ;
        RECT 100.230 140.160 100.490 140.480 ;
        RECT 99.370 137.530 99.970 137.670 ;
        RECT 99.370 135.380 99.510 137.530 ;
        RECT 100.230 137.440 100.490 137.760 ;
        RECT 99.310 135.060 99.570 135.380 ;
        RECT 99.370 134.020 99.510 135.060 ;
        RECT 99.310 133.700 99.570 134.020 ;
        RECT 98.850 130.980 99.110 131.300 ;
        RECT 96.090 129.960 96.350 130.280 ;
        RECT 96.600 128.745 98.140 129.115 ;
        RECT 96.090 127.240 96.350 127.560 ;
        RECT 96.150 119.740 96.290 127.240 ;
        RECT 96.600 123.305 98.140 123.675 ;
        RECT 96.090 119.420 96.350 119.740 ;
        RECT 98.390 118.400 98.650 118.720 ;
        RECT 96.600 117.865 98.140 118.235 ;
        RECT 98.450 117.020 98.590 118.400 ;
        RECT 98.390 116.700 98.650 117.020 ;
        RECT 96.600 112.425 98.140 112.795 ;
        RECT 100.290 111.920 100.430 137.440 ;
        RECT 100.230 111.600 100.490 111.920 ;
        RECT 95.170 111.260 95.430 111.580 ;
        RECT 97.930 110.240 98.190 110.560 ;
        RECT 91.950 109.220 92.210 109.540 ;
        RECT 97.990 108.860 98.130 110.240 ;
        RECT 95.630 108.540 95.890 108.860 ;
        RECT 97.930 108.540 98.190 108.860 ;
        RECT 87.810 108.200 88.070 108.520 ;
        RECT 95.170 107.860 95.430 108.180 ;
        RECT 88.730 107.520 88.990 107.840 ;
        RECT 88.790 106.480 88.930 107.520 ;
        RECT 88.730 106.160 88.990 106.480 ;
        RECT 86.890 105.820 87.150 106.140 ;
        RECT 87.350 105.820 87.610 106.140 ;
        RECT 85.050 103.100 85.310 103.420 ;
        RECT 86.950 103.080 87.090 105.820 ;
        RECT 87.410 103.420 87.550 105.820 ;
        RECT 91.490 105.480 91.750 105.800 ;
        RECT 87.350 103.100 87.610 103.420 ;
        RECT 86.890 102.760 87.150 103.080 ;
        RECT 84.590 102.420 84.850 102.740 ;
        RECT 83.670 102.080 83.930 102.400 ;
        RECT 83.730 100.690 83.870 102.080 ;
        RECT 53.760 99.960 55.810 100.100 ;
        RECT 53.760 98.690 54.040 99.960 ;
        RECT 59.740 98.690 60.020 100.690 ;
        RECT 65.720 98.690 66.000 100.690 ;
        RECT 71.700 98.690 71.980 100.690 ;
        RECT 77.680 98.690 77.960 100.690 ;
        RECT 83.660 98.690 83.940 100.690 ;
        RECT 89.640 100.100 89.920 100.690 ;
        RECT 91.550 100.100 91.690 105.480 ;
        RECT 95.230 104.100 95.370 107.860 ;
        RECT 95.170 103.780 95.430 104.100 ;
        RECT 95.690 100.690 95.830 108.540 ;
        RECT 100.750 107.840 100.890 142.880 ;
        RECT 103.050 138.780 103.190 154.100 ;
        RECT 103.510 138.780 103.650 161.920 ;
        RECT 103.970 160.540 104.110 162.600 ;
        RECT 105.810 160.880 105.950 162.600 ;
        RECT 105.750 160.560 106.010 160.880 ;
        RECT 103.910 160.220 104.170 160.540 ;
        RECT 104.370 154.780 104.630 155.100 ;
        RECT 103.910 153.760 104.170 154.080 ;
        RECT 103.970 152.040 104.110 153.760 ;
        RECT 103.910 151.720 104.170 152.040 ;
        RECT 104.430 151.700 104.570 154.780 ;
        RECT 105.750 153.760 106.010 154.080 ;
        RECT 104.830 151.720 105.090 152.040 ;
        RECT 104.370 151.380 104.630 151.700 ;
        RECT 104.890 150.340 105.030 151.720 ;
        RECT 104.830 150.020 105.090 150.340 ;
        RECT 105.810 149.660 105.950 153.760 ;
        RECT 106.270 149.660 106.410 167.360 ;
        RECT 106.730 162.920 106.870 176.200 ;
        RECT 107.130 171.100 107.390 171.420 ;
        RECT 107.190 168.700 107.330 171.100 ;
        RECT 107.130 168.380 107.390 168.700 ;
        RECT 107.190 162.920 107.330 168.380 ;
        RECT 106.670 162.600 106.930 162.920 ;
        RECT 107.130 162.600 107.390 162.920 ;
        RECT 107.190 161.220 107.330 162.600 ;
        RECT 107.130 160.900 107.390 161.220 ;
        RECT 107.650 160.540 107.790 181.980 ;
        RECT 110.860 180.425 112.400 180.795 ;
        RECT 114.090 179.580 114.230 184.700 ;
        RECT 114.030 179.260 114.290 179.580 ;
        RECT 109.430 178.580 109.690 178.900 ;
        RECT 109.490 177.540 109.630 178.580 ;
        RECT 109.430 177.220 109.690 177.540 ;
        RECT 110.350 176.540 110.610 176.860 ;
        RECT 110.410 173.800 110.550 176.540 ;
        RECT 114.090 176.520 114.230 179.260 ;
        RECT 120.010 176.880 120.270 177.200 ;
        RECT 114.950 176.540 115.210 176.860 ;
        RECT 114.030 176.200 114.290 176.520 ;
        RECT 112.650 175.520 112.910 175.840 ;
        RECT 114.490 175.520 114.750 175.840 ;
        RECT 110.860 174.985 112.400 175.355 ;
        RECT 112.190 173.820 112.450 174.140 ;
        RECT 108.050 173.480 108.310 173.800 ;
        RECT 110.350 173.480 110.610 173.800 ;
        RECT 108.110 168.360 108.250 173.480 ;
        RECT 112.250 171.760 112.390 173.820 ;
        RECT 112.710 173.460 112.850 175.520 ;
        RECT 112.650 173.140 112.910 173.460 ;
        RECT 114.550 172.100 114.690 175.520 ;
        RECT 115.010 174.480 115.150 176.540 ;
        RECT 114.950 174.160 115.210 174.480 ;
        RECT 119.550 173.140 119.810 173.460 ;
        RECT 116.790 172.800 117.050 173.120 ;
        RECT 114.490 171.780 114.750 172.100 ;
        RECT 108.510 171.440 108.770 171.760 ;
        RECT 112.190 171.440 112.450 171.760 ;
        RECT 108.050 168.040 108.310 168.360 ;
        RECT 108.110 166.320 108.250 168.040 ;
        RECT 108.050 166.000 108.310 166.320 ;
        RECT 108.050 160.900 108.310 161.220 ;
        RECT 107.590 160.220 107.850 160.540 ;
        RECT 108.110 157.480 108.250 160.900 ;
        RECT 106.670 157.160 106.930 157.480 ;
        RECT 107.590 157.160 107.850 157.480 ;
        RECT 108.050 157.160 108.310 157.480 ;
        RECT 106.730 155.100 106.870 157.160 ;
        RECT 107.650 155.780 107.790 157.160 ;
        RECT 107.590 155.460 107.850 155.780 ;
        RECT 106.670 154.780 106.930 155.100 ;
        RECT 107.130 154.780 107.390 155.100 ;
        RECT 108.050 154.780 108.310 155.100 ;
        RECT 107.190 152.380 107.330 154.780 ;
        RECT 107.130 152.060 107.390 152.380 ;
        RECT 108.110 151.360 108.250 154.780 ;
        RECT 108.570 152.040 108.710 171.440 ;
        RECT 108.970 171.100 109.230 171.420 ;
        RECT 109.030 167.680 109.170 171.100 ;
        RECT 110.350 170.420 110.610 170.740 ;
        RECT 108.970 167.360 109.230 167.680 ;
        RECT 109.030 165.640 109.170 167.360 ;
        RECT 108.970 165.320 109.230 165.640 ;
        RECT 109.030 154.760 109.170 165.320 ;
        RECT 110.410 165.300 110.550 170.420 ;
        RECT 110.860 169.545 112.400 169.915 ;
        RECT 110.350 164.980 110.610 165.300 ;
        RECT 110.410 160.200 110.550 164.980 ;
        RECT 110.860 164.105 112.400 164.475 ;
        RECT 112.650 161.920 112.910 162.240 ;
        RECT 112.710 160.540 112.850 161.920 ;
        RECT 114.550 161.220 114.690 171.780 ;
        RECT 115.870 164.640 116.130 164.960 ;
        RECT 115.930 162.580 116.070 164.640 ;
        RECT 115.870 162.260 116.130 162.580 ;
        RECT 114.490 160.900 114.750 161.220 ;
        RECT 112.650 160.220 112.910 160.540 ;
        RECT 115.410 160.220 115.670 160.540 ;
        RECT 110.350 159.880 110.610 160.200 ;
        RECT 110.410 157.820 110.550 159.880 ;
        RECT 110.860 158.665 112.400 159.035 ;
        RECT 112.710 157.900 112.850 160.220 ;
        RECT 110.350 157.500 110.610 157.820 ;
        RECT 112.250 157.760 112.850 157.900 ;
        RECT 115.470 157.820 115.610 160.220 ;
        RECT 109.430 157.160 109.690 157.480 ;
        RECT 109.490 155.100 109.630 157.160 ;
        RECT 112.250 157.140 112.390 157.760 ;
        RECT 115.410 157.500 115.670 157.820 ;
        RECT 112.190 156.820 112.450 157.140 ;
        RECT 112.250 155.440 112.390 156.820 ;
        RECT 115.470 155.440 115.610 157.500 ;
        RECT 112.190 155.120 112.450 155.440 ;
        RECT 115.410 155.120 115.670 155.440 ;
        RECT 109.430 154.780 109.690 155.100 ;
        RECT 108.970 154.440 109.230 154.760 ;
        RECT 110.860 153.225 112.400 153.595 ;
        RECT 108.510 151.720 108.770 152.040 ;
        RECT 108.050 151.040 108.310 151.360 ;
        RECT 112.650 151.040 112.910 151.360 ;
        RECT 108.110 150.340 108.250 151.040 ;
        RECT 108.050 150.020 108.310 150.340 ;
        RECT 105.750 149.340 106.010 149.660 ;
        RECT 106.210 149.340 106.470 149.660 ;
        RECT 107.130 149.340 107.390 149.660 ;
        RECT 107.190 147.620 107.330 149.340 ;
        RECT 107.590 148.320 107.850 148.640 ;
        RECT 107.130 147.300 107.390 147.620 ;
        RECT 103.910 146.280 104.170 146.600 ;
        RECT 104.370 146.340 104.630 146.600 ;
        RECT 104.370 146.280 105.490 146.340 ;
        RECT 105.750 146.280 106.010 146.600 ;
        RECT 103.970 143.540 104.110 146.280 ;
        RECT 104.430 146.260 105.490 146.280 ;
        RECT 104.430 146.200 105.550 146.260 ;
        RECT 104.430 143.540 104.570 146.200 ;
        RECT 105.290 145.940 105.550 146.200 ;
        RECT 103.910 143.220 104.170 143.540 ;
        RECT 104.370 143.220 104.630 143.540 ;
        RECT 103.970 141.160 104.110 143.220 ;
        RECT 104.430 142.180 104.570 143.220 ;
        RECT 105.290 142.880 105.550 143.200 ;
        RECT 104.370 141.860 104.630 142.180 ;
        RECT 104.430 141.500 104.570 141.860 ;
        RECT 104.370 141.180 104.630 141.500 ;
        RECT 103.910 140.840 104.170 141.160 ;
        RECT 104.830 140.840 105.090 141.160 ;
        RECT 103.910 140.160 104.170 140.480 ;
        RECT 103.970 139.120 104.110 140.160 ;
        RECT 103.910 138.800 104.170 139.120 ;
        RECT 104.890 138.780 105.030 140.840 ;
        RECT 102.990 138.460 103.250 138.780 ;
        RECT 103.450 138.460 103.710 138.780 ;
        RECT 104.830 138.460 105.090 138.780 ;
        RECT 101.610 137.440 101.870 137.760 ;
        RECT 103.910 137.440 104.170 137.760 ;
        RECT 104.370 137.440 104.630 137.760 ;
        RECT 101.150 134.720 101.410 135.040 ;
        RECT 101.210 133.680 101.350 134.720 ;
        RECT 101.150 133.360 101.410 133.680 ;
        RECT 101.670 131.300 101.810 137.440 ;
        RECT 101.610 130.980 101.870 131.300 ;
        RECT 101.610 129.960 101.870 130.280 ;
        RECT 102.070 129.960 102.330 130.280 ;
        RECT 101.670 127.900 101.810 129.960 ;
        RECT 101.610 127.580 101.870 127.900 ;
        RECT 101.150 124.860 101.410 125.180 ;
        RECT 101.210 120.420 101.350 124.860 ;
        RECT 102.130 124.160 102.270 129.960 ;
        RECT 102.070 123.840 102.330 124.160 ;
        RECT 102.130 123.140 102.270 123.840 ;
        RECT 102.070 122.820 102.330 123.140 ;
        RECT 101.150 120.100 101.410 120.420 ;
        RECT 102.530 118.740 102.790 119.060 ;
        RECT 102.590 117.700 102.730 118.740 ;
        RECT 102.530 117.380 102.790 117.700 ;
        RECT 103.970 111.580 104.110 137.440 ;
        RECT 104.430 128.580 104.570 137.440 ;
        RECT 105.350 134.020 105.490 142.880 ;
        RECT 105.810 141.840 105.950 146.280 ;
        RECT 106.670 142.880 106.930 143.200 ;
        RECT 106.730 142.180 106.870 142.880 ;
        RECT 106.670 141.860 106.930 142.180 ;
        RECT 105.750 141.520 106.010 141.840 ;
        RECT 106.670 141.180 106.930 141.500 ;
        RECT 106.730 138.780 106.870 141.180 ;
        RECT 106.670 138.460 106.930 138.780 ;
        RECT 106.210 134.720 106.470 135.040 ;
        RECT 105.290 133.700 105.550 134.020 ;
        RECT 106.270 133.340 106.410 134.720 ;
        RECT 106.210 133.020 106.470 133.340 ;
        RECT 107.130 133.020 107.390 133.340 ;
        RECT 106.670 130.190 106.930 130.280 ;
        RECT 107.190 130.190 107.330 133.020 ;
        RECT 107.650 131.300 107.790 148.320 ;
        RECT 110.860 147.785 112.400 148.155 ;
        RECT 108.570 146.880 109.630 147.020 ;
        RECT 108.570 141.160 108.710 146.880 ;
        RECT 109.490 146.600 109.630 146.880 ;
        RECT 110.350 146.620 110.610 146.940 ;
        RECT 108.970 146.280 109.230 146.600 ;
        RECT 109.430 146.510 109.690 146.600 ;
        RECT 109.430 146.370 110.090 146.510 ;
        RECT 109.430 146.280 109.690 146.370 ;
        RECT 109.030 144.900 109.170 146.280 ;
        RECT 108.970 144.580 109.230 144.900 ;
        RECT 109.950 144.220 110.090 146.370 ;
        RECT 109.430 143.900 109.690 144.220 ;
        RECT 109.890 143.900 110.150 144.220 ;
        RECT 108.970 141.180 109.230 141.500 ;
        RECT 108.510 140.840 108.770 141.160 ;
        RECT 108.050 140.500 108.310 140.820 ;
        RECT 108.110 136.060 108.250 140.500 ;
        RECT 108.570 138.780 108.710 140.840 ;
        RECT 108.510 138.460 108.770 138.780 ;
        RECT 109.030 138.440 109.170 141.180 ;
        RECT 109.490 139.460 109.630 143.900 ;
        RECT 110.410 141.500 110.550 146.620 ;
        RECT 112.710 146.260 112.850 151.040 ;
        RECT 115.470 149.660 115.610 155.120 ;
        RECT 116.850 155.100 116.990 172.800 ;
        RECT 119.610 172.100 119.750 173.140 ;
        RECT 120.070 172.100 120.210 176.880 ;
        RECT 121.390 176.200 121.650 176.520 ;
        RECT 121.450 173.800 121.590 176.200 ;
        RECT 122.760 174.645 123.040 175.015 ;
        RECT 122.830 173.800 122.970 174.645 ;
        RECT 121.390 173.480 121.650 173.800 ;
        RECT 122.770 173.480 123.030 173.800 ;
        RECT 119.550 171.780 119.810 172.100 ;
        RECT 120.010 171.780 120.270 172.100 ;
        RECT 118.170 168.040 118.430 168.360 ;
        RECT 118.230 166.660 118.370 168.040 ;
        RECT 121.450 168.020 121.590 173.480 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 121.390 167.700 121.650 168.020 ;
        RECT 118.170 166.340 118.430 166.660 ;
        RECT 118.630 165.660 118.890 165.980 ;
        RECT 118.690 161.220 118.830 165.660 ;
        RECT 120.930 164.640 121.190 164.960 ;
        RECT 120.990 163.260 121.130 164.640 ;
        RECT 121.450 163.340 121.590 167.700 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 120.930 162.940 121.190 163.260 ;
        RECT 121.450 163.200 122.510 163.340 ;
        RECT 122.370 162.920 122.510 163.200 ;
        RECT 122.310 162.600 122.570 162.920 ;
        RECT 123.690 162.600 123.950 162.920 ;
        RECT 118.630 160.900 118.890 161.220 ;
        RECT 119.550 160.220 119.810 160.540 ;
        RECT 118.170 159.200 118.430 159.520 ;
        RECT 118.230 157.140 118.370 159.200 ;
        RECT 119.610 158.500 119.750 160.220 ;
        RECT 120.470 159.200 120.730 159.520 ;
        RECT 119.550 158.180 119.810 158.500 ;
        RECT 120.530 157.820 120.670 159.200 ;
        RECT 120.470 157.500 120.730 157.820 ;
        RECT 123.750 157.480 123.890 162.600 ;
        RECT 123.690 157.160 123.950 157.480 ;
        RECT 118.170 156.820 118.430 157.140 ;
        RECT 123.750 156.800 123.890 157.160 ;
        RECT 123.690 156.480 123.950 156.800 ;
        RECT 116.790 154.780 117.050 155.100 ;
        RECT 116.850 152.380 116.990 154.780 ;
        RECT 123.750 152.380 123.890 156.480 ;
        RECT 116.790 152.060 117.050 152.380 ;
        RECT 123.690 152.060 123.950 152.380 ;
        RECT 116.790 151.380 117.050 151.700 ;
        RECT 120.470 151.380 120.730 151.700 ;
        RECT 116.850 150.340 116.990 151.380 ;
        RECT 120.530 150.340 120.670 151.380 ;
        RECT 116.790 150.020 117.050 150.340 ;
        RECT 120.470 150.020 120.730 150.340 ;
        RECT 115.410 149.340 115.670 149.660 ;
        RECT 117.710 149.340 117.970 149.660 ;
        RECT 115.470 146.600 115.610 149.340 ;
        RECT 117.770 147.620 117.910 149.340 ;
        RECT 118.630 148.660 118.890 148.980 ;
        RECT 117.710 147.300 117.970 147.620 ;
        RECT 117.250 146.960 117.510 147.280 ;
        RECT 115.410 146.280 115.670 146.600 ;
        RECT 112.650 145.940 112.910 146.260 ;
        RECT 114.950 143.560 115.210 143.880 ;
        RECT 110.860 142.345 112.400 142.715 ;
        RECT 115.010 141.500 115.150 143.560 ;
        RECT 110.350 141.180 110.610 141.500 ;
        RECT 114.950 141.180 115.210 141.500 ;
        RECT 112.190 140.500 112.450 140.820 ;
        RECT 111.270 140.160 111.530 140.480 ;
        RECT 109.430 139.140 109.690 139.460 ;
        RECT 111.330 139.120 111.470 140.160 ;
        RECT 112.250 139.460 112.390 140.500 ;
        RECT 113.110 140.160 113.370 140.480 ;
        RECT 112.190 139.140 112.450 139.460 ;
        RECT 111.270 138.800 111.530 139.120 ;
        RECT 108.970 138.120 109.230 138.440 ;
        RECT 109.030 136.400 109.170 138.120 ;
        RECT 110.860 136.905 112.400 137.275 ;
        RECT 108.970 136.080 109.230 136.400 ;
        RECT 108.050 135.740 108.310 136.060 ;
        RECT 108.050 134.720 108.310 135.040 ;
        RECT 108.110 133.000 108.250 134.720 ;
        RECT 113.170 133.340 113.310 140.160 ;
        RECT 114.030 137.440 114.290 137.760 ;
        RECT 114.090 135.380 114.230 137.440 ;
        RECT 114.030 135.060 114.290 135.380 ;
        RECT 113.110 133.020 113.370 133.340 ;
        RECT 108.050 132.680 108.310 133.000 ;
        RECT 110.350 132.680 110.610 133.000 ;
        RECT 107.590 130.980 107.850 131.300 ;
        RECT 106.670 130.050 107.330 130.190 ;
        RECT 106.670 129.960 106.930 130.050 ;
        RECT 104.370 128.260 104.630 128.580 ;
        RECT 106.730 127.900 106.870 129.960 ;
        RECT 108.110 129.940 108.250 132.680 ;
        RECT 110.410 131.210 110.550 132.680 ;
        RECT 110.860 131.465 112.400 131.835 ;
        RECT 110.410 131.070 111.010 131.210 ;
        RECT 108.510 129.960 108.770 130.280 ;
        RECT 110.350 130.190 110.610 130.280 ;
        RECT 109.950 130.050 110.610 130.190 ;
        RECT 108.050 129.620 108.310 129.940 ;
        RECT 108.110 128.240 108.250 129.620 ;
        RECT 108.050 127.920 108.310 128.240 ;
        RECT 106.670 127.580 106.930 127.900 ;
        RECT 107.590 127.240 107.850 127.560 ;
        RECT 106.210 126.900 106.470 127.220 ;
        RECT 106.270 125.180 106.410 126.900 ;
        RECT 106.210 124.860 106.470 125.180 ;
        RECT 106.270 122.460 106.410 124.860 ;
        RECT 106.670 123.840 106.930 124.160 ;
        RECT 106.730 122.460 106.870 123.840 ;
        RECT 106.210 122.140 106.470 122.460 ;
        RECT 106.670 122.140 106.930 122.460 ;
        RECT 104.370 121.800 104.630 122.120 ;
        RECT 104.430 120.080 104.570 121.800 ;
        RECT 104.370 119.760 104.630 120.080 ;
        RECT 104.430 119.400 104.570 119.760 ;
        RECT 106.270 119.740 106.410 122.140 ;
        RECT 106.210 119.420 106.470 119.740 ;
        RECT 107.650 119.400 107.790 127.240 ;
        RECT 108.110 122.460 108.250 127.920 ;
        RECT 108.050 122.140 108.310 122.460 ;
        RECT 104.370 119.080 104.630 119.400 ;
        RECT 107.590 119.080 107.850 119.400 ;
        RECT 104.830 118.400 105.090 118.720 ;
        RECT 104.890 117.360 105.030 118.400 ;
        RECT 104.830 117.040 105.090 117.360 ;
        RECT 108.110 117.020 108.250 122.140 ;
        RECT 108.570 119.740 108.710 129.960 ;
        RECT 109.950 127.560 110.090 130.050 ;
        RECT 110.350 129.960 110.610 130.050 ;
        RECT 110.870 127.900 111.010 131.070 ;
        RECT 110.810 127.580 111.070 127.900 ;
        RECT 114.490 127.580 114.750 127.900 ;
        RECT 109.890 127.240 110.150 127.560 ;
        RECT 109.950 124.840 110.090 127.240 ;
        RECT 110.860 126.025 112.400 126.395 ;
        RECT 109.890 124.520 110.150 124.840 ;
        RECT 114.550 123.140 114.690 127.580 ;
        RECT 114.490 122.820 114.750 123.140 ;
        RECT 113.570 122.140 113.830 122.460 ;
        RECT 116.330 122.140 116.590 122.460 ;
        RECT 110.860 120.585 112.400 120.955 ;
        RECT 113.630 119.740 113.770 122.140 ;
        RECT 116.390 120.080 116.530 122.140 ;
        RECT 116.330 119.760 116.590 120.080 ;
        RECT 108.510 119.420 108.770 119.740 ;
        RECT 113.570 119.420 113.830 119.740 ;
        RECT 111.730 118.400 111.990 118.720 ;
        RECT 111.790 117.020 111.930 118.400 ;
        RECT 116.390 117.020 116.530 119.760 ;
        RECT 116.790 118.740 117.050 119.060 ;
        RECT 116.850 117.700 116.990 118.740 ;
        RECT 116.790 117.380 117.050 117.700 ;
        RECT 108.050 116.700 108.310 117.020 ;
        RECT 111.730 116.700 111.990 117.020 ;
        RECT 116.330 116.700 116.590 117.020 ;
        RECT 110.350 116.360 110.610 116.680 ;
        RECT 101.150 111.260 101.410 111.580 ;
        RECT 103.910 111.260 104.170 111.580 ;
        RECT 100.690 107.520 100.950 107.840 ;
        RECT 96.600 106.985 98.140 107.355 ;
        RECT 101.210 103.080 101.350 111.260 ;
        RECT 110.410 110.900 110.550 116.360 ;
        RECT 110.860 115.145 112.400 115.515 ;
        RECT 117.310 113.960 117.450 146.960 ;
        RECT 117.710 146.280 117.970 146.600 ;
        RECT 117.770 141.160 117.910 146.280 ;
        RECT 118.170 145.600 118.430 145.920 ;
        RECT 118.230 144.560 118.370 145.600 ;
        RECT 118.170 144.240 118.430 144.560 ;
        RECT 117.710 140.840 117.970 141.160 ;
        RECT 117.770 138.780 117.910 140.840 ;
        RECT 118.170 140.160 118.430 140.480 ;
        RECT 118.230 139.120 118.370 140.160 ;
        RECT 118.170 138.800 118.430 139.120 ;
        RECT 117.710 138.460 117.970 138.780 ;
        RECT 118.690 124.580 118.830 148.660 ;
        RECT 119.550 146.280 119.810 146.600 ;
        RECT 119.610 142.180 119.750 146.280 ;
        RECT 121.850 145.600 122.110 145.920 ;
        RECT 121.910 144.220 122.050 145.600 ;
        RECT 121.850 143.900 122.110 144.220 ;
        RECT 122.310 143.560 122.570 143.880 ;
        RECT 119.550 141.860 119.810 142.180 ;
        RECT 121.850 140.160 122.110 140.480 ;
        RECT 121.910 138.780 122.050 140.160 ;
        RECT 121.850 138.460 122.110 138.780 ;
        RECT 122.370 138.440 122.510 143.560 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 122.310 138.120 122.570 138.440 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 122.370 135.960 122.510 138.120 ;
        RECT 121.910 135.820 122.510 135.960 ;
        RECT 119.090 135.400 119.350 135.720 ;
        RECT 119.150 134.020 119.290 135.400 ;
        RECT 121.910 135.040 122.050 135.820 ;
        RECT 121.850 134.720 122.110 135.040 ;
        RECT 119.090 133.700 119.350 134.020 ;
        RECT 119.550 127.920 119.810 128.240 ;
        RECT 117.710 124.180 117.970 124.500 ;
        RECT 118.690 124.440 119.290 124.580 ;
        RECT 117.770 123.140 117.910 124.180 ;
        RECT 117.710 122.820 117.970 123.140 ;
        RECT 118.170 121.120 118.430 121.440 ;
        RECT 118.230 117.020 118.370 121.120 ;
        RECT 118.170 116.700 118.430 117.020 ;
        RECT 119.150 113.960 119.290 124.440 ;
        RECT 119.610 123.140 119.750 127.920 ;
        RECT 121.910 127.560 122.050 134.720 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 122.770 127.580 123.030 127.900 ;
        RECT 121.850 127.240 122.110 127.560 ;
        RECT 121.910 125.180 122.050 127.240 ;
        RECT 122.830 125.860 122.970 127.580 ;
        RECT 124.150 126.560 124.410 126.880 ;
        RECT 122.770 125.540 123.030 125.860 ;
        RECT 121.850 124.860 122.110 125.180 ;
        RECT 119.550 122.820 119.810 123.140 ;
        RECT 121.910 119.400 122.050 124.860 ;
        RECT 124.210 124.840 124.350 126.560 ;
        RECT 124.150 124.520 124.410 124.840 ;
        RECT 120.470 119.080 120.730 119.400 ;
        RECT 121.850 119.080 122.110 119.400 ;
        RECT 123.690 119.080 123.950 119.400 ;
        RECT 120.530 117.700 120.670 119.080 ;
        RECT 120.470 117.380 120.730 117.700 ;
        RECT 114.950 113.640 115.210 113.960 ;
        RECT 117.250 113.640 117.510 113.960 ;
        RECT 119.090 113.640 119.350 113.960 ;
        RECT 115.010 111.920 115.150 113.640 ;
        RECT 116.790 113.300 117.050 113.620 ;
        RECT 115.410 112.960 115.670 113.280 ;
        RECT 115.470 111.920 115.610 112.960 ;
        RECT 116.850 111.920 116.990 113.300 ;
        RECT 120.010 112.960 120.270 113.280 ;
        RECT 114.950 111.600 115.210 111.920 ;
        RECT 115.410 111.600 115.670 111.920 ;
        RECT 116.790 111.600 117.050 111.920 ;
        RECT 110.350 110.580 110.610 110.900 ;
        RECT 101.610 110.240 101.870 110.560 ;
        RECT 105.290 110.240 105.550 110.560 ;
        RECT 105.750 110.240 106.010 110.560 ;
        RECT 107.590 110.240 107.850 110.560 ;
        RECT 101.670 106.480 101.810 110.240 ;
        RECT 105.350 106.480 105.490 110.240 ;
        RECT 105.810 108.180 105.950 110.240 ;
        RECT 107.650 108.860 107.790 110.240 ;
        RECT 107.130 108.540 107.390 108.860 ;
        RECT 107.590 108.540 107.850 108.860 ;
        RECT 105.750 107.860 106.010 108.180 ;
        RECT 101.610 106.160 101.870 106.480 ;
        RECT 105.290 106.160 105.550 106.480 ;
        RECT 101.610 105.480 101.870 105.800 ;
        RECT 101.150 102.760 101.410 103.080 ;
        RECT 96.600 101.545 98.140 101.915 ;
        RECT 101.670 100.690 101.810 105.480 ;
        RECT 89.640 99.960 91.690 100.100 ;
        RECT 89.640 98.690 89.920 99.960 ;
        RECT 95.620 98.690 95.900 100.690 ;
        RECT 101.600 98.690 101.880 100.690 ;
        RECT 107.190 100.100 107.330 108.540 ;
        RECT 110.410 108.430 110.550 110.580 ;
        RECT 115.410 110.240 115.670 110.560 ;
        RECT 110.860 109.705 112.400 110.075 ;
        RECT 110.810 108.430 111.070 108.520 ;
        RECT 110.410 108.290 111.070 108.430 ;
        RECT 110.410 106.140 110.550 108.290 ;
        RECT 110.810 108.200 111.070 108.290 ;
        RECT 115.470 106.480 115.610 110.240 ;
        RECT 120.070 108.860 120.210 112.960 ;
        RECT 122.310 109.220 122.570 109.540 ;
        RECT 118.630 108.540 118.890 108.860 ;
        RECT 120.010 108.540 120.270 108.860 ;
        RECT 117.250 107.860 117.510 108.180 ;
        RECT 115.410 106.160 115.670 106.480 ;
        RECT 110.350 105.820 110.610 106.140 ;
        RECT 113.110 105.480 113.370 105.800 ;
        RECT 110.860 104.265 112.400 104.635 ;
        RECT 107.580 100.100 107.860 100.690 ;
        RECT 107.190 99.960 107.860 100.100 ;
        RECT 113.170 100.100 113.310 105.480 ;
        RECT 117.310 104.100 117.450 107.860 ;
        RECT 117.250 103.780 117.510 104.100 ;
        RECT 113.560 100.100 113.840 100.690 ;
        RECT 113.170 99.960 113.840 100.100 ;
        RECT 118.690 100.100 118.830 108.540 ;
        RECT 122.370 106.480 122.510 109.220 ;
        RECT 123.750 108.860 123.890 119.080 ;
        RECT 124.140 114.805 124.420 115.175 ;
        RECT 124.210 113.960 124.350 114.805 ;
        RECT 124.150 113.640 124.410 113.960 ;
        RECT 124.150 110.920 124.410 111.240 ;
        RECT 123.690 108.540 123.950 108.860 ;
        RECT 122.310 106.160 122.570 106.480 ;
        RECT 123.750 106.140 123.890 108.540 ;
        RECT 123.690 105.820 123.950 106.140 ;
        RECT 119.540 100.100 119.820 100.690 ;
        RECT 118.690 99.960 119.820 100.100 ;
        RECT 124.210 100.100 124.350 110.920 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 125.520 100.100 125.800 100.690 ;
        RECT 124.210 99.960 125.800 100.100 ;
        RECT 107.580 98.690 107.860 99.960 ;
        RECT 113.560 98.690 113.840 99.960 ;
        RECT 119.540 98.690 119.820 99.960 ;
        RECT 125.520 98.690 125.800 99.960 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 11.020 215.805 12.600 216.135 ;
        RECT 39.540 215.805 41.120 216.135 ;
        RECT 68.060 215.805 69.640 216.135 ;
        RECT 96.580 215.805 98.160 216.135 ;
        RECT 25.280 213.085 26.860 213.415 ;
        RECT 53.800 213.085 55.380 213.415 ;
        RECT 82.320 213.085 83.900 213.415 ;
        RECT 110.840 213.085 112.420 213.415 ;
        RECT 11.020 210.365 12.600 210.695 ;
        RECT 39.540 210.365 41.120 210.695 ;
        RECT 68.060 210.365 69.640 210.695 ;
        RECT 96.580 210.365 98.160 210.695 ;
        RECT 25.280 207.645 26.860 207.975 ;
        RECT 53.800 207.645 55.380 207.975 ;
        RECT 82.320 207.645 83.900 207.975 ;
        RECT 110.840 207.645 112.420 207.975 ;
        RECT 11.020 204.925 12.600 205.255 ;
        RECT 39.540 204.925 41.120 205.255 ;
        RECT 68.060 204.925 69.640 205.255 ;
        RECT 96.580 204.925 98.160 205.255 ;
        RECT 25.280 202.205 26.860 202.535 ;
        RECT 53.800 202.205 55.380 202.535 ;
        RECT 82.320 202.205 83.900 202.535 ;
        RECT 110.840 202.205 112.420 202.535 ;
        RECT 11.020 199.485 12.600 199.815 ;
        RECT 39.540 199.485 41.120 199.815 ;
        RECT 68.060 199.485 69.640 199.815 ;
        RECT 96.580 199.485 98.160 199.815 ;
        RECT 25.280 196.765 26.860 197.095 ;
        RECT 53.800 196.765 55.380 197.095 ;
        RECT 82.320 196.765 83.900 197.095 ;
        RECT 110.840 196.765 112.420 197.095 ;
        RECT 11.020 194.045 12.600 194.375 ;
        RECT 39.540 194.045 41.120 194.375 ;
        RECT 68.060 194.045 69.640 194.375 ;
        RECT 96.580 194.045 98.160 194.375 ;
        RECT 25.280 191.325 26.860 191.655 ;
        RECT 53.800 191.325 55.380 191.655 ;
        RECT 82.320 191.325 83.900 191.655 ;
        RECT 110.840 191.325 112.420 191.655 ;
        RECT 73.515 189.270 73.845 189.275 ;
        RECT 73.515 189.260 74.100 189.270 ;
        RECT 73.290 188.960 74.100 189.260 ;
        RECT 73.515 188.950 74.100 188.960 ;
        RECT 73.515 188.945 73.845 188.950 ;
        RECT 11.020 188.605 12.600 188.935 ;
        RECT 39.540 188.605 41.120 188.935 ;
        RECT 68.060 188.605 69.640 188.935 ;
        RECT 96.580 188.605 98.160 188.935 ;
        RECT 25.280 185.885 26.860 186.215 ;
        RECT 53.800 185.885 55.380 186.215 ;
        RECT 82.320 185.885 83.900 186.215 ;
        RECT 110.840 185.885 112.420 186.215 ;
        RECT 11.020 183.165 12.600 183.495 ;
        RECT 39.540 183.165 41.120 183.495 ;
        RECT 68.060 183.165 69.640 183.495 ;
        RECT 96.580 183.165 98.160 183.495 ;
        RECT 25.280 180.445 26.860 180.775 ;
        RECT 53.800 180.445 55.380 180.775 ;
        RECT 82.320 180.445 83.900 180.775 ;
        RECT 110.840 180.445 112.420 180.775 ;
        RECT 11.020 177.725 12.600 178.055 ;
        RECT 39.540 177.725 41.120 178.055 ;
        RECT 68.060 177.725 69.640 178.055 ;
        RECT 96.580 177.725 98.160 178.055 ;
        RECT 25.280 175.005 26.860 175.335 ;
        RECT 53.800 175.005 55.380 175.335 ;
        RECT 82.320 175.005 83.900 175.335 ;
        RECT 110.840 175.005 112.420 175.335 ;
        RECT 122.735 174.980 123.065 174.995 ;
        RECT 126.650 174.980 128.650 175.130 ;
        RECT 122.735 174.680 128.650 174.980 ;
        RECT 122.735 174.665 123.065 174.680 ;
        RECT 126.650 174.530 128.650 174.680 ;
        RECT 11.020 172.285 12.600 172.615 ;
        RECT 39.540 172.285 41.120 172.615 ;
        RECT 68.060 172.285 69.640 172.615 ;
        RECT 96.580 172.285 98.160 172.615 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 25.280 169.565 26.860 169.895 ;
        RECT 53.800 169.565 55.380 169.895 ;
        RECT 82.320 169.565 83.900 169.895 ;
        RECT 110.840 169.565 112.420 169.895 ;
        RECT 81.080 167.500 81.460 167.510 ;
        RECT 83.635 167.500 83.965 167.515 ;
        RECT 95.595 167.500 95.925 167.515 ;
        RECT 81.080 167.200 95.925 167.500 ;
        RECT 81.080 167.190 81.460 167.200 ;
        RECT 83.635 167.185 83.965 167.200 ;
        RECT 95.595 167.185 95.925 167.200 ;
        RECT 11.020 166.845 12.600 167.175 ;
        RECT 39.540 166.845 41.120 167.175 ;
        RECT 68.060 166.845 69.640 167.175 ;
        RECT 96.580 166.845 98.160 167.175 ;
        RECT 36.255 164.780 36.585 164.795 ;
        RECT 45.915 164.780 46.245 164.795 ;
        RECT 36.255 164.480 46.245 164.780 ;
        RECT 36.255 164.465 36.585 164.480 ;
        RECT 45.915 164.465 46.245 164.480 ;
        RECT 25.280 164.125 26.860 164.455 ;
        RECT 53.800 164.125 55.380 164.455 ;
        RECT 82.320 164.125 83.900 164.455 ;
        RECT 110.840 164.125 112.420 164.455 ;
        RECT 11.020 161.405 12.600 161.735 ;
        RECT 39.540 161.405 41.120 161.735 ;
        RECT 68.060 161.405 69.640 161.735 ;
        RECT 96.580 161.405 98.160 161.735 ;
        RECT 48.215 160.700 48.545 160.715 ;
        RECT 54.195 160.700 54.525 160.715 ;
        RECT 68.915 160.700 69.245 160.715 ;
        RECT 48.215 160.400 69.245 160.700 ;
        RECT 48.215 160.385 48.545 160.400 ;
        RECT 54.195 160.385 54.525 160.400 ;
        RECT 68.915 160.385 69.245 160.400 ;
        RECT 39.935 159.340 40.265 159.355 ;
        RECT 41.520 159.340 41.900 159.350 ;
        RECT 39.935 159.040 41.900 159.340 ;
        RECT 39.935 159.025 40.265 159.040 ;
        RECT 41.520 159.030 41.900 159.040 ;
        RECT 25.280 158.685 26.860 159.015 ;
        RECT 53.800 158.685 55.380 159.015 ;
        RECT 82.320 158.685 83.900 159.015 ;
        RECT 110.840 158.685 112.420 159.015 ;
        RECT 36.255 157.300 36.585 157.315 ;
        RECT 39.015 157.310 39.345 157.315 ;
        RECT 38.760 157.300 39.345 157.310 ;
        RECT 76.275 157.310 76.605 157.315 ;
        RECT 76.275 157.300 76.860 157.310 ;
        RECT 36.255 157.000 39.750 157.300 ;
        RECT 76.050 157.000 76.860 157.300 ;
        RECT 36.255 156.985 36.585 157.000 ;
        RECT 38.760 156.990 39.345 157.000 ;
        RECT 39.015 156.985 39.345 156.990 ;
        RECT 76.275 156.990 76.860 157.000 ;
        RECT 76.275 156.985 76.605 156.990 ;
        RECT 11.020 155.965 12.600 156.295 ;
        RECT 39.540 155.965 41.120 156.295 ;
        RECT 68.060 155.965 69.640 156.295 ;
        RECT 96.580 155.965 98.160 156.295 ;
        RECT 24.295 154.580 24.625 154.595 ;
        RECT 24.080 154.265 24.625 154.580 ;
        RECT 23.375 153.900 23.705 153.915 ;
        RECT 24.080 153.900 24.380 154.265 ;
        RECT 23.375 153.600 24.380 153.900 ;
        RECT 23.375 153.585 23.705 153.600 ;
        RECT 25.280 153.245 26.860 153.575 ;
        RECT 53.800 153.245 55.380 153.575 ;
        RECT 82.320 153.245 83.900 153.575 ;
        RECT 110.840 153.245 112.420 153.575 ;
        RECT 41.775 151.860 42.105 151.875 ;
        RECT 70.295 151.860 70.625 151.875 ;
        RECT 41.775 151.560 70.625 151.860 ;
        RECT 41.775 151.545 42.105 151.560 ;
        RECT 70.295 151.545 70.625 151.560 ;
        RECT 11.020 150.525 12.600 150.855 ;
        RECT 39.540 150.525 41.120 150.855 ;
        RECT 68.060 150.525 69.640 150.855 ;
        RECT 96.580 150.525 98.160 150.855 ;
        RECT 38.760 149.140 39.140 149.150 ;
        RECT 61.095 149.140 61.425 149.155 ;
        RECT 81.080 149.140 81.460 149.150 ;
        RECT 38.760 148.840 81.460 149.140 ;
        RECT 38.760 148.830 39.140 148.840 ;
        RECT 61.095 148.825 61.425 148.840 ;
        RECT 81.080 148.830 81.460 148.840 ;
        RECT 25.280 147.805 26.860 148.135 ;
        RECT 53.800 147.805 55.380 148.135 ;
        RECT 82.320 147.805 83.900 148.135 ;
        RECT 110.840 147.805 112.420 148.135 ;
        RECT 73.720 147.780 74.100 147.790 ;
        RECT 74.435 147.780 74.765 147.795 ;
        RECT 73.720 147.480 74.765 147.780 ;
        RECT 73.720 147.470 74.100 147.480 ;
        RECT 74.435 147.465 74.765 147.480 ;
        RECT 11.020 145.085 12.600 145.415 ;
        RECT 39.540 145.085 41.120 145.415 ;
        RECT 68.060 145.085 69.640 145.415 ;
        RECT 96.580 145.085 98.160 145.415 ;
        RECT 126.650 145.060 128.650 145.210 ;
        RECT 115.160 144.760 128.650 145.060 ;
        RECT 41.315 144.380 41.645 144.395 ;
        RECT 57.875 144.380 58.205 144.395 ;
        RECT 41.315 144.080 58.205 144.380 ;
        RECT 41.315 144.065 41.645 144.080 ;
        RECT 57.875 144.065 58.205 144.080 ;
        RECT 73.055 144.380 73.385 144.395 ;
        RECT 115.160 144.380 115.460 144.760 ;
        RECT 126.650 144.610 128.650 144.760 ;
        RECT 73.055 144.080 115.460 144.380 ;
        RECT 73.055 144.065 73.385 144.080 ;
        RECT 36.715 143.700 37.045 143.715 ;
        RECT 43.155 143.700 43.485 143.715 ;
        RECT 36.715 143.400 43.485 143.700 ;
        RECT 36.715 143.385 37.045 143.400 ;
        RECT 43.155 143.385 43.485 143.400 ;
        RECT 25.280 142.365 26.860 142.695 ;
        RECT 53.800 142.365 55.380 142.695 ;
        RECT 82.320 142.365 83.900 142.695 ;
        RECT 110.840 142.365 112.420 142.695 ;
        RECT 72.800 140.300 73.180 140.310 ;
        RECT 75.355 140.300 75.685 140.315 ;
        RECT 72.800 140.000 75.685 140.300 ;
        RECT 72.800 139.990 73.180 140.000 ;
        RECT 75.355 139.985 75.685 140.000 ;
        RECT 11.020 139.645 12.600 139.975 ;
        RECT 39.540 139.645 41.120 139.975 ;
        RECT 68.060 139.645 69.640 139.975 ;
        RECT 96.580 139.645 98.160 139.975 ;
        RECT 48.215 138.940 48.545 138.955 ;
        RECT 79.035 138.940 79.365 138.955 ;
        RECT 48.215 138.640 79.365 138.940 ;
        RECT 48.215 138.625 48.545 138.640 ;
        RECT 79.035 138.625 79.365 138.640 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 25.280 136.925 26.860 137.255 ;
        RECT 53.800 136.925 55.380 137.255 ;
        RECT 82.320 136.925 83.900 137.255 ;
        RECT 110.840 136.925 112.420 137.255 ;
        RECT 76.735 135.550 77.065 135.555 ;
        RECT 76.480 135.540 77.065 135.550 ;
        RECT 76.280 135.240 77.065 135.540 ;
        RECT 76.480 135.230 77.065 135.240 ;
        RECT 76.735 135.225 77.065 135.230 ;
        RECT 11.020 134.205 12.600 134.535 ;
        RECT 39.540 134.205 41.120 134.535 ;
        RECT 68.060 134.205 69.640 134.535 ;
        RECT 96.580 134.205 98.160 134.535 ;
        RECT 25.280 131.485 26.860 131.815 ;
        RECT 53.800 131.485 55.380 131.815 ;
        RECT 82.320 131.485 83.900 131.815 ;
        RECT 110.840 131.485 112.420 131.815 ;
        RECT 11.020 128.765 12.600 129.095 ;
        RECT 39.540 128.765 41.120 129.095 ;
        RECT 68.060 128.765 69.640 129.095 ;
        RECT 96.580 128.765 98.160 129.095 ;
        RECT 41.520 128.740 41.900 128.750 ;
        RECT 42.695 128.740 43.025 128.755 ;
        RECT 41.520 128.440 43.025 128.740 ;
        RECT 41.520 128.430 41.900 128.440 ;
        RECT 42.695 128.425 43.025 128.440 ;
        RECT 41.775 128.060 42.105 128.075 ;
        RECT 50.055 128.060 50.385 128.075 ;
        RECT 41.775 127.760 50.385 128.060 ;
        RECT 41.775 127.745 42.105 127.760 ;
        RECT 50.055 127.745 50.385 127.760 ;
        RECT 39.935 127.380 40.265 127.395 ;
        RECT 49.595 127.380 49.925 127.395 ;
        RECT 39.935 127.080 49.925 127.380 ;
        RECT 39.935 127.065 40.265 127.080 ;
        RECT 49.595 127.065 49.925 127.080 ;
        RECT 25.280 126.045 26.860 126.375 ;
        RECT 53.800 126.045 55.380 126.375 ;
        RECT 82.320 126.045 83.900 126.375 ;
        RECT 110.840 126.045 112.420 126.375 ;
        RECT 38.095 125.340 38.425 125.355 ;
        RECT 38.760 125.340 39.140 125.350 ;
        RECT 38.095 125.040 39.140 125.340 ;
        RECT 38.095 125.025 38.425 125.040 ;
        RECT 38.760 125.030 39.140 125.040 ;
        RECT 81.080 125.340 81.460 125.350 ;
        RECT 92.835 125.340 93.165 125.355 ;
        RECT 81.080 125.040 93.165 125.340 ;
        RECT 81.080 125.030 81.460 125.040 ;
        RECT 92.835 125.025 93.165 125.040 ;
        RECT 11.020 123.325 12.600 123.655 ;
        RECT 39.540 123.325 41.120 123.655 ;
        RECT 68.060 123.325 69.640 123.655 ;
        RECT 96.580 123.325 98.160 123.655 ;
        RECT 25.280 120.605 26.860 120.935 ;
        RECT 53.800 120.605 55.380 120.935 ;
        RECT 82.320 120.605 83.900 120.935 ;
        RECT 110.840 120.605 112.420 120.935 ;
        RECT 11.020 117.885 12.600 118.215 ;
        RECT 39.540 117.885 41.120 118.215 ;
        RECT 68.060 117.885 69.640 118.215 ;
        RECT 96.580 117.885 98.160 118.215 ;
        RECT 25.280 115.165 26.860 115.495 ;
        RECT 53.800 115.165 55.380 115.495 ;
        RECT 82.320 115.165 83.900 115.495 ;
        RECT 110.840 115.165 112.420 115.495 ;
        RECT 72.595 115.150 72.925 115.155 ;
        RECT 72.595 115.140 73.180 115.150 ;
        RECT 124.115 115.140 124.445 115.155 ;
        RECT 126.650 115.140 128.650 115.290 ;
        RECT 72.595 114.840 73.380 115.140 ;
        RECT 124.115 114.840 128.650 115.140 ;
        RECT 72.595 114.830 73.180 114.840 ;
        RECT 72.595 114.825 72.925 114.830 ;
        RECT 124.115 114.825 124.445 114.840 ;
        RECT 126.650 114.690 128.650 114.840 ;
        RECT 11.020 112.445 12.600 112.775 ;
        RECT 39.540 112.445 41.120 112.775 ;
        RECT 68.060 112.445 69.640 112.775 ;
        RECT 96.580 112.445 98.160 112.775 ;
        RECT 25.280 109.725 26.860 110.055 ;
        RECT 53.800 109.725 55.380 110.055 ;
        RECT 82.320 109.725 83.900 110.055 ;
        RECT 110.840 109.725 112.420 110.055 ;
        RECT 11.020 107.005 12.600 107.335 ;
        RECT 39.540 107.005 41.120 107.335 ;
        RECT 68.060 107.005 69.640 107.335 ;
        RECT 96.580 107.005 98.160 107.335 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 25.280 104.285 26.860 104.615 ;
        RECT 53.800 104.285 55.380 104.615 ;
        RECT 82.320 104.285 83.900 104.615 ;
        RECT 110.840 104.285 112.420 104.615 ;
        RECT 11.020 101.565 12.600 101.895 ;
        RECT 39.540 101.565 41.120 101.895 ;
        RECT 68.060 101.565 69.640 101.895 ;
        RECT 96.580 101.565 98.160 101.895 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 11.010 101.490 12.610 216.210 ;
        RECT 25.270 101.490 26.870 216.210 ;
        RECT 38.785 156.985 39.115 157.315 ;
        RECT 38.800 149.155 39.100 156.985 ;
        RECT 38.785 148.825 39.115 149.155 ;
        RECT 38.800 125.355 39.100 148.825 ;
        RECT 38.785 125.025 39.115 125.355 ;
        RECT 39.530 101.490 41.130 216.210 ;
        RECT 41.545 159.025 41.875 159.355 ;
        RECT 41.560 128.755 41.860 159.025 ;
        RECT 41.545 128.425 41.875 128.755 ;
        RECT 53.790 101.490 55.390 216.210 ;
        RECT 68.050 101.490 69.650 216.210 ;
        RECT 73.745 188.945 74.075 189.275 ;
        RECT 73.760 147.795 74.060 188.945 ;
        RECT 81.105 167.185 81.435 167.515 ;
        RECT 76.505 156.985 76.835 157.315 ;
        RECT 73.745 147.465 74.075 147.795 ;
        RECT 72.825 139.985 73.155 140.315 ;
        RECT 72.840 115.155 73.140 139.985 ;
        RECT 76.520 135.555 76.820 156.985 ;
        RECT 81.120 149.155 81.420 167.185 ;
        RECT 81.105 148.825 81.435 149.155 ;
        RECT 76.505 135.225 76.835 135.555 ;
        RECT 81.120 125.355 81.420 148.825 ;
        RECT 81.105 125.025 81.435 125.355 ;
        RECT 72.825 114.825 73.155 115.155 ;
        RECT 82.310 101.490 83.910 216.210 ;
        RECT 96.570 101.490 98.170 216.210 ;
        RECT 110.830 101.490 112.430 216.210 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

