VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 27.115 203.925 27.285 204.115 ;
        RECT 28.550 203.975 28.670 204.085 ;
        RECT 29.875 203.925 30.045 204.115 ;
        RECT 30.335 203.925 30.505 204.115 ;
        RECT 31.715 203.925 31.885 204.115 ;
        RECT 35.395 203.925 35.565 204.115 ;
        RECT 38.615 203.925 38.785 204.115 ;
        RECT 39.075 203.925 39.245 204.115 ;
        RECT 41.375 203.925 41.545 204.115 ;
        RECT 41.835 203.925 42.005 204.115 ;
        RECT 43.215 203.925 43.385 204.115 ;
        RECT 44.595 203.925 44.765 204.115 ;
        RECT 45.975 203.925 46.145 204.115 ;
        RECT 47.355 203.925 47.525 204.115 ;
        RECT 49.655 203.970 49.815 204.080 ;
        RECT 50.115 203.925 50.285 204.115 ;
        RECT 52.415 203.925 52.585 204.115 ;
        RECT 52.930 203.975 53.050 204.085 ;
        RECT 53.335 203.925 53.505 204.115 ;
        RECT 54.715 203.925 54.885 204.115 ;
        RECT 56.090 203.925 56.260 204.115 ;
        RECT 58.395 203.925 58.565 204.115 ;
        RECT 58.855 203.925 59.025 204.115 ;
        RECT 61.155 203.925 61.325 204.115 ;
        RECT 63.455 203.925 63.625 204.115 ;
        RECT 26.975 203.115 28.345 203.925 ;
        RECT 28.825 203.015 30.175 203.925 ;
        RECT 30.205 203.015 31.555 203.925 ;
        RECT 31.585 203.015 32.935 203.925 ;
        RECT 32.955 203.115 35.705 203.925 ;
        RECT 35.725 203.055 36.155 203.840 ;
        RECT 36.175 203.115 38.925 203.925 ;
        RECT 38.935 203.145 40.305 203.925 ;
        RECT 40.325 203.015 41.675 203.925 ;
        RECT 41.705 203.015 43.055 203.925 ;
        RECT 43.075 203.145 44.445 203.925 ;
        RECT 44.465 203.015 45.815 203.925 ;
        RECT 45.835 203.145 47.205 203.925 ;
        RECT 47.215 203.145 48.585 203.925 ;
        RECT 48.605 203.055 49.035 203.840 ;
        RECT 49.985 203.015 51.335 203.925 ;
        RECT 51.365 203.015 52.715 203.925 ;
        RECT 53.195 203.145 54.565 203.925 ;
        RECT 54.575 203.145 55.945 203.925 ;
        RECT 55.975 203.015 57.325 203.925 ;
        RECT 57.345 203.015 58.695 203.925 ;
        RECT 58.725 203.015 60.075 203.925 ;
        RECT 60.095 203.145 61.465 203.925 ;
        RECT 61.485 203.055 61.915 203.840 ;
        RECT 61.935 203.245 63.765 203.925 ;
        RECT 63.915 203.895 64.085 204.115 ;
        RECT 67.140 203.925 67.310 204.115 ;
        RECT 70.410 203.975 70.530 204.085 ;
        RECT 74.035 203.925 74.205 204.115 ;
        RECT 74.955 203.925 75.125 204.115 ;
        RECT 85.535 203.925 85.705 204.115 ;
        RECT 86.915 203.925 87.085 204.115 ;
        RECT 88.295 203.970 88.455 204.080 ;
        RECT 88.755 203.925 88.925 204.115 ;
        RECT 95.655 203.925 95.825 204.115 ;
        RECT 96.390 203.925 96.560 204.115 ;
        RECT 109.455 203.925 109.625 204.115 ;
        RECT 109.915 203.925 110.085 204.115 ;
        RECT 111.755 203.970 111.915 204.080 ;
        RECT 113.135 203.925 113.305 204.115 ;
        RECT 66.040 203.895 66.985 203.925 ;
        RECT 63.915 203.695 66.985 203.895 ;
        RECT 63.775 203.215 66.985 203.695 ;
        RECT 63.775 203.015 64.705 203.215 ;
        RECT 66.040 203.015 66.985 203.215 ;
        RECT 66.995 203.015 69.915 203.925 ;
        RECT 70.770 203.245 74.235 203.925 ;
        RECT 70.770 203.015 71.690 203.245 ;
        RECT 74.365 203.055 74.795 203.840 ;
        RECT 74.815 203.245 76.645 203.925 ;
        RECT 76.655 203.245 85.845 203.925 ;
        RECT 76.655 203.015 77.575 203.245 ;
        RECT 80.405 203.025 81.335 203.245 ;
        RECT 85.865 203.015 87.215 203.925 ;
        RECT 87.245 203.055 87.675 203.840 ;
        RECT 88.725 203.245 92.190 203.925 ;
        RECT 91.270 203.015 92.190 203.245 ;
        RECT 92.390 203.245 95.855 203.925 ;
        RECT 95.975 203.245 99.875 203.925 ;
        RECT 92.390 203.015 93.310 203.245 ;
        RECT 95.975 203.015 96.905 203.245 ;
        RECT 100.125 203.055 100.555 203.840 ;
        RECT 100.575 203.245 109.765 203.925 ;
        RECT 100.575 203.015 101.495 203.245 ;
        RECT 104.325 203.025 105.255 203.245 ;
        RECT 109.785 203.015 111.135 203.925 ;
        RECT 112.075 203.115 113.445 203.925 ;
      LAYER nwell ;
        RECT 26.780 199.895 113.640 202.725 ;
      LAYER pwell ;
        RECT 26.975 198.695 28.345 199.505 ;
        RECT 28.815 198.695 30.185 199.475 ;
        RECT 30.205 198.695 31.555 199.605 ;
        RECT 31.585 198.695 32.935 199.605 ;
        RECT 32.965 198.695 34.315 199.605 ;
        RECT 34.335 198.695 35.705 199.475 ;
        RECT 35.725 198.780 36.155 199.565 ;
        RECT 36.635 198.695 38.005 199.475 ;
        RECT 38.015 198.695 39.385 199.475 ;
        RECT 39.395 198.695 42.870 199.605 ;
        RECT 43.085 198.695 44.435 199.605 ;
        RECT 44.465 198.695 45.815 199.605 ;
        RECT 45.835 198.695 47.205 199.475 ;
        RECT 47.225 198.695 48.575 199.605 ;
        RECT 48.690 199.375 49.610 199.605 ;
        RECT 56.785 199.375 57.715 199.595 ;
        RECT 60.545 199.375 61.465 199.605 ;
        RECT 48.690 198.695 52.155 199.375 ;
        RECT 52.275 198.695 61.465 199.375 ;
        RECT 61.485 198.780 61.915 199.565 ;
        RECT 64.590 199.375 65.510 199.605 ;
        RECT 62.045 198.695 65.510 199.375 ;
        RECT 65.615 198.695 68.725 199.605 ;
        RECT 69.320 199.375 70.665 199.605 ;
        RECT 75.185 199.375 76.115 199.595 ;
        RECT 78.945 199.375 79.865 199.605 ;
        RECT 82.530 199.375 83.450 199.605 ;
        RECT 86.210 199.375 87.130 199.605 ;
        RECT 68.835 198.695 70.665 199.375 ;
        RECT 70.675 198.695 79.865 199.375 ;
        RECT 79.985 198.695 83.450 199.375 ;
        RECT 83.665 198.695 87.130 199.375 ;
        RECT 87.245 198.780 87.675 199.565 ;
        RECT 87.705 198.695 89.055 199.605 ;
        RECT 93.585 199.375 94.515 199.595 ;
        RECT 97.345 199.375 98.265 199.605 ;
        RECT 102.785 199.375 103.715 199.595 ;
        RECT 106.545 199.375 107.465 199.605 ;
        RECT 110.130 199.375 111.050 199.605 ;
        RECT 89.075 198.695 98.265 199.375 ;
        RECT 98.275 198.695 107.465 199.375 ;
        RECT 107.585 198.695 111.050 199.375 ;
        RECT 112.075 198.695 113.445 199.505 ;
        RECT 27.115 198.485 27.285 198.695 ;
        RECT 28.495 198.645 28.665 198.675 ;
        RECT 28.495 198.535 28.670 198.645 ;
        RECT 28.495 198.485 28.665 198.535 ;
        RECT 28.955 198.505 29.125 198.695 ;
        RECT 30.335 198.505 30.505 198.695 ;
        RECT 31.715 198.505 31.885 198.695 ;
        RECT 33.095 198.485 33.265 198.675 ;
        RECT 33.555 198.485 33.725 198.675 ;
        RECT 34.015 198.505 34.185 198.695 ;
        RECT 34.475 198.505 34.645 198.695 ;
        RECT 34.935 198.485 35.105 198.675 ;
        RECT 36.370 198.535 36.490 198.645 ;
        RECT 36.775 198.505 36.945 198.695 ;
        RECT 38.155 198.505 38.325 198.695 ;
        RECT 39.540 198.675 39.710 198.695 ;
        RECT 39.535 198.505 39.710 198.675 ;
        RECT 39.535 198.485 39.705 198.505 ;
        RECT 39.995 198.485 40.165 198.675 ;
        RECT 44.135 198.505 44.305 198.695 ;
        RECT 44.590 198.485 44.760 198.675 ;
        RECT 45.055 198.485 45.225 198.675 ;
        RECT 45.515 198.505 45.685 198.695 ;
        RECT 45.975 198.505 46.145 198.695 ;
        RECT 47.355 198.505 47.525 198.695 ;
        RECT 51.955 198.505 52.125 198.695 ;
        RECT 52.415 198.485 52.585 198.695 ;
        RECT 52.930 198.535 53.050 198.645 ;
        RECT 56.555 198.485 56.725 198.675 ;
        RECT 57.015 198.485 57.185 198.675 ;
        RECT 62.075 198.505 62.245 198.695 ;
        RECT 68.515 198.505 68.685 198.695 ;
        RECT 68.975 198.505 69.145 198.695 ;
        RECT 69.430 198.485 69.600 198.675 ;
        RECT 69.895 198.485 70.065 198.675 ;
        RECT 70.815 198.505 70.985 198.695 ;
        RECT 74.035 198.530 74.195 198.640 ;
        RECT 74.955 198.485 75.125 198.675 ;
        RECT 76.335 198.485 76.505 198.675 ;
        RECT 79.555 198.485 79.725 198.675 ;
        RECT 80.015 198.505 80.185 198.695 ;
        RECT 83.235 198.485 83.405 198.675 ;
        RECT 83.695 198.505 83.865 198.695 ;
        RECT 88.755 198.505 88.925 198.695 ;
        RECT 89.215 198.505 89.385 198.695 ;
        RECT 94.735 198.505 94.905 198.675 ;
        RECT 94.735 198.485 94.900 198.505 ;
        RECT 95.470 198.485 95.640 198.675 ;
        RECT 98.415 198.505 98.585 198.695 ;
        RECT 99.795 198.530 99.955 198.640 ;
        RECT 101.175 198.530 101.335 198.640 ;
        RECT 107.615 198.505 107.785 198.695 ;
        RECT 110.375 198.485 110.545 198.675 ;
        RECT 111.755 198.485 111.925 198.675 ;
        RECT 113.135 198.485 113.305 198.695 ;
        RECT 26.975 197.675 28.345 198.485 ;
        RECT 28.465 197.805 31.930 198.485 ;
        RECT 31.010 197.575 31.930 197.805 ;
        RECT 32.045 197.575 33.395 198.485 ;
        RECT 33.425 197.575 34.775 198.485 ;
        RECT 34.905 197.805 38.370 198.485 ;
        RECT 37.450 197.575 38.370 197.805 ;
        RECT 38.475 197.705 39.845 198.485 ;
        RECT 39.855 197.705 41.225 198.485 ;
        RECT 41.430 197.575 44.905 198.485 ;
        RECT 45.025 197.805 48.490 198.485 ;
        RECT 47.570 197.575 48.490 197.805 ;
        RECT 48.605 197.615 49.035 198.400 ;
        RECT 49.150 197.805 52.615 198.485 ;
        RECT 53.290 197.805 56.755 198.485 ;
        RECT 56.875 197.805 67.245 198.485 ;
        RECT 49.150 197.575 50.070 197.805 ;
        RECT 53.290 197.575 54.210 197.805 ;
        RECT 61.385 197.585 62.315 197.805 ;
        RECT 65.035 197.575 67.245 197.805 ;
        RECT 67.455 197.575 69.745 198.485 ;
        RECT 69.755 197.805 73.425 198.485 ;
        RECT 72.495 197.575 73.425 197.805 ;
        RECT 74.365 197.615 74.795 198.400 ;
        RECT 74.825 197.575 76.175 198.485 ;
        RECT 76.295 197.575 79.405 198.485 ;
        RECT 79.525 197.805 82.990 198.485 ;
        RECT 83.095 197.805 92.375 198.485 ;
        RECT 82.070 197.575 82.990 197.805 ;
        RECT 84.455 197.585 85.375 197.805 ;
        RECT 90.040 197.685 92.375 197.805 ;
        RECT 91.455 197.575 92.375 197.685 ;
        RECT 93.065 197.805 94.900 198.485 ;
        RECT 95.055 197.805 98.955 198.485 ;
        RECT 93.065 197.575 93.995 197.805 ;
        RECT 95.055 197.575 95.985 197.805 ;
        RECT 100.125 197.615 100.555 198.400 ;
        RECT 101.495 197.805 110.685 198.485 ;
        RECT 101.495 197.575 102.415 197.805 ;
        RECT 105.245 197.585 106.175 197.805 ;
        RECT 110.705 197.575 112.055 198.485 ;
        RECT 112.075 197.675 113.445 198.485 ;
      LAYER nwell ;
        RECT 26.780 194.455 113.640 197.285 ;
      LAYER pwell ;
        RECT 26.975 193.255 28.345 194.065 ;
        RECT 31.010 193.935 31.930 194.165 ;
        RECT 34.690 193.935 35.610 194.165 ;
        RECT 28.465 193.255 31.930 193.935 ;
        RECT 32.145 193.255 35.610 193.935 ;
        RECT 35.725 193.340 36.155 194.125 ;
        RECT 36.645 193.255 37.995 194.165 ;
        RECT 38.015 193.255 39.385 194.035 ;
        RECT 39.395 193.255 42.870 194.165 ;
        RECT 47.585 193.935 48.515 194.155 ;
        RECT 51.345 193.935 52.265 194.165 ;
        RECT 56.785 193.935 57.715 194.155 ;
        RECT 60.545 193.935 61.465 194.165 ;
        RECT 43.075 193.255 52.265 193.935 ;
        RECT 52.275 193.255 61.465 193.935 ;
        RECT 61.485 193.340 61.915 194.125 ;
        RECT 62.395 193.935 63.740 194.165 ;
        RECT 64.235 193.965 65.180 194.165 ;
        RECT 66.515 193.965 67.445 194.165 ;
        RECT 62.395 193.255 64.225 193.935 ;
        RECT 64.235 193.485 67.445 193.965 ;
        RECT 69.035 193.935 72.035 194.165 ;
        RECT 67.455 193.845 72.035 193.935 ;
        RECT 72.055 193.935 72.975 194.165 ;
        RECT 75.805 193.935 76.735 194.155 ;
        RECT 67.455 193.485 72.045 193.845 ;
        RECT 64.235 193.285 67.305 193.485 ;
        RECT 64.235 193.255 65.180 193.285 ;
        RECT 27.115 193.045 27.285 193.255 ;
        RECT 28.495 193.205 28.665 193.255 ;
        RECT 28.495 193.095 28.670 193.205 ;
        RECT 28.495 193.065 28.665 193.095 ;
        RECT 28.955 193.045 29.125 193.235 ;
        RECT 30.795 193.090 30.955 193.200 ;
        RECT 32.175 193.065 32.345 193.255 ;
        RECT 36.370 193.095 36.490 193.205 ;
        RECT 36.775 193.065 36.945 193.255 ;
        RECT 38.155 193.065 38.325 193.255 ;
        RECT 39.540 193.065 39.710 193.255 ;
        RECT 40.455 193.045 40.625 193.235 ;
        RECT 40.915 193.045 41.085 193.235 ;
        RECT 42.295 193.045 42.465 193.235 ;
        RECT 43.215 193.065 43.385 193.255 ;
        RECT 43.950 193.045 44.120 193.235 ;
        RECT 48.275 193.090 48.435 193.200 ;
        RECT 49.195 193.045 49.365 193.235 ;
        RECT 50.575 193.045 50.745 193.235 ;
        RECT 52.415 193.065 52.585 193.255 ;
        RECT 52.690 193.045 52.860 193.235 ;
        RECT 56.610 193.095 56.730 193.205 ;
        RECT 57.015 193.045 57.185 193.235 ;
        RECT 62.130 193.095 62.250 193.205 ;
        RECT 63.915 193.065 64.085 193.255 ;
        RECT 67.135 193.065 67.305 193.285 ;
        RECT 67.455 193.255 69.025 193.485 ;
        RECT 71.115 193.295 72.045 193.485 ;
        RECT 71.115 193.255 72.035 193.295 ;
        RECT 72.055 193.255 81.245 193.935 ;
        RECT 81.265 193.255 82.615 194.165 ;
        RECT 83.095 193.935 84.025 194.165 ;
        RECT 83.095 193.255 86.995 193.935 ;
        RECT 87.245 193.340 87.675 194.125 ;
        RECT 87.705 193.255 89.055 194.165 ;
        RECT 89.535 193.935 90.465 194.165 ;
        RECT 89.535 193.255 93.435 193.935 ;
        RECT 93.675 193.255 97.150 194.165 ;
        RECT 97.355 193.935 98.285 194.165 ;
        RECT 101.495 193.935 102.425 194.165 ;
        RECT 97.355 193.255 101.255 193.935 ;
        RECT 101.495 193.255 105.395 193.935 ;
        RECT 105.635 193.255 109.110 194.165 ;
        RECT 109.315 193.255 110.685 194.035 ;
        RECT 110.705 193.255 112.055 194.165 ;
        RECT 112.075 193.255 113.445 194.065 ;
        RECT 67.595 193.065 67.765 193.255 ;
        RECT 68.055 193.045 68.225 193.235 ;
        RECT 68.520 193.045 68.690 193.235 ;
        RECT 71.275 193.065 71.445 193.235 ;
        RECT 71.375 193.045 71.445 193.065 ;
        RECT 78.175 193.045 78.345 193.235 ;
        RECT 78.635 193.045 78.805 193.235 ;
        RECT 80.935 193.065 81.105 193.255 ;
        RECT 82.315 193.065 82.485 193.255 ;
        RECT 82.830 193.095 82.950 193.205 ;
        RECT 83.510 193.065 83.680 193.255 ;
        RECT 88.755 193.065 88.925 193.255 ;
        RECT 89.270 193.095 89.390 193.205 ;
        RECT 89.950 193.065 90.120 193.255 ;
        RECT 91.515 193.045 91.685 193.235 ;
        RECT 92.435 193.090 92.595 193.200 ;
        RECT 93.820 193.065 93.990 193.255 ;
        RECT 96.300 193.045 96.470 193.235 ;
        RECT 97.770 193.065 97.940 193.255 ;
        RECT 97.955 193.045 98.125 193.235 ;
        RECT 98.470 193.095 98.590 193.205 ;
        RECT 99.795 193.045 99.965 193.235 ;
        RECT 101.635 193.045 101.805 193.235 ;
        RECT 101.910 193.065 102.080 193.255 ;
        RECT 102.150 193.095 102.270 193.205 ;
        RECT 102.555 193.045 102.725 193.235 ;
        RECT 105.780 193.065 105.950 193.255 ;
        RECT 110.375 193.065 110.545 193.255 ;
        RECT 111.755 193.205 111.925 193.255 ;
        RECT 111.755 193.095 111.930 193.205 ;
        RECT 111.755 193.065 111.925 193.095 ;
        RECT 113.135 193.045 113.305 193.255 ;
        RECT 26.975 192.235 28.345 193.045 ;
        RECT 28.815 192.265 30.185 193.045 ;
        RECT 31.485 192.365 40.765 193.045 ;
        RECT 31.485 192.245 33.820 192.365 ;
        RECT 31.485 192.135 32.405 192.245 ;
        RECT 38.485 192.145 39.405 192.365 ;
        RECT 40.775 192.265 42.145 193.045 ;
        RECT 42.155 192.265 43.525 193.045 ;
        RECT 43.535 192.365 47.435 193.045 ;
        RECT 43.535 192.135 44.465 192.365 ;
        RECT 48.605 192.175 49.035 192.960 ;
        RECT 49.065 192.135 50.415 193.045 ;
        RECT 50.435 192.365 52.265 193.045 ;
        RECT 52.275 192.365 56.175 193.045 ;
        RECT 56.875 192.365 66.065 193.045 ;
        RECT 52.275 192.135 53.205 192.365 ;
        RECT 61.385 192.145 62.315 192.365 ;
        RECT 65.145 192.135 66.065 192.365 ;
        RECT 66.075 192.365 68.365 193.045 ;
        RECT 66.075 192.135 66.995 192.365 ;
        RECT 68.375 192.135 70.985 193.045 ;
        RECT 71.375 192.815 73.645 193.045 ;
        RECT 71.375 192.135 74.130 192.815 ;
        RECT 74.365 192.175 74.795 192.960 ;
        RECT 74.910 192.365 78.375 193.045 ;
        RECT 78.605 192.365 82.070 193.045 ;
        RECT 74.910 192.135 75.830 192.365 ;
        RECT 81.150 192.135 82.070 192.365 ;
        RECT 82.545 192.365 91.825 193.045 ;
        RECT 92.985 192.365 96.885 193.045 ;
        RECT 82.545 192.245 84.880 192.365 ;
        RECT 82.545 192.135 83.465 192.245 ;
        RECT 89.545 192.145 90.465 192.365 ;
        RECT 95.955 192.135 96.885 192.365 ;
        RECT 96.895 192.265 98.265 193.045 ;
        RECT 98.735 192.265 100.105 193.045 ;
        RECT 100.125 192.175 100.555 192.960 ;
        RECT 100.585 192.135 101.935 193.045 ;
        RECT 102.415 192.365 111.605 193.045 ;
        RECT 106.925 192.145 107.855 192.365 ;
        RECT 110.685 192.135 111.605 192.365 ;
        RECT 112.075 192.235 113.445 193.045 ;
      LAYER nwell ;
        RECT 26.780 189.015 113.640 191.845 ;
      LAYER pwell ;
        RECT 26.975 187.815 28.345 188.625 ;
        RECT 28.825 187.815 30.175 188.725 ;
        RECT 30.195 187.815 31.565 188.595 ;
        RECT 34.775 188.495 35.705 188.725 ;
        RECT 31.805 187.815 35.705 188.495 ;
        RECT 35.725 187.900 36.155 188.685 ;
        RECT 36.635 187.815 38.005 188.595 ;
        RECT 38.025 187.815 39.375 188.725 ;
        RECT 39.590 187.815 43.065 188.725 ;
        RECT 43.075 188.495 43.995 188.725 ;
        RECT 46.825 188.495 47.755 188.715 ;
        RECT 43.075 187.815 52.265 188.495 ;
        RECT 52.470 187.815 55.945 188.725 ;
        RECT 55.955 188.495 56.885 188.725 ;
        RECT 55.955 187.815 59.855 188.495 ;
        RECT 60.095 187.815 61.465 188.595 ;
        RECT 61.485 187.900 61.915 188.685 ;
        RECT 62.030 188.495 62.950 188.725 ;
        RECT 62.030 187.815 65.495 188.495 ;
        RECT 65.615 187.815 68.355 188.495 ;
        RECT 68.615 188.045 71.370 188.725 ;
        RECT 74.250 188.495 75.170 188.725 ;
        RECT 77.930 188.495 78.850 188.725 ;
        RECT 82.155 188.495 83.085 188.725 ;
        RECT 86.295 188.495 87.225 188.725 ;
        RECT 68.615 187.815 70.885 188.045 ;
        RECT 71.705 187.815 75.170 188.495 ;
        RECT 75.385 187.815 78.850 188.495 ;
        RECT 79.185 187.815 83.085 188.495 ;
        RECT 83.325 187.815 87.225 188.495 ;
        RECT 87.245 187.900 87.675 188.685 ;
        RECT 87.695 187.815 89.065 188.595 ;
        RECT 89.535 188.495 90.455 188.725 ;
        RECT 93.285 188.495 94.215 188.715 ;
        RECT 89.535 187.815 98.725 188.495 ;
        RECT 98.735 187.815 100.105 188.595 ;
        RECT 100.575 188.495 101.495 188.725 ;
        RECT 104.325 188.495 105.255 188.715 ;
        RECT 100.575 187.815 109.765 188.495 ;
        RECT 109.775 187.815 111.145 188.595 ;
        RECT 112.075 187.815 113.445 188.625 ;
        RECT 27.115 187.605 27.285 187.815 ;
        RECT 28.550 187.655 28.670 187.765 ;
        RECT 29.875 187.625 30.045 187.815 ;
        RECT 30.335 187.625 30.505 187.815 ;
        RECT 35.120 187.625 35.290 187.815 ;
        RECT 36.370 187.655 36.490 187.765 ;
        RECT 36.775 187.625 36.945 187.815 ;
        RECT 37.695 187.605 37.865 187.795 ;
        RECT 38.155 187.625 38.325 187.815 ;
        RECT 42.750 187.625 42.920 187.815 ;
        RECT 46.895 187.605 47.065 187.795 ;
        RECT 47.355 187.605 47.525 187.795 ;
        RECT 49.250 187.655 49.370 187.765 ;
        RECT 49.930 187.605 50.100 187.795 ;
        RECT 51.955 187.625 52.125 187.815 ;
        RECT 53.795 187.605 53.965 187.795 ;
        RECT 55.630 187.625 55.800 187.815 ;
        RECT 56.370 187.625 56.540 187.815 ;
        RECT 58.395 187.605 58.565 187.795 ;
        RECT 59.130 187.605 59.300 187.795 ;
        RECT 60.235 187.625 60.405 187.815 ;
        RECT 63.455 187.650 63.615 187.760 ;
        RECT 65.295 187.605 65.465 187.815 ;
        RECT 65.755 187.625 65.925 187.815 ;
        RECT 68.615 187.795 68.685 187.815 ;
        RECT 68.515 187.625 68.685 187.795 ;
        RECT 71.735 187.625 71.905 187.815 ;
        RECT 68.515 187.605 68.585 187.625 ;
        RECT 73.115 187.605 73.285 187.795 ;
        RECT 74.035 187.650 74.195 187.760 ;
        RECT 75.415 187.625 75.585 187.815 ;
        RECT 76.795 187.605 76.965 187.795 ;
        RECT 77.260 187.605 77.430 187.795 ;
        RECT 82.500 187.625 82.670 187.815 ;
        RECT 86.640 187.625 86.810 187.815 ;
        RECT 88.755 187.625 88.925 187.815 ;
        RECT 89.270 187.655 89.390 187.765 ;
        RECT 89.675 187.605 89.845 187.795 ;
        RECT 90.135 187.605 90.305 187.795 ;
        RECT 93.820 187.605 93.990 187.795 ;
        RECT 97.500 187.605 97.670 187.795 ;
        RECT 98.415 187.625 98.585 187.815 ;
        RECT 99.795 187.625 99.965 187.815 ;
        RECT 100.310 187.655 100.430 187.765 ;
        RECT 104.120 187.605 104.290 187.795 ;
        RECT 108.075 187.605 108.245 187.795 ;
        RECT 109.455 187.625 109.625 187.815 ;
        RECT 110.835 187.625 111.005 187.815 ;
        RECT 111.750 187.605 111.920 187.795 ;
        RECT 113.135 187.605 113.305 187.815 ;
        RECT 26.975 186.795 28.345 187.605 ;
        RECT 28.815 186.925 38.005 187.605 ;
        RECT 38.015 186.925 47.205 187.605 ;
        RECT 28.815 186.695 29.735 186.925 ;
        RECT 32.565 186.705 33.495 186.925 ;
        RECT 38.015 186.695 38.935 186.925 ;
        RECT 41.765 186.705 42.695 186.925 ;
        RECT 47.215 186.825 48.585 187.605 ;
        RECT 48.605 186.735 49.035 187.520 ;
        RECT 49.515 186.925 53.415 187.605 ;
        RECT 49.515 186.695 50.445 186.925 ;
        RECT 53.655 186.825 55.025 187.605 ;
        RECT 55.130 186.925 58.595 187.605 ;
        RECT 58.715 186.925 62.615 187.605 ;
        RECT 63.775 186.925 65.605 187.605 ;
        RECT 66.315 187.375 68.585 187.605 ;
        RECT 68.845 187.565 69.765 187.605 ;
        RECT 55.130 186.695 56.050 186.925 ;
        RECT 58.715 186.695 59.645 186.925 ;
        RECT 63.775 186.695 65.120 186.925 ;
        RECT 65.830 186.695 68.585 187.375 ;
        RECT 68.835 187.375 69.765 187.565 ;
        RECT 71.855 187.375 73.425 187.605 ;
        RECT 68.835 187.015 73.425 187.375 ;
        RECT 68.845 186.925 73.425 187.015 ;
        RECT 68.845 186.695 71.845 186.925 ;
        RECT 74.365 186.735 74.795 187.520 ;
        RECT 74.815 186.925 77.105 187.605 ;
        RECT 74.815 186.695 75.735 186.925 ;
        RECT 77.115 186.695 80.590 187.605 ;
        RECT 80.795 186.925 89.985 187.605 ;
        RECT 90.105 186.925 93.570 187.605 ;
        RECT 80.795 186.695 81.715 186.925 ;
        RECT 84.545 186.705 85.475 186.925 ;
        RECT 92.650 186.695 93.570 186.925 ;
        RECT 93.675 186.695 97.150 187.605 ;
        RECT 97.355 186.695 99.965 187.605 ;
        RECT 100.125 186.735 100.555 187.520 ;
        RECT 100.805 186.925 104.705 187.605 ;
        RECT 103.775 186.695 104.705 186.925 ;
        RECT 104.810 186.925 108.275 187.605 ;
        RECT 104.810 186.695 105.730 186.925 ;
        RECT 108.590 186.695 112.065 187.605 ;
        RECT 112.075 186.795 113.445 187.605 ;
      LAYER nwell ;
        RECT 26.780 183.575 113.640 186.405 ;
      LAYER pwell ;
        RECT 26.975 182.375 28.345 183.185 ;
        RECT 28.825 182.375 30.175 183.285 ;
        RECT 30.205 182.375 31.555 183.285 ;
        RECT 31.575 183.055 32.505 183.285 ;
        RECT 31.575 182.375 35.475 183.055 ;
        RECT 35.725 182.460 36.155 183.245 ;
        RECT 36.635 183.055 37.565 183.285 ;
        RECT 41.235 183.055 42.165 183.285 ;
        RECT 45.375 183.055 46.295 183.285 ;
        RECT 49.125 183.055 50.055 183.275 ;
        RECT 60.535 183.055 61.465 183.285 ;
        RECT 36.635 182.375 40.535 183.055 ;
        RECT 41.235 182.375 45.135 183.055 ;
        RECT 45.375 182.375 54.565 183.055 ;
        RECT 54.585 182.375 57.325 183.055 ;
        RECT 57.565 182.375 61.465 183.055 ;
        RECT 61.485 182.460 61.915 183.245 ;
        RECT 62.030 183.055 62.950 183.285 ;
        RECT 65.710 183.055 66.630 183.285 ;
        RECT 62.030 182.375 65.495 183.055 ;
        RECT 65.710 182.375 69.175 183.055 ;
        RECT 70.410 182.375 73.885 183.285 ;
        RECT 73.895 182.375 77.370 183.285 ;
        RECT 77.575 182.375 81.050 183.285 ;
        RECT 81.810 182.375 85.680 183.285 ;
        RECT 85.865 182.375 87.215 183.285 ;
        RECT 87.245 182.460 87.675 183.245 ;
        RECT 88.810 182.375 92.285 183.285 ;
        RECT 94.950 183.055 95.870 183.285 ;
        RECT 92.405 182.375 95.870 183.055 ;
        RECT 95.985 182.375 97.335 183.285 ;
        RECT 97.365 182.375 98.715 183.285 ;
        RECT 101.850 183.055 102.770 183.285 ;
        RECT 105.530 183.055 106.450 183.285 ;
        RECT 109.210 183.055 110.130 183.285 ;
        RECT 99.305 182.375 102.770 183.055 ;
        RECT 102.985 182.375 106.450 183.055 ;
        RECT 106.665 182.375 110.130 183.055 ;
        RECT 110.695 182.375 112.065 183.155 ;
        RECT 112.075 182.375 113.445 183.185 ;
        RECT 27.115 182.165 27.285 182.375 ;
        RECT 28.550 182.215 28.670 182.325 ;
        RECT 28.955 182.210 29.115 182.320 ;
        RECT 29.875 182.185 30.045 182.375 ;
        RECT 30.335 182.165 30.505 182.375 ;
        RECT 31.990 182.185 32.160 182.375 ;
        RECT 36.370 182.215 36.490 182.325 ;
        RECT 37.050 182.185 37.220 182.375 ;
        RECT 39.535 182.165 39.705 182.355 ;
        RECT 39.995 182.165 40.165 182.355 ;
        RECT 40.970 182.215 41.090 182.325 ;
        RECT 41.375 182.165 41.545 182.355 ;
        RECT 41.650 182.185 41.820 182.375 ;
        RECT 45.060 182.165 45.230 182.355 ;
        RECT 49.195 182.165 49.365 182.355 ;
        RECT 54.255 182.185 54.425 182.375 ;
        RECT 57.015 182.185 57.185 182.375 ;
        RECT 60.880 182.185 61.050 182.375 ;
        RECT 65.295 182.185 65.465 182.375 ;
        RECT 67.135 182.165 67.305 182.355 ;
        RECT 67.650 182.215 67.770 182.325 ;
        RECT 68.055 182.165 68.225 182.355 ;
        RECT 68.975 182.185 69.145 182.375 ;
        RECT 69.895 182.220 70.055 182.330 ;
        RECT 70.815 182.185 70.985 182.355 ;
        RECT 73.570 182.185 73.740 182.375 ;
        RECT 74.040 182.185 74.210 182.375 ;
        RECT 70.915 182.165 70.985 182.185 ;
        RECT 74.955 182.165 75.125 182.355 ;
        RECT 76.850 182.215 76.970 182.325 ;
        RECT 77.720 182.185 77.890 182.375 ;
        RECT 85.535 182.355 85.680 182.375 ;
        RECT 80.660 182.165 80.830 182.355 ;
        RECT 81.400 182.165 81.570 182.355 ;
        RECT 85.075 182.165 85.245 182.355 ;
        RECT 85.535 182.185 85.705 182.355 ;
        RECT 85.995 182.185 86.165 182.375 ;
        RECT 88.295 182.220 88.455 182.330 ;
        RECT 91.970 182.185 92.140 182.375 ;
        RECT 92.435 182.185 92.605 182.375 ;
        RECT 95.655 182.165 95.825 182.355 ;
        RECT 96.390 182.165 96.560 182.355 ;
        RECT 97.035 182.185 97.205 182.375 ;
        RECT 98.415 182.185 98.585 182.375 ;
        RECT 98.930 182.215 99.050 182.325 ;
        RECT 99.335 182.185 99.505 182.375 ;
        RECT 102.095 182.165 102.265 182.355 ;
        RECT 102.555 182.165 102.725 182.355 ;
        RECT 103.015 182.185 103.185 182.375 ;
        RECT 106.695 182.185 106.865 182.375 ;
        RECT 111.755 182.325 111.925 182.375 ;
        RECT 110.430 182.215 110.550 182.325 ;
        RECT 111.755 182.215 111.930 182.325 ;
        RECT 111.755 182.185 111.925 182.215 ;
        RECT 113.135 182.165 113.305 182.375 ;
        RECT 26.975 181.355 28.345 182.165 ;
        RECT 29.285 181.255 30.635 182.165 ;
        RECT 30.655 181.485 39.845 182.165 ;
        RECT 30.655 181.255 31.575 181.485 ;
        RECT 34.405 181.265 35.335 181.485 ;
        RECT 39.865 181.255 41.215 182.165 ;
        RECT 41.345 181.485 44.810 182.165 ;
        RECT 43.890 181.255 44.810 181.485 ;
        RECT 44.915 181.255 48.390 182.165 ;
        RECT 48.605 181.295 49.035 182.080 ;
        RECT 49.055 181.485 58.160 182.165 ;
        RECT 58.255 181.485 67.445 182.165 ;
        RECT 58.255 181.255 59.175 181.485 ;
        RECT 62.005 181.265 62.935 181.485 ;
        RECT 67.915 181.255 70.635 182.165 ;
        RECT 70.915 181.935 73.185 182.165 ;
        RECT 70.915 181.255 73.670 181.935 ;
        RECT 74.365 181.295 74.795 182.080 ;
        RECT 74.815 181.485 76.645 182.165 ;
        RECT 77.345 181.485 81.245 182.165 ;
        RECT 75.300 181.255 76.645 181.485 ;
        RECT 80.315 181.255 81.245 181.485 ;
        RECT 81.255 181.255 84.730 182.165 ;
        RECT 84.935 181.485 94.125 182.165 ;
        RECT 89.445 181.265 90.375 181.485 ;
        RECT 93.205 181.255 94.125 181.485 ;
        RECT 94.135 181.485 95.965 182.165 ;
        RECT 95.975 181.485 99.875 182.165 ;
        RECT 94.135 181.255 95.480 181.485 ;
        RECT 95.975 181.255 96.905 181.485 ;
        RECT 100.125 181.295 100.555 182.080 ;
        RECT 100.575 181.485 102.405 182.165 ;
        RECT 102.415 181.485 111.605 182.165 ;
        RECT 106.925 181.265 107.855 181.485 ;
        RECT 110.685 181.255 111.605 181.485 ;
        RECT 112.075 181.355 113.445 182.165 ;
      LAYER nwell ;
        RECT 26.780 178.135 113.640 180.965 ;
      LAYER pwell ;
        RECT 26.975 176.935 28.345 177.745 ;
        RECT 28.815 176.935 30.185 177.715 ;
        RECT 30.205 176.935 31.555 177.845 ;
        RECT 31.575 177.615 32.505 177.845 ;
        RECT 31.575 176.935 35.475 177.615 ;
        RECT 35.725 177.020 36.155 177.805 ;
        RECT 36.635 176.935 38.005 177.715 ;
        RECT 38.025 176.935 39.375 177.845 ;
        RECT 39.590 176.935 43.065 177.845 ;
        RECT 43.270 176.935 46.745 177.845 ;
        RECT 46.850 177.615 47.770 177.845 ;
        RECT 51.355 177.615 52.700 177.845 ;
        RECT 46.850 176.935 50.315 177.615 ;
        RECT 51.355 176.935 53.185 177.615 ;
        RECT 53.290 176.935 57.160 177.845 ;
        RECT 57.795 176.935 61.270 177.845 ;
        RECT 61.485 177.020 61.915 177.805 ;
        RECT 61.935 176.935 65.410 177.845 ;
        RECT 65.615 176.935 69.090 177.845 ;
        RECT 69.295 177.615 70.640 177.845 ;
        RECT 73.895 177.615 75.240 177.845 ;
        RECT 69.295 176.935 71.125 177.615 ;
        RECT 71.135 176.935 73.875 177.615 ;
        RECT 73.895 176.935 75.725 177.615 ;
        RECT 76.740 176.935 85.845 177.615 ;
        RECT 85.865 176.935 87.215 177.845 ;
        RECT 87.245 177.020 87.675 177.805 ;
        RECT 95.425 177.615 96.355 177.835 ;
        RECT 99.185 177.615 100.105 177.845 ;
        RECT 100.600 177.615 101.945 177.845 ;
        RECT 88.075 176.935 90.500 177.615 ;
        RECT 90.915 176.935 100.105 177.615 ;
        RECT 100.115 176.935 101.945 177.615 ;
        RECT 102.415 177.615 103.335 177.845 ;
        RECT 106.165 177.615 107.095 177.835 ;
        RECT 102.415 176.935 111.605 177.615 ;
        RECT 112.075 176.935 113.445 177.745 ;
        RECT 27.115 176.725 27.285 176.935 ;
        RECT 28.495 176.885 28.665 176.915 ;
        RECT 28.495 176.775 28.670 176.885 ;
        RECT 28.495 176.725 28.665 176.775 ;
        RECT 28.955 176.745 29.125 176.935 ;
        RECT 30.335 176.745 30.505 176.935 ;
        RECT 31.990 176.745 32.160 176.935 ;
        RECT 36.370 176.775 36.490 176.885 ;
        RECT 36.775 176.745 36.945 176.935 ;
        RECT 38.155 176.725 38.325 176.935 ;
        RECT 42.750 176.745 42.920 176.935 ;
        RECT 46.430 176.745 46.600 176.935 ;
        RECT 47.355 176.725 47.525 176.915 ;
        RECT 49.195 176.725 49.365 176.915 ;
        RECT 50.115 176.745 50.285 176.935 ;
        RECT 51.035 176.780 51.195 176.890 ;
        RECT 52.875 176.725 53.045 176.935 ;
        RECT 57.015 176.915 57.160 176.935 ;
        RECT 56.610 176.775 56.730 176.885 ;
        RECT 57.015 176.745 57.185 176.915 ;
        RECT 57.530 176.775 57.650 176.885 ;
        RECT 57.940 176.745 58.110 176.935 ;
        RECT 62.080 176.745 62.250 176.935 ;
        RECT 65.760 176.915 65.930 176.935 ;
        RECT 65.755 176.745 65.930 176.915 ;
        RECT 65.755 176.725 65.925 176.745 ;
        RECT 68.515 176.725 68.685 176.915 ;
        RECT 68.975 176.725 69.145 176.915 ;
        RECT 70.815 176.745 70.985 176.935 ;
        RECT 71.275 176.745 71.445 176.935 ;
        RECT 73.115 176.725 73.285 176.915 ;
        RECT 74.035 176.770 74.195 176.880 ;
        RECT 74.955 176.725 75.125 176.915 ;
        RECT 75.415 176.745 75.585 176.935 ;
        RECT 76.335 176.780 76.495 176.890 ;
        RECT 85.535 176.725 85.705 176.935 ;
        RECT 85.995 176.725 86.165 176.915 ;
        RECT 86.915 176.745 87.085 176.935 ;
        RECT 90.595 176.745 90.765 176.915 ;
        RECT 91.055 176.745 91.225 176.935 ;
        RECT 98.600 176.725 98.770 176.915 ;
        RECT 99.795 176.770 99.955 176.880 ;
        RECT 100.255 176.745 100.425 176.935 ;
        RECT 100.770 176.775 100.890 176.885 ;
        RECT 102.150 176.775 102.270 176.885 ;
        RECT 104.580 176.725 104.750 176.915 ;
        RECT 108.720 176.725 108.890 176.915 ;
        RECT 109.460 176.725 109.630 176.915 ;
        RECT 111.295 176.745 111.465 176.935 ;
        RECT 111.810 176.775 111.930 176.885 ;
        RECT 113.135 176.725 113.305 176.935 ;
        RECT 26.975 175.915 28.345 176.725 ;
        RECT 28.355 176.045 37.635 176.725 ;
        RECT 38.015 176.045 47.205 176.725 ;
        RECT 29.715 175.825 30.635 176.045 ;
        RECT 35.300 175.925 37.635 176.045 ;
        RECT 36.715 175.815 37.635 175.925 ;
        RECT 42.525 175.825 43.455 176.045 ;
        RECT 46.285 175.815 47.205 176.045 ;
        RECT 47.225 175.815 48.575 176.725 ;
        RECT 48.605 175.855 49.035 176.640 ;
        RECT 49.165 176.045 52.630 176.725 ;
        RECT 52.845 176.045 56.310 176.725 ;
        RECT 51.710 175.815 52.630 176.045 ;
        RECT 55.390 175.815 56.310 176.045 ;
        RECT 56.875 176.045 66.065 176.725 ;
        RECT 66.085 176.045 68.825 176.725 ;
        RECT 68.835 176.045 70.665 176.725 ;
        RECT 56.875 175.815 57.795 176.045 ;
        RECT 60.625 175.825 61.555 176.045 ;
        RECT 69.320 175.815 70.665 176.045 ;
        RECT 70.705 175.815 73.425 176.725 ;
        RECT 74.365 175.855 74.795 176.640 ;
        RECT 74.825 175.815 76.175 176.725 ;
        RECT 76.565 176.045 85.845 176.725 ;
        RECT 85.855 176.045 94.960 176.725 ;
        RECT 95.285 176.045 99.185 176.725 ;
        RECT 76.565 175.925 78.900 176.045 ;
        RECT 76.565 175.815 77.485 175.925 ;
        RECT 83.565 175.825 84.485 176.045 ;
        RECT 98.255 175.815 99.185 176.045 ;
        RECT 100.125 175.855 100.555 176.640 ;
        RECT 101.265 176.045 105.165 176.725 ;
        RECT 105.405 176.045 109.305 176.725 ;
        RECT 104.235 175.815 105.165 176.045 ;
        RECT 108.375 175.815 109.305 176.045 ;
        RECT 109.315 175.815 111.925 176.725 ;
        RECT 112.075 175.915 113.445 176.725 ;
      LAYER nwell ;
        RECT 26.780 172.695 113.640 175.525 ;
      LAYER pwell ;
        RECT 29.495 172.315 30.445 172.405 ;
        RECT 26.975 171.495 28.345 172.305 ;
        RECT 28.515 171.495 30.445 172.315 ;
        RECT 31.575 172.175 32.505 172.405 ;
        RECT 31.575 171.495 35.475 172.175 ;
        RECT 35.725 171.580 36.155 172.365 ;
        RECT 36.270 171.495 40.140 172.405 ;
        RECT 44.825 172.175 45.755 172.395 ;
        RECT 48.585 172.175 49.505 172.405 ;
        RECT 54.025 172.175 54.955 172.395 ;
        RECT 57.785 172.175 58.705 172.405 ;
        RECT 40.315 171.495 49.505 172.175 ;
        RECT 49.515 171.495 58.705 172.175 ;
        RECT 58.855 171.495 61.465 172.405 ;
        RECT 61.485 171.580 61.915 172.365 ;
        RECT 61.935 172.175 62.855 172.405 ;
        RECT 65.685 172.175 66.615 172.395 ;
        RECT 75.185 172.295 76.105 172.405 ;
        RECT 75.185 172.175 77.520 172.295 ;
        RECT 82.185 172.175 83.105 172.395 ;
        RECT 84.960 172.175 86.305 172.405 ;
        RECT 61.935 171.495 71.125 172.175 ;
        RECT 71.145 171.495 73.885 172.175 ;
        RECT 75.185 171.495 84.465 172.175 ;
        RECT 84.475 171.495 86.305 172.175 ;
        RECT 87.245 171.580 87.675 172.365 ;
        RECT 88.065 172.295 88.985 172.405 ;
        RECT 88.065 172.175 90.400 172.295 ;
        RECT 95.065 172.175 95.985 172.395 ;
        RECT 100.555 172.175 101.485 172.405 ;
        RECT 88.065 171.495 97.345 172.175 ;
        RECT 97.585 171.495 101.485 172.175 ;
        RECT 101.495 172.175 102.415 172.405 ;
        RECT 105.245 172.175 106.175 172.395 ;
        RECT 101.495 171.495 110.685 172.175 ;
        RECT 110.705 171.495 112.055 172.405 ;
        RECT 112.075 171.495 113.445 172.305 ;
        RECT 27.115 171.285 27.285 171.495 ;
        RECT 28.515 171.475 28.665 171.495 ;
        RECT 28.495 171.285 28.665 171.475 ;
        RECT 31.255 171.340 31.415 171.450 ;
        RECT 31.990 171.305 32.160 171.495 ;
        RECT 39.995 171.475 40.140 171.495 ;
        RECT 39.995 171.305 40.165 171.475 ;
        RECT 40.455 171.305 40.625 171.495 ;
        RECT 46.895 171.285 47.065 171.475 ;
        RECT 47.355 171.285 47.525 171.475 ;
        RECT 49.470 171.285 49.640 171.475 ;
        RECT 49.655 171.305 49.825 171.495 ;
        RECT 53.610 171.285 53.780 171.475 ;
        RECT 57.750 171.285 57.920 171.475 ;
        RECT 61.150 171.305 61.320 171.495 ;
        RECT 65.020 171.285 65.190 171.475 ;
        RECT 68.975 171.285 69.145 171.475 ;
        RECT 70.815 171.305 70.985 171.495 ;
        RECT 71.730 171.285 71.900 171.475 ;
        RECT 73.575 171.285 73.745 171.495 ;
        RECT 74.090 171.335 74.210 171.445 ;
        RECT 74.495 171.340 74.655 171.450 ;
        RECT 75.875 171.285 76.045 171.475 ;
        RECT 79.740 171.285 79.910 171.475 ;
        RECT 81.395 171.285 81.565 171.475 ;
        RECT 84.155 171.305 84.325 171.495 ;
        RECT 84.615 171.305 84.785 171.495 ;
        RECT 86.915 171.340 87.075 171.450 ;
        RECT 91.055 171.285 91.225 171.475 ;
        RECT 94.920 171.285 95.090 171.475 ;
        RECT 96.115 171.330 96.275 171.440 ;
        RECT 96.580 171.285 96.750 171.475 ;
        RECT 97.035 171.305 97.205 171.495 ;
        RECT 100.720 171.285 100.890 171.475 ;
        RECT 100.900 171.305 101.070 171.495 ;
        RECT 107.615 171.285 107.785 171.475 ;
        RECT 110.375 171.305 110.545 171.495 ;
        RECT 111.290 171.285 111.460 171.475 ;
        RECT 111.755 171.445 111.925 171.495 ;
        RECT 111.755 171.335 111.930 171.445 ;
        RECT 111.755 171.305 111.925 171.335 ;
        RECT 113.135 171.285 113.305 171.495 ;
        RECT 26.975 170.475 28.345 171.285 ;
        RECT 28.355 170.605 37.635 171.285 ;
        RECT 38.100 170.605 47.205 171.285 ;
        RECT 29.715 170.385 30.635 170.605 ;
        RECT 35.300 170.485 37.635 170.605 ;
        RECT 47.215 170.505 48.585 171.285 ;
        RECT 36.715 170.375 37.635 170.485 ;
        RECT 48.605 170.415 49.035 171.200 ;
        RECT 49.055 170.605 52.955 171.285 ;
        RECT 53.195 170.605 57.095 171.285 ;
        RECT 57.335 170.605 61.235 171.285 ;
        RECT 61.705 170.605 65.605 171.285 ;
        RECT 49.055 170.375 49.985 170.605 ;
        RECT 53.195 170.375 54.125 170.605 ;
        RECT 57.335 170.375 58.265 170.605 ;
        RECT 64.675 170.375 65.605 170.605 ;
        RECT 65.710 170.605 69.175 171.285 ;
        RECT 65.710 170.375 66.630 170.605 ;
        RECT 69.435 170.375 72.045 171.285 ;
        RECT 72.055 170.605 73.885 171.285 ;
        RECT 72.055 170.375 73.400 170.605 ;
        RECT 74.365 170.415 74.795 171.200 ;
        RECT 74.815 170.505 76.185 171.285 ;
        RECT 76.425 170.605 80.325 171.285 ;
        RECT 79.395 170.375 80.325 170.605 ;
        RECT 80.345 170.375 81.695 171.285 ;
        RECT 82.085 170.605 91.365 171.285 ;
        RECT 91.605 170.605 95.505 171.285 ;
        RECT 82.085 170.485 84.420 170.605 ;
        RECT 82.085 170.375 83.005 170.485 ;
        RECT 89.085 170.385 90.005 170.605 ;
        RECT 94.575 170.375 95.505 170.605 ;
        RECT 96.435 170.375 99.910 171.285 ;
        RECT 100.125 170.415 100.555 171.200 ;
        RECT 100.575 170.375 104.050 171.285 ;
        RECT 104.350 170.605 107.815 171.285 ;
        RECT 104.350 170.375 105.270 170.605 ;
        RECT 108.130 170.375 111.605 171.285 ;
        RECT 112.075 170.475 113.445 171.285 ;
      LAYER nwell ;
        RECT 26.780 167.255 113.640 170.085 ;
      LAYER pwell ;
        RECT 30.415 166.875 31.365 166.965 ;
        RECT 26.975 166.055 28.345 166.865 ;
        RECT 29.435 166.055 31.365 166.875 ;
        RECT 31.575 166.735 32.505 166.965 ;
        RECT 31.575 166.055 35.475 166.735 ;
        RECT 35.725 166.140 36.155 166.925 ;
        RECT 36.635 166.055 38.005 166.835 ;
        RECT 38.210 166.055 41.685 166.965 ;
        RECT 42.065 166.855 42.985 166.965 ;
        RECT 42.065 166.735 44.400 166.855 ;
        RECT 49.065 166.735 49.985 166.955 ;
        RECT 51.355 166.735 52.285 166.965 ;
        RECT 42.065 166.055 51.345 166.735 ;
        RECT 51.355 166.055 55.255 166.735 ;
        RECT 56.415 166.055 57.785 166.835 ;
        RECT 57.795 166.055 61.270 166.965 ;
        RECT 61.485 166.140 61.915 166.925 ;
        RECT 61.935 166.055 65.410 166.965 ;
        RECT 66.075 166.055 68.685 166.965 ;
        RECT 69.030 166.055 72.505 166.965 ;
        RECT 72.515 166.055 75.990 166.965 ;
        RECT 76.565 166.855 77.485 166.965 ;
        RECT 76.565 166.735 78.900 166.855 ;
        RECT 83.565 166.735 84.485 166.955 ;
        RECT 76.565 166.055 85.845 166.735 ;
        RECT 85.855 166.055 87.225 166.835 ;
        RECT 87.245 166.140 87.675 166.925 ;
        RECT 90.895 166.735 91.825 166.965 ;
        RECT 87.925 166.055 91.825 166.735 ;
        RECT 91.930 166.735 92.850 166.965 ;
        RECT 91.930 166.055 95.395 166.735 ;
        RECT 95.515 166.055 98.990 166.965 ;
        RECT 99.655 166.055 102.265 166.965 ;
        RECT 102.415 166.735 103.335 166.965 ;
        RECT 106.165 166.735 107.095 166.955 ;
        RECT 102.415 166.055 111.605 166.735 ;
        RECT 112.075 166.055 113.445 166.865 ;
        RECT 27.115 165.845 27.285 166.055 ;
        RECT 29.435 166.035 29.585 166.055 ;
        RECT 28.955 165.900 29.115 166.010 ;
        RECT 29.415 165.865 29.585 166.035 ;
        RECT 31.990 165.865 32.160 166.055 ;
        RECT 36.370 165.895 36.490 166.005 ;
        RECT 36.775 165.865 36.945 166.055 ;
        RECT 37.695 165.845 37.865 166.035 ;
        RECT 39.075 165.845 39.245 166.035 ;
        RECT 39.995 165.890 40.155 166.000 ;
        RECT 40.730 165.845 40.900 166.035 ;
        RECT 41.370 165.865 41.540 166.055 ;
        RECT 44.650 165.895 44.770 166.005 ;
        RECT 45.055 165.845 45.225 166.035 ;
        RECT 49.195 165.865 49.365 166.035 ;
        RECT 51.035 165.865 51.205 166.055 ;
        RECT 49.215 165.845 49.365 165.865 ;
        RECT 51.500 165.845 51.670 166.035 ;
        RECT 51.770 165.865 51.940 166.055 ;
        RECT 56.095 165.900 56.255 166.010 ;
        RECT 56.555 165.865 56.725 166.055 ;
        RECT 57.940 165.865 58.110 166.055 ;
        RECT 58.390 165.845 58.560 166.035 ;
        RECT 58.910 165.895 59.030 166.005 ;
        RECT 62.080 165.865 62.250 166.055 ;
        RECT 65.810 165.895 65.930 166.005 ;
        RECT 66.220 165.865 66.390 166.055 ;
        RECT 68.515 165.845 68.685 166.035 ;
        RECT 70.355 165.845 70.525 166.035 ;
        RECT 70.820 165.845 70.990 166.035 ;
        RECT 72.190 165.865 72.360 166.055 ;
        RECT 72.660 165.865 72.830 166.055 ;
        RECT 76.335 165.845 76.505 166.035 ;
        RECT 77.715 165.845 77.885 166.035 ;
        RECT 81.580 165.845 81.750 166.035 ;
        RECT 82.315 165.845 82.485 166.035 ;
        RECT 84.155 165.890 84.315 166.000 ;
        RECT 84.615 165.845 84.785 166.035 ;
        RECT 85.535 165.865 85.705 166.055 ;
        RECT 85.995 165.845 86.165 166.035 ;
        RECT 86.915 165.865 87.085 166.055 ;
        RECT 26.975 165.035 28.345 165.845 ;
        RECT 28.725 165.165 38.005 165.845 ;
        RECT 28.725 165.045 31.060 165.165 ;
        RECT 28.725 164.935 29.645 165.045 ;
        RECT 35.725 164.945 36.645 165.165 ;
        RECT 38.015 165.065 39.385 165.845 ;
        RECT 40.315 165.165 44.215 165.845 ;
        RECT 45.025 165.165 48.490 165.845 ;
        RECT 40.315 164.935 41.245 165.165 ;
        RECT 47.570 164.935 48.490 165.165 ;
        RECT 48.605 164.975 49.035 165.760 ;
        RECT 49.215 165.025 51.145 165.845 ;
        RECT 50.195 164.935 51.145 165.025 ;
        RECT 51.355 164.935 54.830 165.845 ;
        RECT 55.230 164.935 58.705 165.845 ;
        RECT 59.545 165.165 68.825 165.845 ;
        RECT 68.835 165.165 70.665 165.845 ;
        RECT 59.545 165.045 61.880 165.165 ;
        RECT 59.545 164.935 60.465 165.045 ;
        RECT 66.545 164.945 67.465 165.165 ;
        RECT 68.835 164.935 70.180 165.165 ;
        RECT 70.675 164.935 74.150 165.845 ;
        RECT 74.365 164.975 74.795 165.760 ;
        RECT 74.815 165.165 76.645 165.845 ;
        RECT 74.815 164.935 76.160 165.165 ;
        RECT 76.665 164.935 78.015 165.845 ;
        RECT 78.265 165.165 82.165 165.845 ;
        RECT 81.235 164.935 82.165 165.165 ;
        RECT 82.175 165.065 83.545 165.845 ;
        RECT 84.485 164.935 85.835 165.845 ;
        RECT 85.855 165.065 87.225 165.845 ;
        RECT 87.235 165.815 88.180 165.845 ;
        RECT 89.670 165.815 89.840 166.035 ;
        RECT 90.140 165.845 90.310 166.035 ;
        RECT 91.240 165.865 91.410 166.055 ;
        RECT 93.820 165.845 93.990 166.035 ;
        RECT 95.195 165.865 95.365 166.055 ;
        RECT 95.660 165.865 95.830 166.055 ;
        RECT 99.800 166.035 99.970 166.055 ;
        RECT 99.390 165.895 99.510 166.005 ;
        RECT 99.790 165.865 99.970 166.035 ;
        RECT 87.235 165.135 89.985 165.815 ;
        RECT 87.235 164.935 88.180 165.135 ;
        RECT 89.995 164.935 93.470 165.845 ;
        RECT 93.675 164.935 97.150 165.845 ;
        RECT 97.355 165.815 98.300 165.845 ;
        RECT 99.790 165.815 99.960 165.865 ;
        RECT 101.635 165.845 101.805 166.035 ;
        RECT 102.150 165.895 102.270 166.005 ;
        RECT 111.295 165.865 111.465 166.055 ;
        RECT 111.755 166.005 111.925 166.035 ;
        RECT 111.755 165.895 111.930 166.005 ;
        RECT 111.755 165.845 111.925 165.895 ;
        RECT 113.135 165.845 113.305 166.055 ;
        RECT 97.355 165.135 100.105 165.815 ;
        RECT 97.355 164.935 98.300 165.135 ;
        RECT 100.125 164.975 100.555 165.760 ;
        RECT 100.575 165.065 101.945 165.845 ;
        RECT 102.785 165.165 112.065 165.845 ;
        RECT 102.785 165.045 105.120 165.165 ;
        RECT 102.785 164.935 103.705 165.045 ;
        RECT 109.785 164.945 110.705 165.165 ;
        RECT 112.075 165.035 113.445 165.845 ;
      LAYER nwell ;
        RECT 26.780 161.815 113.640 164.645 ;
      LAYER pwell ;
        RECT 30.415 161.435 31.365 161.525 ;
        RECT 26.975 160.615 28.345 161.425 ;
        RECT 29.435 160.615 31.365 161.435 ;
        RECT 34.775 161.295 35.705 161.525 ;
        RECT 31.805 160.615 35.705 161.295 ;
        RECT 35.725 160.700 36.155 161.485 ;
        RECT 37.535 161.295 38.455 161.515 ;
        RECT 44.535 161.415 45.455 161.525 ;
        RECT 43.120 161.295 45.455 161.415 ;
        RECT 36.175 160.615 45.455 161.295 ;
        RECT 45.835 160.615 49.310 161.525 ;
        RECT 49.975 160.615 53.450 161.525 ;
        RECT 53.665 160.615 55.015 161.525 ;
        RECT 55.965 160.615 57.315 161.525 ;
        RECT 57.335 160.615 60.810 161.525 ;
        RECT 61.485 160.700 61.915 161.485 ;
        RECT 62.020 160.615 71.125 161.295 ;
        RECT 72.055 160.615 74.775 161.525 ;
        RECT 74.815 160.615 78.290 161.525 ;
        RECT 78.965 160.615 80.315 161.525 ;
        RECT 80.345 160.615 81.695 161.525 ;
        RECT 81.725 160.615 83.075 161.525 ;
        RECT 86.295 161.295 87.225 161.525 ;
        RECT 83.325 160.615 87.225 161.295 ;
        RECT 87.245 160.700 87.675 161.485 ;
        RECT 87.705 160.615 89.055 161.525 ;
        RECT 92.650 161.295 93.570 161.525 ;
        RECT 90.105 160.615 93.570 161.295 ;
        RECT 93.675 160.615 97.150 161.525 ;
        RECT 98.010 160.615 101.485 161.525 ;
        RECT 104.695 161.295 105.625 161.525 ;
        RECT 108.835 161.295 109.765 161.525 ;
        RECT 101.725 160.615 105.625 161.295 ;
        RECT 105.865 160.615 109.765 161.295 ;
        RECT 109.775 160.615 111.145 161.395 ;
        RECT 112.075 160.615 113.445 161.425 ;
        RECT 27.115 160.405 27.285 160.615 ;
        RECT 29.435 160.595 29.585 160.615 ;
        RECT 28.955 160.460 29.115 160.570 ;
        RECT 29.415 160.425 29.585 160.595 ;
        RECT 26.975 159.595 28.345 160.405 ;
        RECT 28.355 160.375 29.300 160.405 ;
        RECT 30.790 160.375 30.960 160.595 ;
        RECT 31.115 160.375 32.060 160.405 ;
        RECT 33.550 160.375 33.720 160.595 ;
        RECT 35.120 160.425 35.290 160.615 ;
        RECT 36.315 160.425 36.485 160.615 ;
        RECT 37.235 160.405 37.405 160.595 ;
        RECT 37.700 160.405 37.870 160.595 ;
        RECT 41.380 160.405 41.550 160.595 ;
        RECT 45.060 160.405 45.230 160.595 ;
        RECT 45.980 160.425 46.150 160.615 ;
        RECT 49.195 160.405 49.365 160.595 ;
        RECT 49.710 160.455 49.830 160.565 ;
        RECT 50.120 160.425 50.290 160.615 ;
        RECT 53.795 160.425 53.965 160.615 ;
        RECT 55.635 160.460 55.795 160.570 ;
        RECT 56.095 160.425 56.265 160.615 ;
        RECT 57.480 160.425 57.650 160.615 ;
        RECT 61.210 160.455 61.330 160.565 ;
        RECT 62.260 160.405 62.430 160.595 ;
        RECT 63.455 160.450 63.615 160.560 ;
        RECT 63.915 160.405 64.085 160.595 ;
        RECT 66.675 160.405 66.845 160.595 ;
        RECT 69.435 160.405 69.605 160.595 ;
        RECT 69.895 160.405 70.065 160.595 ;
        RECT 70.815 160.425 70.985 160.615 ;
        RECT 71.735 160.405 71.905 160.595 ;
        RECT 72.195 160.425 72.365 160.615 ;
        RECT 74.960 160.425 75.130 160.615 ;
        RECT 75.875 160.405 76.045 160.595 ;
        RECT 76.335 160.405 76.505 160.595 ;
        RECT 78.690 160.455 78.810 160.565 ;
        RECT 79.095 160.425 79.265 160.615 ;
        RECT 81.395 160.425 81.565 160.615 ;
        RECT 81.855 160.425 82.025 160.615 ;
        RECT 86.640 160.425 86.810 160.615 ;
        RECT 86.915 160.405 87.085 160.595 ;
        RECT 87.375 160.405 87.545 160.595 ;
        RECT 87.835 160.425 88.005 160.615 ;
        RECT 89.675 160.460 89.835 160.570 ;
        RECT 90.135 160.425 90.305 160.615 ;
        RECT 93.820 160.425 93.990 160.615 ;
        RECT 101.170 160.595 101.340 160.615 ;
        RECT 96.580 160.405 96.750 160.595 ;
        RECT 97.550 160.455 97.670 160.565 ;
        RECT 100.770 160.455 100.890 160.565 ;
        RECT 101.170 160.425 101.345 160.595 ;
        RECT 102.610 160.455 102.730 160.565 ;
        RECT 105.040 160.425 105.210 160.615 ;
        RECT 101.175 160.405 101.345 160.425 ;
        RECT 106.420 160.405 106.590 160.595 ;
        RECT 107.155 160.405 107.325 160.595 ;
        RECT 109.180 160.425 109.350 160.615 ;
        RECT 109.915 160.425 110.085 160.615 ;
        RECT 111.755 160.405 111.925 160.595 ;
        RECT 113.135 160.405 113.305 160.615 ;
        RECT 28.355 159.695 31.105 160.375 ;
        RECT 31.115 159.695 33.865 160.375 ;
        RECT 33.970 159.725 37.435 160.405 ;
        RECT 28.355 159.495 29.300 159.695 ;
        RECT 31.115 159.495 32.060 159.695 ;
        RECT 33.970 159.495 34.890 159.725 ;
        RECT 37.555 159.495 41.030 160.405 ;
        RECT 41.235 159.495 44.710 160.405 ;
        RECT 44.915 159.495 48.390 160.405 ;
        RECT 48.605 159.535 49.035 160.320 ;
        RECT 49.055 159.725 58.335 160.405 ;
        RECT 58.945 159.725 62.845 160.405 ;
        RECT 50.415 159.505 51.335 159.725 ;
        RECT 56.000 159.605 58.335 159.725 ;
        RECT 57.415 159.495 58.335 159.605 ;
        RECT 61.915 159.495 62.845 159.725 ;
        RECT 63.775 159.625 65.145 160.405 ;
        RECT 65.155 159.725 66.985 160.405 ;
        RECT 67.005 159.725 69.745 160.405 ;
        RECT 69.755 159.725 71.585 160.405 ;
        RECT 71.595 159.725 74.335 160.405 ;
        RECT 65.155 159.495 66.500 159.725 ;
        RECT 70.240 159.495 71.585 159.725 ;
        RECT 74.365 159.535 74.795 160.320 ;
        RECT 74.815 159.625 76.185 160.405 ;
        RECT 76.195 159.625 77.565 160.405 ;
        RECT 77.945 159.725 87.225 160.405 ;
        RECT 87.235 159.725 96.425 160.405 ;
        RECT 77.945 159.605 80.280 159.725 ;
        RECT 77.945 159.495 78.865 159.605 ;
        RECT 84.945 159.505 85.865 159.725 ;
        RECT 91.745 159.505 92.675 159.725 ;
        RECT 95.505 159.495 96.425 159.725 ;
        RECT 96.435 159.495 99.910 160.405 ;
        RECT 100.125 159.535 100.555 160.320 ;
        RECT 101.045 159.495 102.395 160.405 ;
        RECT 103.105 159.725 107.005 160.405 ;
        RECT 107.125 159.725 110.590 160.405 ;
        RECT 106.075 159.495 107.005 159.725 ;
        RECT 109.670 159.495 110.590 159.725 ;
        RECT 110.705 159.495 112.055 160.405 ;
        RECT 112.075 159.595 113.445 160.405 ;
      LAYER nwell ;
        RECT 26.780 156.375 113.640 159.205 ;
      LAYER pwell ;
        RECT 29.495 155.995 30.445 156.085 ;
        RECT 26.975 155.175 28.345 155.985 ;
        RECT 28.515 155.175 30.445 155.995 ;
        RECT 30.655 155.855 31.585 156.085 ;
        RECT 30.655 155.175 34.555 155.855 ;
        RECT 35.725 155.260 36.155 156.045 ;
        RECT 36.175 155.885 37.120 156.085 ;
        RECT 38.935 155.885 39.880 156.085 ;
        RECT 41.695 155.885 42.640 156.085 ;
        RECT 36.175 155.205 38.925 155.885 ;
        RECT 38.935 155.205 41.685 155.885 ;
        RECT 41.695 155.205 44.445 155.885 ;
        RECT 36.175 155.175 37.120 155.205 ;
        RECT 27.115 154.965 27.285 155.175 ;
        RECT 28.515 155.155 28.665 155.175 ;
        RECT 28.495 154.985 28.665 155.155 ;
        RECT 31.070 154.985 31.240 155.175 ;
        RECT 35.395 155.020 35.555 155.130 ;
        RECT 37.695 154.965 37.865 155.155 ;
        RECT 38.610 154.985 38.780 155.205 ;
        RECT 38.935 155.175 39.880 155.205 ;
        RECT 40.455 154.965 40.625 155.155 ;
        RECT 41.190 154.965 41.360 155.155 ;
        RECT 41.370 154.985 41.540 155.205 ;
        RECT 41.695 155.175 42.640 155.205 ;
        RECT 44.130 154.985 44.300 155.205 ;
        RECT 44.455 155.175 47.930 156.085 ;
        RECT 48.135 155.175 51.610 156.085 ;
        RECT 51.815 155.175 53.185 155.955 ;
        RECT 53.195 155.855 54.125 156.085 ;
        RECT 53.195 155.175 57.095 155.855 ;
        RECT 58.255 155.175 61.465 156.085 ;
        RECT 61.485 155.260 61.915 156.045 ;
        RECT 65.595 155.855 66.525 156.085 ;
        RECT 62.625 155.175 66.525 155.855 ;
        RECT 66.545 155.175 67.895 156.085 ;
        RECT 69.320 155.855 70.665 156.085 ;
        RECT 71.160 155.855 72.505 156.085 ;
        RECT 68.835 155.175 70.665 155.855 ;
        RECT 70.675 155.175 72.505 155.855 ;
        RECT 72.975 155.885 73.920 156.085 ;
        RECT 72.975 155.205 75.725 155.885 ;
        RECT 72.975 155.175 73.920 155.205 ;
        RECT 44.600 154.985 44.770 155.175 ;
        RECT 45.515 155.010 45.675 155.120 ;
        RECT 26.975 154.155 28.345 154.965 ;
        RECT 28.725 154.285 38.005 154.965 ;
        RECT 38.025 154.285 40.765 154.965 ;
        RECT 40.775 154.285 44.675 154.965 ;
        RECT 45.980 154.935 46.150 155.155 ;
        RECT 48.280 154.985 48.450 155.175 ;
        RECT 51.035 154.985 51.205 155.155 ;
        RECT 52.875 154.985 53.045 155.175 ;
        RECT 53.610 154.985 53.780 155.175 ;
        RECT 57.935 155.020 58.095 155.130 ;
        RECT 58.395 154.985 58.565 155.175 ;
        RECT 51.035 154.965 51.185 154.985 ;
        RECT 60.695 154.965 60.865 155.155 ;
        RECT 61.615 155.010 61.775 155.120 ;
        RECT 62.130 155.015 62.250 155.125 ;
        RECT 65.940 154.985 66.110 155.175 ;
        RECT 67.595 154.985 67.765 155.175 ;
        RECT 68.515 155.020 68.675 155.130 ;
        RECT 68.975 154.985 69.145 155.175 ;
        RECT 70.815 154.965 70.985 155.175 ;
        RECT 71.330 155.015 71.450 155.125 ;
        RECT 72.710 155.015 72.830 155.125 ;
        RECT 47.640 154.935 48.585 154.965 ;
        RECT 28.725 154.165 31.060 154.285 ;
        RECT 28.725 154.055 29.645 154.165 ;
        RECT 35.725 154.065 36.645 154.285 ;
        RECT 40.775 154.055 41.705 154.285 ;
        RECT 45.835 154.255 48.585 154.935 ;
        RECT 47.640 154.055 48.585 154.255 ;
        RECT 48.605 154.095 49.035 154.880 ;
        RECT 49.255 154.145 51.185 154.965 ;
        RECT 51.725 154.285 61.005 154.965 ;
        RECT 61.935 154.285 71.125 154.965 ;
        RECT 71.595 154.935 72.540 154.965 ;
        RECT 74.030 154.935 74.200 155.155 ;
        RECT 74.960 154.965 75.130 155.155 ;
        RECT 75.410 154.985 75.580 155.205 ;
        RECT 75.735 155.175 79.210 156.085 ;
        RECT 82.615 155.855 83.545 156.085 ;
        RECT 79.645 155.175 83.545 155.855 ;
        RECT 83.650 155.855 84.570 156.085 ;
        RECT 83.650 155.175 87.115 155.855 ;
        RECT 87.245 155.260 87.675 156.045 ;
        RECT 88.155 155.885 89.100 156.085 ;
        RECT 92.720 155.885 93.665 156.085 ;
        RECT 88.155 155.205 90.905 155.885 ;
        RECT 90.915 155.205 93.665 155.885 ;
        RECT 88.155 155.175 89.100 155.205 ;
        RECT 75.880 154.985 76.050 155.175 ;
        RECT 82.960 154.985 83.130 155.175 ;
        RECT 86.915 154.985 87.085 155.175 ;
        RECT 87.835 155.125 88.005 155.155 ;
        RECT 87.835 155.015 88.010 155.125 ;
        RECT 87.835 154.965 88.005 155.015 ;
        RECT 89.215 154.965 89.385 155.155 ;
        RECT 51.725 154.165 54.060 154.285 ;
        RECT 49.255 154.055 50.205 154.145 ;
        RECT 51.725 154.055 52.645 154.165 ;
        RECT 58.725 154.065 59.645 154.285 ;
        RECT 61.935 154.055 62.855 154.285 ;
        RECT 65.685 154.065 66.615 154.285 ;
        RECT 71.595 154.255 74.345 154.935 ;
        RECT 71.595 154.055 72.540 154.255 ;
        RECT 74.365 154.095 74.795 154.880 ;
        RECT 74.815 154.055 78.290 154.965 ;
        RECT 78.865 154.285 88.145 154.965 ;
        RECT 78.865 154.165 81.200 154.285 ;
        RECT 78.865 154.055 79.785 154.165 ;
        RECT 85.865 154.065 86.785 154.285 ;
        RECT 88.155 154.185 89.525 154.965 ;
        RECT 89.680 154.935 89.850 155.155 ;
        RECT 90.590 154.985 90.760 155.205 ;
        RECT 91.060 154.985 91.230 155.205 ;
        RECT 92.720 155.175 93.665 155.205 ;
        RECT 93.675 155.175 97.150 156.085 ;
        RECT 97.355 155.175 100.830 156.085 ;
        RECT 101.045 155.175 102.395 156.085 ;
        RECT 102.785 155.975 103.705 156.085 ;
        RECT 102.785 155.855 105.120 155.975 ;
        RECT 109.785 155.855 110.705 156.075 ;
        RECT 102.785 155.175 112.065 155.855 ;
        RECT 112.075 155.175 113.445 155.985 ;
        RECT 92.440 154.965 92.610 155.155 ;
        RECT 93.820 154.985 93.990 155.175 ;
        RECT 97.500 154.985 97.670 155.175 ;
        RECT 99.520 154.965 99.690 155.155 ;
        RECT 100.770 155.015 100.890 155.125 ;
        RECT 101.175 154.965 101.345 155.175 ;
        RECT 111.755 154.965 111.925 155.175 ;
        RECT 113.135 154.965 113.305 155.175 ;
        RECT 91.340 154.935 92.285 154.965 ;
        RECT 89.535 154.255 92.285 154.935 ;
        RECT 91.340 154.055 92.285 154.255 ;
        RECT 92.295 154.055 95.770 154.965 ;
        RECT 96.205 154.285 100.105 154.965 ;
        RECT 99.175 154.055 100.105 154.285 ;
        RECT 100.125 154.095 100.555 154.880 ;
        RECT 101.035 154.185 102.405 154.965 ;
        RECT 102.785 154.285 112.065 154.965 ;
        RECT 102.785 154.165 105.120 154.285 ;
        RECT 102.785 154.055 103.705 154.165 ;
        RECT 109.785 154.065 110.705 154.285 ;
        RECT 112.075 154.155 113.445 154.965 ;
      LAYER nwell ;
        RECT 26.780 150.935 113.640 153.765 ;
      LAYER pwell ;
        RECT 30.415 150.555 31.365 150.645 ;
        RECT 26.975 149.735 28.345 150.545 ;
        RECT 29.435 149.735 31.365 150.555 ;
        RECT 31.575 150.415 32.505 150.645 ;
        RECT 31.575 149.735 35.475 150.415 ;
        RECT 35.725 149.820 36.155 150.605 ;
        RECT 37.535 150.415 38.455 150.635 ;
        RECT 44.535 150.535 45.455 150.645 ;
        RECT 43.120 150.415 45.455 150.535 ;
        RECT 36.175 149.735 45.455 150.415 ;
        RECT 45.845 149.735 47.195 150.645 ;
        RECT 49.480 150.445 50.425 150.645 ;
        RECT 47.675 149.765 50.425 150.445 ;
        RECT 53.090 150.415 54.010 150.645 ;
        RECT 27.115 149.525 27.285 149.735 ;
        RECT 29.435 149.715 29.585 149.735 ;
        RECT 28.955 149.580 29.115 149.690 ;
        RECT 29.415 149.545 29.585 149.715 ;
        RECT 31.990 149.545 32.160 149.735 ;
        RECT 36.315 149.545 36.485 149.735 ;
        RECT 37.695 149.525 37.865 149.715 ;
        RECT 45.975 149.545 46.145 149.735 ;
        RECT 46.895 149.525 47.065 149.715 ;
        RECT 47.355 149.685 47.525 149.715 ;
        RECT 47.355 149.575 47.530 149.685 ;
        RECT 47.355 149.525 47.525 149.575 ;
        RECT 47.820 149.545 47.990 149.765 ;
        RECT 49.480 149.735 50.425 149.765 ;
        RECT 50.545 149.735 54.010 150.415 ;
        RECT 54.115 149.735 57.590 150.645 ;
        RECT 60.450 150.415 61.370 150.645 ;
        RECT 57.905 149.735 61.370 150.415 ;
        RECT 61.485 149.820 61.915 150.605 ;
        RECT 63.225 150.535 64.145 150.645 ;
        RECT 63.225 150.415 65.560 150.535 ;
        RECT 70.225 150.415 71.145 150.635 ;
        RECT 63.225 149.735 72.505 150.415 ;
        RECT 72.525 149.735 73.875 150.645 ;
        RECT 73.895 149.735 75.265 150.515 ;
        RECT 75.275 149.735 78.025 150.545 ;
        RECT 78.035 149.735 79.405 150.515 ;
        RECT 79.415 150.415 80.345 150.645 ;
        RECT 79.415 149.735 83.315 150.415 ;
        RECT 83.565 149.735 84.915 150.645 ;
        RECT 84.935 149.735 86.305 150.515 ;
        RECT 87.245 149.820 87.675 150.605 ;
        RECT 89.755 150.555 90.705 150.645 ;
        RECT 88.775 149.735 90.705 150.555 ;
        RECT 94.115 150.415 95.045 150.645 ;
        RECT 91.145 149.735 95.045 150.415 ;
        RECT 95.055 150.445 96.000 150.645 ;
        RECT 98.015 150.555 98.965 150.645 ;
        RECT 95.055 149.765 97.805 150.445 ;
        RECT 95.055 149.735 96.000 149.765 ;
        RECT 49.250 149.575 49.370 149.685 ;
        RECT 26.975 148.715 28.345 149.525 ;
        RECT 28.725 148.845 38.005 149.525 ;
        RECT 38.100 148.845 47.205 149.525 ;
        RECT 28.725 148.725 31.060 148.845 ;
        RECT 28.725 148.615 29.645 148.725 ;
        RECT 35.725 148.625 36.645 148.845 ;
        RECT 47.215 148.745 48.585 149.525 ;
        RECT 49.660 149.495 49.830 149.715 ;
        RECT 50.575 149.545 50.745 149.735 ;
        RECT 52.420 149.525 52.590 149.715 ;
        RECT 54.260 149.545 54.430 149.735 ;
        RECT 56.100 149.525 56.270 149.715 ;
        RECT 57.935 149.545 58.105 149.735 ;
        RECT 59.830 149.575 59.950 149.685 ;
        RECT 60.240 149.525 60.410 149.715 ;
        RECT 62.535 149.580 62.695 149.690 ;
        RECT 67.320 149.525 67.490 149.715 ;
        RECT 69.435 149.525 69.605 149.715 ;
        RECT 69.895 149.525 70.065 149.715 ;
        RECT 72.195 149.545 72.365 149.735 ;
        RECT 72.655 149.545 72.825 149.735 ;
        RECT 51.320 149.495 52.265 149.525 ;
        RECT 48.605 148.655 49.035 149.440 ;
        RECT 49.515 148.815 52.265 149.495 ;
        RECT 51.320 148.615 52.265 148.815 ;
        RECT 52.275 148.615 55.750 149.525 ;
        RECT 55.955 148.615 59.430 149.525 ;
        RECT 60.095 148.615 63.570 149.525 ;
        RECT 64.005 148.845 67.905 149.525 ;
        RECT 67.915 148.845 69.745 149.525 ;
        RECT 69.755 148.845 71.585 149.525 ;
        RECT 71.595 149.495 72.540 149.525 ;
        RECT 74.030 149.495 74.200 149.715 ;
        RECT 74.955 149.685 75.125 149.735 ;
        RECT 74.955 149.575 75.130 149.685 ;
        RECT 74.955 149.545 75.125 149.575 ;
        RECT 75.420 149.525 75.590 149.715 ;
        RECT 77.715 149.545 77.885 149.735 ;
        RECT 78.175 149.545 78.345 149.735 ;
        RECT 79.830 149.545 80.000 149.735 ;
        RECT 84.615 149.545 84.785 149.735 ;
        RECT 85.075 149.545 85.245 149.735 ;
        RECT 88.775 149.715 88.925 149.735 ;
        RECT 86.915 149.580 87.075 149.690 ;
        RECT 88.295 149.525 88.465 149.715 ;
        RECT 88.755 149.545 88.925 149.715 ;
        RECT 94.460 149.545 94.630 149.735 ;
        RECT 97.490 149.545 97.660 149.765 ;
        RECT 98.015 149.735 99.945 150.555 ;
        RECT 100.125 149.735 101.475 150.645 ;
        RECT 104.695 150.415 105.625 150.645 ;
        RECT 101.725 149.735 105.625 150.415 ;
        RECT 106.555 149.735 107.925 150.515 ;
        RECT 108.395 149.735 109.765 150.515 ;
        RECT 109.775 149.735 111.145 150.515 ;
        RECT 112.075 149.735 113.445 150.545 ;
        RECT 99.795 149.715 99.945 149.735 ;
        RECT 97.955 149.525 98.125 149.715 ;
        RECT 98.415 149.525 98.585 149.715 ;
        RECT 99.795 149.685 99.965 149.715 ;
        RECT 99.795 149.575 99.970 149.685 ;
        RECT 99.795 149.545 99.965 149.575 ;
        RECT 100.255 149.545 100.425 149.735 ;
        RECT 100.770 149.575 100.890 149.685 ;
        RECT 105.040 149.545 105.210 149.735 ;
        RECT 106.235 149.580 106.395 149.690 ;
        RECT 106.695 149.545 106.865 149.735 ;
        RECT 108.130 149.575 108.250 149.685 ;
        RECT 108.535 149.545 108.705 149.735 ;
        RECT 109.915 149.545 110.085 149.735 ;
        RECT 110.375 149.525 110.545 149.715 ;
        RECT 110.835 149.525 111.005 149.715 ;
        RECT 111.755 149.580 111.915 149.690 ;
        RECT 113.135 149.525 113.305 149.735 ;
        RECT 66.975 148.615 67.905 148.845 ;
        RECT 71.595 148.815 74.345 149.495 ;
        RECT 71.595 148.615 72.540 148.815 ;
        RECT 74.365 148.655 74.795 149.440 ;
        RECT 75.275 148.615 78.750 149.525 ;
        RECT 79.325 148.845 88.605 149.525 ;
        RECT 88.985 148.845 98.265 149.525 ;
        RECT 79.325 148.725 81.660 148.845 ;
        RECT 79.325 148.615 80.245 148.725 ;
        RECT 86.325 148.625 87.245 148.845 ;
        RECT 88.985 148.725 91.320 148.845 ;
        RECT 88.985 148.615 89.905 148.725 ;
        RECT 95.985 148.625 96.905 148.845 ;
        RECT 98.285 148.615 99.635 149.525 ;
        RECT 100.125 148.655 100.555 149.440 ;
        RECT 101.405 148.845 110.685 149.525 ;
        RECT 101.405 148.725 103.740 148.845 ;
        RECT 101.405 148.615 102.325 148.725 ;
        RECT 108.405 148.625 109.325 148.845 ;
        RECT 110.705 148.615 112.055 149.525 ;
        RECT 112.075 148.715 113.445 149.525 ;
      LAYER nwell ;
        RECT 26.780 145.495 113.640 148.325 ;
      LAYER pwell ;
        RECT 30.415 145.115 31.365 145.205 ;
        RECT 26.975 144.295 28.345 145.105 ;
        RECT 29.435 144.295 31.365 145.115 ;
        RECT 31.575 144.975 32.505 145.205 ;
        RECT 31.575 144.295 35.475 144.975 ;
        RECT 35.725 144.380 36.155 145.165 ;
        RECT 39.375 144.975 40.305 145.205 ;
        RECT 36.405 144.295 40.305 144.975 ;
        RECT 40.685 145.095 41.605 145.205 ;
        RECT 40.685 144.975 43.020 145.095 ;
        RECT 47.685 144.975 48.605 145.195 ;
        RECT 53.175 144.975 54.105 145.205 ;
        RECT 40.685 144.295 49.965 144.975 ;
        RECT 50.205 144.295 54.105 144.975 ;
        RECT 54.310 144.295 57.785 145.205 ;
        RECT 57.795 144.295 61.270 145.205 ;
        RECT 61.485 144.380 61.915 145.165 ;
        RECT 62.865 144.295 64.215 145.205 ;
        RECT 67.435 144.975 68.365 145.205 ;
        RECT 69.975 145.115 70.925 145.205 ;
        RECT 64.465 144.295 68.365 144.975 ;
        RECT 68.995 144.295 70.925 145.115 ;
        RECT 73.895 145.005 74.840 145.205 ;
        RECT 71.135 144.295 73.875 144.975 ;
        RECT 73.895 144.325 76.645 145.005 ;
        RECT 73.895 144.295 74.840 144.325 ;
        RECT 27.115 144.085 27.285 144.295 ;
        RECT 29.435 144.275 29.585 144.295 ;
        RECT 28.955 144.130 29.115 144.250 ;
        RECT 29.415 144.105 29.585 144.275 ;
        RECT 31.990 144.105 32.160 144.295 ;
        RECT 38.615 144.085 38.785 144.275 ;
        RECT 39.720 144.105 39.890 144.295 ;
        RECT 48.275 144.085 48.445 144.275 ;
        RECT 49.250 144.135 49.370 144.245 ;
        RECT 49.655 144.105 49.825 144.295 ;
        RECT 53.520 144.105 53.690 144.295 ;
        RECT 55.170 144.105 55.340 144.275 ;
        RECT 56.555 144.085 56.725 144.275 ;
        RECT 57.070 144.135 57.190 144.245 ;
        RECT 57.470 144.105 57.640 144.295 ;
        RECT 57.940 144.105 58.110 144.295 ;
        RECT 60.880 144.085 61.050 144.275 ;
        RECT 62.535 144.085 62.705 144.275 ;
        RECT 62.995 144.105 63.165 144.295 ;
        RECT 67.780 144.105 67.950 144.295 ;
        RECT 68.995 144.275 69.145 144.295 ;
        RECT 68.570 144.135 68.690 144.245 ;
        RECT 68.975 144.105 69.145 144.275 ;
        RECT 71.275 144.105 71.445 144.295 ;
        RECT 72.195 144.085 72.365 144.275 ;
        RECT 73.575 144.085 73.745 144.275 ;
        RECT 74.090 144.135 74.210 144.245 ;
        RECT 76.330 144.105 76.500 144.325 ;
        RECT 76.655 144.295 80.130 145.205 ;
        RECT 83.995 144.975 84.925 145.205 ;
        RECT 81.025 144.295 84.925 144.975 ;
        RECT 84.935 144.295 86.305 145.075 ;
        RECT 87.245 144.380 87.675 145.165 ;
        RECT 90.895 144.975 91.825 145.205 ;
        RECT 87.925 144.295 91.825 144.975 ;
        RECT 91.845 144.295 93.195 145.205 ;
        RECT 93.415 145.115 94.365 145.205 ;
        RECT 96.655 145.115 97.605 145.205 ;
        RECT 93.415 144.295 95.345 145.115 ;
        RECT 76.800 144.105 76.970 144.295 ;
        RECT 77.715 144.085 77.885 144.275 ;
        RECT 80.530 144.135 80.650 144.245 ;
        RECT 81.580 144.085 81.750 144.275 ;
        RECT 84.155 144.105 84.325 144.275 ;
        RECT 84.340 144.105 84.510 144.295 ;
        RECT 85.075 144.105 85.245 144.295 ;
        RECT 86.915 144.140 87.075 144.250 ;
        RECT 91.240 144.105 91.410 144.295 ;
        RECT 91.975 144.105 92.145 144.295 ;
        RECT 95.195 144.275 95.345 144.295 ;
        RECT 95.675 144.295 97.605 145.115 ;
        RECT 98.475 145.115 99.425 145.205 ;
        RECT 100.775 145.115 101.725 145.205 ;
        RECT 98.475 144.295 100.405 145.115 ;
        RECT 100.775 144.295 102.705 145.115 ;
        RECT 102.885 144.295 104.235 145.205 ;
        RECT 104.265 144.295 105.615 145.205 ;
        RECT 106.555 144.295 107.925 145.075 ;
        RECT 107.945 144.295 109.295 145.205 ;
        RECT 109.315 144.295 110.685 145.075 ;
        RECT 110.695 144.295 112.065 145.075 ;
        RECT 112.075 144.295 113.445 145.105 ;
        RECT 95.675 144.275 95.825 144.295 ;
        RECT 100.255 144.275 100.405 144.295 ;
        RECT 102.555 144.275 102.705 144.295 ;
        RECT 84.155 144.085 84.305 144.105 ;
        RECT 93.355 144.085 93.525 144.275 ;
        RECT 93.815 144.085 93.985 144.275 ;
        RECT 95.195 144.105 95.365 144.275 ;
        RECT 95.655 144.105 95.825 144.275 ;
        RECT 98.010 144.135 98.130 144.245 ;
        RECT 99.520 144.085 99.690 144.275 ;
        RECT 100.255 144.105 100.425 144.275 ;
        RECT 101.635 144.085 101.805 144.275 ;
        RECT 102.555 144.105 102.725 144.275 ;
        RECT 103.015 144.105 103.185 144.295 ;
        RECT 104.395 144.105 104.565 144.295 ;
        RECT 106.235 144.140 106.395 144.250 ;
        RECT 106.695 144.105 106.865 144.295 ;
        RECT 108.995 144.105 109.165 144.295 ;
        RECT 109.455 144.105 109.625 144.295 ;
        RECT 111.295 144.085 111.465 144.275 ;
        RECT 111.755 144.245 111.925 144.295 ;
        RECT 111.755 144.135 111.930 144.245 ;
        RECT 111.755 144.105 111.925 144.135 ;
        RECT 113.135 144.085 113.305 144.295 ;
        RECT 26.975 143.275 28.345 144.085 ;
        RECT 29.645 143.405 38.925 144.085 ;
        RECT 39.305 143.405 48.585 144.085 ;
        RECT 29.645 143.285 31.980 143.405 ;
        RECT 29.645 143.175 30.565 143.285 ;
        RECT 36.645 143.185 37.565 143.405 ;
        RECT 39.305 143.285 41.640 143.405 ;
        RECT 39.305 143.175 40.225 143.285 ;
        RECT 46.305 143.185 47.225 143.405 ;
        RECT 48.605 143.215 49.035 144.000 ;
        RECT 50.595 143.405 54.545 144.085 ;
        RECT 55.495 143.305 56.865 144.085 ;
        RECT 57.565 143.405 61.465 144.085 ;
        RECT 60.535 143.175 61.465 143.405 ;
        RECT 61.475 143.275 62.845 144.085 ;
        RECT 63.225 143.405 72.505 144.085 ;
        RECT 63.225 143.285 65.560 143.405 ;
        RECT 63.225 143.175 64.145 143.285 ;
        RECT 70.225 143.185 71.145 143.405 ;
        RECT 72.515 143.305 73.885 144.085 ;
        RECT 74.365 143.215 74.795 144.000 ;
        RECT 74.815 143.175 77.975 144.085 ;
        RECT 78.265 143.405 82.165 144.085 ;
        RECT 81.235 143.175 82.165 143.405 ;
        RECT 82.375 143.265 84.305 144.085 ;
        RECT 84.560 143.405 93.665 144.085 ;
        RECT 93.675 143.305 95.045 144.085 ;
        RECT 96.205 143.405 100.105 144.085 ;
        RECT 82.375 143.175 83.325 143.265 ;
        RECT 99.175 143.175 100.105 143.405 ;
        RECT 100.125 143.215 100.555 144.000 ;
        RECT 100.575 143.305 101.945 144.085 ;
        RECT 102.325 143.405 111.605 144.085 ;
        RECT 102.325 143.285 104.660 143.405 ;
        RECT 102.325 143.175 103.245 143.285 ;
        RECT 109.325 143.185 110.245 143.405 ;
        RECT 112.075 143.275 113.445 144.085 ;
      LAYER nwell ;
        RECT 26.780 140.055 113.640 142.885 ;
      LAYER pwell ;
        RECT 30.415 139.675 31.365 139.765 ;
        RECT 26.975 138.855 28.345 139.665 ;
        RECT 29.435 138.855 31.365 139.675 ;
        RECT 31.575 139.535 32.505 139.765 ;
        RECT 31.575 138.855 35.475 139.535 ;
        RECT 35.725 138.940 36.155 139.725 ;
        RECT 36.175 138.855 39.335 139.765 ;
        RECT 39.765 139.655 40.685 139.765 ;
        RECT 39.765 139.535 42.100 139.655 ;
        RECT 46.765 139.535 47.685 139.755 ;
        RECT 60.060 139.565 61.005 139.765 ;
        RECT 39.765 138.855 49.045 139.535 ;
        RECT 49.055 138.855 58.160 139.535 ;
        RECT 58.255 138.885 61.005 139.565 ;
        RECT 61.485 138.940 61.915 139.725 ;
        RECT 27.115 138.645 27.285 138.855 ;
        RECT 29.435 138.835 29.585 138.855 ;
        RECT 28.955 138.700 29.115 138.810 ;
        RECT 29.415 138.665 29.585 138.835 ;
        RECT 31.990 138.665 32.160 138.855 ;
        RECT 38.615 138.645 38.785 138.835 ;
        RECT 39.075 138.645 39.245 138.855 ;
        RECT 48.735 138.665 48.905 138.855 ;
        RECT 49.195 138.645 49.365 138.855 ;
        RECT 58.400 138.665 58.570 138.885 ;
        RECT 60.060 138.855 61.005 138.885 ;
        RECT 61.945 138.855 63.295 139.765 ;
        RECT 66.515 139.535 67.445 139.765 ;
        RECT 77.945 139.655 78.865 139.765 ;
        RECT 77.945 139.535 80.280 139.655 ;
        RECT 84.945 139.535 85.865 139.755 ;
        RECT 63.545 138.855 67.445 139.535 ;
        RECT 68.375 138.855 77.480 139.535 ;
        RECT 77.945 138.855 87.225 139.535 ;
        RECT 87.245 138.940 87.675 139.725 ;
        RECT 88.065 139.655 88.985 139.765 ;
        RECT 88.065 139.535 90.400 139.655 ;
        RECT 95.065 139.535 95.985 139.755 ;
        RECT 101.015 139.535 101.945 139.765 ;
        RECT 88.065 138.855 97.345 139.535 ;
        RECT 98.045 138.855 101.945 139.535 ;
        RECT 102.325 139.655 103.245 139.765 ;
        RECT 102.325 139.535 104.660 139.655 ;
        RECT 109.325 139.535 110.245 139.755 ;
        RECT 102.325 138.855 111.605 139.535 ;
        RECT 112.075 138.855 113.445 139.665 ;
        RECT 58.910 138.695 59.030 138.805 ;
        RECT 59.315 138.645 59.485 138.835 ;
        RECT 61.210 138.695 61.330 138.805 ;
        RECT 62.075 138.665 62.245 138.855 ;
        RECT 66.860 138.665 67.030 138.855 ;
        RECT 68.055 138.700 68.215 138.810 ;
        RECT 68.515 138.665 68.685 138.855 ;
        RECT 69.895 138.645 70.065 138.835 ;
        RECT 70.410 138.695 70.530 138.805 ;
        RECT 70.815 138.665 70.985 138.835 ;
        RECT 70.835 138.645 70.985 138.665 ;
        RECT 74.035 138.645 74.205 138.835 ;
        RECT 78.360 138.645 78.530 138.835 ;
        RECT 80.935 138.665 81.105 138.835 ;
        RECT 83.235 138.665 83.405 138.835 ;
        RECT 84.155 138.690 84.315 138.800 ;
        RECT 86.915 138.665 87.085 138.855 ;
        RECT 80.935 138.645 81.085 138.665 ;
        RECT 83.235 138.645 83.385 138.665 ;
        RECT 88.020 138.645 88.190 138.835 ;
        RECT 89.675 138.645 89.845 138.835 ;
        RECT 90.135 138.645 90.305 138.835 ;
        RECT 91.570 138.695 91.690 138.805 ;
        RECT 95.380 138.645 95.550 138.835 ;
        RECT 97.035 138.665 97.205 138.855 ;
        RECT 97.550 138.695 97.670 138.805 ;
        RECT 99.520 138.645 99.690 138.835 ;
        RECT 101.360 138.665 101.530 138.855 ;
        RECT 109.915 138.645 110.085 138.835 ;
        RECT 111.295 138.645 111.465 138.855 ;
        RECT 111.810 138.695 111.930 138.805 ;
        RECT 113.135 138.645 113.305 138.855 ;
        RECT 26.975 137.835 28.345 138.645 ;
        RECT 28.555 137.965 38.925 138.645 ;
        RECT 38.935 137.965 48.215 138.645 ;
        RECT 28.555 137.735 30.765 137.965 ;
        RECT 33.485 137.745 34.415 137.965 ;
        RECT 40.295 137.745 41.215 137.965 ;
        RECT 45.880 137.845 48.215 137.965 ;
        RECT 47.295 137.735 48.215 137.845 ;
        RECT 48.605 137.775 49.035 138.560 ;
        RECT 49.055 137.965 58.335 138.645 ;
        RECT 50.415 137.745 51.335 137.965 ;
        RECT 56.000 137.845 58.335 137.965 ;
        RECT 59.175 137.865 60.545 138.645 ;
        RECT 60.925 137.965 70.205 138.645 ;
        RECT 57.415 137.735 58.335 137.845 ;
        RECT 60.925 137.845 63.260 137.965 ;
        RECT 60.925 137.735 61.845 137.845 ;
        RECT 67.925 137.745 68.845 137.965 ;
        RECT 70.835 137.825 72.765 138.645 ;
        RECT 72.975 137.865 74.345 138.645 ;
        RECT 71.815 137.735 72.765 137.825 ;
        RECT 74.365 137.775 74.795 138.560 ;
        RECT 75.045 137.965 78.945 138.645 ;
        RECT 78.015 137.735 78.945 137.965 ;
        RECT 79.155 137.825 81.085 138.645 ;
        RECT 81.455 137.825 83.385 138.645 ;
        RECT 84.705 137.965 88.605 138.645 ;
        RECT 79.155 137.735 80.105 137.825 ;
        RECT 81.455 137.735 82.405 137.825 ;
        RECT 87.675 137.735 88.605 137.965 ;
        RECT 88.625 137.735 89.975 138.645 ;
        RECT 90.005 137.735 91.355 138.645 ;
        RECT 92.065 137.965 95.965 138.645 ;
        RECT 96.205 137.965 100.105 138.645 ;
        RECT 95.035 137.735 95.965 137.965 ;
        RECT 99.175 137.735 100.105 137.965 ;
        RECT 100.125 137.775 100.555 138.560 ;
        RECT 100.945 137.965 110.225 138.645 ;
        RECT 100.945 137.845 103.280 137.965 ;
        RECT 100.945 137.735 101.865 137.845 ;
        RECT 107.945 137.745 108.865 137.965 ;
        RECT 110.235 137.865 111.605 138.645 ;
        RECT 112.075 137.835 113.445 138.645 ;
      LAYER nwell ;
        RECT 26.780 134.615 113.640 137.445 ;
      LAYER pwell ;
        RECT 26.975 133.415 28.345 134.225 ;
        RECT 28.355 133.415 29.725 134.195 ;
        RECT 29.745 133.415 31.095 134.325 ;
        RECT 34.315 134.095 35.245 134.325 ;
        RECT 31.345 133.415 35.245 134.095 ;
        RECT 35.725 133.500 36.155 134.285 ;
        RECT 36.315 133.415 38.925 134.325 ;
        RECT 40.295 134.095 41.215 134.315 ;
        RECT 47.295 134.215 48.215 134.325 ;
        RECT 45.880 134.095 48.215 134.215 ;
        RECT 38.935 133.415 48.215 134.095 ;
        RECT 48.965 134.215 49.885 134.325 ;
        RECT 48.965 134.095 51.300 134.215 ;
        RECT 55.965 134.095 56.885 134.315 ;
        RECT 58.255 134.125 59.200 134.325 ;
        RECT 48.965 133.415 58.245 134.095 ;
        RECT 58.255 133.445 61.005 134.125 ;
        RECT 61.485 133.500 61.915 134.285 ;
        RECT 62.305 134.215 63.225 134.325 ;
        RECT 62.305 134.095 64.640 134.215 ;
        RECT 69.305 134.095 70.225 134.315 ;
        RECT 71.965 134.215 72.885 134.325 ;
        RECT 71.965 134.095 74.300 134.215 ;
        RECT 78.965 134.095 79.885 134.315 ;
        RECT 81.255 134.095 82.185 134.325 ;
        RECT 58.255 133.415 59.200 133.445 ;
        RECT 27.115 133.205 27.285 133.415 ;
        RECT 28.495 133.205 28.665 133.415 ;
        RECT 29.875 133.225 30.045 133.415 ;
        RECT 34.660 133.225 34.830 133.415 ;
        RECT 35.450 133.255 35.570 133.365 ;
        RECT 38.610 133.225 38.780 133.415 ;
        RECT 39.075 133.225 39.245 133.415 ;
        RECT 39.995 133.205 40.165 133.395 ;
        RECT 40.730 133.205 40.900 133.395 ;
        RECT 44.870 133.205 45.040 133.395 ;
        RECT 52.600 133.205 52.770 133.395 ;
        RECT 57.935 133.225 58.105 133.415 ;
        RECT 60.690 133.225 60.860 133.445 ;
        RECT 62.305 133.415 71.585 134.095 ;
        RECT 71.965 133.415 81.245 134.095 ;
        RECT 81.255 133.415 85.155 134.095 ;
        RECT 85.395 133.415 86.765 134.195 ;
        RECT 87.245 133.500 87.675 134.285 ;
        RECT 88.065 134.215 88.985 134.325 ;
        RECT 88.065 134.095 90.400 134.215 ;
        RECT 95.065 134.095 95.985 134.315 ;
        RECT 97.725 134.215 98.645 134.325 ;
        RECT 97.725 134.095 100.060 134.215 ;
        RECT 104.725 134.095 105.645 134.315 ;
        RECT 88.065 133.415 97.345 134.095 ;
        RECT 97.725 133.415 107.005 134.095 ;
        RECT 107.025 133.415 108.375 134.325 ;
        RECT 108.855 133.415 110.685 134.225 ;
        RECT 110.695 133.415 112.065 134.195 ;
        RECT 112.075 133.415 113.445 134.225 ;
        RECT 61.210 133.255 61.330 133.365 ;
        RECT 62.535 133.205 62.705 133.395 ;
        RECT 66.400 133.205 66.570 133.395 ;
        RECT 67.135 133.205 67.305 133.395 ;
        RECT 68.570 133.255 68.690 133.365 ;
        RECT 71.275 133.205 71.445 133.415 ;
        RECT 71.735 133.205 71.905 133.395 ;
        RECT 73.115 133.205 73.285 133.395 ;
        RECT 74.955 133.205 75.125 133.395 ;
        RECT 80.935 133.225 81.105 133.415 ;
        RECT 81.670 133.225 81.840 133.415 ;
        RECT 86.455 133.225 86.625 133.415 ;
        RECT 86.970 133.255 87.090 133.365 ;
        RECT 93.815 133.205 93.985 133.395 ;
        RECT 94.275 133.205 94.445 133.395 ;
        RECT 95.710 133.255 95.830 133.365 ;
        RECT 97.035 133.225 97.205 133.415 ;
        RECT 99.520 133.205 99.690 133.395 ;
        RECT 100.715 133.205 100.885 133.395 ;
        RECT 102.555 133.250 102.715 133.360 ;
        RECT 103.015 133.205 103.185 133.395 ;
        RECT 104.855 133.250 105.015 133.360 ;
        RECT 105.315 133.205 105.485 133.395 ;
        RECT 106.695 133.205 106.865 133.415 ;
        RECT 107.155 133.225 107.325 133.415 ;
        RECT 108.590 133.360 108.710 133.365 ;
        RECT 108.535 133.255 108.710 133.360 ;
        RECT 108.535 133.250 108.695 133.255 ;
        RECT 109.915 133.205 110.085 133.395 ;
        RECT 110.375 133.205 110.545 133.415 ;
        RECT 111.745 133.365 111.915 133.415 ;
        RECT 111.745 133.255 111.930 133.365 ;
        RECT 111.745 133.225 111.915 133.255 ;
        RECT 113.135 133.205 113.305 133.415 ;
        RECT 26.975 132.395 28.345 133.205 ;
        RECT 28.355 132.425 29.725 133.205 ;
        RECT 29.935 132.525 40.305 133.205 ;
        RECT 40.315 132.525 44.215 133.205 ;
        RECT 44.455 132.525 48.355 133.205 ;
        RECT 29.935 132.295 32.145 132.525 ;
        RECT 34.865 132.305 35.795 132.525 ;
        RECT 40.315 132.295 41.245 132.525 ;
        RECT 44.455 132.295 45.385 132.525 ;
        RECT 48.605 132.335 49.035 133.120 ;
        RECT 49.285 132.525 53.185 133.205 ;
        RECT 52.255 132.295 53.185 132.525 ;
        RECT 53.565 132.525 62.845 133.205 ;
        RECT 63.085 132.525 66.985 133.205 ;
        RECT 53.565 132.405 55.900 132.525 ;
        RECT 53.565 132.295 54.485 132.405 ;
        RECT 60.565 132.305 61.485 132.525 ;
        RECT 66.055 132.295 66.985 132.525 ;
        RECT 66.995 132.425 68.365 133.205 ;
        RECT 68.835 132.395 71.585 133.205 ;
        RECT 71.605 132.295 72.955 133.205 ;
        RECT 72.985 132.295 74.335 133.205 ;
        RECT 74.365 132.335 74.795 133.120 ;
        RECT 74.815 132.525 84.095 133.205 ;
        RECT 76.175 132.305 77.095 132.525 ;
        RECT 81.760 132.405 84.095 132.525 ;
        RECT 83.175 132.295 84.095 132.405 ;
        RECT 84.845 132.525 94.125 133.205 ;
        RECT 84.845 132.405 87.180 132.525 ;
        RECT 84.845 132.295 85.765 132.405 ;
        RECT 91.845 132.305 92.765 132.525 ;
        RECT 94.135 132.425 95.505 133.205 ;
        RECT 96.205 132.525 100.105 133.205 ;
        RECT 99.175 132.295 100.105 132.525 ;
        RECT 100.125 132.335 100.555 133.120 ;
        RECT 100.575 132.425 101.945 133.205 ;
        RECT 102.885 132.295 104.235 133.205 ;
        RECT 105.175 132.425 106.545 133.205 ;
        RECT 106.565 132.295 107.915 133.205 ;
        RECT 108.855 132.425 110.225 133.205 ;
        RECT 110.245 132.295 111.595 133.205 ;
        RECT 112.075 132.395 113.445 133.205 ;
      LAYER nwell ;
        RECT 26.780 129.175 113.640 132.005 ;
      LAYER pwell ;
        RECT 26.975 127.975 28.345 128.785 ;
        RECT 28.355 127.975 29.725 128.755 ;
        RECT 29.745 127.975 31.095 128.885 ;
        RECT 31.585 127.975 32.935 128.885 ;
        RECT 33.875 127.975 35.245 128.755 ;
        RECT 35.725 128.060 36.155 128.845 ;
        RECT 37.105 127.975 38.455 128.885 ;
        RECT 38.475 127.975 39.845 128.755 ;
        RECT 39.865 127.975 41.215 128.885 ;
        RECT 41.235 127.975 42.605 128.755 ;
        RECT 42.815 128.655 45.025 128.885 ;
        RECT 47.745 128.655 48.675 128.875 ;
        RECT 42.815 127.975 53.185 128.655 ;
        RECT 54.125 127.975 55.475 128.885 ;
        RECT 59.395 128.795 60.345 128.885 ;
        RECT 55.495 127.975 56.865 128.755 ;
        RECT 56.875 127.975 58.245 128.755 ;
        RECT 58.415 127.975 60.345 128.795 ;
        RECT 61.485 128.060 61.915 128.845 ;
        RECT 62.395 127.975 64.225 128.785 ;
        RECT 64.245 127.975 65.595 128.885 ;
        RECT 65.615 127.975 69.285 128.785 ;
        RECT 69.295 127.975 74.805 128.785 ;
        RECT 74.815 127.975 76.185 128.755 ;
        RECT 76.195 127.975 77.565 128.755 ;
        RECT 77.575 127.975 78.945 128.755 ;
        RECT 78.955 127.975 81.565 128.885 ;
        RECT 81.715 127.975 85.385 128.785 ;
        RECT 85.405 127.975 86.755 128.885 ;
        RECT 87.245 128.060 87.675 128.845 ;
        RECT 88.615 127.975 89.985 128.755 ;
        RECT 90.005 127.975 91.355 128.885 ;
        RECT 91.845 127.975 93.195 128.885 ;
        RECT 93.215 127.975 94.585 128.755 ;
        RECT 94.595 127.975 95.965 128.755 ;
        RECT 95.985 127.975 97.335 128.885 ;
        RECT 98.275 127.975 99.645 128.755 ;
        RECT 100.125 127.975 101.475 128.885 ;
        RECT 106.005 128.655 106.935 128.875 ;
        RECT 109.655 128.655 111.865 128.885 ;
        RECT 101.495 127.975 111.865 128.655 ;
        RECT 112.075 127.975 113.445 128.785 ;
        RECT 27.115 127.765 27.285 127.975 ;
        RECT 28.495 127.925 28.665 127.975 ;
        RECT 28.495 127.815 28.670 127.925 ;
        RECT 28.495 127.785 28.665 127.815 ;
        RECT 29.875 127.765 30.045 127.975 ;
        RECT 30.335 127.765 30.505 127.955 ;
        RECT 31.310 127.815 31.430 127.925 ;
        RECT 31.715 127.785 31.885 127.975 ;
        RECT 32.635 127.765 32.805 127.955 ;
        RECT 33.095 127.765 33.265 127.955 ;
        RECT 33.555 127.820 33.715 127.930 ;
        RECT 34.015 127.785 34.185 127.975 ;
        RECT 34.475 127.765 34.645 127.955 ;
        RECT 35.450 127.815 35.570 127.925 ;
        RECT 35.855 127.765 36.025 127.955 ;
        RECT 36.775 127.820 36.935 127.930 ;
        RECT 37.235 127.765 37.405 127.975 ;
        RECT 38.615 127.785 38.785 127.975 ;
        RECT 39.995 127.785 40.165 127.975 ;
        RECT 42.295 127.785 42.465 127.975 ;
        RECT 48.275 127.810 48.435 127.920 ;
        RECT 49.250 127.815 49.370 127.925 ;
        RECT 51.950 127.765 52.120 127.955 ;
        RECT 52.875 127.785 53.045 127.975 ;
        RECT 53.795 127.820 53.955 127.930 ;
        RECT 54.255 127.765 54.425 127.975 ;
        RECT 54.715 127.765 54.885 127.955 ;
        RECT 55.635 127.785 55.805 127.975 ;
        RECT 56.095 127.765 56.265 127.955 ;
        RECT 57.015 127.785 57.185 127.975 ;
        RECT 58.415 127.955 58.565 127.975 ;
        RECT 58.395 127.785 58.565 127.955 ;
        RECT 61.155 127.820 61.315 127.930 ;
        RECT 62.130 127.815 62.250 127.925 ;
        RECT 63.915 127.785 64.085 127.975 ;
        RECT 65.295 127.785 65.465 127.975 ;
        RECT 66.675 127.765 66.845 127.955 ;
        RECT 68.055 127.765 68.225 127.955 ;
        RECT 68.975 127.785 69.145 127.975 ;
        RECT 69.435 127.765 69.605 127.955 ;
        RECT 70.870 127.815 70.990 127.925 ;
        RECT 72.655 127.765 72.825 127.955 ;
        RECT 73.115 127.765 73.285 127.955 ;
        RECT 74.495 127.785 74.665 127.975 ;
        RECT 74.955 127.765 75.125 127.975 ;
        RECT 76.335 127.785 76.505 127.975 ;
        RECT 78.635 127.785 78.805 127.975 ;
        RECT 79.100 127.785 79.270 127.975 ;
        RECT 85.075 127.785 85.245 127.975 ;
        RECT 85.535 127.785 85.705 127.975 ;
        RECT 85.995 127.810 86.155 127.920 ;
        RECT 86.455 127.765 86.625 127.955 ;
        RECT 86.970 127.815 87.090 127.925 ;
        RECT 88.295 127.820 88.455 127.930 ;
        RECT 88.755 127.785 88.925 127.975 ;
        RECT 90.135 127.785 90.305 127.975 ;
        RECT 91.570 127.815 91.690 127.925 ;
        RECT 92.895 127.785 93.065 127.975 ;
        RECT 93.355 127.785 93.525 127.975 ;
        RECT 94.735 127.785 94.905 127.975 ;
        RECT 97.035 127.785 97.205 127.975 ;
        RECT 97.955 127.765 98.125 127.955 ;
        RECT 98.415 127.785 98.585 127.975 ;
        RECT 99.335 127.765 99.505 127.955 ;
        RECT 99.850 127.815 99.970 127.925 ;
        RECT 100.255 127.785 100.425 127.975 ;
        RECT 101.175 127.810 101.335 127.920 ;
        RECT 101.635 127.765 101.805 127.975 ;
        RECT 113.135 127.765 113.305 127.975 ;
        RECT 26.975 126.955 28.345 127.765 ;
        RECT 28.825 126.855 30.175 127.765 ;
        RECT 30.195 126.985 31.565 127.765 ;
        RECT 31.575 126.955 32.945 127.765 ;
        RECT 32.955 126.985 34.325 127.765 ;
        RECT 34.335 126.985 35.705 127.765 ;
        RECT 35.715 126.985 37.085 127.765 ;
        RECT 37.095 127.085 47.465 127.765 ;
        RECT 41.605 126.865 42.535 127.085 ;
        RECT 45.255 126.855 47.465 127.085 ;
        RECT 48.605 126.895 49.035 127.680 ;
        RECT 49.655 126.855 52.265 127.765 ;
        RECT 53.205 126.855 54.555 127.765 ;
        RECT 54.575 126.985 55.945 127.765 ;
        RECT 55.955 127.085 66.325 127.765 ;
        RECT 60.465 126.865 61.395 127.085 ;
        RECT 64.115 126.855 66.325 127.085 ;
        RECT 66.535 126.985 67.905 127.765 ;
        RECT 67.925 126.855 69.275 127.765 ;
        RECT 69.295 126.985 70.665 127.765 ;
        RECT 71.135 126.955 72.965 127.765 ;
        RECT 72.975 126.985 74.345 127.765 ;
        RECT 74.365 126.895 74.795 127.680 ;
        RECT 74.815 127.085 85.185 127.765 ;
        RECT 79.325 126.865 80.255 127.085 ;
        RECT 82.975 126.855 85.185 127.085 ;
        RECT 86.315 126.985 87.685 127.765 ;
        RECT 87.895 127.085 98.265 127.765 ;
        RECT 87.895 126.855 90.105 127.085 ;
        RECT 92.825 126.865 93.755 127.085 ;
        RECT 98.275 126.985 99.645 127.765 ;
        RECT 100.125 126.895 100.555 127.680 ;
        RECT 101.495 127.085 111.865 127.765 ;
        RECT 106.005 126.865 106.935 127.085 ;
        RECT 109.655 126.855 111.865 127.085 ;
        RECT 112.075 126.955 113.445 127.765 ;
      LAYER nwell ;
        RECT 26.780 123.735 113.640 126.565 ;
      LAYER pwell ;
        RECT 26.975 122.535 28.345 123.345 ;
        RECT 28.365 122.535 29.715 123.445 ;
        RECT 29.735 122.535 31.565 123.345 ;
        RECT 31.585 122.535 32.935 123.445 ;
        RECT 32.965 122.535 34.315 123.445 ;
        RECT 34.345 122.535 35.695 123.445 ;
        RECT 35.725 122.620 36.155 123.405 ;
        RECT 36.185 122.535 37.535 123.445 ;
        RECT 37.555 122.535 38.925 123.315 ;
        RECT 38.945 122.535 40.295 123.445 ;
        RECT 44.825 123.215 45.755 123.435 ;
        RECT 48.475 123.215 50.685 123.445 ;
        RECT 40.315 122.535 50.685 123.215 ;
        RECT 51.095 123.215 53.305 123.445 ;
        RECT 56.025 123.215 56.955 123.435 ;
        RECT 51.095 122.535 61.465 123.215 ;
        RECT 61.485 122.620 61.915 123.405 ;
        RECT 62.135 123.215 64.345 123.445 ;
        RECT 67.065 123.215 67.995 123.435 ;
        RECT 72.715 123.215 74.925 123.445 ;
        RECT 77.645 123.215 78.575 123.435 ;
        RECT 62.135 122.535 72.505 123.215 ;
        RECT 72.715 122.535 83.085 123.215 ;
        RECT 83.105 122.535 84.455 123.445 ;
        RECT 84.485 122.535 85.835 123.445 ;
        RECT 85.865 122.535 87.215 123.445 ;
        RECT 87.245 122.620 87.675 123.405 ;
        RECT 87.895 123.215 90.105 123.445 ;
        RECT 92.825 123.215 93.755 123.435 ;
        RECT 98.475 123.215 100.685 123.445 ;
        RECT 103.405 123.215 104.335 123.435 ;
        RECT 87.895 122.535 98.265 123.215 ;
        RECT 98.475 122.535 108.845 123.215 ;
        RECT 108.865 122.535 110.215 123.445 ;
        RECT 110.235 122.535 111.605 123.315 ;
        RECT 112.075 122.535 113.445 123.345 ;
        RECT 27.115 122.325 27.285 122.535 ;
        RECT 29.415 122.345 29.585 122.535 ;
        RECT 29.875 122.325 30.045 122.515 ;
        RECT 31.255 122.345 31.425 122.535 ;
        RECT 32.635 122.345 32.805 122.535 ;
        RECT 33.095 122.345 33.265 122.535 ;
        RECT 34.475 122.345 34.645 122.535 ;
        RECT 35.395 122.325 35.565 122.515 ;
        RECT 36.315 122.345 36.485 122.535 ;
        RECT 37.695 122.345 37.865 122.535 ;
        RECT 39.075 122.345 39.245 122.535 ;
        RECT 40.455 122.345 40.625 122.535 ;
        RECT 46.435 122.325 46.605 122.515 ;
        RECT 46.950 122.375 47.070 122.485 ;
        RECT 48.275 122.325 48.445 122.515 ;
        RECT 49.655 122.370 49.815 122.480 ;
        RECT 50.115 122.325 50.285 122.515 ;
        RECT 52.875 122.325 53.045 122.515 ;
        RECT 54.255 122.325 54.425 122.515 ;
        RECT 55.175 122.370 55.335 122.480 ;
        RECT 56.555 122.325 56.725 122.515 ;
        RECT 57.070 122.375 57.190 122.485 ;
        RECT 59.775 122.325 59.945 122.515 ;
        RECT 60.235 122.325 60.405 122.515 ;
        RECT 61.155 122.345 61.325 122.535 ;
        RECT 62.130 122.375 62.250 122.485 ;
        RECT 62.535 122.325 62.705 122.515 ;
        RECT 72.195 122.345 72.365 122.535 ;
        RECT 74.035 122.325 74.205 122.515 ;
        RECT 75.010 122.375 75.130 122.485 ;
        RECT 76.335 122.325 76.505 122.515 ;
        RECT 76.795 122.325 76.965 122.515 ;
        RECT 82.775 122.345 82.945 122.535 ;
        RECT 84.155 122.345 84.325 122.535 ;
        RECT 85.535 122.345 85.705 122.535 ;
        RECT 86.915 122.345 87.085 122.535 ;
        RECT 87.835 122.325 88.005 122.515 ;
        RECT 89.270 122.375 89.390 122.485 ;
        RECT 97.955 122.345 98.125 122.535 ;
        RECT 99.795 122.325 99.965 122.515 ;
        RECT 101.175 122.370 101.335 122.480 ;
        RECT 108.535 122.345 108.705 122.535 ;
        RECT 109.915 122.345 110.085 122.535 ;
        RECT 111.295 122.345 111.465 122.535 ;
        RECT 111.755 122.485 111.925 122.515 ;
        RECT 111.755 122.375 111.930 122.485 ;
        RECT 111.755 122.325 111.925 122.375 ;
        RECT 113.135 122.325 113.305 122.535 ;
        RECT 26.975 121.515 28.345 122.325 ;
        RECT 28.355 121.515 30.185 122.325 ;
        RECT 30.195 121.515 35.705 122.325 ;
        RECT 35.725 121.455 36.155 122.240 ;
        RECT 36.375 121.645 46.745 122.325 ;
        RECT 36.375 121.415 38.585 121.645 ;
        RECT 41.305 121.425 42.235 121.645 ;
        RECT 47.225 121.415 48.575 122.325 ;
        RECT 48.605 121.455 49.035 122.240 ;
        RECT 49.975 121.545 51.345 122.325 ;
        RECT 51.355 121.515 53.185 122.325 ;
        RECT 53.195 121.545 54.565 122.325 ;
        RECT 55.505 121.415 56.855 122.325 ;
        RECT 57.335 121.515 60.085 122.325 ;
        RECT 60.105 121.415 61.455 122.325 ;
        RECT 61.485 121.455 61.915 122.240 ;
        RECT 62.405 121.415 63.755 122.325 ;
        RECT 63.975 121.645 74.345 122.325 ;
        RECT 63.975 121.415 66.185 121.645 ;
        RECT 68.905 121.425 69.835 121.645 ;
        RECT 74.365 121.455 74.795 122.240 ;
        RECT 75.285 121.415 76.635 122.325 ;
        RECT 76.655 121.645 87.025 122.325 ;
        RECT 81.165 121.425 82.095 121.645 ;
        RECT 84.815 121.415 87.025 121.645 ;
        RECT 87.245 121.455 87.675 122.240 ;
        RECT 87.705 121.415 89.055 122.325 ;
        RECT 89.735 121.645 100.105 122.325 ;
        RECT 89.735 121.415 91.945 121.645 ;
        RECT 94.665 121.425 95.595 121.645 ;
        RECT 100.125 121.455 100.555 122.240 ;
        RECT 101.695 121.645 112.065 122.325 ;
        RECT 101.695 121.415 103.905 121.645 ;
        RECT 106.625 121.425 107.555 121.645 ;
        RECT 112.075 121.515 113.445 122.325 ;
      LAYER nwell ;
        RECT 26.780 119.520 113.640 121.125 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 26.970 203.945 113.450 204.115 ;
        RECT 27.055 203.195 28.265 203.945 ;
        RECT 27.055 202.655 27.575 203.195 ;
        RECT 28.955 203.125 29.165 203.945 ;
        RECT 29.335 203.145 29.665 203.775 ;
        RECT 27.745 202.485 28.265 203.025 ;
        RECT 29.335 202.545 29.585 203.145 ;
        RECT 29.835 203.125 30.065 203.945 ;
        RECT 30.315 203.125 30.545 203.945 ;
        RECT 30.715 203.145 31.045 203.775 ;
        RECT 29.755 202.705 30.085 202.955 ;
        RECT 30.295 202.705 30.625 202.955 ;
        RECT 30.795 202.545 31.045 203.145 ;
        RECT 31.215 203.125 31.425 203.945 ;
        RECT 31.695 203.125 31.925 203.945 ;
        RECT 32.095 203.145 32.425 203.775 ;
        RECT 31.675 202.705 32.005 202.955 ;
        RECT 32.175 202.545 32.425 203.145 ;
        RECT 32.595 203.125 32.805 203.945 ;
        RECT 33.035 203.175 35.625 203.945 ;
        RECT 35.795 203.220 36.085 203.945 ;
        RECT 36.255 203.175 38.845 203.945 ;
        RECT 39.105 203.395 39.275 203.775 ;
        RECT 39.455 203.565 39.785 203.945 ;
        RECT 39.105 203.225 39.770 203.395 ;
        RECT 39.965 203.270 40.225 203.775 ;
        RECT 27.055 201.395 28.265 202.485 ;
        RECT 28.955 201.395 29.165 202.535 ;
        RECT 29.335 201.565 29.665 202.545 ;
        RECT 29.835 201.395 30.065 202.535 ;
        RECT 30.315 201.395 30.545 202.535 ;
        RECT 30.715 201.565 31.045 202.545 ;
        RECT 31.215 201.395 31.425 202.535 ;
        RECT 31.695 201.395 31.925 202.535 ;
        RECT 32.095 201.565 32.425 202.545 ;
        RECT 32.595 201.395 32.805 202.535 ;
        RECT 33.035 202.485 34.245 203.005 ;
        RECT 34.415 202.655 35.625 203.175 ;
        RECT 33.035 201.395 35.625 202.485 ;
        RECT 35.795 201.395 36.085 202.560 ;
        RECT 36.255 202.485 37.465 203.005 ;
        RECT 37.635 202.655 38.845 203.175 ;
        RECT 39.035 202.675 39.365 203.045 ;
        RECT 39.600 202.970 39.770 203.225 ;
        RECT 39.600 202.640 39.885 202.970 ;
        RECT 39.600 202.495 39.770 202.640 ;
        RECT 36.255 201.395 38.845 202.485 ;
        RECT 39.105 202.325 39.770 202.495 ;
        RECT 40.055 202.470 40.225 203.270 ;
        RECT 40.455 203.125 40.665 203.945 ;
        RECT 40.835 203.145 41.165 203.775 ;
        RECT 40.835 202.545 41.085 203.145 ;
        RECT 41.335 203.125 41.565 203.945 ;
        RECT 41.815 203.125 42.045 203.945 ;
        RECT 42.215 203.145 42.545 203.775 ;
        RECT 41.255 202.705 41.585 202.955 ;
        RECT 41.795 202.705 42.125 202.955 ;
        RECT 42.295 202.545 42.545 203.145 ;
        RECT 42.715 203.125 42.925 203.945 ;
        RECT 43.245 203.395 43.415 203.775 ;
        RECT 43.595 203.565 43.925 203.945 ;
        RECT 43.245 203.225 43.910 203.395 ;
        RECT 44.105 203.270 44.365 203.775 ;
        RECT 43.175 202.675 43.505 203.045 ;
        RECT 43.740 202.970 43.910 203.225 ;
        RECT 39.105 201.565 39.275 202.325 ;
        RECT 39.455 201.395 39.785 202.155 ;
        RECT 39.955 201.565 40.225 202.470 ;
        RECT 40.455 201.395 40.665 202.535 ;
        RECT 40.835 201.565 41.165 202.545 ;
        RECT 41.335 201.395 41.565 202.535 ;
        RECT 41.815 201.395 42.045 202.535 ;
        RECT 42.215 201.565 42.545 202.545 ;
        RECT 43.740 202.640 44.025 202.970 ;
        RECT 42.715 201.395 42.925 202.535 ;
        RECT 43.740 202.495 43.910 202.640 ;
        RECT 43.245 202.325 43.910 202.495 ;
        RECT 44.195 202.470 44.365 203.270 ;
        RECT 44.575 203.125 44.805 203.945 ;
        RECT 44.975 203.145 45.305 203.775 ;
        RECT 44.555 202.705 44.885 202.955 ;
        RECT 45.055 202.545 45.305 203.145 ;
        RECT 45.475 203.125 45.685 203.945 ;
        RECT 46.005 203.395 46.175 203.775 ;
        RECT 46.355 203.565 46.685 203.945 ;
        RECT 46.005 203.225 46.670 203.395 ;
        RECT 46.865 203.270 47.125 203.775 ;
        RECT 45.935 202.675 46.265 203.045 ;
        RECT 46.500 202.970 46.670 203.225 ;
        RECT 43.245 201.565 43.415 202.325 ;
        RECT 43.595 201.395 43.925 202.155 ;
        RECT 44.095 201.565 44.365 202.470 ;
        RECT 44.575 201.395 44.805 202.535 ;
        RECT 44.975 201.565 45.305 202.545 ;
        RECT 46.500 202.640 46.785 202.970 ;
        RECT 45.475 201.395 45.685 202.535 ;
        RECT 46.500 202.495 46.670 202.640 ;
        RECT 46.005 202.325 46.670 202.495 ;
        RECT 46.955 202.470 47.125 203.270 ;
        RECT 47.385 203.395 47.555 203.775 ;
        RECT 47.735 203.565 48.065 203.945 ;
        RECT 47.385 203.225 48.050 203.395 ;
        RECT 48.245 203.270 48.505 203.775 ;
        RECT 47.315 202.675 47.645 203.045 ;
        RECT 47.880 202.970 48.050 203.225 ;
        RECT 47.880 202.640 48.165 202.970 ;
        RECT 47.880 202.495 48.050 202.640 ;
        RECT 46.005 201.565 46.175 202.325 ;
        RECT 46.355 201.395 46.685 202.155 ;
        RECT 46.855 201.565 47.125 202.470 ;
        RECT 47.385 202.325 48.050 202.495 ;
        RECT 48.335 202.470 48.505 203.270 ;
        RECT 48.675 203.220 48.965 203.945 ;
        RECT 50.095 203.125 50.325 203.945 ;
        RECT 50.495 203.145 50.825 203.775 ;
        RECT 50.075 202.705 50.405 202.955 ;
        RECT 47.385 201.565 47.555 202.325 ;
        RECT 47.735 201.395 48.065 202.155 ;
        RECT 48.235 201.565 48.505 202.470 ;
        RECT 48.675 201.395 48.965 202.560 ;
        RECT 50.575 202.545 50.825 203.145 ;
        RECT 50.995 203.125 51.205 203.945 ;
        RECT 51.495 203.125 51.705 203.945 ;
        RECT 51.875 203.145 52.205 203.775 ;
        RECT 50.095 201.395 50.325 202.535 ;
        RECT 50.495 201.565 50.825 202.545 ;
        RECT 51.875 202.545 52.125 203.145 ;
        RECT 52.375 203.125 52.605 203.945 ;
        RECT 53.365 203.395 53.535 203.775 ;
        RECT 53.715 203.565 54.045 203.945 ;
        RECT 53.365 203.225 54.030 203.395 ;
        RECT 54.225 203.270 54.485 203.775 ;
        RECT 52.295 202.705 52.625 202.955 ;
        RECT 53.295 202.675 53.625 203.045 ;
        RECT 53.860 202.970 54.030 203.225 ;
        RECT 53.860 202.640 54.145 202.970 ;
        RECT 50.995 201.395 51.205 202.535 ;
        RECT 51.495 201.395 51.705 202.535 ;
        RECT 51.875 201.565 52.205 202.545 ;
        RECT 52.375 201.395 52.605 202.535 ;
        RECT 53.860 202.495 54.030 202.640 ;
        RECT 53.365 202.325 54.030 202.495 ;
        RECT 54.315 202.470 54.485 203.270 ;
        RECT 54.745 203.395 54.915 203.775 ;
        RECT 55.095 203.565 55.425 203.945 ;
        RECT 54.745 203.225 55.410 203.395 ;
        RECT 55.605 203.270 55.865 203.775 ;
        RECT 54.675 202.675 55.005 203.045 ;
        RECT 55.240 202.970 55.410 203.225 ;
        RECT 55.240 202.640 55.525 202.970 ;
        RECT 55.240 202.495 55.410 202.640 ;
        RECT 53.365 201.565 53.535 202.325 ;
        RECT 53.715 201.395 54.045 202.155 ;
        RECT 54.215 201.565 54.485 202.470 ;
        RECT 54.745 202.325 55.410 202.495 ;
        RECT 55.695 202.470 55.865 203.270 ;
        RECT 56.035 203.145 56.345 203.945 ;
        RECT 56.550 203.145 57.245 203.775 ;
        RECT 56.045 202.705 56.380 202.975 ;
        RECT 56.550 202.545 56.720 203.145 ;
        RECT 57.475 203.125 57.685 203.945 ;
        RECT 57.855 203.145 58.185 203.775 ;
        RECT 56.890 202.705 57.225 202.955 ;
        RECT 57.855 202.545 58.105 203.145 ;
        RECT 58.355 203.125 58.585 203.945 ;
        RECT 58.835 203.125 59.065 203.945 ;
        RECT 59.235 203.145 59.565 203.775 ;
        RECT 58.275 202.705 58.605 202.955 ;
        RECT 58.815 202.705 59.145 202.955 ;
        RECT 59.315 202.545 59.565 203.145 ;
        RECT 59.735 203.125 59.945 203.945 ;
        RECT 60.175 203.270 60.435 203.775 ;
        RECT 60.615 203.565 60.945 203.945 ;
        RECT 61.125 203.395 61.295 203.775 ;
        RECT 54.745 201.565 54.915 202.325 ;
        RECT 55.095 201.395 55.425 202.155 ;
        RECT 55.595 201.565 55.865 202.470 ;
        RECT 56.035 201.395 56.315 202.535 ;
        RECT 56.485 201.565 56.815 202.545 ;
        RECT 56.985 201.395 57.245 202.535 ;
        RECT 57.475 201.395 57.685 202.535 ;
        RECT 57.855 201.565 58.185 202.545 ;
        RECT 58.355 201.395 58.585 202.535 ;
        RECT 58.835 201.395 59.065 202.535 ;
        RECT 59.235 201.565 59.565 202.545 ;
        RECT 59.735 201.395 59.945 202.535 ;
        RECT 60.175 202.470 60.345 203.270 ;
        RECT 60.630 203.225 61.295 203.395 ;
        RECT 60.630 202.970 60.800 203.225 ;
        RECT 61.555 203.220 61.845 203.945 ;
        RECT 62.020 203.545 62.355 203.945 ;
        RECT 62.525 203.375 62.730 203.775 ;
        RECT 62.940 203.465 63.215 203.945 ;
        RECT 63.425 203.445 63.685 203.775 ;
        RECT 62.045 203.205 62.730 203.375 ;
        RECT 60.515 202.640 60.800 202.970 ;
        RECT 61.035 202.675 61.365 203.045 ;
        RECT 60.630 202.495 60.800 202.640 ;
        RECT 60.175 201.565 60.445 202.470 ;
        RECT 60.630 202.325 61.295 202.495 ;
        RECT 60.615 201.395 60.945 202.155 ;
        RECT 61.125 201.565 61.295 202.325 ;
        RECT 61.555 201.395 61.845 202.560 ;
        RECT 62.045 202.175 62.385 203.205 ;
        RECT 62.555 202.535 62.805 203.035 ;
        RECT 62.985 202.705 63.345 203.285 ;
        RECT 63.515 202.535 63.685 203.445 ;
        RECT 63.855 203.125 64.115 203.945 ;
        RECT 64.285 203.125 64.615 203.545 ;
        RECT 64.795 203.375 65.055 203.775 ;
        RECT 65.225 203.545 65.555 203.945 ;
        RECT 65.725 203.375 65.895 203.725 ;
        RECT 66.065 203.545 66.440 203.945 ;
        RECT 64.795 203.205 66.460 203.375 ;
        RECT 66.630 203.270 66.905 203.615 ;
        RECT 64.365 203.035 64.615 203.125 ;
        RECT 66.290 203.035 66.460 203.205 ;
        RECT 63.860 202.705 64.195 202.955 ;
        RECT 64.365 202.705 65.080 203.035 ;
        RECT 65.295 202.705 66.120 203.035 ;
        RECT 66.290 202.705 66.565 203.035 ;
        RECT 62.555 202.365 63.685 202.535 ;
        RECT 62.045 202.000 62.710 202.175 ;
        RECT 62.020 201.395 62.355 201.820 ;
        RECT 62.525 201.595 62.710 202.000 ;
        RECT 62.915 201.395 63.245 202.175 ;
        RECT 63.415 201.595 63.685 202.365 ;
        RECT 63.855 201.395 64.115 202.535 ;
        RECT 64.365 202.145 64.535 202.705 ;
        RECT 64.795 202.245 65.125 202.535 ;
        RECT 65.295 202.415 65.540 202.705 ;
        RECT 66.290 202.535 66.460 202.705 ;
        RECT 66.735 202.535 66.905 203.270 ;
        RECT 65.800 202.365 66.460 202.535 ;
        RECT 65.800 202.245 65.970 202.365 ;
        RECT 64.795 202.075 65.970 202.245 ;
        RECT 64.355 201.575 65.970 201.905 ;
        RECT 66.140 201.395 66.420 202.195 ;
        RECT 66.630 201.565 66.905 202.535 ;
        RECT 67.085 203.220 67.415 203.730 ;
        RECT 67.585 203.545 67.915 203.945 ;
        RECT 68.965 203.375 69.295 203.715 ;
        RECT 69.465 203.545 69.795 203.945 ;
        RECT 67.085 202.455 67.275 203.220 ;
        RECT 67.585 203.205 69.950 203.375 ;
        RECT 67.585 203.035 67.755 203.205 ;
        RECT 67.445 202.705 67.755 203.035 ;
        RECT 67.925 202.705 68.230 203.035 ;
        RECT 67.085 201.605 67.415 202.455 ;
        RECT 67.585 201.395 67.835 202.535 ;
        RECT 68.015 202.375 68.230 202.705 ;
        RECT 68.405 202.375 68.690 203.035 ;
        RECT 68.885 202.375 69.150 203.035 ;
        RECT 69.365 202.375 69.610 203.035 ;
        RECT 69.780 202.205 69.950 203.205 ;
        RECT 68.025 202.035 69.315 202.205 ;
        RECT 68.025 201.615 68.275 202.035 ;
        RECT 68.505 201.395 68.835 201.865 ;
        RECT 69.065 201.615 69.315 202.035 ;
        RECT 69.495 202.035 69.950 202.205 ;
        RECT 70.755 203.205 71.140 203.775 ;
        RECT 71.310 203.485 71.635 203.945 ;
        RECT 72.155 203.315 72.435 203.775 ;
        RECT 70.755 202.535 71.035 203.205 ;
        RECT 71.310 203.145 72.435 203.315 ;
        RECT 71.310 203.035 71.760 203.145 ;
        RECT 71.205 202.705 71.760 203.035 ;
        RECT 72.625 202.975 73.025 203.775 ;
        RECT 73.425 203.485 73.695 203.945 ;
        RECT 73.865 203.315 74.150 203.775 ;
        RECT 69.495 201.605 69.825 202.035 ;
        RECT 70.755 201.565 71.140 202.535 ;
        RECT 71.310 202.245 71.760 202.705 ;
        RECT 71.930 202.415 73.025 202.975 ;
        RECT 71.310 202.025 72.435 202.245 ;
        RECT 71.310 201.395 71.635 201.855 ;
        RECT 72.155 201.565 72.435 202.025 ;
        RECT 72.625 201.565 73.025 202.415 ;
        RECT 73.195 203.145 74.150 203.315 ;
        RECT 74.435 203.220 74.725 203.945 ;
        RECT 74.895 203.445 75.155 203.775 ;
        RECT 75.365 203.465 75.640 203.945 ;
        RECT 73.195 202.245 73.405 203.145 ;
        RECT 73.575 202.415 74.265 202.975 ;
        RECT 73.195 202.025 74.150 202.245 ;
        RECT 73.425 201.395 73.695 201.855 ;
        RECT 73.865 201.565 74.150 202.025 ;
        RECT 74.435 201.395 74.725 202.560 ;
        RECT 74.895 202.535 75.065 203.445 ;
        RECT 75.850 203.375 76.055 203.775 ;
        RECT 76.225 203.545 76.560 203.945 ;
        RECT 75.235 202.705 75.595 203.285 ;
        RECT 75.850 203.205 76.535 203.375 ;
        RECT 75.775 202.535 76.025 203.035 ;
        RECT 74.895 202.365 76.025 202.535 ;
        RECT 74.895 201.595 75.165 202.365 ;
        RECT 76.195 202.175 76.535 203.205 ;
        RECT 75.335 201.395 75.665 202.175 ;
        RECT 75.870 202.000 76.535 202.175 ;
        RECT 76.740 203.235 76.995 203.765 ;
        RECT 77.165 203.485 77.470 203.945 ;
        RECT 77.715 203.565 78.785 203.735 ;
        RECT 76.740 202.585 76.950 203.235 ;
        RECT 77.715 203.210 78.035 203.565 ;
        RECT 77.710 203.035 78.035 203.210 ;
        RECT 77.120 202.735 78.035 203.035 ;
        RECT 78.205 202.995 78.445 203.395 ;
        RECT 78.615 203.335 78.785 203.565 ;
        RECT 78.955 203.505 79.145 203.945 ;
        RECT 79.315 203.495 80.265 203.775 ;
        RECT 80.485 203.585 80.835 203.755 ;
        RECT 78.615 203.165 79.145 203.335 ;
        RECT 77.120 202.705 77.860 202.735 ;
        RECT 75.870 201.595 76.055 202.000 ;
        RECT 76.225 201.395 76.560 201.820 ;
        RECT 76.740 201.705 76.995 202.585 ;
        RECT 77.165 201.395 77.470 202.535 ;
        RECT 77.690 202.115 77.860 202.705 ;
        RECT 78.205 202.625 78.745 202.995 ;
        RECT 78.925 202.885 79.145 203.165 ;
        RECT 79.315 202.715 79.485 203.495 ;
        RECT 79.080 202.545 79.485 202.715 ;
        RECT 79.655 202.705 80.005 203.325 ;
        RECT 79.080 202.455 79.250 202.545 ;
        RECT 80.175 202.535 80.385 203.325 ;
        RECT 78.030 202.285 79.250 202.455 ;
        RECT 79.710 202.375 80.385 202.535 ;
        RECT 77.690 201.945 78.490 202.115 ;
        RECT 77.810 201.395 78.140 201.775 ;
        RECT 78.320 201.655 78.490 201.945 ;
        RECT 79.080 201.905 79.250 202.285 ;
        RECT 79.420 202.365 80.385 202.375 ;
        RECT 80.575 203.195 80.835 203.585 ;
        RECT 81.045 203.485 81.375 203.945 ;
        RECT 82.250 203.555 83.105 203.725 ;
        RECT 83.310 203.555 83.805 203.725 ;
        RECT 83.975 203.585 84.305 203.945 ;
        RECT 80.575 202.505 80.745 203.195 ;
        RECT 80.915 202.845 81.085 203.025 ;
        RECT 81.255 203.015 82.045 203.265 ;
        RECT 82.250 202.845 82.420 203.555 ;
        RECT 82.590 203.045 82.945 203.265 ;
        RECT 80.915 202.675 82.605 202.845 ;
        RECT 79.420 202.075 79.880 202.365 ;
        RECT 80.575 202.335 82.075 202.505 ;
        RECT 80.575 202.195 80.745 202.335 ;
        RECT 80.185 202.025 80.745 202.195 ;
        RECT 78.660 201.395 78.910 201.855 ;
        RECT 79.080 201.565 79.950 201.905 ;
        RECT 80.185 201.565 80.355 202.025 ;
        RECT 81.190 201.995 82.265 202.165 ;
        RECT 80.525 201.395 80.895 201.855 ;
        RECT 81.190 201.655 81.360 201.995 ;
        RECT 81.530 201.395 81.860 201.825 ;
        RECT 82.095 201.655 82.265 201.995 ;
        RECT 82.435 201.895 82.605 202.675 ;
        RECT 82.775 202.455 82.945 203.045 ;
        RECT 83.115 202.645 83.465 203.265 ;
        RECT 82.775 202.065 83.240 202.455 ;
        RECT 83.635 202.195 83.805 203.555 ;
        RECT 83.975 202.365 84.435 203.415 ;
        RECT 83.410 202.025 83.805 202.195 ;
        RECT 83.410 201.895 83.580 202.025 ;
        RECT 82.435 201.565 83.115 201.895 ;
        RECT 83.330 201.565 83.580 201.895 ;
        RECT 83.750 201.395 84.000 201.855 ;
        RECT 84.170 201.580 84.495 202.365 ;
        RECT 84.665 201.565 84.835 203.685 ;
        RECT 85.005 203.565 85.335 203.945 ;
        RECT 85.505 203.395 85.760 203.685 ;
        RECT 85.010 203.225 85.760 203.395 ;
        RECT 85.010 202.235 85.240 203.225 ;
        RECT 85.995 203.125 86.205 203.945 ;
        RECT 86.375 203.145 86.705 203.775 ;
        RECT 85.410 202.405 85.760 203.055 ;
        RECT 86.375 202.545 86.625 203.145 ;
        RECT 86.875 203.125 87.105 203.945 ;
        RECT 87.315 203.220 87.605 203.945 ;
        RECT 88.810 203.315 89.095 203.775 ;
        RECT 89.265 203.485 89.535 203.945 ;
        RECT 88.810 203.145 89.765 203.315 ;
        RECT 86.795 202.705 87.125 202.955 ;
        RECT 85.010 202.065 85.760 202.235 ;
        RECT 85.005 201.395 85.335 201.895 ;
        RECT 85.505 201.565 85.760 202.065 ;
        RECT 85.995 201.395 86.205 202.535 ;
        RECT 86.375 201.565 86.705 202.545 ;
        RECT 86.875 201.395 87.105 202.535 ;
        RECT 87.315 201.395 87.605 202.560 ;
        RECT 88.695 202.415 89.385 202.975 ;
        RECT 89.555 202.245 89.765 203.145 ;
        RECT 88.810 202.025 89.765 202.245 ;
        RECT 89.935 202.975 90.335 203.775 ;
        RECT 90.525 203.315 90.805 203.775 ;
        RECT 91.325 203.485 91.650 203.945 ;
        RECT 90.525 203.145 91.650 203.315 ;
        RECT 91.820 203.205 92.205 203.775 ;
        RECT 91.200 203.035 91.650 203.145 ;
        RECT 89.935 202.415 91.030 202.975 ;
        RECT 91.200 202.705 91.755 203.035 ;
        RECT 88.810 201.565 89.095 202.025 ;
        RECT 89.265 201.395 89.535 201.855 ;
        RECT 89.935 201.565 90.335 202.415 ;
        RECT 91.200 202.245 91.650 202.705 ;
        RECT 91.925 202.535 92.205 203.205 ;
        RECT 90.525 202.025 91.650 202.245 ;
        RECT 90.525 201.565 90.805 202.025 ;
        RECT 91.325 201.395 91.650 201.855 ;
        RECT 91.820 201.565 92.205 202.535 ;
        RECT 92.375 203.205 92.760 203.775 ;
        RECT 92.930 203.485 93.255 203.945 ;
        RECT 93.775 203.315 94.055 203.775 ;
        RECT 92.375 202.535 92.655 203.205 ;
        RECT 92.930 203.145 94.055 203.315 ;
        RECT 92.930 203.035 93.380 203.145 ;
        RECT 92.825 202.705 93.380 203.035 ;
        RECT 94.245 202.975 94.645 203.775 ;
        RECT 95.045 203.485 95.315 203.945 ;
        RECT 95.485 203.315 95.770 203.775 ;
        RECT 92.375 201.565 92.760 202.535 ;
        RECT 92.930 202.245 93.380 202.705 ;
        RECT 93.550 202.415 94.645 202.975 ;
        RECT 92.930 202.025 94.055 202.245 ;
        RECT 92.930 201.395 93.255 201.855 ;
        RECT 93.775 201.565 94.055 202.025 ;
        RECT 94.245 201.565 94.645 202.415 ;
        RECT 94.815 203.145 95.770 203.315 ;
        RECT 96.060 203.205 96.315 203.775 ;
        RECT 96.485 203.545 96.815 203.945 ;
        RECT 97.240 203.410 97.770 203.775 ;
        RECT 97.240 203.375 97.415 203.410 ;
        RECT 96.485 203.205 97.415 203.375 ;
        RECT 94.815 202.245 95.025 203.145 ;
        RECT 95.195 202.415 95.885 202.975 ;
        RECT 96.060 202.535 96.230 203.205 ;
        RECT 96.485 203.035 96.655 203.205 ;
        RECT 96.400 202.705 96.655 203.035 ;
        RECT 96.880 202.705 97.075 203.035 ;
        RECT 94.815 202.025 95.770 202.245 ;
        RECT 95.045 201.395 95.315 201.855 ;
        RECT 95.485 201.565 95.770 202.025 ;
        RECT 96.060 201.565 96.395 202.535 ;
        RECT 96.565 201.395 96.735 202.535 ;
        RECT 96.905 201.735 97.075 202.705 ;
        RECT 97.245 202.075 97.415 203.205 ;
        RECT 97.585 202.415 97.755 203.215 ;
        RECT 97.960 202.925 98.235 203.775 ;
        RECT 97.955 202.755 98.235 202.925 ;
        RECT 97.960 202.615 98.235 202.755 ;
        RECT 98.405 202.415 98.595 203.775 ;
        RECT 98.775 203.410 99.285 203.945 ;
        RECT 99.505 203.135 99.750 203.740 ;
        RECT 100.195 203.220 100.485 203.945 ;
        RECT 100.660 203.235 100.915 203.765 ;
        RECT 101.085 203.485 101.390 203.945 ;
        RECT 101.635 203.565 102.705 203.735 ;
        RECT 98.795 202.965 100.025 203.135 ;
        RECT 97.585 202.245 98.595 202.415 ;
        RECT 98.765 202.400 99.515 202.590 ;
        RECT 97.245 201.905 98.370 202.075 ;
        RECT 98.765 201.735 98.935 202.400 ;
        RECT 99.685 202.155 100.025 202.965 ;
        RECT 100.660 202.585 100.870 203.235 ;
        RECT 101.635 203.210 101.955 203.565 ;
        RECT 101.630 203.035 101.955 203.210 ;
        RECT 101.040 202.735 101.955 203.035 ;
        RECT 102.125 202.995 102.365 203.395 ;
        RECT 102.535 203.335 102.705 203.565 ;
        RECT 102.875 203.505 103.065 203.945 ;
        RECT 103.235 203.495 104.185 203.775 ;
        RECT 104.405 203.585 104.755 203.755 ;
        RECT 102.535 203.165 103.065 203.335 ;
        RECT 101.040 202.705 101.780 202.735 ;
        RECT 96.905 201.565 98.935 201.735 ;
        RECT 99.105 201.395 99.275 202.155 ;
        RECT 99.510 201.745 100.025 202.155 ;
        RECT 100.195 201.395 100.485 202.560 ;
        RECT 100.660 201.705 100.915 202.585 ;
        RECT 101.085 201.395 101.390 202.535 ;
        RECT 101.610 202.115 101.780 202.705 ;
        RECT 102.125 202.625 102.665 202.995 ;
        RECT 102.845 202.885 103.065 203.165 ;
        RECT 103.235 202.715 103.405 203.495 ;
        RECT 103.000 202.545 103.405 202.715 ;
        RECT 103.575 202.705 103.925 203.325 ;
        RECT 103.000 202.455 103.170 202.545 ;
        RECT 104.095 202.535 104.305 203.325 ;
        RECT 101.950 202.285 103.170 202.455 ;
        RECT 103.630 202.375 104.305 202.535 ;
        RECT 101.610 201.945 102.410 202.115 ;
        RECT 101.730 201.395 102.060 201.775 ;
        RECT 102.240 201.655 102.410 201.945 ;
        RECT 103.000 201.905 103.170 202.285 ;
        RECT 103.340 202.365 104.305 202.375 ;
        RECT 104.495 203.195 104.755 203.585 ;
        RECT 104.965 203.485 105.295 203.945 ;
        RECT 106.170 203.555 107.025 203.725 ;
        RECT 107.230 203.555 107.725 203.725 ;
        RECT 107.895 203.585 108.225 203.945 ;
        RECT 104.495 202.505 104.665 203.195 ;
        RECT 104.835 202.845 105.005 203.025 ;
        RECT 105.175 203.015 105.965 203.265 ;
        RECT 106.170 202.845 106.340 203.555 ;
        RECT 106.510 203.045 106.865 203.265 ;
        RECT 104.835 202.675 106.525 202.845 ;
        RECT 103.340 202.075 103.800 202.365 ;
        RECT 104.495 202.335 105.995 202.505 ;
        RECT 104.495 202.195 104.665 202.335 ;
        RECT 104.105 202.025 104.665 202.195 ;
        RECT 102.580 201.395 102.830 201.855 ;
        RECT 103.000 201.565 103.870 201.905 ;
        RECT 104.105 201.565 104.275 202.025 ;
        RECT 105.110 201.995 106.185 202.165 ;
        RECT 104.445 201.395 104.815 201.855 ;
        RECT 105.110 201.655 105.280 201.995 ;
        RECT 105.450 201.395 105.780 201.825 ;
        RECT 106.015 201.655 106.185 201.995 ;
        RECT 106.355 201.895 106.525 202.675 ;
        RECT 106.695 202.455 106.865 203.045 ;
        RECT 107.035 202.645 107.385 203.265 ;
        RECT 106.695 202.065 107.160 202.455 ;
        RECT 107.555 202.195 107.725 203.555 ;
        RECT 107.895 202.365 108.355 203.415 ;
        RECT 107.330 202.025 107.725 202.195 ;
        RECT 107.330 201.895 107.500 202.025 ;
        RECT 106.355 201.565 107.035 201.895 ;
        RECT 107.250 201.565 107.500 201.895 ;
        RECT 107.670 201.395 107.920 201.855 ;
        RECT 108.090 201.580 108.415 202.365 ;
        RECT 108.585 201.565 108.755 203.685 ;
        RECT 108.925 203.565 109.255 203.945 ;
        RECT 109.425 203.395 109.680 203.685 ;
        RECT 108.930 203.225 109.680 203.395 ;
        RECT 108.930 202.235 109.160 203.225 ;
        RECT 109.895 203.125 110.125 203.945 ;
        RECT 110.295 203.145 110.625 203.775 ;
        RECT 109.330 202.405 109.680 203.055 ;
        RECT 109.875 202.705 110.205 202.955 ;
        RECT 110.375 202.545 110.625 203.145 ;
        RECT 110.795 203.125 111.005 203.945 ;
        RECT 112.155 203.195 113.365 203.945 ;
        RECT 108.930 202.065 109.680 202.235 ;
        RECT 108.925 201.395 109.255 201.895 ;
        RECT 109.425 201.565 109.680 202.065 ;
        RECT 109.895 201.395 110.125 202.535 ;
        RECT 110.295 201.565 110.625 202.545 ;
        RECT 110.795 201.395 111.005 202.535 ;
        RECT 112.155 202.485 112.675 203.025 ;
        RECT 112.845 202.655 113.365 203.195 ;
        RECT 112.155 201.395 113.365 202.485 ;
        RECT 26.970 201.225 113.450 201.395 ;
        RECT 27.055 200.135 28.265 201.225 ;
        RECT 27.055 199.425 27.575 199.965 ;
        RECT 27.745 199.595 28.265 200.135 ;
        RECT 28.985 200.295 29.155 201.055 ;
        RECT 29.335 200.465 29.665 201.225 ;
        RECT 28.985 200.125 29.650 200.295 ;
        RECT 29.835 200.150 30.105 201.055 ;
        RECT 29.480 199.980 29.650 200.125 ;
        RECT 28.915 199.575 29.245 199.945 ;
        RECT 29.480 199.650 29.765 199.980 ;
        RECT 27.055 198.675 28.265 199.425 ;
        RECT 29.480 199.395 29.650 199.650 ;
        RECT 28.985 199.225 29.650 199.395 ;
        RECT 29.935 199.350 30.105 200.150 ;
        RECT 30.315 200.085 30.545 201.225 ;
        RECT 30.715 200.075 31.045 201.055 ;
        RECT 31.215 200.085 31.425 201.225 ;
        RECT 31.695 200.085 31.925 201.225 ;
        RECT 32.095 200.075 32.425 201.055 ;
        RECT 32.595 200.085 32.805 201.225 ;
        RECT 33.095 200.085 33.305 201.225 ;
        RECT 30.295 199.665 30.625 199.915 ;
        RECT 28.985 198.845 29.155 199.225 ;
        RECT 29.335 198.675 29.665 199.055 ;
        RECT 29.845 198.845 30.105 199.350 ;
        RECT 30.315 198.675 30.545 199.495 ;
        RECT 30.795 199.475 31.045 200.075 ;
        RECT 31.675 199.665 32.005 199.915 ;
        RECT 30.715 198.845 31.045 199.475 ;
        RECT 31.215 198.675 31.425 199.495 ;
        RECT 31.695 198.675 31.925 199.495 ;
        RECT 32.175 199.475 32.425 200.075 ;
        RECT 33.475 200.075 33.805 201.055 ;
        RECT 33.975 200.085 34.205 201.225 ;
        RECT 34.505 200.295 34.675 201.055 ;
        RECT 34.855 200.465 35.185 201.225 ;
        RECT 34.505 200.125 35.170 200.295 ;
        RECT 35.355 200.150 35.625 201.055 ;
        RECT 32.095 198.845 32.425 199.475 ;
        RECT 32.595 198.675 32.805 199.495 ;
        RECT 33.095 198.675 33.305 199.495 ;
        RECT 33.475 199.475 33.725 200.075 ;
        RECT 35.000 199.980 35.170 200.125 ;
        RECT 33.895 199.665 34.225 199.915 ;
        RECT 34.435 199.575 34.765 199.945 ;
        RECT 35.000 199.650 35.285 199.980 ;
        RECT 33.475 198.845 33.805 199.475 ;
        RECT 33.975 198.675 34.205 199.495 ;
        RECT 35.000 199.395 35.170 199.650 ;
        RECT 34.505 199.225 35.170 199.395 ;
        RECT 35.455 199.350 35.625 200.150 ;
        RECT 35.795 200.060 36.085 201.225 ;
        RECT 36.805 200.295 36.975 201.055 ;
        RECT 37.155 200.465 37.485 201.225 ;
        RECT 36.805 200.125 37.470 200.295 ;
        RECT 37.655 200.150 37.925 201.055 ;
        RECT 37.300 199.980 37.470 200.125 ;
        RECT 36.735 199.575 37.065 199.945 ;
        RECT 37.300 199.650 37.585 199.980 ;
        RECT 34.505 198.845 34.675 199.225 ;
        RECT 34.855 198.675 35.185 199.055 ;
        RECT 35.365 198.845 35.625 199.350 ;
        RECT 35.795 198.675 36.085 199.400 ;
        RECT 37.300 199.395 37.470 199.650 ;
        RECT 36.805 199.225 37.470 199.395 ;
        RECT 37.755 199.350 37.925 200.150 ;
        RECT 38.185 200.295 38.355 201.055 ;
        RECT 38.535 200.465 38.865 201.225 ;
        RECT 38.185 200.125 38.850 200.295 ;
        RECT 39.035 200.150 39.305 201.055 ;
        RECT 38.680 199.980 38.850 200.125 ;
        RECT 38.115 199.575 38.445 199.945 ;
        RECT 38.680 199.650 38.965 199.980 ;
        RECT 38.680 199.395 38.850 199.650 ;
        RECT 36.805 198.845 36.975 199.225 ;
        RECT 37.155 198.675 37.485 199.055 ;
        RECT 37.665 198.845 37.925 199.350 ;
        RECT 38.185 199.225 38.850 199.395 ;
        RECT 39.135 199.350 39.305 200.150 ;
        RECT 38.185 198.845 38.355 199.225 ;
        RECT 38.535 198.675 38.865 199.055 ;
        RECT 39.045 198.845 39.305 199.350 ;
        RECT 39.475 200.085 39.815 201.055 ;
        RECT 39.985 200.085 40.155 201.225 ;
        RECT 40.425 200.425 40.675 201.225 ;
        RECT 41.320 200.255 41.650 201.055 ;
        RECT 41.950 200.425 42.280 201.225 ;
        RECT 42.450 200.255 42.780 201.055 ;
        RECT 40.345 200.085 42.780 200.255 ;
        RECT 43.215 200.085 43.425 201.225 ;
        RECT 39.475 199.475 39.650 200.085 ;
        RECT 40.345 199.835 40.515 200.085 ;
        RECT 39.820 199.665 40.515 199.835 ;
        RECT 40.690 199.665 41.110 199.865 ;
        RECT 41.280 199.665 41.610 199.865 ;
        RECT 41.780 199.665 42.110 199.865 ;
        RECT 39.475 198.845 39.815 199.475 ;
        RECT 39.985 198.675 40.235 199.475 ;
        RECT 40.425 199.325 41.650 199.495 ;
        RECT 40.425 198.845 40.755 199.325 ;
        RECT 40.925 198.675 41.150 199.135 ;
        RECT 41.320 198.845 41.650 199.325 ;
        RECT 42.280 199.455 42.450 200.085 ;
        RECT 43.595 200.075 43.925 201.055 ;
        RECT 44.095 200.085 44.325 201.225 ;
        RECT 44.595 200.085 44.805 201.225 ;
        RECT 44.975 200.075 45.305 201.055 ;
        RECT 45.475 200.085 45.705 201.225 ;
        RECT 46.005 200.295 46.175 201.055 ;
        RECT 46.355 200.465 46.685 201.225 ;
        RECT 46.005 200.125 46.670 200.295 ;
        RECT 46.855 200.150 47.125 201.055 ;
        RECT 42.635 199.665 42.985 199.915 ;
        RECT 42.280 198.845 42.780 199.455 ;
        RECT 43.215 198.675 43.425 199.495 ;
        RECT 43.595 199.475 43.845 200.075 ;
        RECT 44.015 199.665 44.345 199.915 ;
        RECT 43.595 198.845 43.925 199.475 ;
        RECT 44.095 198.675 44.325 199.495 ;
        RECT 44.595 198.675 44.805 199.495 ;
        RECT 44.975 199.475 45.225 200.075 ;
        RECT 46.500 199.980 46.670 200.125 ;
        RECT 45.395 199.665 45.725 199.915 ;
        RECT 45.935 199.575 46.265 199.945 ;
        RECT 46.500 199.650 46.785 199.980 ;
        RECT 44.975 198.845 45.305 199.475 ;
        RECT 45.475 198.675 45.705 199.495 ;
        RECT 46.500 199.395 46.670 199.650 ;
        RECT 46.005 199.225 46.670 199.395 ;
        RECT 46.955 199.350 47.125 200.150 ;
        RECT 47.335 200.085 47.565 201.225 ;
        RECT 47.735 200.075 48.065 201.055 ;
        RECT 48.235 200.085 48.445 201.225 ;
        RECT 48.675 200.085 49.060 201.055 ;
        RECT 49.230 200.765 49.555 201.225 ;
        RECT 50.075 200.595 50.355 201.055 ;
        RECT 49.230 200.375 50.355 200.595 ;
        RECT 47.315 199.665 47.645 199.915 ;
        RECT 46.005 198.845 46.175 199.225 ;
        RECT 46.355 198.675 46.685 199.055 ;
        RECT 46.865 198.845 47.125 199.350 ;
        RECT 47.335 198.675 47.565 199.495 ;
        RECT 47.815 199.475 48.065 200.075 ;
        RECT 47.735 198.845 48.065 199.475 ;
        RECT 48.235 198.675 48.445 199.495 ;
        RECT 48.675 199.415 48.955 200.085 ;
        RECT 49.230 199.915 49.680 200.375 ;
        RECT 50.545 200.205 50.945 201.055 ;
        RECT 51.345 200.765 51.615 201.225 ;
        RECT 51.785 200.595 52.070 201.055 ;
        RECT 49.125 199.585 49.680 199.915 ;
        RECT 49.850 199.645 50.945 200.205 ;
        RECT 49.230 199.475 49.680 199.585 ;
        RECT 48.675 198.845 49.060 199.415 ;
        RECT 49.230 199.305 50.355 199.475 ;
        RECT 49.230 198.675 49.555 199.135 ;
        RECT 50.075 198.845 50.355 199.305 ;
        RECT 50.545 198.845 50.945 199.645 ;
        RECT 51.115 200.375 52.070 200.595 ;
        RECT 52.360 200.555 52.615 201.055 ;
        RECT 52.785 200.725 53.115 201.225 ;
        RECT 52.360 200.385 53.110 200.555 ;
        RECT 51.115 199.475 51.325 200.375 ;
        RECT 51.495 199.645 52.185 200.205 ;
        RECT 52.360 199.565 52.710 200.215 ;
        RECT 51.115 199.305 52.070 199.475 ;
        RECT 52.880 199.395 53.110 200.385 ;
        RECT 51.345 198.675 51.615 199.135 ;
        RECT 51.785 198.845 52.070 199.305 ;
        RECT 52.360 199.225 53.110 199.395 ;
        RECT 52.360 198.935 52.615 199.225 ;
        RECT 52.785 198.675 53.115 199.055 ;
        RECT 53.285 198.935 53.455 201.055 ;
        RECT 53.625 200.255 53.950 201.040 ;
        RECT 54.120 200.765 54.370 201.225 ;
        RECT 54.540 200.725 54.790 201.055 ;
        RECT 55.005 200.725 55.685 201.055 ;
        RECT 54.540 200.595 54.710 200.725 ;
        RECT 54.315 200.425 54.710 200.595 ;
        RECT 53.685 199.205 54.145 200.255 ;
        RECT 54.315 199.065 54.485 200.425 ;
        RECT 54.880 200.165 55.345 200.555 ;
        RECT 54.655 199.355 55.005 199.975 ;
        RECT 55.175 199.575 55.345 200.165 ;
        RECT 55.515 199.945 55.685 200.725 ;
        RECT 55.855 200.625 56.025 200.965 ;
        RECT 56.260 200.795 56.590 201.225 ;
        RECT 56.760 200.625 56.930 200.965 ;
        RECT 57.225 200.765 57.595 201.225 ;
        RECT 55.855 200.455 56.930 200.625 ;
        RECT 57.765 200.595 57.935 201.055 ;
        RECT 58.170 200.715 59.040 201.055 ;
        RECT 59.210 200.765 59.460 201.225 ;
        RECT 57.375 200.425 57.935 200.595 ;
        RECT 57.375 200.285 57.545 200.425 ;
        RECT 56.045 200.115 57.545 200.285 ;
        RECT 58.240 200.255 58.700 200.545 ;
        RECT 55.515 199.775 57.205 199.945 ;
        RECT 55.175 199.355 55.530 199.575 ;
        RECT 55.700 199.065 55.870 199.775 ;
        RECT 56.075 199.355 56.865 199.605 ;
        RECT 57.035 199.595 57.205 199.775 ;
        RECT 57.375 199.425 57.545 200.115 ;
        RECT 53.815 198.675 54.145 199.035 ;
        RECT 54.315 198.895 54.810 199.065 ;
        RECT 55.015 198.895 55.870 199.065 ;
        RECT 56.745 198.675 57.075 199.135 ;
        RECT 57.285 199.035 57.545 199.425 ;
        RECT 57.735 200.245 58.700 200.255 ;
        RECT 58.870 200.335 59.040 200.715 ;
        RECT 59.630 200.675 59.800 200.965 ;
        RECT 59.980 200.845 60.310 201.225 ;
        RECT 59.630 200.505 60.430 200.675 ;
        RECT 57.735 200.085 58.410 200.245 ;
        RECT 58.870 200.165 60.090 200.335 ;
        RECT 57.735 199.295 57.945 200.085 ;
        RECT 58.870 200.075 59.040 200.165 ;
        RECT 58.115 199.295 58.465 199.915 ;
        RECT 58.635 199.905 59.040 200.075 ;
        RECT 58.635 199.125 58.805 199.905 ;
        RECT 58.975 199.455 59.195 199.735 ;
        RECT 59.375 199.625 59.915 199.995 ;
        RECT 60.260 199.915 60.430 200.505 ;
        RECT 60.650 200.085 60.955 201.225 ;
        RECT 61.125 200.035 61.380 200.915 ;
        RECT 61.555 200.060 61.845 201.225 ;
        RECT 62.130 200.595 62.415 201.055 ;
        RECT 62.585 200.765 62.855 201.225 ;
        RECT 62.130 200.375 63.085 200.595 ;
        RECT 60.260 199.885 61.000 199.915 ;
        RECT 58.975 199.285 59.505 199.455 ;
        RECT 57.285 198.865 57.635 199.035 ;
        RECT 57.855 198.845 58.805 199.125 ;
        RECT 58.975 198.675 59.165 199.115 ;
        RECT 59.335 199.055 59.505 199.285 ;
        RECT 59.675 199.225 59.915 199.625 ;
        RECT 60.085 199.585 61.000 199.885 ;
        RECT 60.085 199.410 60.410 199.585 ;
        RECT 60.085 199.055 60.405 199.410 ;
        RECT 61.170 199.385 61.380 200.035 ;
        RECT 62.015 199.645 62.705 200.205 ;
        RECT 62.875 199.475 63.085 200.375 ;
        RECT 59.335 198.885 60.405 199.055 ;
        RECT 60.650 198.675 60.955 199.135 ;
        RECT 61.125 198.855 61.380 199.385 ;
        RECT 61.555 198.675 61.845 199.400 ;
        RECT 62.130 199.305 63.085 199.475 ;
        RECT 63.255 200.205 63.655 201.055 ;
        RECT 63.845 200.595 64.125 201.055 ;
        RECT 64.645 200.765 64.970 201.225 ;
        RECT 63.845 200.375 64.970 200.595 ;
        RECT 63.255 199.645 64.350 200.205 ;
        RECT 64.520 199.915 64.970 200.375 ;
        RECT 65.140 200.085 65.525 201.055 ;
        RECT 65.715 200.715 66.015 201.225 ;
        RECT 66.185 200.715 66.565 200.885 ;
        RECT 67.145 200.715 67.775 201.225 ;
        RECT 66.185 200.545 66.355 200.715 ;
        RECT 67.945 200.545 68.275 201.055 ;
        RECT 68.445 200.715 68.745 201.225 ;
        RECT 62.130 198.845 62.415 199.305 ;
        RECT 62.585 198.675 62.855 199.135 ;
        RECT 63.255 198.845 63.655 199.645 ;
        RECT 64.520 199.585 65.075 199.915 ;
        RECT 64.520 199.475 64.970 199.585 ;
        RECT 63.845 199.305 64.970 199.475 ;
        RECT 65.245 199.415 65.525 200.085 ;
        RECT 63.845 198.845 64.125 199.305 ;
        RECT 64.645 198.675 64.970 199.135 ;
        RECT 65.140 198.845 65.525 199.415 ;
        RECT 65.695 200.345 66.355 200.545 ;
        RECT 66.525 200.375 68.745 200.545 ;
        RECT 65.695 199.415 65.865 200.345 ;
        RECT 66.525 200.175 66.695 200.375 ;
        RECT 66.035 200.005 66.695 200.175 ;
        RECT 66.865 200.035 68.405 200.205 ;
        RECT 66.035 199.585 66.205 200.005 ;
        RECT 66.865 199.835 67.035 200.035 ;
        RECT 66.435 199.665 67.035 199.835 ;
        RECT 67.205 199.665 67.900 199.865 ;
        RECT 68.160 199.585 68.405 200.035 ;
        RECT 66.525 199.415 67.435 199.495 ;
        RECT 65.695 198.935 66.015 199.415 ;
        RECT 66.185 199.325 67.435 199.415 ;
        RECT 66.185 199.245 66.695 199.325 ;
        RECT 66.185 198.845 66.415 199.245 ;
        RECT 66.585 198.675 66.935 199.065 ;
        RECT 67.105 198.845 67.435 199.325 ;
        RECT 67.605 198.675 67.775 199.495 ;
        RECT 68.575 199.415 68.745 200.375 ;
        RECT 69.005 200.295 69.175 201.055 ;
        RECT 69.390 200.465 69.720 201.225 ;
        RECT 69.005 200.125 69.720 200.295 ;
        RECT 69.890 200.150 70.145 201.055 ;
        RECT 68.915 199.575 69.270 199.945 ;
        RECT 69.550 199.915 69.720 200.125 ;
        RECT 69.550 199.585 69.805 199.915 ;
        RECT 68.280 198.870 68.745 199.415 ;
        RECT 69.550 199.395 69.720 199.585 ;
        RECT 69.975 199.420 70.145 200.150 ;
        RECT 70.320 200.075 70.580 201.225 ;
        RECT 70.760 200.555 71.015 201.055 ;
        RECT 71.185 200.725 71.515 201.225 ;
        RECT 70.760 200.385 71.510 200.555 ;
        RECT 70.760 199.565 71.110 200.215 ;
        RECT 69.005 199.225 69.720 199.395 ;
        RECT 69.005 198.845 69.175 199.225 ;
        RECT 69.390 198.675 69.720 199.055 ;
        RECT 69.890 198.845 70.145 199.420 ;
        RECT 70.320 198.675 70.580 199.515 ;
        RECT 71.280 199.395 71.510 200.385 ;
        RECT 70.760 199.225 71.510 199.395 ;
        RECT 70.760 198.935 71.015 199.225 ;
        RECT 71.185 198.675 71.515 199.055 ;
        RECT 71.685 198.935 71.855 201.055 ;
        RECT 72.025 200.255 72.350 201.040 ;
        RECT 72.520 200.765 72.770 201.225 ;
        RECT 72.940 200.725 73.190 201.055 ;
        RECT 73.405 200.725 74.085 201.055 ;
        RECT 72.940 200.595 73.110 200.725 ;
        RECT 72.715 200.425 73.110 200.595 ;
        RECT 72.085 199.205 72.545 200.255 ;
        RECT 72.715 199.065 72.885 200.425 ;
        RECT 73.280 200.165 73.745 200.555 ;
        RECT 73.055 199.355 73.405 199.975 ;
        RECT 73.575 199.575 73.745 200.165 ;
        RECT 73.915 199.945 74.085 200.725 ;
        RECT 74.255 200.625 74.425 200.965 ;
        RECT 74.660 200.795 74.990 201.225 ;
        RECT 75.160 200.625 75.330 200.965 ;
        RECT 75.625 200.765 75.995 201.225 ;
        RECT 74.255 200.455 75.330 200.625 ;
        RECT 76.165 200.595 76.335 201.055 ;
        RECT 76.570 200.715 77.440 201.055 ;
        RECT 77.610 200.765 77.860 201.225 ;
        RECT 75.775 200.425 76.335 200.595 ;
        RECT 75.775 200.285 75.945 200.425 ;
        RECT 74.445 200.115 75.945 200.285 ;
        RECT 76.640 200.255 77.100 200.545 ;
        RECT 73.915 199.775 75.605 199.945 ;
        RECT 73.575 199.355 73.930 199.575 ;
        RECT 74.100 199.065 74.270 199.775 ;
        RECT 74.475 199.355 75.265 199.605 ;
        RECT 75.435 199.595 75.605 199.775 ;
        RECT 75.775 199.425 75.945 200.115 ;
        RECT 72.215 198.675 72.545 199.035 ;
        RECT 72.715 198.895 73.210 199.065 ;
        RECT 73.415 198.895 74.270 199.065 ;
        RECT 75.145 198.675 75.475 199.135 ;
        RECT 75.685 199.035 75.945 199.425 ;
        RECT 76.135 200.245 77.100 200.255 ;
        RECT 77.270 200.335 77.440 200.715 ;
        RECT 78.030 200.675 78.200 200.965 ;
        RECT 78.380 200.845 78.710 201.225 ;
        RECT 78.030 200.505 78.830 200.675 ;
        RECT 76.135 200.085 76.810 200.245 ;
        RECT 77.270 200.165 78.490 200.335 ;
        RECT 76.135 199.295 76.345 200.085 ;
        RECT 77.270 200.075 77.440 200.165 ;
        RECT 76.515 199.295 76.865 199.915 ;
        RECT 77.035 199.905 77.440 200.075 ;
        RECT 77.035 199.125 77.205 199.905 ;
        RECT 77.375 199.455 77.595 199.735 ;
        RECT 77.775 199.625 78.315 199.995 ;
        RECT 78.660 199.915 78.830 200.505 ;
        RECT 79.050 200.085 79.355 201.225 ;
        RECT 79.525 200.035 79.780 200.915 ;
        RECT 80.070 200.595 80.355 201.055 ;
        RECT 80.525 200.765 80.795 201.225 ;
        RECT 80.070 200.375 81.025 200.595 ;
        RECT 78.660 199.885 79.400 199.915 ;
        RECT 77.375 199.285 77.905 199.455 ;
        RECT 75.685 198.865 76.035 199.035 ;
        RECT 76.255 198.845 77.205 199.125 ;
        RECT 77.375 198.675 77.565 199.115 ;
        RECT 77.735 199.055 77.905 199.285 ;
        RECT 78.075 199.225 78.315 199.625 ;
        RECT 78.485 199.585 79.400 199.885 ;
        RECT 78.485 199.410 78.810 199.585 ;
        RECT 78.485 199.055 78.805 199.410 ;
        RECT 79.570 199.385 79.780 200.035 ;
        RECT 79.955 199.645 80.645 200.205 ;
        RECT 80.815 199.475 81.025 200.375 ;
        RECT 77.735 198.885 78.805 199.055 ;
        RECT 79.050 198.675 79.355 199.135 ;
        RECT 79.525 198.855 79.780 199.385 ;
        RECT 80.070 199.305 81.025 199.475 ;
        RECT 81.195 200.205 81.595 201.055 ;
        RECT 81.785 200.595 82.065 201.055 ;
        RECT 82.585 200.765 82.910 201.225 ;
        RECT 81.785 200.375 82.910 200.595 ;
        RECT 81.195 199.645 82.290 200.205 ;
        RECT 82.460 199.915 82.910 200.375 ;
        RECT 83.080 200.085 83.465 201.055 ;
        RECT 83.750 200.595 84.035 201.055 ;
        RECT 84.205 200.765 84.475 201.225 ;
        RECT 83.750 200.375 84.705 200.595 ;
        RECT 80.070 198.845 80.355 199.305 ;
        RECT 80.525 198.675 80.795 199.135 ;
        RECT 81.195 198.845 81.595 199.645 ;
        RECT 82.460 199.585 83.015 199.915 ;
        RECT 82.460 199.475 82.910 199.585 ;
        RECT 81.785 199.305 82.910 199.475 ;
        RECT 83.185 199.415 83.465 200.085 ;
        RECT 83.635 199.645 84.325 200.205 ;
        RECT 84.495 199.475 84.705 200.375 ;
        RECT 81.785 198.845 82.065 199.305 ;
        RECT 82.585 198.675 82.910 199.135 ;
        RECT 83.080 198.845 83.465 199.415 ;
        RECT 83.750 199.305 84.705 199.475 ;
        RECT 84.875 200.205 85.275 201.055 ;
        RECT 85.465 200.595 85.745 201.055 ;
        RECT 86.265 200.765 86.590 201.225 ;
        RECT 85.465 200.375 86.590 200.595 ;
        RECT 84.875 199.645 85.970 200.205 ;
        RECT 86.140 199.915 86.590 200.375 ;
        RECT 86.760 200.085 87.145 201.055 ;
        RECT 83.750 198.845 84.035 199.305 ;
        RECT 84.205 198.675 84.475 199.135 ;
        RECT 84.875 198.845 85.275 199.645 ;
        RECT 86.140 199.585 86.695 199.915 ;
        RECT 86.140 199.475 86.590 199.585 ;
        RECT 85.465 199.305 86.590 199.475 ;
        RECT 86.865 199.415 87.145 200.085 ;
        RECT 87.315 200.060 87.605 201.225 ;
        RECT 87.835 200.085 88.045 201.225 ;
        RECT 88.215 200.075 88.545 201.055 ;
        RECT 88.715 200.085 88.945 201.225 ;
        RECT 89.160 200.555 89.415 201.055 ;
        RECT 89.585 200.725 89.915 201.225 ;
        RECT 89.160 200.385 89.910 200.555 ;
        RECT 85.465 198.845 85.745 199.305 ;
        RECT 86.265 198.675 86.590 199.135 ;
        RECT 86.760 198.845 87.145 199.415 ;
        RECT 87.315 198.675 87.605 199.400 ;
        RECT 87.835 198.675 88.045 199.495 ;
        RECT 88.215 199.475 88.465 200.075 ;
        RECT 88.635 199.665 88.965 199.915 ;
        RECT 89.160 199.565 89.510 200.215 ;
        RECT 88.215 198.845 88.545 199.475 ;
        RECT 88.715 198.675 88.945 199.495 ;
        RECT 89.680 199.395 89.910 200.385 ;
        RECT 89.160 199.225 89.910 199.395 ;
        RECT 89.160 198.935 89.415 199.225 ;
        RECT 89.585 198.675 89.915 199.055 ;
        RECT 90.085 198.935 90.255 201.055 ;
        RECT 90.425 200.255 90.750 201.040 ;
        RECT 90.920 200.765 91.170 201.225 ;
        RECT 91.340 200.725 91.590 201.055 ;
        RECT 91.805 200.725 92.485 201.055 ;
        RECT 91.340 200.595 91.510 200.725 ;
        RECT 91.115 200.425 91.510 200.595 ;
        RECT 90.485 199.205 90.945 200.255 ;
        RECT 91.115 199.065 91.285 200.425 ;
        RECT 91.680 200.165 92.145 200.555 ;
        RECT 91.455 199.355 91.805 199.975 ;
        RECT 91.975 199.575 92.145 200.165 ;
        RECT 92.315 199.945 92.485 200.725 ;
        RECT 92.655 200.625 92.825 200.965 ;
        RECT 93.060 200.795 93.390 201.225 ;
        RECT 93.560 200.625 93.730 200.965 ;
        RECT 94.025 200.765 94.395 201.225 ;
        RECT 92.655 200.455 93.730 200.625 ;
        RECT 94.565 200.595 94.735 201.055 ;
        RECT 94.970 200.715 95.840 201.055 ;
        RECT 96.010 200.765 96.260 201.225 ;
        RECT 94.175 200.425 94.735 200.595 ;
        RECT 94.175 200.285 94.345 200.425 ;
        RECT 92.845 200.115 94.345 200.285 ;
        RECT 95.040 200.255 95.500 200.545 ;
        RECT 92.315 199.775 94.005 199.945 ;
        RECT 91.975 199.355 92.330 199.575 ;
        RECT 92.500 199.065 92.670 199.775 ;
        RECT 92.875 199.355 93.665 199.605 ;
        RECT 93.835 199.595 94.005 199.775 ;
        RECT 94.175 199.425 94.345 200.115 ;
        RECT 90.615 198.675 90.945 199.035 ;
        RECT 91.115 198.895 91.610 199.065 ;
        RECT 91.815 198.895 92.670 199.065 ;
        RECT 93.545 198.675 93.875 199.135 ;
        RECT 94.085 199.035 94.345 199.425 ;
        RECT 94.535 200.245 95.500 200.255 ;
        RECT 95.670 200.335 95.840 200.715 ;
        RECT 96.430 200.675 96.600 200.965 ;
        RECT 96.780 200.845 97.110 201.225 ;
        RECT 96.430 200.505 97.230 200.675 ;
        RECT 94.535 200.085 95.210 200.245 ;
        RECT 95.670 200.165 96.890 200.335 ;
        RECT 94.535 199.295 94.745 200.085 ;
        RECT 95.670 200.075 95.840 200.165 ;
        RECT 94.915 199.295 95.265 199.915 ;
        RECT 95.435 199.905 95.840 200.075 ;
        RECT 95.435 199.125 95.605 199.905 ;
        RECT 95.775 199.455 95.995 199.735 ;
        RECT 96.175 199.625 96.715 199.995 ;
        RECT 97.060 199.915 97.230 200.505 ;
        RECT 97.450 200.085 97.755 201.225 ;
        RECT 97.925 200.035 98.180 200.915 ;
        RECT 98.360 200.555 98.615 201.055 ;
        RECT 98.785 200.725 99.115 201.225 ;
        RECT 98.360 200.385 99.110 200.555 ;
        RECT 97.060 199.885 97.800 199.915 ;
        RECT 95.775 199.285 96.305 199.455 ;
        RECT 94.085 198.865 94.435 199.035 ;
        RECT 94.655 198.845 95.605 199.125 ;
        RECT 95.775 198.675 95.965 199.115 ;
        RECT 96.135 199.055 96.305 199.285 ;
        RECT 96.475 199.225 96.715 199.625 ;
        RECT 96.885 199.585 97.800 199.885 ;
        RECT 96.885 199.410 97.210 199.585 ;
        RECT 96.885 199.055 97.205 199.410 ;
        RECT 97.970 199.385 98.180 200.035 ;
        RECT 98.360 199.565 98.710 200.215 ;
        RECT 98.880 199.395 99.110 200.385 ;
        RECT 96.135 198.885 97.205 199.055 ;
        RECT 97.450 198.675 97.755 199.135 ;
        RECT 97.925 198.855 98.180 199.385 ;
        RECT 98.360 199.225 99.110 199.395 ;
        RECT 98.360 198.935 98.615 199.225 ;
        RECT 98.785 198.675 99.115 199.055 ;
        RECT 99.285 198.935 99.455 201.055 ;
        RECT 99.625 200.255 99.950 201.040 ;
        RECT 100.120 200.765 100.370 201.225 ;
        RECT 100.540 200.725 100.790 201.055 ;
        RECT 101.005 200.725 101.685 201.055 ;
        RECT 100.540 200.595 100.710 200.725 ;
        RECT 100.315 200.425 100.710 200.595 ;
        RECT 99.685 199.205 100.145 200.255 ;
        RECT 100.315 199.065 100.485 200.425 ;
        RECT 100.880 200.165 101.345 200.555 ;
        RECT 100.655 199.355 101.005 199.975 ;
        RECT 101.175 199.575 101.345 200.165 ;
        RECT 101.515 199.945 101.685 200.725 ;
        RECT 101.855 200.625 102.025 200.965 ;
        RECT 102.260 200.795 102.590 201.225 ;
        RECT 102.760 200.625 102.930 200.965 ;
        RECT 103.225 200.765 103.595 201.225 ;
        RECT 101.855 200.455 102.930 200.625 ;
        RECT 103.765 200.595 103.935 201.055 ;
        RECT 104.170 200.715 105.040 201.055 ;
        RECT 105.210 200.765 105.460 201.225 ;
        RECT 103.375 200.425 103.935 200.595 ;
        RECT 103.375 200.285 103.545 200.425 ;
        RECT 102.045 200.115 103.545 200.285 ;
        RECT 104.240 200.255 104.700 200.545 ;
        RECT 101.515 199.775 103.205 199.945 ;
        RECT 101.175 199.355 101.530 199.575 ;
        RECT 101.700 199.065 101.870 199.775 ;
        RECT 102.075 199.355 102.865 199.605 ;
        RECT 103.035 199.595 103.205 199.775 ;
        RECT 103.375 199.425 103.545 200.115 ;
        RECT 99.815 198.675 100.145 199.035 ;
        RECT 100.315 198.895 100.810 199.065 ;
        RECT 101.015 198.895 101.870 199.065 ;
        RECT 102.745 198.675 103.075 199.135 ;
        RECT 103.285 199.035 103.545 199.425 ;
        RECT 103.735 200.245 104.700 200.255 ;
        RECT 104.870 200.335 105.040 200.715 ;
        RECT 105.630 200.675 105.800 200.965 ;
        RECT 105.980 200.845 106.310 201.225 ;
        RECT 105.630 200.505 106.430 200.675 ;
        RECT 103.735 200.085 104.410 200.245 ;
        RECT 104.870 200.165 106.090 200.335 ;
        RECT 103.735 199.295 103.945 200.085 ;
        RECT 104.870 200.075 105.040 200.165 ;
        RECT 104.115 199.295 104.465 199.915 ;
        RECT 104.635 199.905 105.040 200.075 ;
        RECT 104.635 199.125 104.805 199.905 ;
        RECT 104.975 199.455 105.195 199.735 ;
        RECT 105.375 199.625 105.915 199.995 ;
        RECT 106.260 199.915 106.430 200.505 ;
        RECT 106.650 200.085 106.955 201.225 ;
        RECT 107.125 200.035 107.380 200.915 ;
        RECT 107.670 200.595 107.955 201.055 ;
        RECT 108.125 200.765 108.395 201.225 ;
        RECT 107.670 200.375 108.625 200.595 ;
        RECT 106.260 199.885 107.000 199.915 ;
        RECT 104.975 199.285 105.505 199.455 ;
        RECT 103.285 198.865 103.635 199.035 ;
        RECT 103.855 198.845 104.805 199.125 ;
        RECT 104.975 198.675 105.165 199.115 ;
        RECT 105.335 199.055 105.505 199.285 ;
        RECT 105.675 199.225 105.915 199.625 ;
        RECT 106.085 199.585 107.000 199.885 ;
        RECT 106.085 199.410 106.410 199.585 ;
        RECT 106.085 199.055 106.405 199.410 ;
        RECT 107.170 199.385 107.380 200.035 ;
        RECT 107.555 199.645 108.245 200.205 ;
        RECT 108.415 199.475 108.625 200.375 ;
        RECT 105.335 198.885 106.405 199.055 ;
        RECT 106.650 198.675 106.955 199.135 ;
        RECT 107.125 198.855 107.380 199.385 ;
        RECT 107.670 199.305 108.625 199.475 ;
        RECT 108.795 200.205 109.195 201.055 ;
        RECT 109.385 200.595 109.665 201.055 ;
        RECT 110.185 200.765 110.510 201.225 ;
        RECT 109.385 200.375 110.510 200.595 ;
        RECT 108.795 199.645 109.890 200.205 ;
        RECT 110.060 199.915 110.510 200.375 ;
        RECT 110.680 200.085 111.065 201.055 ;
        RECT 107.670 198.845 107.955 199.305 ;
        RECT 108.125 198.675 108.395 199.135 ;
        RECT 108.795 198.845 109.195 199.645 ;
        RECT 110.060 199.585 110.615 199.915 ;
        RECT 110.060 199.475 110.510 199.585 ;
        RECT 109.385 199.305 110.510 199.475 ;
        RECT 110.785 199.415 111.065 200.085 ;
        RECT 112.155 200.135 113.365 201.225 ;
        RECT 112.155 199.595 112.675 200.135 ;
        RECT 112.845 199.425 113.365 199.965 ;
        RECT 109.385 198.845 109.665 199.305 ;
        RECT 110.185 198.675 110.510 199.135 ;
        RECT 110.680 198.845 111.065 199.415 ;
        RECT 112.155 198.675 113.365 199.425 ;
        RECT 26.970 198.505 113.450 198.675 ;
        RECT 27.055 197.755 28.265 198.505 ;
        RECT 28.550 197.875 28.835 198.335 ;
        RECT 29.005 198.045 29.275 198.505 ;
        RECT 27.055 197.215 27.575 197.755 ;
        RECT 28.550 197.705 29.505 197.875 ;
        RECT 27.745 197.045 28.265 197.585 ;
        RECT 27.055 195.955 28.265 197.045 ;
        RECT 28.435 196.975 29.125 197.535 ;
        RECT 29.295 196.805 29.505 197.705 ;
        RECT 28.550 196.585 29.505 196.805 ;
        RECT 29.675 197.535 30.075 198.335 ;
        RECT 30.265 197.875 30.545 198.335 ;
        RECT 31.065 198.045 31.390 198.505 ;
        RECT 30.265 197.705 31.390 197.875 ;
        RECT 31.560 197.765 31.945 198.335 ;
        RECT 30.940 197.595 31.390 197.705 ;
        RECT 29.675 196.975 30.770 197.535 ;
        RECT 30.940 197.265 31.495 197.595 ;
        RECT 28.550 196.125 28.835 196.585 ;
        RECT 29.005 195.955 29.275 196.415 ;
        RECT 29.675 196.125 30.075 196.975 ;
        RECT 30.940 196.805 31.390 197.265 ;
        RECT 31.665 197.095 31.945 197.765 ;
        RECT 32.175 197.685 32.385 198.505 ;
        RECT 32.555 197.705 32.885 198.335 ;
        RECT 32.555 197.105 32.805 197.705 ;
        RECT 33.055 197.685 33.285 198.505 ;
        RECT 33.535 197.685 33.765 198.505 ;
        RECT 33.935 197.705 34.265 198.335 ;
        RECT 32.975 197.265 33.305 197.515 ;
        RECT 33.515 197.265 33.845 197.515 ;
        RECT 34.015 197.105 34.265 197.705 ;
        RECT 34.435 197.685 34.645 198.505 ;
        RECT 34.990 197.875 35.275 198.335 ;
        RECT 35.445 198.045 35.715 198.505 ;
        RECT 34.990 197.705 35.945 197.875 ;
        RECT 30.265 196.585 31.390 196.805 ;
        RECT 30.265 196.125 30.545 196.585 ;
        RECT 31.065 195.955 31.390 196.415 ;
        RECT 31.560 196.125 31.945 197.095 ;
        RECT 32.175 195.955 32.385 197.095 ;
        RECT 32.555 196.125 32.885 197.105 ;
        RECT 33.055 195.955 33.285 197.095 ;
        RECT 33.535 195.955 33.765 197.095 ;
        RECT 33.935 196.125 34.265 197.105 ;
        RECT 34.435 195.955 34.645 197.095 ;
        RECT 34.875 196.975 35.565 197.535 ;
        RECT 35.735 196.805 35.945 197.705 ;
        RECT 34.990 196.585 35.945 196.805 ;
        RECT 36.115 197.535 36.515 198.335 ;
        RECT 36.705 197.875 36.985 198.335 ;
        RECT 37.505 198.045 37.830 198.505 ;
        RECT 36.705 197.705 37.830 197.875 ;
        RECT 38.000 197.765 38.385 198.335 ;
        RECT 37.380 197.595 37.830 197.705 ;
        RECT 36.115 196.975 37.210 197.535 ;
        RECT 37.380 197.265 37.935 197.595 ;
        RECT 34.990 196.125 35.275 196.585 ;
        RECT 35.445 195.955 35.715 196.415 ;
        RECT 36.115 196.125 36.515 196.975 ;
        RECT 37.380 196.805 37.830 197.265 ;
        RECT 38.105 197.095 38.385 197.765 ;
        RECT 36.705 196.585 37.830 196.805 ;
        RECT 36.705 196.125 36.985 196.585 ;
        RECT 37.505 195.955 37.830 196.415 ;
        RECT 38.000 196.125 38.385 197.095 ;
        RECT 38.555 197.830 38.815 198.335 ;
        RECT 38.995 198.125 39.325 198.505 ;
        RECT 39.505 197.955 39.675 198.335 ;
        RECT 38.555 197.030 38.725 197.830 ;
        RECT 39.010 197.785 39.675 197.955 ;
        RECT 40.025 197.955 40.195 198.335 ;
        RECT 40.375 198.125 40.705 198.505 ;
        RECT 40.025 197.785 40.690 197.955 ;
        RECT 40.885 197.830 41.145 198.335 ;
        RECT 39.010 197.530 39.180 197.785 ;
        RECT 38.895 197.200 39.180 197.530 ;
        RECT 39.415 197.235 39.745 197.605 ;
        RECT 39.955 197.235 40.285 197.605 ;
        RECT 40.520 197.530 40.690 197.785 ;
        RECT 39.010 197.055 39.180 197.200 ;
        RECT 40.520 197.200 40.805 197.530 ;
        RECT 40.520 197.055 40.690 197.200 ;
        RECT 38.555 196.125 38.825 197.030 ;
        RECT 39.010 196.885 39.675 197.055 ;
        RECT 38.995 195.955 39.325 196.715 ;
        RECT 39.505 196.125 39.675 196.885 ;
        RECT 40.025 196.885 40.690 197.055 ;
        RECT 40.975 197.030 41.145 197.830 ;
        RECT 41.520 197.725 42.020 198.335 ;
        RECT 41.315 197.265 41.665 197.515 ;
        RECT 41.850 197.095 42.020 197.725 ;
        RECT 42.650 197.855 42.980 198.335 ;
        RECT 43.150 198.045 43.375 198.505 ;
        RECT 43.545 197.855 43.875 198.335 ;
        RECT 42.650 197.685 43.875 197.855 ;
        RECT 44.065 197.705 44.315 198.505 ;
        RECT 44.485 197.705 44.825 198.335 ;
        RECT 45.110 197.875 45.395 198.335 ;
        RECT 45.565 198.045 45.835 198.505 ;
        RECT 45.110 197.705 46.065 197.875 ;
        RECT 42.190 197.315 42.520 197.515 ;
        RECT 42.690 197.315 43.020 197.515 ;
        RECT 43.190 197.315 43.610 197.515 ;
        RECT 43.785 197.345 44.480 197.515 ;
        RECT 43.785 197.095 43.955 197.345 ;
        RECT 44.650 197.145 44.825 197.705 ;
        RECT 44.595 197.095 44.825 197.145 ;
        RECT 40.025 196.125 40.195 196.885 ;
        RECT 40.375 195.955 40.705 196.715 ;
        RECT 40.875 196.125 41.145 197.030 ;
        RECT 41.520 196.925 43.955 197.095 ;
        RECT 41.520 196.125 41.850 196.925 ;
        RECT 42.020 195.955 42.350 196.755 ;
        RECT 42.650 196.125 42.980 196.925 ;
        RECT 43.625 195.955 43.875 196.755 ;
        RECT 44.145 195.955 44.315 197.095 ;
        RECT 44.485 196.125 44.825 197.095 ;
        RECT 44.995 196.975 45.685 197.535 ;
        RECT 45.855 196.805 46.065 197.705 ;
        RECT 45.110 196.585 46.065 196.805 ;
        RECT 46.235 197.535 46.635 198.335 ;
        RECT 46.825 197.875 47.105 198.335 ;
        RECT 47.625 198.045 47.950 198.505 ;
        RECT 46.825 197.705 47.950 197.875 ;
        RECT 48.120 197.765 48.505 198.335 ;
        RECT 48.675 197.780 48.965 198.505 ;
        RECT 47.500 197.595 47.950 197.705 ;
        RECT 46.235 196.975 47.330 197.535 ;
        RECT 47.500 197.265 48.055 197.595 ;
        RECT 45.110 196.125 45.395 196.585 ;
        RECT 45.565 195.955 45.835 196.415 ;
        RECT 46.235 196.125 46.635 196.975 ;
        RECT 47.500 196.805 47.950 197.265 ;
        RECT 48.225 197.095 48.505 197.765 ;
        RECT 49.135 197.765 49.520 198.335 ;
        RECT 49.690 198.045 50.015 198.505 ;
        RECT 50.535 197.875 50.815 198.335 ;
        RECT 46.825 196.585 47.950 196.805 ;
        RECT 46.825 196.125 47.105 196.585 ;
        RECT 47.625 195.955 47.950 196.415 ;
        RECT 48.120 196.125 48.505 197.095 ;
        RECT 48.675 195.955 48.965 197.120 ;
        RECT 49.135 197.095 49.415 197.765 ;
        RECT 49.690 197.705 50.815 197.875 ;
        RECT 49.690 197.595 50.140 197.705 ;
        RECT 49.585 197.265 50.140 197.595 ;
        RECT 51.005 197.535 51.405 198.335 ;
        RECT 51.805 198.045 52.075 198.505 ;
        RECT 52.245 197.875 52.530 198.335 ;
        RECT 49.135 196.125 49.520 197.095 ;
        RECT 49.690 196.805 50.140 197.265 ;
        RECT 50.310 196.975 51.405 197.535 ;
        RECT 49.690 196.585 50.815 196.805 ;
        RECT 49.690 195.955 50.015 196.415 ;
        RECT 50.535 196.125 50.815 196.585 ;
        RECT 51.005 196.125 51.405 196.975 ;
        RECT 51.575 197.705 52.530 197.875 ;
        RECT 53.275 197.765 53.660 198.335 ;
        RECT 53.830 198.045 54.155 198.505 ;
        RECT 54.675 197.875 54.955 198.335 ;
        RECT 51.575 196.805 51.785 197.705 ;
        RECT 51.955 196.975 52.645 197.535 ;
        RECT 53.275 197.095 53.555 197.765 ;
        RECT 53.830 197.705 54.955 197.875 ;
        RECT 53.830 197.595 54.280 197.705 ;
        RECT 53.725 197.265 54.280 197.595 ;
        RECT 55.145 197.535 55.545 198.335 ;
        RECT 55.945 198.045 56.215 198.505 ;
        RECT 56.385 197.875 56.670 198.335 ;
        RECT 51.575 196.585 52.530 196.805 ;
        RECT 51.805 195.955 52.075 196.415 ;
        RECT 52.245 196.125 52.530 196.585 ;
        RECT 53.275 196.125 53.660 197.095 ;
        RECT 53.830 196.805 54.280 197.265 ;
        RECT 54.450 196.975 55.545 197.535 ;
        RECT 53.830 196.585 54.955 196.805 ;
        RECT 53.830 195.955 54.155 196.415 ;
        RECT 54.675 196.125 54.955 196.585 ;
        RECT 55.145 196.125 55.545 196.975 ;
        RECT 55.715 197.705 56.670 197.875 ;
        RECT 56.960 197.955 57.215 198.245 ;
        RECT 57.385 198.125 57.715 198.505 ;
        RECT 56.960 197.785 57.710 197.955 ;
        RECT 55.715 196.805 55.925 197.705 ;
        RECT 56.095 196.975 56.785 197.535 ;
        RECT 56.960 196.965 57.310 197.615 ;
        RECT 55.715 196.585 56.670 196.805 ;
        RECT 57.480 196.795 57.710 197.785 ;
        RECT 55.945 195.955 56.215 196.415 ;
        RECT 56.385 196.125 56.670 196.585 ;
        RECT 56.960 196.625 57.710 196.795 ;
        RECT 56.960 196.125 57.215 196.625 ;
        RECT 57.385 195.955 57.715 196.455 ;
        RECT 57.885 196.125 58.055 198.245 ;
        RECT 58.415 198.145 58.745 198.505 ;
        RECT 58.915 198.115 59.410 198.285 ;
        RECT 59.615 198.115 60.470 198.285 ;
        RECT 58.285 196.925 58.745 197.975 ;
        RECT 58.225 196.140 58.550 196.925 ;
        RECT 58.915 196.755 59.085 198.115 ;
        RECT 59.255 197.205 59.605 197.825 ;
        RECT 59.775 197.605 60.130 197.825 ;
        RECT 59.775 197.015 59.945 197.605 ;
        RECT 60.300 197.405 60.470 198.115 ;
        RECT 61.345 198.045 61.675 198.505 ;
        RECT 61.885 198.145 62.235 198.315 ;
        RECT 60.675 197.575 61.465 197.825 ;
        RECT 61.885 197.755 62.145 198.145 ;
        RECT 62.455 198.055 63.405 198.335 ;
        RECT 63.575 198.065 63.765 198.505 ;
        RECT 63.935 198.125 65.005 198.295 ;
        RECT 61.635 197.405 61.805 197.585 ;
        RECT 58.915 196.585 59.310 196.755 ;
        RECT 59.480 196.625 59.945 197.015 ;
        RECT 60.115 197.235 61.805 197.405 ;
        RECT 59.140 196.455 59.310 196.585 ;
        RECT 60.115 196.455 60.285 197.235 ;
        RECT 61.975 197.065 62.145 197.755 ;
        RECT 60.645 196.895 62.145 197.065 ;
        RECT 62.335 197.095 62.545 197.885 ;
        RECT 62.715 197.265 63.065 197.885 ;
        RECT 63.235 197.275 63.405 198.055 ;
        RECT 63.935 197.895 64.105 198.125 ;
        RECT 63.575 197.725 64.105 197.895 ;
        RECT 63.575 197.445 63.795 197.725 ;
        RECT 64.275 197.555 64.515 197.955 ;
        RECT 63.235 197.105 63.640 197.275 ;
        RECT 63.975 197.185 64.515 197.555 ;
        RECT 64.685 197.770 65.005 198.125 ;
        RECT 64.685 197.515 65.010 197.770 ;
        RECT 65.205 197.695 65.375 198.505 ;
        RECT 65.545 197.855 65.875 198.335 ;
        RECT 66.045 198.035 66.215 198.505 ;
        RECT 66.385 197.855 66.715 198.335 ;
        RECT 66.885 198.035 67.055 198.505 ;
        RECT 65.545 197.685 67.310 197.855 ;
        RECT 67.535 197.765 68.230 198.335 ;
        RECT 68.400 197.765 68.750 198.290 ;
        RECT 64.685 197.305 66.715 197.515 ;
        RECT 64.685 197.295 65.030 197.305 ;
        RECT 62.335 196.935 63.010 197.095 ;
        RECT 63.470 197.015 63.640 197.105 ;
        RECT 62.335 196.925 63.300 196.935 ;
        RECT 61.975 196.755 62.145 196.895 ;
        RECT 58.720 195.955 58.970 196.415 ;
        RECT 59.140 196.125 59.390 196.455 ;
        RECT 59.605 196.125 60.285 196.455 ;
        RECT 60.455 196.555 61.530 196.725 ;
        RECT 61.975 196.585 62.535 196.755 ;
        RECT 62.840 196.635 63.300 196.925 ;
        RECT 63.470 196.845 64.690 197.015 ;
        RECT 60.455 196.215 60.625 196.555 ;
        RECT 60.860 195.955 61.190 196.385 ;
        RECT 61.360 196.215 61.530 196.555 ;
        RECT 61.825 195.955 62.195 196.415 ;
        RECT 62.365 196.125 62.535 196.585 ;
        RECT 63.470 196.465 63.640 196.845 ;
        RECT 64.860 196.675 65.030 197.295 ;
        RECT 66.900 197.135 67.310 197.685 ;
        RECT 62.770 196.125 63.640 196.465 ;
        RECT 64.230 196.505 65.030 196.675 ;
        RECT 63.810 195.955 64.060 196.415 ;
        RECT 64.230 196.215 64.400 196.505 ;
        RECT 64.580 195.955 64.910 196.335 ;
        RECT 65.205 195.955 65.375 197.015 ;
        RECT 65.585 196.965 67.310 197.135 ;
        RECT 65.585 196.125 65.875 196.965 ;
        RECT 66.045 195.955 66.215 196.795 ;
        RECT 66.425 196.125 66.675 196.965 ;
        RECT 67.535 196.925 67.775 197.595 ;
        RECT 67.955 197.095 68.125 197.765 ;
        RECT 68.400 197.595 68.605 197.765 ;
        RECT 68.940 197.595 69.155 198.290 ;
        RECT 69.325 197.765 69.660 198.505 ;
        RECT 69.920 197.935 70.095 198.335 ;
        RECT 70.265 198.125 70.595 198.505 ;
        RECT 70.840 198.005 71.070 198.335 ;
        RECT 69.920 197.765 70.550 197.935 ;
        RECT 70.380 197.595 70.550 197.765 ;
        RECT 68.295 197.265 68.605 197.595 ;
        RECT 68.775 197.265 69.155 197.595 ;
        RECT 69.355 197.265 69.640 197.595 ;
        RECT 67.955 196.925 69.235 197.095 ;
        RECT 66.885 195.955 67.055 196.795 ;
        RECT 67.555 195.955 67.835 196.755 ;
        RECT 68.035 196.125 68.365 196.925 ;
        RECT 68.565 195.955 68.735 196.755 ;
        RECT 68.905 196.125 69.235 196.925 ;
        RECT 69.405 195.955 69.665 197.095 ;
        RECT 69.835 196.915 70.200 197.595 ;
        RECT 70.380 197.265 70.730 197.595 ;
        RECT 70.380 196.745 70.550 197.265 ;
        RECT 69.920 196.575 70.550 196.745 ;
        RECT 70.900 196.715 71.070 198.005 ;
        RECT 71.270 196.895 71.550 198.170 ;
        RECT 71.775 197.485 72.045 198.170 ;
        RECT 72.505 198.125 72.835 198.505 ;
        RECT 73.005 198.250 73.340 198.295 ;
        RECT 71.735 197.315 72.045 197.485 ;
        RECT 71.775 196.895 72.045 197.315 ;
        RECT 72.235 196.895 72.575 197.925 ;
        RECT 73.005 197.785 73.345 198.250 ;
        RECT 72.745 197.265 73.005 197.595 ;
        RECT 72.745 196.715 72.915 197.265 ;
        RECT 73.175 197.095 73.345 197.785 ;
        RECT 74.435 197.780 74.725 198.505 ;
        RECT 74.935 197.685 75.165 198.505 ;
        RECT 75.335 197.705 75.665 198.335 ;
        RECT 74.915 197.265 75.245 197.515 ;
        RECT 69.920 196.125 70.095 196.575 ;
        RECT 70.900 196.545 72.915 196.715 ;
        RECT 70.265 195.955 70.595 196.395 ;
        RECT 70.900 196.125 71.070 196.545 ;
        RECT 71.305 195.955 71.975 196.365 ;
        RECT 72.190 196.125 72.360 196.545 ;
        RECT 72.560 195.955 72.890 196.365 ;
        RECT 73.085 196.125 73.345 197.095 ;
        RECT 74.435 195.955 74.725 197.120 ;
        RECT 75.415 197.105 75.665 197.705 ;
        RECT 75.835 197.685 76.045 198.505 ;
        RECT 76.275 197.765 76.740 198.310 ;
        RECT 74.935 195.955 75.165 197.095 ;
        RECT 75.335 196.125 75.665 197.105 ;
        RECT 75.835 195.955 76.045 197.095 ;
        RECT 76.275 196.805 76.445 197.765 ;
        RECT 77.245 197.685 77.415 198.505 ;
        RECT 77.585 197.855 77.915 198.335 ;
        RECT 78.085 198.115 78.435 198.505 ;
        RECT 78.605 197.935 78.835 198.335 ;
        RECT 78.325 197.855 78.835 197.935 ;
        RECT 77.585 197.765 78.835 197.855 ;
        RECT 79.005 197.765 79.325 198.245 ;
        RECT 77.585 197.685 78.495 197.765 ;
        RECT 76.615 197.145 76.860 197.595 ;
        RECT 77.120 197.315 77.815 197.515 ;
        RECT 77.985 197.345 78.585 197.515 ;
        RECT 77.985 197.145 78.155 197.345 ;
        RECT 78.815 197.175 78.985 197.595 ;
        RECT 76.615 196.975 78.155 197.145 ;
        RECT 78.325 197.005 78.985 197.175 ;
        RECT 78.325 196.805 78.495 197.005 ;
        RECT 79.155 196.835 79.325 197.765 ;
        RECT 79.610 197.875 79.895 198.335 ;
        RECT 80.065 198.045 80.335 198.505 ;
        RECT 79.610 197.705 80.565 197.875 ;
        RECT 79.495 196.975 80.185 197.535 ;
        RECT 76.275 196.635 78.495 196.805 ;
        RECT 78.665 196.635 79.325 196.835 ;
        RECT 80.355 196.805 80.565 197.705 ;
        RECT 76.275 195.955 76.575 196.465 ;
        RECT 76.745 196.125 77.075 196.635 ;
        RECT 78.665 196.465 78.835 196.635 ;
        RECT 79.610 196.585 80.565 196.805 ;
        RECT 80.735 197.535 81.135 198.335 ;
        RECT 81.325 197.875 81.605 198.335 ;
        RECT 82.125 198.045 82.450 198.505 ;
        RECT 81.325 197.705 82.450 197.875 ;
        RECT 82.620 197.765 83.005 198.335 ;
        RECT 83.265 197.955 83.435 198.245 ;
        RECT 83.605 198.125 83.935 198.505 ;
        RECT 83.265 197.785 83.930 197.955 ;
        RECT 82.000 197.595 82.450 197.705 ;
        RECT 80.735 196.975 81.830 197.535 ;
        RECT 82.000 197.265 82.555 197.595 ;
        RECT 77.245 195.955 77.875 196.465 ;
        RECT 78.455 196.295 78.835 196.465 ;
        RECT 79.005 195.955 79.305 196.465 ;
        RECT 79.610 196.125 79.895 196.585 ;
        RECT 80.065 195.955 80.335 196.415 ;
        RECT 80.735 196.125 81.135 196.975 ;
        RECT 82.000 196.805 82.450 197.265 ;
        RECT 82.725 197.095 83.005 197.765 ;
        RECT 81.325 196.585 82.450 196.805 ;
        RECT 81.325 196.125 81.605 196.585 ;
        RECT 82.125 195.955 82.450 196.415 ;
        RECT 82.620 196.125 83.005 197.095 ;
        RECT 83.180 196.965 83.530 197.615 ;
        RECT 83.700 196.795 83.930 197.785 ;
        RECT 83.265 196.625 83.930 196.795 ;
        RECT 83.265 196.125 83.435 196.625 ;
        RECT 83.605 195.955 83.935 196.455 ;
        RECT 84.105 196.125 84.330 198.245 ;
        RECT 84.545 198.125 84.875 198.505 ;
        RECT 85.045 197.955 85.215 198.285 ;
        RECT 85.515 198.125 86.530 198.325 ;
        RECT 84.520 197.765 85.215 197.955 ;
        RECT 84.520 196.795 84.690 197.765 ;
        RECT 84.860 196.965 85.270 197.585 ;
        RECT 85.440 197.015 85.660 197.885 ;
        RECT 85.840 197.575 86.190 197.945 ;
        RECT 86.360 197.395 86.530 198.125 ;
        RECT 86.700 198.065 87.110 198.505 ;
        RECT 87.400 197.865 87.650 198.295 ;
        RECT 87.850 198.045 88.170 198.505 ;
        RECT 88.730 198.115 89.580 198.285 ;
        RECT 86.700 197.525 87.110 197.855 ;
        RECT 87.400 197.525 87.820 197.865 ;
        RECT 86.110 197.355 86.530 197.395 ;
        RECT 86.110 197.185 87.460 197.355 ;
        RECT 84.520 196.625 85.215 196.795 ;
        RECT 85.440 196.635 85.940 197.015 ;
        RECT 84.545 195.955 84.875 196.455 ;
        RECT 85.045 196.125 85.215 196.625 ;
        RECT 86.110 196.340 86.280 197.185 ;
        RECT 87.210 197.025 87.460 197.185 ;
        RECT 86.450 196.755 86.700 197.015 ;
        RECT 87.630 196.755 87.820 197.525 ;
        RECT 86.450 196.505 87.820 196.755 ;
        RECT 87.990 197.695 89.240 197.865 ;
        RECT 87.990 196.935 88.160 197.695 ;
        RECT 88.910 197.575 89.240 197.695 ;
        RECT 88.330 197.115 88.510 197.525 ;
        RECT 89.410 197.355 89.580 198.115 ;
        RECT 89.780 198.025 90.440 198.505 ;
        RECT 90.620 197.910 90.940 198.240 ;
        RECT 89.770 197.585 90.430 197.855 ;
        RECT 89.770 197.525 90.100 197.585 ;
        RECT 90.250 197.355 90.580 197.415 ;
        RECT 88.680 197.185 90.580 197.355 ;
        RECT 87.990 196.625 88.510 196.935 ;
        RECT 88.680 196.675 88.850 197.185 ;
        RECT 90.750 197.015 90.940 197.910 ;
        RECT 89.020 196.845 90.940 197.015 ;
        RECT 90.620 196.825 90.940 196.845 ;
        RECT 91.140 197.595 91.390 198.245 ;
        RECT 91.570 198.045 91.855 198.505 ;
        RECT 92.035 197.795 92.290 198.325 ;
        RECT 91.140 197.265 91.940 197.595 ;
        RECT 88.680 196.505 89.890 196.675 ;
        RECT 85.450 196.170 86.280 196.340 ;
        RECT 86.520 195.955 86.900 196.335 ;
        RECT 87.080 196.215 87.250 196.505 ;
        RECT 88.680 196.425 88.850 196.505 ;
        RECT 87.420 195.955 87.750 196.335 ;
        RECT 88.220 196.175 88.850 196.425 ;
        RECT 89.030 195.955 89.450 196.335 ;
        RECT 89.650 196.215 89.890 196.505 ;
        RECT 90.120 195.955 90.450 196.645 ;
        RECT 90.620 196.215 90.790 196.825 ;
        RECT 91.140 196.675 91.390 197.265 ;
        RECT 92.110 196.935 92.290 197.795 ;
        RECT 92.035 196.805 92.290 196.935 ;
        RECT 92.870 197.765 93.485 198.335 ;
        RECT 93.655 197.995 93.870 198.505 ;
        RECT 94.100 197.995 94.380 198.325 ;
        RECT 94.560 197.995 94.800 198.505 ;
        RECT 91.060 196.165 91.390 196.675 ;
        RECT 91.570 195.955 91.855 196.755 ;
        RECT 92.035 196.635 92.375 196.805 ;
        RECT 92.870 196.745 93.185 197.765 ;
        RECT 93.355 197.095 93.525 197.595 ;
        RECT 93.775 197.265 94.040 197.825 ;
        RECT 94.210 197.095 94.380 197.995 ;
        RECT 94.550 197.265 94.905 197.825 ;
        RECT 95.140 197.765 95.395 198.335 ;
        RECT 95.565 198.105 95.895 198.505 ;
        RECT 96.320 197.970 96.850 198.335 ;
        RECT 97.040 198.165 97.315 198.335 ;
        RECT 97.035 197.995 97.315 198.165 ;
        RECT 96.320 197.935 96.495 197.970 ;
        RECT 95.565 197.765 96.495 197.935 ;
        RECT 95.140 197.095 95.310 197.765 ;
        RECT 95.565 197.595 95.735 197.765 ;
        RECT 95.480 197.265 95.735 197.595 ;
        RECT 95.960 197.265 96.155 197.595 ;
        RECT 93.355 196.925 94.780 197.095 ;
        RECT 92.035 196.265 92.290 196.635 ;
        RECT 92.870 196.125 93.405 196.745 ;
        RECT 93.575 195.955 93.905 196.755 ;
        RECT 94.390 196.750 94.780 196.925 ;
        RECT 95.140 196.125 95.475 197.095 ;
        RECT 95.645 195.955 95.815 197.095 ;
        RECT 95.985 196.295 96.155 197.265 ;
        RECT 96.325 196.635 96.495 197.765 ;
        RECT 96.665 196.975 96.835 197.775 ;
        RECT 97.040 197.175 97.315 197.995 ;
        RECT 97.485 196.975 97.675 198.335 ;
        RECT 97.855 197.970 98.365 198.505 ;
        RECT 98.585 197.695 98.830 198.300 ;
        RECT 100.195 197.780 100.485 198.505 ;
        RECT 101.580 197.795 101.835 198.325 ;
        RECT 102.005 198.045 102.310 198.505 ;
        RECT 102.555 198.125 103.625 198.295 ;
        RECT 97.875 197.525 99.105 197.695 ;
        RECT 96.665 196.805 97.675 196.975 ;
        RECT 97.845 196.960 98.595 197.150 ;
        RECT 96.325 196.465 97.450 196.635 ;
        RECT 97.845 196.295 98.015 196.960 ;
        RECT 98.765 196.715 99.105 197.525 ;
        RECT 101.580 197.145 101.790 197.795 ;
        RECT 102.555 197.770 102.875 198.125 ;
        RECT 102.550 197.595 102.875 197.770 ;
        RECT 101.960 197.295 102.875 197.595 ;
        RECT 103.045 197.555 103.285 197.955 ;
        RECT 103.455 197.895 103.625 198.125 ;
        RECT 103.795 198.065 103.985 198.505 ;
        RECT 104.155 198.055 105.105 198.335 ;
        RECT 105.325 198.145 105.675 198.315 ;
        RECT 103.455 197.725 103.985 197.895 ;
        RECT 101.960 197.265 102.700 197.295 ;
        RECT 95.985 196.125 98.015 196.295 ;
        RECT 98.185 195.955 98.355 196.715 ;
        RECT 98.590 196.305 99.105 196.715 ;
        RECT 100.195 195.955 100.485 197.120 ;
        RECT 101.580 196.265 101.835 197.145 ;
        RECT 102.005 195.955 102.310 197.095 ;
        RECT 102.530 196.675 102.700 197.265 ;
        RECT 103.045 197.185 103.585 197.555 ;
        RECT 103.765 197.445 103.985 197.725 ;
        RECT 104.155 197.275 104.325 198.055 ;
        RECT 103.920 197.105 104.325 197.275 ;
        RECT 104.495 197.265 104.845 197.885 ;
        RECT 103.920 197.015 104.090 197.105 ;
        RECT 105.015 197.095 105.225 197.885 ;
        RECT 102.870 196.845 104.090 197.015 ;
        RECT 104.550 196.935 105.225 197.095 ;
        RECT 102.530 196.505 103.330 196.675 ;
        RECT 102.650 195.955 102.980 196.335 ;
        RECT 103.160 196.215 103.330 196.505 ;
        RECT 103.920 196.465 104.090 196.845 ;
        RECT 104.260 196.925 105.225 196.935 ;
        RECT 105.415 197.755 105.675 198.145 ;
        RECT 105.885 198.045 106.215 198.505 ;
        RECT 107.090 198.115 107.945 198.285 ;
        RECT 108.150 198.115 108.645 198.285 ;
        RECT 108.815 198.145 109.145 198.505 ;
        RECT 105.415 197.065 105.585 197.755 ;
        RECT 105.755 197.405 105.925 197.585 ;
        RECT 106.095 197.575 106.885 197.825 ;
        RECT 107.090 197.405 107.260 198.115 ;
        RECT 107.430 197.605 107.785 197.825 ;
        RECT 105.755 197.235 107.445 197.405 ;
        RECT 104.260 196.635 104.720 196.925 ;
        RECT 105.415 196.895 106.915 197.065 ;
        RECT 105.415 196.755 105.585 196.895 ;
        RECT 105.025 196.585 105.585 196.755 ;
        RECT 103.500 195.955 103.750 196.415 ;
        RECT 103.920 196.125 104.790 196.465 ;
        RECT 105.025 196.125 105.195 196.585 ;
        RECT 106.030 196.555 107.105 196.725 ;
        RECT 105.365 195.955 105.735 196.415 ;
        RECT 106.030 196.215 106.200 196.555 ;
        RECT 106.370 195.955 106.700 196.385 ;
        RECT 106.935 196.215 107.105 196.555 ;
        RECT 107.275 196.455 107.445 197.235 ;
        RECT 107.615 197.015 107.785 197.605 ;
        RECT 107.955 197.205 108.305 197.825 ;
        RECT 107.615 196.625 108.080 197.015 ;
        RECT 108.475 196.755 108.645 198.115 ;
        RECT 108.815 196.925 109.275 197.975 ;
        RECT 108.250 196.585 108.645 196.755 ;
        RECT 108.250 196.455 108.420 196.585 ;
        RECT 107.275 196.125 107.955 196.455 ;
        RECT 108.170 196.125 108.420 196.455 ;
        RECT 108.590 195.955 108.840 196.415 ;
        RECT 109.010 196.140 109.335 196.925 ;
        RECT 109.505 196.125 109.675 198.245 ;
        RECT 109.845 198.125 110.175 198.505 ;
        RECT 110.345 197.955 110.600 198.245 ;
        RECT 109.850 197.785 110.600 197.955 ;
        RECT 109.850 196.795 110.080 197.785 ;
        RECT 110.835 197.685 111.045 198.505 ;
        RECT 111.215 197.705 111.545 198.335 ;
        RECT 110.250 196.965 110.600 197.615 ;
        RECT 111.215 197.105 111.465 197.705 ;
        RECT 111.715 197.685 111.945 198.505 ;
        RECT 112.155 197.755 113.365 198.505 ;
        RECT 111.635 197.265 111.965 197.515 ;
        RECT 109.850 196.625 110.600 196.795 ;
        RECT 109.845 195.955 110.175 196.455 ;
        RECT 110.345 196.125 110.600 196.625 ;
        RECT 110.835 195.955 111.045 197.095 ;
        RECT 111.215 196.125 111.545 197.105 ;
        RECT 111.715 195.955 111.945 197.095 ;
        RECT 112.155 197.045 112.675 197.585 ;
        RECT 112.845 197.215 113.365 197.755 ;
        RECT 112.155 195.955 113.365 197.045 ;
        RECT 26.970 195.785 113.450 195.955 ;
        RECT 27.055 194.695 28.265 195.785 ;
        RECT 28.550 195.155 28.835 195.615 ;
        RECT 29.005 195.325 29.275 195.785 ;
        RECT 28.550 194.935 29.505 195.155 ;
        RECT 27.055 193.985 27.575 194.525 ;
        RECT 27.745 194.155 28.265 194.695 ;
        RECT 28.435 194.205 29.125 194.765 ;
        RECT 29.295 194.035 29.505 194.935 ;
        RECT 27.055 193.235 28.265 193.985 ;
        RECT 28.550 193.865 29.505 194.035 ;
        RECT 29.675 194.765 30.075 195.615 ;
        RECT 30.265 195.155 30.545 195.615 ;
        RECT 31.065 195.325 31.390 195.785 ;
        RECT 30.265 194.935 31.390 195.155 ;
        RECT 29.675 194.205 30.770 194.765 ;
        RECT 30.940 194.475 31.390 194.935 ;
        RECT 31.560 194.645 31.945 195.615 ;
        RECT 32.230 195.155 32.515 195.615 ;
        RECT 32.685 195.325 32.955 195.785 ;
        RECT 32.230 194.935 33.185 195.155 ;
        RECT 28.550 193.405 28.835 193.865 ;
        RECT 29.005 193.235 29.275 193.695 ;
        RECT 29.675 193.405 30.075 194.205 ;
        RECT 30.940 194.145 31.495 194.475 ;
        RECT 30.940 194.035 31.390 194.145 ;
        RECT 30.265 193.865 31.390 194.035 ;
        RECT 31.665 193.975 31.945 194.645 ;
        RECT 32.115 194.205 32.805 194.765 ;
        RECT 32.975 194.035 33.185 194.935 ;
        RECT 30.265 193.405 30.545 193.865 ;
        RECT 31.065 193.235 31.390 193.695 ;
        RECT 31.560 193.405 31.945 193.975 ;
        RECT 32.230 193.865 33.185 194.035 ;
        RECT 33.355 194.765 33.755 195.615 ;
        RECT 33.945 195.155 34.225 195.615 ;
        RECT 34.745 195.325 35.070 195.785 ;
        RECT 33.945 194.935 35.070 195.155 ;
        RECT 33.355 194.205 34.450 194.765 ;
        RECT 34.620 194.475 35.070 194.935 ;
        RECT 35.240 194.645 35.625 195.615 ;
        RECT 32.230 193.405 32.515 193.865 ;
        RECT 32.685 193.235 32.955 193.695 ;
        RECT 33.355 193.405 33.755 194.205 ;
        RECT 34.620 194.145 35.175 194.475 ;
        RECT 34.620 194.035 35.070 194.145 ;
        RECT 33.945 193.865 35.070 194.035 ;
        RECT 35.345 193.975 35.625 194.645 ;
        RECT 35.795 194.620 36.085 195.785 ;
        RECT 36.755 194.645 36.985 195.785 ;
        RECT 37.155 194.635 37.485 195.615 ;
        RECT 37.655 194.645 37.865 195.785 ;
        RECT 38.185 194.855 38.355 195.615 ;
        RECT 38.535 195.025 38.865 195.785 ;
        RECT 38.185 194.685 38.850 194.855 ;
        RECT 39.035 194.710 39.305 195.615 ;
        RECT 36.735 194.225 37.065 194.475 ;
        RECT 33.945 193.405 34.225 193.865 ;
        RECT 34.745 193.235 35.070 193.695 ;
        RECT 35.240 193.405 35.625 193.975 ;
        RECT 35.795 193.235 36.085 193.960 ;
        RECT 36.755 193.235 36.985 194.055 ;
        RECT 37.235 194.035 37.485 194.635 ;
        RECT 38.680 194.540 38.850 194.685 ;
        RECT 38.115 194.135 38.445 194.505 ;
        RECT 38.680 194.210 38.965 194.540 ;
        RECT 37.155 193.405 37.485 194.035 ;
        RECT 37.655 193.235 37.865 194.055 ;
        RECT 38.680 193.955 38.850 194.210 ;
        RECT 38.185 193.785 38.850 193.955 ;
        RECT 39.135 193.910 39.305 194.710 ;
        RECT 38.185 193.405 38.355 193.785 ;
        RECT 38.535 193.235 38.865 193.615 ;
        RECT 39.045 193.405 39.305 193.910 ;
        RECT 39.475 194.645 39.815 195.615 ;
        RECT 39.985 194.645 40.155 195.785 ;
        RECT 40.425 194.985 40.675 195.785 ;
        RECT 41.320 194.815 41.650 195.615 ;
        RECT 41.950 194.985 42.280 195.785 ;
        RECT 42.450 194.815 42.780 195.615 ;
        RECT 43.160 195.115 43.415 195.615 ;
        RECT 43.585 195.285 43.915 195.785 ;
        RECT 43.160 194.945 43.910 195.115 ;
        RECT 40.345 194.645 42.780 194.815 ;
        RECT 39.475 194.035 39.650 194.645 ;
        RECT 40.345 194.395 40.515 194.645 ;
        RECT 39.820 194.225 40.515 194.395 ;
        RECT 40.690 194.225 41.110 194.425 ;
        RECT 41.280 194.225 41.610 194.425 ;
        RECT 41.780 194.225 42.110 194.425 ;
        RECT 39.475 193.405 39.815 194.035 ;
        RECT 39.985 193.235 40.235 194.035 ;
        RECT 40.425 193.885 41.650 194.055 ;
        RECT 40.425 193.405 40.755 193.885 ;
        RECT 40.925 193.235 41.150 193.695 ;
        RECT 41.320 193.405 41.650 193.885 ;
        RECT 42.280 194.015 42.450 194.645 ;
        RECT 42.635 194.225 42.985 194.475 ;
        RECT 43.160 194.125 43.510 194.775 ;
        RECT 42.280 193.405 42.780 194.015 ;
        RECT 43.680 193.955 43.910 194.945 ;
        RECT 43.160 193.785 43.910 193.955 ;
        RECT 43.160 193.495 43.415 193.785 ;
        RECT 43.585 193.235 43.915 193.615 ;
        RECT 44.085 193.495 44.255 195.615 ;
        RECT 44.425 194.815 44.750 195.600 ;
        RECT 44.920 195.325 45.170 195.785 ;
        RECT 45.340 195.285 45.590 195.615 ;
        RECT 45.805 195.285 46.485 195.615 ;
        RECT 45.340 195.155 45.510 195.285 ;
        RECT 45.115 194.985 45.510 195.155 ;
        RECT 44.485 193.765 44.945 194.815 ;
        RECT 45.115 193.625 45.285 194.985 ;
        RECT 45.680 194.725 46.145 195.115 ;
        RECT 45.455 193.915 45.805 194.535 ;
        RECT 45.975 194.135 46.145 194.725 ;
        RECT 46.315 194.505 46.485 195.285 ;
        RECT 46.655 195.185 46.825 195.525 ;
        RECT 47.060 195.355 47.390 195.785 ;
        RECT 47.560 195.185 47.730 195.525 ;
        RECT 48.025 195.325 48.395 195.785 ;
        RECT 46.655 195.015 47.730 195.185 ;
        RECT 48.565 195.155 48.735 195.615 ;
        RECT 48.970 195.275 49.840 195.615 ;
        RECT 50.010 195.325 50.260 195.785 ;
        RECT 48.175 194.985 48.735 195.155 ;
        RECT 48.175 194.845 48.345 194.985 ;
        RECT 46.845 194.675 48.345 194.845 ;
        RECT 49.040 194.815 49.500 195.105 ;
        RECT 46.315 194.335 48.005 194.505 ;
        RECT 45.975 193.915 46.330 194.135 ;
        RECT 46.500 193.625 46.670 194.335 ;
        RECT 46.875 193.915 47.665 194.165 ;
        RECT 47.835 194.155 48.005 194.335 ;
        RECT 48.175 193.985 48.345 194.675 ;
        RECT 44.615 193.235 44.945 193.595 ;
        RECT 45.115 193.455 45.610 193.625 ;
        RECT 45.815 193.455 46.670 193.625 ;
        RECT 47.545 193.235 47.875 193.695 ;
        RECT 48.085 193.595 48.345 193.985 ;
        RECT 48.535 194.805 49.500 194.815 ;
        RECT 49.670 194.895 49.840 195.275 ;
        RECT 50.430 195.235 50.600 195.525 ;
        RECT 50.780 195.405 51.110 195.785 ;
        RECT 50.430 195.065 51.230 195.235 ;
        RECT 48.535 194.645 49.210 194.805 ;
        RECT 49.670 194.725 50.890 194.895 ;
        RECT 48.535 193.855 48.745 194.645 ;
        RECT 49.670 194.635 49.840 194.725 ;
        RECT 48.915 193.855 49.265 194.475 ;
        RECT 49.435 194.465 49.840 194.635 ;
        RECT 49.435 193.685 49.605 194.465 ;
        RECT 49.775 194.015 49.995 194.295 ;
        RECT 50.175 194.185 50.715 194.555 ;
        RECT 51.060 194.475 51.230 195.065 ;
        RECT 51.450 194.645 51.755 195.785 ;
        RECT 51.925 194.595 52.180 195.475 ;
        RECT 52.360 195.115 52.615 195.615 ;
        RECT 52.785 195.285 53.115 195.785 ;
        RECT 52.360 194.945 53.110 195.115 ;
        RECT 51.060 194.445 51.800 194.475 ;
        RECT 49.775 193.845 50.305 194.015 ;
        RECT 48.085 193.425 48.435 193.595 ;
        RECT 48.655 193.405 49.605 193.685 ;
        RECT 49.775 193.235 49.965 193.675 ;
        RECT 50.135 193.615 50.305 193.845 ;
        RECT 50.475 193.785 50.715 194.185 ;
        RECT 50.885 194.145 51.800 194.445 ;
        RECT 50.885 193.970 51.210 194.145 ;
        RECT 50.885 193.615 51.205 193.970 ;
        RECT 51.970 193.945 52.180 194.595 ;
        RECT 52.360 194.125 52.710 194.775 ;
        RECT 52.880 193.955 53.110 194.945 ;
        RECT 50.135 193.445 51.205 193.615 ;
        RECT 51.450 193.235 51.755 193.695 ;
        RECT 51.925 193.415 52.180 193.945 ;
        RECT 52.360 193.785 53.110 193.955 ;
        RECT 52.360 193.495 52.615 193.785 ;
        RECT 52.785 193.235 53.115 193.615 ;
        RECT 53.285 193.495 53.455 195.615 ;
        RECT 53.625 194.815 53.950 195.600 ;
        RECT 54.120 195.325 54.370 195.785 ;
        RECT 54.540 195.285 54.790 195.615 ;
        RECT 55.005 195.285 55.685 195.615 ;
        RECT 54.540 195.155 54.710 195.285 ;
        RECT 54.315 194.985 54.710 195.155 ;
        RECT 53.685 193.765 54.145 194.815 ;
        RECT 54.315 193.625 54.485 194.985 ;
        RECT 54.880 194.725 55.345 195.115 ;
        RECT 54.655 193.915 55.005 194.535 ;
        RECT 55.175 194.135 55.345 194.725 ;
        RECT 55.515 194.505 55.685 195.285 ;
        RECT 55.855 195.185 56.025 195.525 ;
        RECT 56.260 195.355 56.590 195.785 ;
        RECT 56.760 195.185 56.930 195.525 ;
        RECT 57.225 195.325 57.595 195.785 ;
        RECT 55.855 195.015 56.930 195.185 ;
        RECT 57.765 195.155 57.935 195.615 ;
        RECT 58.170 195.275 59.040 195.615 ;
        RECT 59.210 195.325 59.460 195.785 ;
        RECT 57.375 194.985 57.935 195.155 ;
        RECT 57.375 194.845 57.545 194.985 ;
        RECT 56.045 194.675 57.545 194.845 ;
        RECT 58.240 194.815 58.700 195.105 ;
        RECT 55.515 194.335 57.205 194.505 ;
        RECT 55.175 193.915 55.530 194.135 ;
        RECT 55.700 193.625 55.870 194.335 ;
        RECT 56.075 193.915 56.865 194.165 ;
        RECT 57.035 194.155 57.205 194.335 ;
        RECT 57.375 193.985 57.545 194.675 ;
        RECT 53.815 193.235 54.145 193.595 ;
        RECT 54.315 193.455 54.810 193.625 ;
        RECT 55.015 193.455 55.870 193.625 ;
        RECT 56.745 193.235 57.075 193.695 ;
        RECT 57.285 193.595 57.545 193.985 ;
        RECT 57.735 194.805 58.700 194.815 ;
        RECT 58.870 194.895 59.040 195.275 ;
        RECT 59.630 195.235 59.800 195.525 ;
        RECT 59.980 195.405 60.310 195.785 ;
        RECT 59.630 195.065 60.430 195.235 ;
        RECT 57.735 194.645 58.410 194.805 ;
        RECT 58.870 194.725 60.090 194.895 ;
        RECT 57.735 193.855 57.945 194.645 ;
        RECT 58.870 194.635 59.040 194.725 ;
        RECT 58.115 193.855 58.465 194.475 ;
        RECT 58.635 194.465 59.040 194.635 ;
        RECT 58.635 193.685 58.805 194.465 ;
        RECT 58.975 194.015 59.195 194.295 ;
        RECT 59.375 194.185 59.915 194.555 ;
        RECT 60.260 194.475 60.430 195.065 ;
        RECT 60.650 194.645 60.955 195.785 ;
        RECT 61.125 194.595 61.380 195.475 ;
        RECT 61.555 194.620 61.845 195.785 ;
        RECT 62.480 194.635 62.740 195.785 ;
        RECT 62.915 194.710 63.170 195.615 ;
        RECT 63.340 195.025 63.670 195.785 ;
        RECT 63.885 194.855 64.055 195.615 ;
        RECT 60.260 194.445 61.000 194.475 ;
        RECT 58.975 193.845 59.505 194.015 ;
        RECT 57.285 193.425 57.635 193.595 ;
        RECT 57.855 193.405 58.805 193.685 ;
        RECT 58.975 193.235 59.165 193.675 ;
        RECT 59.335 193.615 59.505 193.845 ;
        RECT 59.675 193.785 59.915 194.185 ;
        RECT 60.085 194.145 61.000 194.445 ;
        RECT 60.085 193.970 60.410 194.145 ;
        RECT 60.085 193.615 60.405 193.970 ;
        RECT 61.170 193.945 61.380 194.595 ;
        RECT 59.335 193.445 60.405 193.615 ;
        RECT 60.650 193.235 60.955 193.695 ;
        RECT 61.125 193.415 61.380 193.945 ;
        RECT 61.555 193.235 61.845 193.960 ;
        RECT 62.480 193.235 62.740 194.075 ;
        RECT 62.915 193.980 63.085 194.710 ;
        RECT 63.340 194.685 64.055 194.855 ;
        RECT 63.340 194.475 63.510 194.685 ;
        RECT 64.315 194.645 64.590 195.615 ;
        RECT 64.800 194.985 65.080 195.785 ;
        RECT 65.250 195.275 66.865 195.605 ;
        RECT 65.250 194.935 66.425 195.105 ;
        RECT 65.250 194.815 65.420 194.935 ;
        RECT 64.760 194.645 65.420 194.815 ;
        RECT 63.255 194.145 63.510 194.475 ;
        RECT 62.915 193.405 63.170 193.980 ;
        RECT 63.340 193.955 63.510 194.145 ;
        RECT 63.790 194.135 64.145 194.505 ;
        RECT 63.340 193.785 64.055 193.955 ;
        RECT 63.340 193.235 63.670 193.615 ;
        RECT 63.885 193.405 64.055 193.785 ;
        RECT 64.315 193.910 64.485 194.645 ;
        RECT 64.760 194.475 64.930 194.645 ;
        RECT 65.680 194.475 65.925 194.765 ;
        RECT 66.095 194.645 66.425 194.935 ;
        RECT 66.685 194.475 66.855 195.035 ;
        RECT 67.105 194.645 67.365 195.785 ;
        RECT 67.535 195.285 67.795 195.615 ;
        RECT 68.105 195.405 68.435 195.785 ;
        RECT 67.535 194.605 67.705 195.285 ;
        RECT 68.675 195.235 68.865 195.615 ;
        RECT 69.115 195.405 69.445 195.785 ;
        RECT 69.655 195.235 69.825 195.615 ;
        RECT 70.020 195.405 70.350 195.785 ;
        RECT 70.610 195.235 70.780 195.615 ;
        RECT 71.205 195.405 71.535 195.785 ;
        RECT 67.875 194.775 68.225 195.105 ;
        RECT 68.675 195.065 69.415 195.235 ;
        RECT 68.495 194.725 69.075 194.895 ;
        RECT 68.495 194.605 68.665 194.725 ;
        RECT 64.655 194.145 64.930 194.475 ;
        RECT 65.100 194.145 65.925 194.475 ;
        RECT 66.140 194.145 66.855 194.475 ;
        RECT 67.025 194.225 67.360 194.475 ;
        RECT 67.535 194.435 68.665 194.605 ;
        RECT 69.245 194.555 69.415 195.065 ;
        RECT 64.760 193.975 64.930 194.145 ;
        RECT 66.605 194.055 66.855 194.145 ;
        RECT 64.315 193.565 64.590 193.910 ;
        RECT 64.760 193.805 66.425 193.975 ;
        RECT 64.780 193.235 65.155 193.635 ;
        RECT 65.325 193.455 65.495 193.805 ;
        RECT 65.665 193.235 65.995 193.635 ;
        RECT 66.165 193.405 66.425 193.805 ;
        RECT 66.605 193.635 66.935 194.055 ;
        RECT 67.105 193.235 67.365 194.055 ;
        RECT 67.535 193.735 67.705 194.435 ;
        RECT 68.845 194.385 69.415 194.555 ;
        RECT 69.585 195.065 71.535 195.235 ;
        RECT 68.055 194.095 68.675 194.265 ;
        RECT 68.055 193.915 68.265 194.095 ;
        RECT 68.845 193.905 69.015 194.385 ;
        RECT 69.585 194.075 69.755 195.065 ;
        RECT 70.345 194.475 70.530 194.785 ;
        RECT 70.800 194.475 70.995 194.785 ;
        RECT 67.535 193.405 67.795 193.735 ;
        RECT 68.105 193.235 68.435 193.615 ;
        RECT 68.615 193.575 69.015 193.905 ;
        RECT 69.205 193.745 69.755 194.075 ;
        RECT 69.925 193.575 70.095 194.475 ;
        RECT 68.615 193.405 70.095 193.575 ;
        RECT 70.345 194.145 70.575 194.475 ;
        RECT 70.800 194.145 71.055 194.475 ;
        RECT 71.365 194.145 71.535 195.065 ;
        RECT 70.345 193.565 70.530 194.145 ;
        RECT 70.800 193.570 70.995 194.145 ;
        RECT 71.205 193.235 71.535 193.615 ;
        RECT 71.705 193.405 71.965 195.615 ;
        RECT 72.140 194.595 72.395 195.475 ;
        RECT 72.565 194.645 72.870 195.785 ;
        RECT 73.210 195.405 73.540 195.785 ;
        RECT 73.720 195.235 73.890 195.525 ;
        RECT 74.060 195.325 74.310 195.785 ;
        RECT 73.090 195.065 73.890 195.235 ;
        RECT 74.480 195.275 75.350 195.615 ;
        RECT 72.140 193.945 72.350 194.595 ;
        RECT 73.090 194.475 73.260 195.065 ;
        RECT 74.480 194.895 74.650 195.275 ;
        RECT 75.585 195.155 75.755 195.615 ;
        RECT 75.925 195.325 76.295 195.785 ;
        RECT 76.590 195.185 76.760 195.525 ;
        RECT 76.930 195.355 77.260 195.785 ;
        RECT 77.495 195.185 77.665 195.525 ;
        RECT 73.430 194.725 74.650 194.895 ;
        RECT 74.820 194.815 75.280 195.105 ;
        RECT 75.585 194.985 76.145 195.155 ;
        RECT 76.590 195.015 77.665 195.185 ;
        RECT 77.835 195.285 78.515 195.615 ;
        RECT 78.730 195.285 78.980 195.615 ;
        RECT 79.150 195.325 79.400 195.785 ;
        RECT 75.975 194.845 76.145 194.985 ;
        RECT 74.820 194.805 75.785 194.815 ;
        RECT 74.480 194.635 74.650 194.725 ;
        RECT 75.110 194.645 75.785 194.805 ;
        RECT 72.520 194.445 73.260 194.475 ;
        RECT 72.520 194.145 73.435 194.445 ;
        RECT 73.110 193.970 73.435 194.145 ;
        RECT 72.140 193.415 72.395 193.945 ;
        RECT 72.565 193.235 72.870 193.695 ;
        RECT 73.115 193.615 73.435 193.970 ;
        RECT 73.605 194.185 74.145 194.555 ;
        RECT 74.480 194.465 74.885 194.635 ;
        RECT 73.605 193.785 73.845 194.185 ;
        RECT 74.325 194.015 74.545 194.295 ;
        RECT 74.015 193.845 74.545 194.015 ;
        RECT 74.015 193.615 74.185 193.845 ;
        RECT 74.715 193.685 74.885 194.465 ;
        RECT 75.055 193.855 75.405 194.475 ;
        RECT 75.575 193.855 75.785 194.645 ;
        RECT 75.975 194.675 77.475 194.845 ;
        RECT 75.975 193.985 76.145 194.675 ;
        RECT 77.835 194.505 78.005 195.285 ;
        RECT 78.810 195.155 78.980 195.285 ;
        RECT 76.315 194.335 78.005 194.505 ;
        RECT 78.175 194.725 78.640 195.115 ;
        RECT 78.810 194.985 79.205 195.155 ;
        RECT 76.315 194.155 76.485 194.335 ;
        RECT 73.115 193.445 74.185 193.615 ;
        RECT 74.355 193.235 74.545 193.675 ;
        RECT 74.715 193.405 75.665 193.685 ;
        RECT 75.975 193.595 76.235 193.985 ;
        RECT 76.655 193.915 77.445 194.165 ;
        RECT 75.885 193.425 76.235 193.595 ;
        RECT 76.445 193.235 76.775 193.695 ;
        RECT 77.650 193.625 77.820 194.335 ;
        RECT 78.175 194.135 78.345 194.725 ;
        RECT 77.990 193.915 78.345 194.135 ;
        RECT 78.515 193.915 78.865 194.535 ;
        RECT 79.035 193.625 79.205 194.985 ;
        RECT 79.570 194.815 79.895 195.600 ;
        RECT 79.375 193.765 79.835 194.815 ;
        RECT 77.650 193.455 78.505 193.625 ;
        RECT 78.710 193.455 79.205 193.625 ;
        RECT 79.375 193.235 79.705 193.595 ;
        RECT 80.065 193.495 80.235 195.615 ;
        RECT 80.405 195.285 80.735 195.785 ;
        RECT 80.905 195.115 81.160 195.615 ;
        RECT 80.410 194.945 81.160 195.115 ;
        RECT 80.410 193.955 80.640 194.945 ;
        RECT 80.810 194.125 81.160 194.775 ;
        RECT 81.395 194.645 81.605 195.785 ;
        RECT 81.775 194.635 82.105 195.615 ;
        RECT 82.275 194.645 82.505 195.785 ;
        RECT 83.180 194.645 83.515 195.615 ;
        RECT 83.685 194.645 83.855 195.785 ;
        RECT 84.025 195.445 86.055 195.615 ;
        RECT 80.410 193.785 81.160 193.955 ;
        RECT 80.405 193.235 80.735 193.615 ;
        RECT 80.905 193.495 81.160 193.785 ;
        RECT 81.395 193.235 81.605 194.055 ;
        RECT 81.775 194.035 82.025 194.635 ;
        RECT 82.195 194.225 82.525 194.475 ;
        RECT 81.775 193.405 82.105 194.035 ;
        RECT 82.275 193.235 82.505 194.055 ;
        RECT 83.180 193.975 83.350 194.645 ;
        RECT 84.025 194.475 84.195 195.445 ;
        RECT 83.520 194.145 83.775 194.475 ;
        RECT 84.000 194.145 84.195 194.475 ;
        RECT 84.365 195.105 85.490 195.275 ;
        RECT 83.605 193.975 83.775 194.145 ;
        RECT 84.365 193.975 84.535 195.105 ;
        RECT 83.180 193.405 83.435 193.975 ;
        RECT 83.605 193.805 84.535 193.975 ;
        RECT 84.705 194.765 85.715 194.935 ;
        RECT 84.705 193.965 84.875 194.765 ;
        RECT 84.360 193.770 84.535 193.805 ;
        RECT 83.605 193.235 83.935 193.635 ;
        RECT 84.360 193.405 84.890 193.770 ;
        RECT 85.080 193.745 85.355 194.565 ;
        RECT 85.075 193.575 85.355 193.745 ;
        RECT 85.080 193.405 85.355 193.575 ;
        RECT 85.525 193.405 85.715 194.765 ;
        RECT 85.885 194.780 86.055 195.445 ;
        RECT 86.225 195.025 86.395 195.785 ;
        RECT 86.630 195.025 87.145 195.435 ;
        RECT 85.885 194.590 86.635 194.780 ;
        RECT 86.805 194.215 87.145 195.025 ;
        RECT 87.315 194.620 87.605 195.785 ;
        RECT 87.835 194.645 88.045 195.785 ;
        RECT 88.215 194.635 88.545 195.615 ;
        RECT 88.715 194.645 88.945 195.785 ;
        RECT 89.620 194.645 89.955 195.615 ;
        RECT 90.125 194.645 90.295 195.785 ;
        RECT 90.465 195.445 92.495 195.615 ;
        RECT 85.915 194.045 87.145 194.215 ;
        RECT 85.895 193.235 86.405 193.770 ;
        RECT 86.625 193.440 86.870 194.045 ;
        RECT 87.315 193.235 87.605 193.960 ;
        RECT 87.835 193.235 88.045 194.055 ;
        RECT 88.215 194.035 88.465 194.635 ;
        RECT 88.635 194.225 88.965 194.475 ;
        RECT 88.215 193.405 88.545 194.035 ;
        RECT 88.715 193.235 88.945 194.055 ;
        RECT 89.620 193.975 89.790 194.645 ;
        RECT 90.465 194.475 90.635 195.445 ;
        RECT 89.960 194.145 90.215 194.475 ;
        RECT 90.440 194.145 90.635 194.475 ;
        RECT 90.805 195.105 91.930 195.275 ;
        RECT 90.045 193.975 90.215 194.145 ;
        RECT 90.805 193.975 90.975 195.105 ;
        RECT 89.620 193.405 89.875 193.975 ;
        RECT 90.045 193.805 90.975 193.975 ;
        RECT 91.145 194.765 92.155 194.935 ;
        RECT 91.145 193.965 91.315 194.765 ;
        RECT 91.520 194.425 91.795 194.565 ;
        RECT 91.515 194.255 91.795 194.425 ;
        RECT 90.800 193.770 90.975 193.805 ;
        RECT 90.045 193.235 90.375 193.635 ;
        RECT 90.800 193.405 91.330 193.770 ;
        RECT 91.520 193.405 91.795 194.255 ;
        RECT 91.965 193.405 92.155 194.765 ;
        RECT 92.325 194.780 92.495 195.445 ;
        RECT 92.665 195.025 92.835 195.785 ;
        RECT 93.070 195.025 93.585 195.435 ;
        RECT 92.325 194.590 93.075 194.780 ;
        RECT 93.245 194.215 93.585 195.025 ;
        RECT 92.355 194.045 93.585 194.215 ;
        RECT 93.755 194.645 94.095 195.615 ;
        RECT 94.265 194.645 94.435 195.785 ;
        RECT 94.705 194.985 94.955 195.785 ;
        RECT 95.600 194.815 95.930 195.615 ;
        RECT 96.230 194.985 96.560 195.785 ;
        RECT 96.730 194.815 97.060 195.615 ;
        RECT 94.625 194.645 97.060 194.815 ;
        RECT 97.440 194.645 97.775 195.615 ;
        RECT 97.945 194.645 98.115 195.785 ;
        RECT 98.285 195.445 100.315 195.615 ;
        RECT 92.335 193.235 92.845 193.770 ;
        RECT 93.065 193.440 93.310 194.045 ;
        RECT 93.755 194.035 93.930 194.645 ;
        RECT 94.625 194.395 94.795 194.645 ;
        RECT 94.100 194.225 94.795 194.395 ;
        RECT 94.970 194.225 95.390 194.425 ;
        RECT 95.560 194.225 95.890 194.425 ;
        RECT 96.060 194.225 96.390 194.425 ;
        RECT 93.755 193.405 94.095 194.035 ;
        RECT 94.265 193.235 94.515 194.035 ;
        RECT 94.705 193.885 95.930 194.055 ;
        RECT 94.705 193.405 95.035 193.885 ;
        RECT 95.205 193.235 95.430 193.695 ;
        RECT 95.600 193.405 95.930 193.885 ;
        RECT 96.560 194.015 96.730 194.645 ;
        RECT 96.915 194.225 97.265 194.475 ;
        RECT 96.560 193.405 97.060 194.015 ;
        RECT 97.440 193.975 97.610 194.645 ;
        RECT 98.285 194.475 98.455 195.445 ;
        RECT 97.780 194.145 98.035 194.475 ;
        RECT 98.260 194.145 98.455 194.475 ;
        RECT 98.625 195.105 99.750 195.275 ;
        RECT 97.865 193.975 98.035 194.145 ;
        RECT 98.625 193.975 98.795 195.105 ;
        RECT 97.440 193.405 97.695 193.975 ;
        RECT 97.865 193.805 98.795 193.975 ;
        RECT 98.965 194.765 99.975 194.935 ;
        RECT 98.965 193.965 99.135 194.765 ;
        RECT 99.340 194.425 99.615 194.565 ;
        RECT 99.335 194.255 99.615 194.425 ;
        RECT 98.620 193.770 98.795 193.805 ;
        RECT 97.865 193.235 98.195 193.635 ;
        RECT 98.620 193.405 99.150 193.770 ;
        RECT 99.340 193.405 99.615 194.255 ;
        RECT 99.785 193.405 99.975 194.765 ;
        RECT 100.145 194.780 100.315 195.445 ;
        RECT 100.485 195.025 100.655 195.785 ;
        RECT 100.890 195.025 101.405 195.435 ;
        RECT 100.145 194.590 100.895 194.780 ;
        RECT 101.065 194.215 101.405 195.025 ;
        RECT 100.175 194.045 101.405 194.215 ;
        RECT 101.580 194.645 101.915 195.615 ;
        RECT 102.085 194.645 102.255 195.785 ;
        RECT 102.425 195.445 104.455 195.615 ;
        RECT 100.155 193.235 100.665 193.770 ;
        RECT 100.885 193.440 101.130 194.045 ;
        RECT 101.580 193.975 101.750 194.645 ;
        RECT 102.425 194.475 102.595 195.445 ;
        RECT 101.920 194.145 102.175 194.475 ;
        RECT 102.400 194.145 102.595 194.475 ;
        RECT 102.765 195.105 103.890 195.275 ;
        RECT 102.005 193.975 102.175 194.145 ;
        RECT 102.765 193.975 102.935 195.105 ;
        RECT 101.580 193.405 101.835 193.975 ;
        RECT 102.005 193.805 102.935 193.975 ;
        RECT 103.105 194.765 104.115 194.935 ;
        RECT 103.105 193.965 103.275 194.765 ;
        RECT 102.760 193.770 102.935 193.805 ;
        RECT 102.005 193.235 102.335 193.635 ;
        RECT 102.760 193.405 103.290 193.770 ;
        RECT 103.480 193.745 103.755 194.565 ;
        RECT 103.475 193.575 103.755 193.745 ;
        RECT 103.480 193.405 103.755 193.575 ;
        RECT 103.925 193.405 104.115 194.765 ;
        RECT 104.285 194.780 104.455 195.445 ;
        RECT 104.625 195.025 104.795 195.785 ;
        RECT 105.030 195.025 105.545 195.435 ;
        RECT 104.285 194.590 105.035 194.780 ;
        RECT 105.205 194.215 105.545 195.025 ;
        RECT 104.315 194.045 105.545 194.215 ;
        RECT 105.715 194.645 106.055 195.615 ;
        RECT 106.225 194.645 106.395 195.785 ;
        RECT 106.665 194.985 106.915 195.785 ;
        RECT 107.560 194.815 107.890 195.615 ;
        RECT 108.190 194.985 108.520 195.785 ;
        RECT 108.690 194.815 109.020 195.615 ;
        RECT 106.585 194.645 109.020 194.815 ;
        RECT 109.395 194.710 109.665 195.615 ;
        RECT 109.835 195.025 110.165 195.785 ;
        RECT 110.345 194.855 110.515 195.615 ;
        RECT 104.295 193.235 104.805 193.770 ;
        RECT 105.025 193.440 105.270 194.045 ;
        RECT 105.715 194.035 105.890 194.645 ;
        RECT 106.585 194.395 106.755 194.645 ;
        RECT 106.060 194.225 106.755 194.395 ;
        RECT 106.930 194.225 107.350 194.425 ;
        RECT 107.520 194.225 107.850 194.425 ;
        RECT 108.020 194.225 108.350 194.425 ;
        RECT 105.715 193.405 106.055 194.035 ;
        RECT 106.225 193.235 106.475 194.035 ;
        RECT 106.665 193.885 107.890 194.055 ;
        RECT 106.665 193.405 106.995 193.885 ;
        RECT 107.165 193.235 107.390 193.695 ;
        RECT 107.560 193.405 107.890 193.885 ;
        RECT 108.520 194.015 108.690 194.645 ;
        RECT 108.875 194.225 109.225 194.475 ;
        RECT 108.520 193.405 109.020 194.015 ;
        RECT 109.395 193.910 109.565 194.710 ;
        RECT 109.850 194.685 110.515 194.855 ;
        RECT 109.850 194.540 110.020 194.685 ;
        RECT 110.835 194.645 111.045 195.785 ;
        RECT 109.735 194.210 110.020 194.540 ;
        RECT 111.215 194.635 111.545 195.615 ;
        RECT 111.715 194.645 111.945 195.785 ;
        RECT 112.155 194.695 113.365 195.785 ;
        RECT 109.850 193.955 110.020 194.210 ;
        RECT 110.255 194.135 110.585 194.505 ;
        RECT 109.395 193.405 109.655 193.910 ;
        RECT 109.850 193.785 110.515 193.955 ;
        RECT 109.835 193.235 110.165 193.615 ;
        RECT 110.345 193.405 110.515 193.785 ;
        RECT 110.835 193.235 111.045 194.055 ;
        RECT 111.215 194.035 111.465 194.635 ;
        RECT 111.635 194.225 111.965 194.475 ;
        RECT 112.155 194.155 112.675 194.695 ;
        RECT 111.215 193.405 111.545 194.035 ;
        RECT 111.715 193.235 111.945 194.055 ;
        RECT 112.845 193.985 113.365 194.525 ;
        RECT 112.155 193.235 113.365 193.985 ;
        RECT 26.970 193.065 113.450 193.235 ;
        RECT 27.055 192.315 28.265 193.065 ;
        RECT 28.985 192.515 29.155 192.895 ;
        RECT 29.335 192.685 29.665 193.065 ;
        RECT 28.985 192.345 29.650 192.515 ;
        RECT 29.845 192.390 30.105 192.895 ;
        RECT 27.055 191.775 27.575 192.315 ;
        RECT 27.745 191.605 28.265 192.145 ;
        RECT 28.915 191.795 29.245 192.165 ;
        RECT 29.480 192.090 29.650 192.345 ;
        RECT 29.480 191.760 29.765 192.090 ;
        RECT 29.480 191.615 29.650 191.760 ;
        RECT 27.055 190.515 28.265 191.605 ;
        RECT 28.985 191.445 29.650 191.615 ;
        RECT 29.935 191.590 30.105 192.390 ;
        RECT 28.985 190.685 29.155 191.445 ;
        RECT 29.335 190.515 29.665 191.275 ;
        RECT 29.835 190.685 30.105 191.590 ;
        RECT 31.570 192.355 31.825 192.885 ;
        RECT 32.005 192.605 32.290 193.065 ;
        RECT 31.570 191.495 31.750 192.355 ;
        RECT 32.470 192.155 32.720 192.805 ;
        RECT 31.920 191.825 32.720 192.155 ;
        RECT 31.570 191.025 31.825 191.495 ;
        RECT 31.485 190.855 31.825 191.025 ;
        RECT 31.570 190.825 31.825 190.855 ;
        RECT 32.005 190.515 32.290 191.315 ;
        RECT 32.470 191.235 32.720 191.825 ;
        RECT 32.920 192.470 33.240 192.800 ;
        RECT 33.420 192.585 34.080 193.065 ;
        RECT 34.280 192.675 35.130 192.845 ;
        RECT 32.920 191.575 33.110 192.470 ;
        RECT 33.430 192.145 34.090 192.415 ;
        RECT 33.760 192.085 34.090 192.145 ;
        RECT 33.280 191.915 33.610 191.975 ;
        RECT 34.280 191.915 34.450 192.675 ;
        RECT 35.690 192.605 36.010 193.065 ;
        RECT 36.210 192.425 36.460 192.855 ;
        RECT 36.750 192.625 37.160 193.065 ;
        RECT 37.330 192.685 38.345 192.885 ;
        RECT 34.620 192.255 35.870 192.425 ;
        RECT 34.620 192.135 34.950 192.255 ;
        RECT 33.280 191.745 35.180 191.915 ;
        RECT 32.920 191.405 34.840 191.575 ;
        RECT 32.920 191.385 33.240 191.405 ;
        RECT 32.470 190.725 32.800 191.235 ;
        RECT 33.070 190.775 33.240 191.385 ;
        RECT 35.010 191.235 35.180 191.745 ;
        RECT 35.350 191.675 35.530 192.085 ;
        RECT 35.700 191.495 35.870 192.255 ;
        RECT 33.410 190.515 33.740 191.205 ;
        RECT 33.970 191.065 35.180 191.235 ;
        RECT 35.350 191.185 35.870 191.495 ;
        RECT 36.040 192.085 36.460 192.425 ;
        RECT 36.750 192.085 37.160 192.415 ;
        RECT 36.040 191.315 36.230 192.085 ;
        RECT 37.330 191.955 37.500 192.685 ;
        RECT 38.645 192.515 38.815 192.845 ;
        RECT 38.985 192.685 39.315 193.065 ;
        RECT 37.670 192.135 38.020 192.505 ;
        RECT 37.330 191.915 37.750 191.955 ;
        RECT 36.400 191.745 37.750 191.915 ;
        RECT 36.400 191.585 36.650 191.745 ;
        RECT 37.160 191.315 37.410 191.575 ;
        RECT 36.040 191.065 37.410 191.315 ;
        RECT 33.970 190.775 34.210 191.065 ;
        RECT 35.010 190.985 35.180 191.065 ;
        RECT 34.410 190.515 34.830 190.895 ;
        RECT 35.010 190.735 35.640 190.985 ;
        RECT 36.110 190.515 36.440 190.895 ;
        RECT 36.610 190.775 36.780 191.065 ;
        RECT 37.580 190.900 37.750 191.745 ;
        RECT 38.200 191.575 38.420 192.445 ;
        RECT 38.645 192.325 39.340 192.515 ;
        RECT 37.920 191.195 38.420 191.575 ;
        RECT 38.590 191.525 39.000 192.145 ;
        RECT 39.170 191.355 39.340 192.325 ;
        RECT 38.645 191.185 39.340 191.355 ;
        RECT 36.960 190.515 37.340 190.895 ;
        RECT 37.580 190.730 38.410 190.900 ;
        RECT 38.645 190.685 38.815 191.185 ;
        RECT 38.985 190.515 39.315 191.015 ;
        RECT 39.530 190.685 39.755 192.805 ;
        RECT 39.925 192.685 40.255 193.065 ;
        RECT 40.425 192.515 40.595 192.805 ;
        RECT 39.930 192.345 40.595 192.515 ;
        RECT 40.945 192.515 41.115 192.895 ;
        RECT 41.295 192.685 41.625 193.065 ;
        RECT 40.945 192.345 41.610 192.515 ;
        RECT 41.805 192.390 42.065 192.895 ;
        RECT 39.930 191.355 40.160 192.345 ;
        RECT 40.330 191.525 40.680 192.175 ;
        RECT 40.875 191.795 41.205 192.165 ;
        RECT 41.440 192.090 41.610 192.345 ;
        RECT 41.440 191.760 41.725 192.090 ;
        RECT 41.440 191.615 41.610 191.760 ;
        RECT 40.945 191.445 41.610 191.615 ;
        RECT 41.895 191.590 42.065 192.390 ;
        RECT 42.325 192.515 42.495 192.895 ;
        RECT 42.675 192.685 43.005 193.065 ;
        RECT 42.325 192.345 42.990 192.515 ;
        RECT 43.185 192.390 43.445 192.895 ;
        RECT 42.255 191.795 42.585 192.165 ;
        RECT 42.820 192.090 42.990 192.345 ;
        RECT 42.820 191.760 43.105 192.090 ;
        RECT 42.820 191.615 42.990 191.760 ;
        RECT 39.930 191.185 40.595 191.355 ;
        RECT 39.925 190.515 40.255 191.015 ;
        RECT 40.425 190.685 40.595 191.185 ;
        RECT 40.945 190.685 41.115 191.445 ;
        RECT 41.295 190.515 41.625 191.275 ;
        RECT 41.795 190.685 42.065 191.590 ;
        RECT 42.325 191.445 42.990 191.615 ;
        RECT 43.275 191.590 43.445 192.390 ;
        RECT 42.325 190.685 42.495 191.445 ;
        RECT 42.675 190.515 43.005 191.275 ;
        RECT 43.175 190.685 43.445 191.590 ;
        RECT 43.620 192.325 43.875 192.895 ;
        RECT 44.045 192.665 44.375 193.065 ;
        RECT 44.800 192.530 45.330 192.895 ;
        RECT 44.800 192.495 44.975 192.530 ;
        RECT 44.045 192.325 44.975 192.495 ;
        RECT 43.620 191.655 43.790 192.325 ;
        RECT 44.045 192.155 44.215 192.325 ;
        RECT 43.960 191.825 44.215 192.155 ;
        RECT 44.440 191.825 44.635 192.155 ;
        RECT 43.620 190.685 43.955 191.655 ;
        RECT 44.125 190.515 44.295 191.655 ;
        RECT 44.465 190.855 44.635 191.825 ;
        RECT 44.805 191.195 44.975 192.325 ;
        RECT 45.145 191.535 45.315 192.335 ;
        RECT 45.520 192.045 45.795 192.895 ;
        RECT 45.515 191.875 45.795 192.045 ;
        RECT 45.520 191.735 45.795 191.875 ;
        RECT 45.965 191.535 46.155 192.895 ;
        RECT 46.335 192.530 46.845 193.065 ;
        RECT 47.065 192.255 47.310 192.860 ;
        RECT 48.675 192.340 48.965 193.065 ;
        RECT 46.355 192.085 47.585 192.255 ;
        RECT 49.175 192.245 49.405 193.065 ;
        RECT 49.575 192.265 49.905 192.895 ;
        RECT 45.145 191.365 46.155 191.535 ;
        RECT 46.325 191.520 47.075 191.710 ;
        RECT 44.805 191.025 45.930 191.195 ;
        RECT 46.325 190.855 46.495 191.520 ;
        RECT 47.245 191.275 47.585 192.085 ;
        RECT 49.155 191.825 49.485 192.075 ;
        RECT 44.465 190.685 46.495 190.855 ;
        RECT 46.665 190.515 46.835 191.275 ;
        RECT 47.070 190.865 47.585 191.275 ;
        RECT 48.675 190.515 48.965 191.680 ;
        RECT 49.655 191.665 49.905 192.265 ;
        RECT 50.075 192.245 50.285 193.065 ;
        RECT 50.515 192.565 50.775 192.895 ;
        RECT 50.985 192.585 51.260 193.065 ;
        RECT 49.175 190.515 49.405 191.655 ;
        RECT 49.575 190.685 49.905 191.665 ;
        RECT 50.515 191.655 50.685 192.565 ;
        RECT 51.470 192.495 51.675 192.895 ;
        RECT 51.845 192.665 52.180 193.065 ;
        RECT 50.855 191.825 51.215 192.405 ;
        RECT 51.470 192.325 52.155 192.495 ;
        RECT 51.395 191.655 51.645 192.155 ;
        RECT 50.075 190.515 50.285 191.655 ;
        RECT 50.515 191.485 51.645 191.655 ;
        RECT 50.515 190.715 50.785 191.485 ;
        RECT 51.815 191.295 52.155 192.325 ;
        RECT 50.955 190.515 51.285 191.295 ;
        RECT 51.490 191.120 52.155 191.295 ;
        RECT 52.360 192.325 52.615 192.895 ;
        RECT 52.785 192.665 53.115 193.065 ;
        RECT 53.540 192.530 54.070 192.895 ;
        RECT 54.260 192.725 54.535 192.895 ;
        RECT 54.255 192.555 54.535 192.725 ;
        RECT 53.540 192.495 53.715 192.530 ;
        RECT 52.785 192.325 53.715 192.495 ;
        RECT 52.360 191.655 52.530 192.325 ;
        RECT 52.785 192.155 52.955 192.325 ;
        RECT 52.700 191.825 52.955 192.155 ;
        RECT 53.180 191.825 53.375 192.155 ;
        RECT 51.490 190.715 51.675 191.120 ;
        RECT 51.845 190.515 52.180 190.940 ;
        RECT 52.360 190.685 52.695 191.655 ;
        RECT 52.865 190.515 53.035 191.655 ;
        RECT 53.205 190.855 53.375 191.825 ;
        RECT 53.545 191.195 53.715 192.325 ;
        RECT 53.885 191.535 54.055 192.335 ;
        RECT 54.260 191.735 54.535 192.555 ;
        RECT 54.705 191.535 54.895 192.895 ;
        RECT 55.075 192.530 55.585 193.065 ;
        RECT 55.805 192.255 56.050 192.860 ;
        RECT 56.960 192.515 57.215 192.805 ;
        RECT 57.385 192.685 57.715 193.065 ;
        RECT 56.960 192.345 57.710 192.515 ;
        RECT 55.095 192.085 56.325 192.255 ;
        RECT 53.885 191.365 54.895 191.535 ;
        RECT 55.065 191.520 55.815 191.710 ;
        RECT 53.545 191.025 54.670 191.195 ;
        RECT 55.065 190.855 55.235 191.520 ;
        RECT 55.985 191.275 56.325 192.085 ;
        RECT 56.960 191.525 57.310 192.175 ;
        RECT 57.480 191.355 57.710 192.345 ;
        RECT 53.205 190.685 55.235 190.855 ;
        RECT 55.405 190.515 55.575 191.275 ;
        RECT 55.810 190.865 56.325 191.275 ;
        RECT 56.960 191.185 57.710 191.355 ;
        RECT 56.960 190.685 57.215 191.185 ;
        RECT 57.385 190.515 57.715 191.015 ;
        RECT 57.885 190.685 58.055 192.805 ;
        RECT 58.415 192.705 58.745 193.065 ;
        RECT 58.915 192.675 59.410 192.845 ;
        RECT 59.615 192.675 60.470 192.845 ;
        RECT 58.285 191.485 58.745 192.535 ;
        RECT 58.225 190.700 58.550 191.485 ;
        RECT 58.915 191.315 59.085 192.675 ;
        RECT 59.255 191.765 59.605 192.385 ;
        RECT 59.775 192.165 60.130 192.385 ;
        RECT 59.775 191.575 59.945 192.165 ;
        RECT 60.300 191.965 60.470 192.675 ;
        RECT 61.345 192.605 61.675 193.065 ;
        RECT 61.885 192.705 62.235 192.875 ;
        RECT 60.675 192.135 61.465 192.385 ;
        RECT 61.885 192.315 62.145 192.705 ;
        RECT 62.455 192.615 63.405 192.895 ;
        RECT 63.575 192.625 63.765 193.065 ;
        RECT 63.935 192.685 65.005 192.855 ;
        RECT 61.635 191.965 61.805 192.145 ;
        RECT 58.915 191.145 59.310 191.315 ;
        RECT 59.480 191.185 59.945 191.575 ;
        RECT 60.115 191.795 61.805 191.965 ;
        RECT 59.140 191.015 59.310 191.145 ;
        RECT 60.115 191.015 60.285 191.795 ;
        RECT 61.975 191.625 62.145 192.315 ;
        RECT 60.645 191.455 62.145 191.625 ;
        RECT 62.335 191.655 62.545 192.445 ;
        RECT 62.715 191.825 63.065 192.445 ;
        RECT 63.235 191.835 63.405 192.615 ;
        RECT 63.935 192.455 64.105 192.685 ;
        RECT 63.575 192.285 64.105 192.455 ;
        RECT 63.575 192.005 63.795 192.285 ;
        RECT 64.275 192.115 64.515 192.515 ;
        RECT 63.235 191.665 63.640 191.835 ;
        RECT 63.975 191.745 64.515 192.115 ;
        RECT 64.685 192.330 65.005 192.685 ;
        RECT 65.250 192.605 65.555 193.065 ;
        RECT 65.725 192.355 65.980 192.885 ;
        RECT 64.685 192.155 65.010 192.330 ;
        RECT 64.685 191.855 65.600 192.155 ;
        RECT 64.860 191.825 65.600 191.855 ;
        RECT 62.335 191.495 63.010 191.655 ;
        RECT 63.470 191.575 63.640 191.665 ;
        RECT 62.335 191.485 63.300 191.495 ;
        RECT 61.975 191.315 62.145 191.455 ;
        RECT 58.720 190.515 58.970 190.975 ;
        RECT 59.140 190.685 59.390 191.015 ;
        RECT 59.605 190.685 60.285 191.015 ;
        RECT 60.455 191.115 61.530 191.285 ;
        RECT 61.975 191.145 62.535 191.315 ;
        RECT 62.840 191.195 63.300 191.485 ;
        RECT 63.470 191.405 64.690 191.575 ;
        RECT 60.455 190.775 60.625 191.115 ;
        RECT 60.860 190.515 61.190 190.945 ;
        RECT 61.360 190.775 61.530 191.115 ;
        RECT 61.825 190.515 62.195 190.975 ;
        RECT 62.365 190.685 62.535 191.145 ;
        RECT 63.470 191.025 63.640 191.405 ;
        RECT 64.860 191.235 65.030 191.825 ;
        RECT 65.770 191.705 65.980 192.355 ;
        RECT 62.770 190.685 63.640 191.025 ;
        RECT 64.230 191.065 65.030 191.235 ;
        RECT 63.810 190.515 64.060 190.975 ;
        RECT 64.230 190.775 64.400 191.065 ;
        RECT 64.580 190.515 64.910 190.895 ;
        RECT 65.250 190.515 65.555 191.655 ;
        RECT 65.725 190.825 65.980 191.705 ;
        RECT 66.155 192.415 66.415 192.895 ;
        RECT 66.585 192.525 66.835 193.065 ;
        RECT 66.155 191.385 66.325 192.415 ;
        RECT 67.005 192.360 67.225 192.845 ;
        RECT 66.495 191.765 66.725 192.160 ;
        RECT 66.895 191.935 67.225 192.360 ;
        RECT 67.395 192.685 68.285 192.855 ;
        RECT 67.395 191.960 67.565 192.685 ;
        RECT 67.735 192.130 68.285 192.515 ;
        RECT 68.545 192.415 68.715 192.895 ;
        RECT 68.895 192.585 69.135 193.065 ;
        RECT 69.385 192.415 69.555 192.895 ;
        RECT 69.725 192.585 70.055 193.065 ;
        RECT 70.225 192.415 70.395 192.895 ;
        RECT 68.545 192.245 69.180 192.415 ;
        RECT 69.385 192.245 70.395 192.415 ;
        RECT 70.565 192.265 70.895 193.065 ;
        RECT 71.485 192.670 71.815 193.065 ;
        RECT 71.985 192.495 72.185 192.850 ;
        RECT 72.355 192.665 72.685 193.065 ;
        RECT 72.855 192.495 73.055 192.840 ;
        RECT 71.215 192.325 73.055 192.495 ;
        RECT 73.225 192.325 73.555 193.065 ;
        RECT 73.790 192.495 73.960 192.745 ;
        RECT 73.790 192.325 74.265 192.495 ;
        RECT 74.435 192.340 74.725 193.065 ;
        RECT 69.010 192.075 69.180 192.245 ;
        RECT 69.895 192.215 70.395 192.245 ;
        RECT 67.395 191.890 68.285 191.960 ;
        RECT 67.390 191.865 68.285 191.890 ;
        RECT 67.380 191.850 68.285 191.865 ;
        RECT 67.375 191.835 68.285 191.850 ;
        RECT 68.460 191.835 68.840 192.075 ;
        RECT 69.010 191.905 69.510 192.075 ;
        RECT 67.365 191.830 68.285 191.835 ;
        RECT 67.360 191.820 68.285 191.830 ;
        RECT 67.355 191.810 68.285 191.820 ;
        RECT 67.345 191.805 68.285 191.810 ;
        RECT 67.335 191.795 68.285 191.805 ;
        RECT 67.325 191.790 68.285 191.795 ;
        RECT 67.325 191.785 67.660 191.790 ;
        RECT 67.310 191.780 67.660 191.785 ;
        RECT 67.295 191.770 67.660 191.780 ;
        RECT 67.270 191.765 67.660 191.770 ;
        RECT 66.495 191.760 67.660 191.765 ;
        RECT 66.495 191.725 67.630 191.760 ;
        RECT 66.495 191.700 67.595 191.725 ;
        RECT 66.495 191.670 67.565 191.700 ;
        RECT 66.495 191.640 67.545 191.670 ;
        RECT 66.495 191.610 67.525 191.640 ;
        RECT 66.495 191.600 67.455 191.610 ;
        RECT 66.495 191.590 67.430 191.600 ;
        RECT 66.495 191.575 67.410 191.590 ;
        RECT 66.495 191.560 67.390 191.575 ;
        RECT 66.600 191.550 67.385 191.560 ;
        RECT 66.600 191.515 67.370 191.550 ;
        RECT 66.155 190.685 66.430 191.385 ;
        RECT 66.600 191.265 67.355 191.515 ;
        RECT 67.525 191.195 67.855 191.440 ;
        RECT 68.025 191.340 68.285 191.790 ;
        RECT 69.010 191.665 69.180 191.905 ;
        RECT 69.900 191.705 70.395 192.215 ;
        RECT 68.465 191.495 69.180 191.665 ;
        RECT 69.385 191.535 70.395 191.705 ;
        RECT 67.670 191.170 67.855 191.195 ;
        RECT 67.670 191.070 68.285 191.170 ;
        RECT 66.600 190.515 66.855 191.060 ;
        RECT 67.025 190.685 67.505 191.025 ;
        RECT 67.680 190.515 68.285 191.070 ;
        RECT 68.465 190.685 68.795 191.495 ;
        RECT 68.965 190.515 69.205 191.315 ;
        RECT 69.385 190.685 69.555 191.535 ;
        RECT 69.725 190.515 70.055 191.315 ;
        RECT 70.225 190.685 70.395 191.535 ;
        RECT 70.565 190.515 70.895 191.665 ;
        RECT 71.215 190.700 71.475 192.325 ;
        RECT 71.655 191.355 71.875 192.155 ;
        RECT 72.115 191.535 72.415 192.155 ;
        RECT 72.585 191.535 72.915 192.155 ;
        RECT 73.085 191.535 73.405 192.155 ;
        RECT 73.575 191.535 73.925 192.155 ;
        RECT 74.095 191.355 74.265 192.325 ;
        RECT 74.895 192.325 75.280 192.895 ;
        RECT 75.450 192.605 75.775 193.065 ;
        RECT 76.295 192.435 76.575 192.895 ;
        RECT 71.655 191.145 74.265 191.355 ;
        RECT 73.225 190.515 73.555 190.965 ;
        RECT 74.435 190.515 74.725 191.680 ;
        RECT 74.895 191.655 75.175 192.325 ;
        RECT 75.450 192.265 76.575 192.435 ;
        RECT 75.450 192.155 75.900 192.265 ;
        RECT 75.345 191.825 75.900 192.155 ;
        RECT 76.765 192.095 77.165 192.895 ;
        RECT 77.565 192.605 77.835 193.065 ;
        RECT 78.005 192.435 78.290 192.895 ;
        RECT 74.895 190.685 75.280 191.655 ;
        RECT 75.450 191.365 75.900 191.825 ;
        RECT 76.070 191.535 77.165 192.095 ;
        RECT 75.450 191.145 76.575 191.365 ;
        RECT 75.450 190.515 75.775 190.975 ;
        RECT 76.295 190.685 76.575 191.145 ;
        RECT 76.765 190.685 77.165 191.535 ;
        RECT 77.335 192.265 78.290 192.435 ;
        RECT 78.690 192.435 78.975 192.895 ;
        RECT 79.145 192.605 79.415 193.065 ;
        RECT 78.690 192.265 79.645 192.435 ;
        RECT 77.335 191.365 77.545 192.265 ;
        RECT 77.715 191.535 78.405 192.095 ;
        RECT 78.575 191.535 79.265 192.095 ;
        RECT 79.435 191.365 79.645 192.265 ;
        RECT 77.335 191.145 78.290 191.365 ;
        RECT 77.565 190.515 77.835 190.975 ;
        RECT 78.005 190.685 78.290 191.145 ;
        RECT 78.690 191.145 79.645 191.365 ;
        RECT 79.815 192.095 80.215 192.895 ;
        RECT 80.405 192.435 80.685 192.895 ;
        RECT 81.205 192.605 81.530 193.065 ;
        RECT 80.405 192.265 81.530 192.435 ;
        RECT 81.700 192.325 82.085 192.895 ;
        RECT 81.080 192.155 81.530 192.265 ;
        RECT 79.815 191.535 80.910 192.095 ;
        RECT 81.080 191.825 81.635 192.155 ;
        RECT 78.690 190.685 78.975 191.145 ;
        RECT 79.145 190.515 79.415 190.975 ;
        RECT 79.815 190.685 80.215 191.535 ;
        RECT 81.080 191.365 81.530 191.825 ;
        RECT 81.805 191.655 82.085 192.325 ;
        RECT 80.405 191.145 81.530 191.365 ;
        RECT 80.405 190.685 80.685 191.145 ;
        RECT 81.205 190.515 81.530 190.975 ;
        RECT 81.700 190.685 82.085 191.655 ;
        RECT 82.630 192.355 82.885 192.885 ;
        RECT 83.065 192.605 83.350 193.065 ;
        RECT 82.630 191.495 82.810 192.355 ;
        RECT 83.530 192.155 83.780 192.805 ;
        RECT 82.980 191.825 83.780 192.155 ;
        RECT 82.630 191.025 82.885 191.495 ;
        RECT 82.545 190.855 82.885 191.025 ;
        RECT 82.630 190.825 82.885 190.855 ;
        RECT 83.065 190.515 83.350 191.315 ;
        RECT 83.530 191.235 83.780 191.825 ;
        RECT 83.980 192.470 84.300 192.800 ;
        RECT 84.480 192.585 85.140 193.065 ;
        RECT 85.340 192.675 86.190 192.845 ;
        RECT 83.980 191.575 84.170 192.470 ;
        RECT 84.490 192.145 85.150 192.415 ;
        RECT 84.820 192.085 85.150 192.145 ;
        RECT 84.340 191.915 84.670 191.975 ;
        RECT 85.340 191.915 85.510 192.675 ;
        RECT 86.750 192.605 87.070 193.065 ;
        RECT 87.270 192.425 87.520 192.855 ;
        RECT 87.810 192.625 88.220 193.065 ;
        RECT 88.390 192.685 89.405 192.885 ;
        RECT 85.680 192.255 86.930 192.425 ;
        RECT 85.680 192.135 86.010 192.255 ;
        RECT 84.340 191.745 86.240 191.915 ;
        RECT 83.980 191.405 85.900 191.575 ;
        RECT 83.980 191.385 84.300 191.405 ;
        RECT 83.530 190.725 83.860 191.235 ;
        RECT 84.130 190.775 84.300 191.385 ;
        RECT 86.070 191.235 86.240 191.745 ;
        RECT 86.410 191.675 86.590 192.085 ;
        RECT 86.760 191.495 86.930 192.255 ;
        RECT 84.470 190.515 84.800 191.205 ;
        RECT 85.030 191.065 86.240 191.235 ;
        RECT 86.410 191.185 86.930 191.495 ;
        RECT 87.100 192.085 87.520 192.425 ;
        RECT 87.810 192.085 88.220 192.415 ;
        RECT 87.100 191.315 87.290 192.085 ;
        RECT 88.390 191.955 88.560 192.685 ;
        RECT 89.705 192.515 89.875 192.845 ;
        RECT 90.045 192.685 90.375 193.065 ;
        RECT 88.730 192.135 89.080 192.505 ;
        RECT 88.390 191.915 88.810 191.955 ;
        RECT 87.460 191.745 88.810 191.915 ;
        RECT 87.460 191.585 87.710 191.745 ;
        RECT 88.220 191.315 88.470 191.575 ;
        RECT 87.100 191.065 88.470 191.315 ;
        RECT 85.030 190.775 85.270 191.065 ;
        RECT 86.070 190.985 86.240 191.065 ;
        RECT 85.470 190.515 85.890 190.895 ;
        RECT 86.070 190.735 86.700 190.985 ;
        RECT 87.170 190.515 87.500 190.895 ;
        RECT 87.670 190.775 87.840 191.065 ;
        RECT 88.640 190.900 88.810 191.745 ;
        RECT 89.260 191.575 89.480 192.445 ;
        RECT 89.705 192.325 90.400 192.515 ;
        RECT 88.980 191.195 89.480 191.575 ;
        RECT 89.650 191.525 90.060 192.145 ;
        RECT 90.230 191.355 90.400 192.325 ;
        RECT 89.705 191.185 90.400 191.355 ;
        RECT 88.020 190.515 88.400 190.895 ;
        RECT 88.640 190.730 89.470 190.900 ;
        RECT 89.705 190.685 89.875 191.185 ;
        RECT 90.045 190.515 90.375 191.015 ;
        RECT 90.590 190.685 90.815 192.805 ;
        RECT 90.985 192.685 91.315 193.065 ;
        RECT 91.485 192.515 91.655 192.805 ;
        RECT 90.990 192.345 91.655 192.515 ;
        RECT 90.990 191.355 91.220 192.345 ;
        RECT 93.110 192.255 93.355 192.860 ;
        RECT 93.575 192.530 94.085 193.065 ;
        RECT 91.390 191.525 91.740 192.175 ;
        RECT 92.835 192.085 94.065 192.255 ;
        RECT 90.990 191.185 91.655 191.355 ;
        RECT 90.985 190.515 91.315 191.015 ;
        RECT 91.485 190.685 91.655 191.185 ;
        RECT 92.835 191.275 93.175 192.085 ;
        RECT 93.345 191.520 94.095 191.710 ;
        RECT 92.835 190.865 93.350 191.275 ;
        RECT 93.585 190.515 93.755 191.275 ;
        RECT 93.925 190.855 94.095 191.520 ;
        RECT 94.265 191.535 94.455 192.895 ;
        RECT 94.625 192.045 94.900 192.895 ;
        RECT 95.090 192.530 95.620 192.895 ;
        RECT 96.045 192.665 96.375 193.065 ;
        RECT 95.445 192.495 95.620 192.530 ;
        RECT 94.625 191.875 94.905 192.045 ;
        RECT 94.625 191.735 94.900 191.875 ;
        RECT 95.105 191.535 95.275 192.335 ;
        RECT 94.265 191.365 95.275 191.535 ;
        RECT 95.445 192.325 96.375 192.495 ;
        RECT 96.545 192.325 96.800 192.895 ;
        RECT 95.445 191.195 95.615 192.325 ;
        RECT 96.205 192.155 96.375 192.325 ;
        RECT 94.490 191.025 95.615 191.195 ;
        RECT 95.785 191.825 95.980 192.155 ;
        RECT 96.205 191.825 96.460 192.155 ;
        RECT 95.785 190.855 95.955 191.825 ;
        RECT 96.630 191.655 96.800 192.325 ;
        RECT 93.925 190.685 95.955 190.855 ;
        RECT 96.125 190.515 96.295 191.655 ;
        RECT 96.465 190.685 96.800 191.655 ;
        RECT 96.975 192.390 97.235 192.895 ;
        RECT 97.415 192.685 97.745 193.065 ;
        RECT 97.925 192.515 98.095 192.895 ;
        RECT 96.975 191.590 97.145 192.390 ;
        RECT 97.430 192.345 98.095 192.515 ;
        RECT 98.815 192.390 99.075 192.895 ;
        RECT 99.255 192.685 99.585 193.065 ;
        RECT 99.765 192.515 99.935 192.895 ;
        RECT 97.430 192.090 97.600 192.345 ;
        RECT 97.315 191.760 97.600 192.090 ;
        RECT 97.835 191.795 98.165 192.165 ;
        RECT 97.430 191.615 97.600 191.760 ;
        RECT 96.975 190.685 97.245 191.590 ;
        RECT 97.430 191.445 98.095 191.615 ;
        RECT 97.415 190.515 97.745 191.275 ;
        RECT 97.925 190.685 98.095 191.445 ;
        RECT 98.815 191.590 98.985 192.390 ;
        RECT 99.270 192.345 99.935 192.515 ;
        RECT 99.270 192.090 99.440 192.345 ;
        RECT 100.195 192.340 100.485 193.065 ;
        RECT 100.715 192.245 100.925 193.065 ;
        RECT 101.095 192.265 101.425 192.895 ;
        RECT 99.155 191.760 99.440 192.090 ;
        RECT 99.675 191.795 100.005 192.165 ;
        RECT 99.270 191.615 99.440 191.760 ;
        RECT 98.815 190.685 99.085 191.590 ;
        RECT 99.270 191.445 99.935 191.615 ;
        RECT 99.255 190.515 99.585 191.275 ;
        RECT 99.765 190.685 99.935 191.445 ;
        RECT 100.195 190.515 100.485 191.680 ;
        RECT 101.095 191.665 101.345 192.265 ;
        RECT 101.595 192.245 101.825 193.065 ;
        RECT 102.500 192.515 102.755 192.805 ;
        RECT 102.925 192.685 103.255 193.065 ;
        RECT 102.500 192.345 103.250 192.515 ;
        RECT 101.515 191.825 101.845 192.075 ;
        RECT 100.715 190.515 100.925 191.655 ;
        RECT 101.095 190.685 101.425 191.665 ;
        RECT 101.595 190.515 101.825 191.655 ;
        RECT 102.500 191.525 102.850 192.175 ;
        RECT 103.020 191.355 103.250 192.345 ;
        RECT 102.500 191.185 103.250 191.355 ;
        RECT 102.500 190.685 102.755 191.185 ;
        RECT 102.925 190.515 103.255 191.015 ;
        RECT 103.425 190.685 103.595 192.805 ;
        RECT 103.955 192.705 104.285 193.065 ;
        RECT 104.455 192.675 104.950 192.845 ;
        RECT 105.155 192.675 106.010 192.845 ;
        RECT 103.825 191.485 104.285 192.535 ;
        RECT 103.765 190.700 104.090 191.485 ;
        RECT 104.455 191.315 104.625 192.675 ;
        RECT 104.795 191.765 105.145 192.385 ;
        RECT 105.315 192.165 105.670 192.385 ;
        RECT 105.315 191.575 105.485 192.165 ;
        RECT 105.840 191.965 106.010 192.675 ;
        RECT 106.885 192.605 107.215 193.065 ;
        RECT 107.425 192.705 107.775 192.875 ;
        RECT 106.215 192.135 107.005 192.385 ;
        RECT 107.425 192.315 107.685 192.705 ;
        RECT 107.995 192.615 108.945 192.895 ;
        RECT 109.115 192.625 109.305 193.065 ;
        RECT 109.475 192.685 110.545 192.855 ;
        RECT 107.175 191.965 107.345 192.145 ;
        RECT 104.455 191.145 104.850 191.315 ;
        RECT 105.020 191.185 105.485 191.575 ;
        RECT 105.655 191.795 107.345 191.965 ;
        RECT 104.680 191.015 104.850 191.145 ;
        RECT 105.655 191.015 105.825 191.795 ;
        RECT 107.515 191.625 107.685 192.315 ;
        RECT 106.185 191.455 107.685 191.625 ;
        RECT 107.875 191.655 108.085 192.445 ;
        RECT 108.255 191.825 108.605 192.445 ;
        RECT 108.775 191.835 108.945 192.615 ;
        RECT 109.475 192.455 109.645 192.685 ;
        RECT 109.115 192.285 109.645 192.455 ;
        RECT 109.115 192.005 109.335 192.285 ;
        RECT 109.815 192.115 110.055 192.515 ;
        RECT 108.775 191.665 109.180 191.835 ;
        RECT 109.515 191.745 110.055 192.115 ;
        RECT 110.225 192.330 110.545 192.685 ;
        RECT 110.790 192.605 111.095 193.065 ;
        RECT 111.265 192.355 111.520 192.885 ;
        RECT 110.225 192.155 110.550 192.330 ;
        RECT 110.225 191.855 111.140 192.155 ;
        RECT 110.400 191.825 111.140 191.855 ;
        RECT 107.875 191.495 108.550 191.655 ;
        RECT 109.010 191.575 109.180 191.665 ;
        RECT 107.875 191.485 108.840 191.495 ;
        RECT 107.515 191.315 107.685 191.455 ;
        RECT 104.260 190.515 104.510 190.975 ;
        RECT 104.680 190.685 104.930 191.015 ;
        RECT 105.145 190.685 105.825 191.015 ;
        RECT 105.995 191.115 107.070 191.285 ;
        RECT 107.515 191.145 108.075 191.315 ;
        RECT 108.380 191.195 108.840 191.485 ;
        RECT 109.010 191.405 110.230 191.575 ;
        RECT 105.995 190.775 106.165 191.115 ;
        RECT 106.400 190.515 106.730 190.945 ;
        RECT 106.900 190.775 107.070 191.115 ;
        RECT 107.365 190.515 107.735 190.975 ;
        RECT 107.905 190.685 108.075 191.145 ;
        RECT 109.010 191.025 109.180 191.405 ;
        RECT 110.400 191.235 110.570 191.825 ;
        RECT 111.310 191.705 111.520 192.355 ;
        RECT 112.155 192.315 113.365 193.065 ;
        RECT 108.310 190.685 109.180 191.025 ;
        RECT 109.770 191.065 110.570 191.235 ;
        RECT 109.350 190.515 109.600 190.975 ;
        RECT 109.770 190.775 109.940 191.065 ;
        RECT 110.120 190.515 110.450 190.895 ;
        RECT 110.790 190.515 111.095 191.655 ;
        RECT 111.265 190.825 111.520 191.705 ;
        RECT 112.155 191.605 112.675 192.145 ;
        RECT 112.845 191.775 113.365 192.315 ;
        RECT 112.155 190.515 113.365 191.605 ;
        RECT 26.970 190.345 113.450 190.515 ;
        RECT 27.055 189.255 28.265 190.345 ;
        RECT 27.055 188.545 27.575 189.085 ;
        RECT 27.745 188.715 28.265 189.255 ;
        RECT 28.955 189.205 29.165 190.345 ;
        RECT 29.335 189.195 29.665 190.175 ;
        RECT 29.835 189.205 30.065 190.345 ;
        RECT 30.365 189.415 30.535 190.175 ;
        RECT 30.715 189.585 31.045 190.345 ;
        RECT 30.365 189.245 31.030 189.415 ;
        RECT 31.215 189.270 31.485 190.175 ;
        RECT 27.055 187.795 28.265 188.545 ;
        RECT 28.955 187.795 29.165 188.615 ;
        RECT 29.335 188.595 29.585 189.195 ;
        RECT 30.860 189.100 31.030 189.245 ;
        RECT 29.755 188.785 30.085 189.035 ;
        RECT 30.295 188.695 30.625 189.065 ;
        RECT 30.860 188.770 31.145 189.100 ;
        RECT 29.335 187.965 29.665 188.595 ;
        RECT 29.835 187.795 30.065 188.615 ;
        RECT 30.860 188.515 31.030 188.770 ;
        RECT 30.365 188.345 31.030 188.515 ;
        RECT 31.315 188.470 31.485 189.270 ;
        RECT 31.655 189.585 32.170 189.995 ;
        RECT 32.405 189.585 32.575 190.345 ;
        RECT 32.745 190.005 34.775 190.175 ;
        RECT 31.655 188.775 31.995 189.585 ;
        RECT 32.745 189.340 32.915 190.005 ;
        RECT 33.310 189.665 34.435 189.835 ;
        RECT 32.165 189.150 32.915 189.340 ;
        RECT 33.085 189.325 34.095 189.495 ;
        RECT 31.655 188.605 32.885 188.775 ;
        RECT 30.365 187.965 30.535 188.345 ;
        RECT 30.715 187.795 31.045 188.175 ;
        RECT 31.225 187.965 31.485 188.470 ;
        RECT 31.930 188.000 32.175 188.605 ;
        RECT 32.395 187.795 32.905 188.330 ;
        RECT 33.085 187.965 33.275 189.325 ;
        RECT 33.445 188.985 33.720 189.125 ;
        RECT 33.445 188.815 33.725 188.985 ;
        RECT 33.445 187.965 33.720 188.815 ;
        RECT 33.925 188.525 34.095 189.325 ;
        RECT 34.265 188.535 34.435 189.665 ;
        RECT 34.605 189.035 34.775 190.005 ;
        RECT 34.945 189.205 35.115 190.345 ;
        RECT 35.285 189.205 35.620 190.175 ;
        RECT 34.605 188.705 34.800 189.035 ;
        RECT 35.025 188.705 35.280 189.035 ;
        RECT 35.025 188.535 35.195 188.705 ;
        RECT 35.450 188.535 35.620 189.205 ;
        RECT 35.795 189.180 36.085 190.345 ;
        RECT 36.805 189.415 36.975 190.175 ;
        RECT 37.155 189.585 37.485 190.345 ;
        RECT 36.805 189.245 37.470 189.415 ;
        RECT 37.655 189.270 37.925 190.175 ;
        RECT 37.300 189.100 37.470 189.245 ;
        RECT 36.735 188.695 37.065 189.065 ;
        RECT 37.300 188.770 37.585 189.100 ;
        RECT 34.265 188.365 35.195 188.535 ;
        RECT 34.265 188.330 34.440 188.365 ;
        RECT 33.910 187.965 34.440 188.330 ;
        RECT 34.865 187.795 35.195 188.195 ;
        RECT 35.365 187.965 35.620 188.535 ;
        RECT 35.795 187.795 36.085 188.520 ;
        RECT 37.300 188.515 37.470 188.770 ;
        RECT 36.805 188.345 37.470 188.515 ;
        RECT 37.755 188.470 37.925 189.270 ;
        RECT 38.135 189.205 38.365 190.345 ;
        RECT 38.535 189.195 38.865 190.175 ;
        RECT 39.035 189.205 39.245 190.345 ;
        RECT 39.680 189.375 40.010 190.175 ;
        RECT 40.180 189.545 40.510 190.345 ;
        RECT 40.810 189.375 41.140 190.175 ;
        RECT 41.785 189.545 42.035 190.345 ;
        RECT 39.680 189.205 42.115 189.375 ;
        RECT 42.305 189.205 42.475 190.345 ;
        RECT 42.645 189.205 42.985 190.175 ;
        RECT 38.115 188.785 38.445 189.035 ;
        RECT 36.805 187.965 36.975 188.345 ;
        RECT 37.155 187.795 37.485 188.175 ;
        RECT 37.665 187.965 37.925 188.470 ;
        RECT 38.135 187.795 38.365 188.615 ;
        RECT 38.615 188.595 38.865 189.195 ;
        RECT 39.475 188.785 39.825 189.035 ;
        RECT 38.535 187.965 38.865 188.595 ;
        RECT 39.035 187.795 39.245 188.615 ;
        RECT 40.010 188.575 40.180 189.205 ;
        RECT 40.350 188.785 40.680 188.985 ;
        RECT 40.850 188.785 41.180 188.985 ;
        RECT 41.350 188.785 41.770 188.985 ;
        RECT 41.945 188.955 42.115 189.205 ;
        RECT 41.945 188.785 42.640 188.955 ;
        RECT 39.680 187.965 40.180 188.575 ;
        RECT 40.810 188.445 42.035 188.615 ;
        RECT 42.810 188.595 42.985 189.205 ;
        RECT 40.810 187.965 41.140 188.445 ;
        RECT 41.310 187.795 41.535 188.255 ;
        RECT 41.705 187.965 42.035 188.445 ;
        RECT 42.225 187.795 42.475 188.595 ;
        RECT 42.645 187.965 42.985 188.595 ;
        RECT 43.160 189.155 43.415 190.035 ;
        RECT 43.585 189.205 43.890 190.345 ;
        RECT 44.230 189.965 44.560 190.345 ;
        RECT 44.740 189.795 44.910 190.085 ;
        RECT 45.080 189.885 45.330 190.345 ;
        RECT 44.110 189.625 44.910 189.795 ;
        RECT 45.500 189.835 46.370 190.175 ;
        RECT 43.160 188.505 43.370 189.155 ;
        RECT 44.110 189.035 44.280 189.625 ;
        RECT 45.500 189.455 45.670 189.835 ;
        RECT 46.605 189.715 46.775 190.175 ;
        RECT 46.945 189.885 47.315 190.345 ;
        RECT 47.610 189.745 47.780 190.085 ;
        RECT 47.950 189.915 48.280 190.345 ;
        RECT 48.515 189.745 48.685 190.085 ;
        RECT 44.450 189.285 45.670 189.455 ;
        RECT 45.840 189.375 46.300 189.665 ;
        RECT 46.605 189.545 47.165 189.715 ;
        RECT 47.610 189.575 48.685 189.745 ;
        RECT 48.855 189.845 49.535 190.175 ;
        RECT 49.750 189.845 50.000 190.175 ;
        RECT 50.170 189.885 50.420 190.345 ;
        RECT 46.995 189.405 47.165 189.545 ;
        RECT 45.840 189.365 46.805 189.375 ;
        RECT 45.500 189.195 45.670 189.285 ;
        RECT 46.130 189.205 46.805 189.365 ;
        RECT 43.540 189.005 44.280 189.035 ;
        RECT 43.540 188.705 44.455 189.005 ;
        RECT 44.130 188.530 44.455 188.705 ;
        RECT 43.160 187.975 43.415 188.505 ;
        RECT 43.585 187.795 43.890 188.255 ;
        RECT 44.135 188.175 44.455 188.530 ;
        RECT 44.625 188.745 45.165 189.115 ;
        RECT 45.500 189.025 45.905 189.195 ;
        RECT 44.625 188.345 44.865 188.745 ;
        RECT 45.345 188.575 45.565 188.855 ;
        RECT 45.035 188.405 45.565 188.575 ;
        RECT 45.035 188.175 45.205 188.405 ;
        RECT 45.735 188.245 45.905 189.025 ;
        RECT 46.075 188.415 46.425 189.035 ;
        RECT 46.595 188.415 46.805 189.205 ;
        RECT 46.995 189.235 48.495 189.405 ;
        RECT 46.995 188.545 47.165 189.235 ;
        RECT 48.855 189.065 49.025 189.845 ;
        RECT 49.830 189.715 50.000 189.845 ;
        RECT 47.335 188.895 49.025 189.065 ;
        RECT 49.195 189.285 49.660 189.675 ;
        RECT 49.830 189.545 50.225 189.715 ;
        RECT 47.335 188.715 47.505 188.895 ;
        RECT 44.135 188.005 45.205 188.175 ;
        RECT 45.375 187.795 45.565 188.235 ;
        RECT 45.735 187.965 46.685 188.245 ;
        RECT 46.995 188.155 47.255 188.545 ;
        RECT 47.675 188.475 48.465 188.725 ;
        RECT 46.905 187.985 47.255 188.155 ;
        RECT 47.465 187.795 47.795 188.255 ;
        RECT 48.670 188.185 48.840 188.895 ;
        RECT 49.195 188.695 49.365 189.285 ;
        RECT 49.010 188.475 49.365 188.695 ;
        RECT 49.535 188.475 49.885 189.095 ;
        RECT 50.055 188.185 50.225 189.545 ;
        RECT 50.590 189.375 50.915 190.160 ;
        RECT 50.395 188.325 50.855 189.375 ;
        RECT 48.670 188.015 49.525 188.185 ;
        RECT 49.730 188.015 50.225 188.185 ;
        RECT 50.395 187.795 50.725 188.155 ;
        RECT 51.085 188.055 51.255 190.175 ;
        RECT 51.425 189.845 51.755 190.345 ;
        RECT 51.925 189.675 52.180 190.175 ;
        RECT 51.430 189.505 52.180 189.675 ;
        RECT 51.430 188.515 51.660 189.505 ;
        RECT 52.560 189.375 52.890 190.175 ;
        RECT 53.060 189.545 53.390 190.345 ;
        RECT 53.690 189.375 54.020 190.175 ;
        RECT 54.665 189.545 54.915 190.345 ;
        RECT 51.830 188.685 52.180 189.335 ;
        RECT 52.560 189.205 54.995 189.375 ;
        RECT 55.185 189.205 55.355 190.345 ;
        RECT 55.525 189.205 55.865 190.175 ;
        RECT 52.355 188.785 52.705 189.035 ;
        RECT 52.890 188.575 53.060 189.205 ;
        RECT 53.230 188.785 53.560 188.985 ;
        RECT 53.730 188.785 54.060 188.985 ;
        RECT 54.230 188.785 54.650 188.985 ;
        RECT 54.825 188.955 54.995 189.205 ;
        RECT 54.825 188.785 55.520 188.955 ;
        RECT 51.430 188.345 52.180 188.515 ;
        RECT 51.425 187.795 51.755 188.175 ;
        RECT 51.925 188.055 52.180 188.345 ;
        RECT 52.560 187.965 53.060 188.575 ;
        RECT 53.690 188.445 54.915 188.615 ;
        RECT 55.690 188.595 55.865 189.205 ;
        RECT 53.690 187.965 54.020 188.445 ;
        RECT 54.190 187.795 54.415 188.255 ;
        RECT 54.585 187.965 54.915 188.445 ;
        RECT 55.105 187.795 55.355 188.595 ;
        RECT 55.525 187.965 55.865 188.595 ;
        RECT 56.040 189.205 56.375 190.175 ;
        RECT 56.545 189.205 56.715 190.345 ;
        RECT 56.885 190.005 58.915 190.175 ;
        RECT 56.040 188.535 56.210 189.205 ;
        RECT 56.885 189.035 57.055 190.005 ;
        RECT 56.380 188.705 56.635 189.035 ;
        RECT 56.860 188.705 57.055 189.035 ;
        RECT 57.225 189.665 58.350 189.835 ;
        RECT 56.465 188.535 56.635 188.705 ;
        RECT 57.225 188.535 57.395 189.665 ;
        RECT 56.040 187.965 56.295 188.535 ;
        RECT 56.465 188.365 57.395 188.535 ;
        RECT 57.565 189.325 58.575 189.495 ;
        RECT 57.565 188.525 57.735 189.325 ;
        RECT 57.940 188.645 58.215 189.125 ;
        RECT 57.935 188.475 58.215 188.645 ;
        RECT 57.220 188.330 57.395 188.365 ;
        RECT 56.465 187.795 56.795 188.195 ;
        RECT 57.220 187.965 57.750 188.330 ;
        RECT 57.940 187.965 58.215 188.475 ;
        RECT 58.385 187.965 58.575 189.325 ;
        RECT 58.745 189.340 58.915 190.005 ;
        RECT 59.085 189.585 59.255 190.345 ;
        RECT 59.490 189.585 60.005 189.995 ;
        RECT 58.745 189.150 59.495 189.340 ;
        RECT 59.665 188.775 60.005 189.585 ;
        RECT 60.265 189.415 60.435 190.175 ;
        RECT 60.615 189.585 60.945 190.345 ;
        RECT 60.265 189.245 60.930 189.415 ;
        RECT 61.115 189.270 61.385 190.175 ;
        RECT 60.760 189.100 60.930 189.245 ;
        RECT 58.775 188.605 60.005 188.775 ;
        RECT 60.195 188.695 60.525 189.065 ;
        RECT 60.760 188.770 61.045 189.100 ;
        RECT 58.755 187.795 59.265 188.330 ;
        RECT 59.485 188.000 59.730 188.605 ;
        RECT 60.760 188.515 60.930 188.770 ;
        RECT 60.265 188.345 60.930 188.515 ;
        RECT 61.215 188.470 61.385 189.270 ;
        RECT 61.555 189.180 61.845 190.345 ;
        RECT 62.015 189.205 62.400 190.175 ;
        RECT 62.570 189.885 62.895 190.345 ;
        RECT 63.415 189.715 63.695 190.175 ;
        RECT 62.570 189.495 63.695 189.715 ;
        RECT 62.015 188.535 62.295 189.205 ;
        RECT 62.570 189.035 63.020 189.495 ;
        RECT 63.885 189.325 64.285 190.175 ;
        RECT 64.685 189.885 64.955 190.345 ;
        RECT 65.125 189.715 65.410 190.175 ;
        RECT 62.465 188.705 63.020 189.035 ;
        RECT 63.190 188.765 64.285 189.325 ;
        RECT 62.570 188.595 63.020 188.705 ;
        RECT 60.265 187.965 60.435 188.345 ;
        RECT 60.615 187.795 60.945 188.175 ;
        RECT 61.125 187.965 61.385 188.470 ;
        RECT 61.555 187.795 61.845 188.520 ;
        RECT 62.015 187.965 62.400 188.535 ;
        RECT 62.570 188.425 63.695 188.595 ;
        RECT 62.570 187.795 62.895 188.255 ;
        RECT 63.415 187.965 63.695 188.425 ;
        RECT 63.885 187.965 64.285 188.765 ;
        RECT 64.455 189.495 65.410 189.715 ;
        RECT 64.455 188.595 64.665 189.495 ;
        RECT 65.695 189.375 66.005 190.175 ;
        RECT 66.175 189.545 66.485 190.345 ;
        RECT 66.655 189.715 66.915 190.175 ;
        RECT 67.085 189.885 67.340 190.345 ;
        RECT 67.515 189.715 67.775 190.175 ;
        RECT 66.655 189.545 67.775 189.715 ;
        RECT 64.835 188.765 65.525 189.325 ;
        RECT 65.695 189.205 66.725 189.375 ;
        RECT 64.455 188.425 65.410 188.595 ;
        RECT 64.685 187.795 64.955 188.255 ;
        RECT 65.125 187.965 65.410 188.425 ;
        RECT 65.695 188.295 65.865 189.205 ;
        RECT 66.035 188.465 66.385 189.035 ;
        RECT 66.555 188.955 66.725 189.205 ;
        RECT 67.515 189.295 67.775 189.545 ;
        RECT 67.945 189.475 68.230 190.345 ;
        RECT 67.515 189.125 68.270 189.295 ;
        RECT 66.555 188.785 67.695 188.955 ;
        RECT 67.865 188.615 68.270 189.125 ;
        RECT 66.620 188.445 68.270 188.615 ;
        RECT 68.455 188.535 68.715 190.160 ;
        RECT 70.465 189.895 70.795 190.345 ;
        RECT 71.790 189.715 72.075 190.175 ;
        RECT 72.245 189.885 72.515 190.345 ;
        RECT 68.895 189.505 71.505 189.715 ;
        RECT 68.895 188.705 69.115 189.505 ;
        RECT 69.355 188.705 69.655 189.325 ;
        RECT 69.825 188.705 70.155 189.325 ;
        RECT 70.325 188.705 70.645 189.325 ;
        RECT 70.815 188.705 71.165 189.325 ;
        RECT 71.335 188.535 71.505 189.505 ;
        RECT 71.790 189.495 72.745 189.715 ;
        RECT 71.675 188.765 72.365 189.325 ;
        RECT 72.535 188.595 72.745 189.495 ;
        RECT 65.695 187.965 65.995 188.295 ;
        RECT 66.165 187.795 66.440 188.275 ;
        RECT 66.620 188.055 66.915 188.445 ;
        RECT 67.085 187.795 67.340 188.275 ;
        RECT 67.515 188.055 67.775 188.445 ;
        RECT 68.455 188.365 70.295 188.535 ;
        RECT 67.945 187.795 68.225 188.275 ;
        RECT 68.725 187.795 69.055 188.190 ;
        RECT 69.225 188.010 69.425 188.365 ;
        RECT 69.595 187.795 69.925 188.195 ;
        RECT 70.095 188.020 70.295 188.365 ;
        RECT 70.465 187.795 70.795 188.535 ;
        RECT 71.030 188.365 71.505 188.535 ;
        RECT 71.790 188.425 72.745 188.595 ;
        RECT 72.915 189.325 73.315 190.175 ;
        RECT 73.505 189.715 73.785 190.175 ;
        RECT 74.305 189.885 74.630 190.345 ;
        RECT 73.505 189.495 74.630 189.715 ;
        RECT 72.915 188.765 74.010 189.325 ;
        RECT 74.180 189.035 74.630 189.495 ;
        RECT 74.800 189.205 75.185 190.175 ;
        RECT 75.470 189.715 75.755 190.175 ;
        RECT 75.925 189.885 76.195 190.345 ;
        RECT 75.470 189.495 76.425 189.715 ;
        RECT 71.030 188.115 71.200 188.365 ;
        RECT 71.790 187.965 72.075 188.425 ;
        RECT 72.245 187.795 72.515 188.255 ;
        RECT 72.915 187.965 73.315 188.765 ;
        RECT 74.180 188.705 74.735 189.035 ;
        RECT 74.180 188.595 74.630 188.705 ;
        RECT 73.505 188.425 74.630 188.595 ;
        RECT 74.905 188.535 75.185 189.205 ;
        RECT 75.355 188.765 76.045 189.325 ;
        RECT 76.215 188.595 76.425 189.495 ;
        RECT 73.505 187.965 73.785 188.425 ;
        RECT 74.305 187.795 74.630 188.255 ;
        RECT 74.800 187.965 75.185 188.535 ;
        RECT 75.470 188.425 76.425 188.595 ;
        RECT 76.595 189.325 76.995 190.175 ;
        RECT 77.185 189.715 77.465 190.175 ;
        RECT 77.985 189.885 78.310 190.345 ;
        RECT 77.185 189.495 78.310 189.715 ;
        RECT 76.595 188.765 77.690 189.325 ;
        RECT 77.860 189.035 78.310 189.495 ;
        RECT 78.480 189.205 78.865 190.175 ;
        RECT 75.470 187.965 75.755 188.425 ;
        RECT 75.925 187.795 76.195 188.255 ;
        RECT 76.595 187.965 76.995 188.765 ;
        RECT 77.860 188.705 78.415 189.035 ;
        RECT 77.860 188.595 78.310 188.705 ;
        RECT 77.185 188.425 78.310 188.595 ;
        RECT 78.585 188.535 78.865 189.205 ;
        RECT 79.035 189.585 79.550 189.995 ;
        RECT 79.785 189.585 79.955 190.345 ;
        RECT 80.125 190.005 82.155 190.175 ;
        RECT 79.035 188.775 79.375 189.585 ;
        RECT 80.125 189.340 80.295 190.005 ;
        RECT 80.690 189.665 81.815 189.835 ;
        RECT 79.545 189.150 80.295 189.340 ;
        RECT 80.465 189.325 81.475 189.495 ;
        RECT 79.035 188.605 80.265 188.775 ;
        RECT 77.185 187.965 77.465 188.425 ;
        RECT 77.985 187.795 78.310 188.255 ;
        RECT 78.480 187.965 78.865 188.535 ;
        RECT 79.310 188.000 79.555 188.605 ;
        RECT 79.775 187.795 80.285 188.330 ;
        RECT 80.465 187.965 80.655 189.325 ;
        RECT 80.825 188.985 81.100 189.125 ;
        RECT 80.825 188.815 81.105 188.985 ;
        RECT 80.825 187.965 81.100 188.815 ;
        RECT 81.305 188.525 81.475 189.325 ;
        RECT 81.645 188.535 81.815 189.665 ;
        RECT 81.985 189.035 82.155 190.005 ;
        RECT 82.325 189.205 82.495 190.345 ;
        RECT 82.665 189.205 83.000 190.175 ;
        RECT 81.985 188.705 82.180 189.035 ;
        RECT 82.405 188.705 82.660 189.035 ;
        RECT 82.405 188.535 82.575 188.705 ;
        RECT 82.830 188.535 83.000 189.205 ;
        RECT 83.175 189.585 83.690 189.995 ;
        RECT 83.925 189.585 84.095 190.345 ;
        RECT 84.265 190.005 86.295 190.175 ;
        RECT 83.175 188.775 83.515 189.585 ;
        RECT 84.265 189.340 84.435 190.005 ;
        RECT 84.830 189.665 85.955 189.835 ;
        RECT 83.685 189.150 84.435 189.340 ;
        RECT 84.605 189.325 85.615 189.495 ;
        RECT 83.175 188.605 84.405 188.775 ;
        RECT 81.645 188.365 82.575 188.535 ;
        RECT 81.645 188.330 81.820 188.365 ;
        RECT 81.290 187.965 81.820 188.330 ;
        RECT 82.245 187.795 82.575 188.195 ;
        RECT 82.745 187.965 83.000 188.535 ;
        RECT 83.450 188.000 83.695 188.605 ;
        RECT 83.915 187.795 84.425 188.330 ;
        RECT 84.605 187.965 84.795 189.325 ;
        RECT 84.965 188.305 85.240 189.125 ;
        RECT 85.445 188.525 85.615 189.325 ;
        RECT 85.785 188.535 85.955 189.665 ;
        RECT 86.125 189.035 86.295 190.005 ;
        RECT 86.465 189.205 86.635 190.345 ;
        RECT 86.805 189.205 87.140 190.175 ;
        RECT 86.125 188.705 86.320 189.035 ;
        RECT 86.545 188.705 86.800 189.035 ;
        RECT 86.545 188.535 86.715 188.705 ;
        RECT 86.970 188.535 87.140 189.205 ;
        RECT 87.315 189.180 87.605 190.345 ;
        RECT 87.775 189.270 88.045 190.175 ;
        RECT 88.215 189.585 88.545 190.345 ;
        RECT 88.725 189.415 88.895 190.175 ;
        RECT 85.785 188.365 86.715 188.535 ;
        RECT 85.785 188.330 85.960 188.365 ;
        RECT 84.965 188.135 85.245 188.305 ;
        RECT 84.965 187.965 85.240 188.135 ;
        RECT 85.430 187.965 85.960 188.330 ;
        RECT 86.385 187.795 86.715 188.195 ;
        RECT 86.885 187.965 87.140 188.535 ;
        RECT 87.315 187.795 87.605 188.520 ;
        RECT 87.775 188.470 87.945 189.270 ;
        RECT 88.230 189.245 88.895 189.415 ;
        RECT 88.230 189.100 88.400 189.245 ;
        RECT 88.115 188.770 88.400 189.100 ;
        RECT 89.620 189.155 89.875 190.035 ;
        RECT 90.045 189.205 90.350 190.345 ;
        RECT 90.690 189.965 91.020 190.345 ;
        RECT 91.200 189.795 91.370 190.085 ;
        RECT 91.540 189.885 91.790 190.345 ;
        RECT 90.570 189.625 91.370 189.795 ;
        RECT 91.960 189.835 92.830 190.175 ;
        RECT 88.230 188.515 88.400 188.770 ;
        RECT 88.635 188.695 88.965 189.065 ;
        RECT 87.775 187.965 88.035 188.470 ;
        RECT 88.230 188.345 88.895 188.515 ;
        RECT 88.215 187.795 88.545 188.175 ;
        RECT 88.725 187.965 88.895 188.345 ;
        RECT 89.620 188.505 89.830 189.155 ;
        RECT 90.570 189.035 90.740 189.625 ;
        RECT 91.960 189.455 92.130 189.835 ;
        RECT 93.065 189.715 93.235 190.175 ;
        RECT 93.405 189.885 93.775 190.345 ;
        RECT 94.070 189.745 94.240 190.085 ;
        RECT 94.410 189.915 94.740 190.345 ;
        RECT 94.975 189.745 95.145 190.085 ;
        RECT 90.910 189.285 92.130 189.455 ;
        RECT 92.300 189.375 92.760 189.665 ;
        RECT 93.065 189.545 93.625 189.715 ;
        RECT 94.070 189.575 95.145 189.745 ;
        RECT 95.315 189.845 95.995 190.175 ;
        RECT 96.210 189.845 96.460 190.175 ;
        RECT 96.630 189.885 96.880 190.345 ;
        RECT 93.455 189.405 93.625 189.545 ;
        RECT 92.300 189.365 93.265 189.375 ;
        RECT 91.960 189.195 92.130 189.285 ;
        RECT 92.590 189.205 93.265 189.365 ;
        RECT 90.000 189.005 90.740 189.035 ;
        RECT 90.000 188.705 90.915 189.005 ;
        RECT 90.590 188.530 90.915 188.705 ;
        RECT 89.620 187.975 89.875 188.505 ;
        RECT 90.045 187.795 90.350 188.255 ;
        RECT 90.595 188.175 90.915 188.530 ;
        RECT 91.085 188.745 91.625 189.115 ;
        RECT 91.960 189.025 92.365 189.195 ;
        RECT 91.085 188.345 91.325 188.745 ;
        RECT 91.805 188.575 92.025 188.855 ;
        RECT 91.495 188.405 92.025 188.575 ;
        RECT 91.495 188.175 91.665 188.405 ;
        RECT 92.195 188.245 92.365 189.025 ;
        RECT 92.535 188.415 92.885 189.035 ;
        RECT 93.055 188.415 93.265 189.205 ;
        RECT 93.455 189.235 94.955 189.405 ;
        RECT 93.455 188.545 93.625 189.235 ;
        RECT 95.315 189.065 95.485 189.845 ;
        RECT 96.290 189.715 96.460 189.845 ;
        RECT 93.795 188.895 95.485 189.065 ;
        RECT 95.655 189.285 96.120 189.675 ;
        RECT 96.290 189.545 96.685 189.715 ;
        RECT 93.795 188.715 93.965 188.895 ;
        RECT 90.595 188.005 91.665 188.175 ;
        RECT 91.835 187.795 92.025 188.235 ;
        RECT 92.195 187.965 93.145 188.245 ;
        RECT 93.455 188.155 93.715 188.545 ;
        RECT 94.135 188.475 94.925 188.725 ;
        RECT 93.365 187.985 93.715 188.155 ;
        RECT 93.925 187.795 94.255 188.255 ;
        RECT 95.130 188.185 95.300 188.895 ;
        RECT 95.655 188.695 95.825 189.285 ;
        RECT 95.470 188.475 95.825 188.695 ;
        RECT 95.995 188.475 96.345 189.095 ;
        RECT 96.515 188.185 96.685 189.545 ;
        RECT 97.050 189.375 97.375 190.160 ;
        RECT 96.855 188.325 97.315 189.375 ;
        RECT 95.130 188.015 95.985 188.185 ;
        RECT 96.190 188.015 96.685 188.185 ;
        RECT 96.855 187.795 97.185 188.155 ;
        RECT 97.545 188.055 97.715 190.175 ;
        RECT 97.885 189.845 98.215 190.345 ;
        RECT 98.385 189.675 98.640 190.175 ;
        RECT 97.890 189.505 98.640 189.675 ;
        RECT 97.890 188.515 98.120 189.505 ;
        RECT 98.290 188.685 98.640 189.335 ;
        RECT 98.815 189.270 99.085 190.175 ;
        RECT 99.255 189.585 99.585 190.345 ;
        RECT 99.765 189.415 99.935 190.175 ;
        RECT 97.890 188.345 98.640 188.515 ;
        RECT 97.885 187.795 98.215 188.175 ;
        RECT 98.385 188.055 98.640 188.345 ;
        RECT 98.815 188.470 98.985 189.270 ;
        RECT 99.270 189.245 99.935 189.415 ;
        RECT 99.270 189.100 99.440 189.245 ;
        RECT 99.155 188.770 99.440 189.100 ;
        RECT 100.660 189.155 100.915 190.035 ;
        RECT 101.085 189.205 101.390 190.345 ;
        RECT 101.730 189.965 102.060 190.345 ;
        RECT 102.240 189.795 102.410 190.085 ;
        RECT 102.580 189.885 102.830 190.345 ;
        RECT 101.610 189.625 102.410 189.795 ;
        RECT 103.000 189.835 103.870 190.175 ;
        RECT 99.270 188.515 99.440 188.770 ;
        RECT 99.675 188.695 100.005 189.065 ;
        RECT 98.815 187.965 99.075 188.470 ;
        RECT 99.270 188.345 99.935 188.515 ;
        RECT 99.255 187.795 99.585 188.175 ;
        RECT 99.765 187.965 99.935 188.345 ;
        RECT 100.660 188.505 100.870 189.155 ;
        RECT 101.610 189.035 101.780 189.625 ;
        RECT 103.000 189.455 103.170 189.835 ;
        RECT 104.105 189.715 104.275 190.175 ;
        RECT 104.445 189.885 104.815 190.345 ;
        RECT 105.110 189.745 105.280 190.085 ;
        RECT 105.450 189.915 105.780 190.345 ;
        RECT 106.015 189.745 106.185 190.085 ;
        RECT 101.950 189.285 103.170 189.455 ;
        RECT 103.340 189.375 103.800 189.665 ;
        RECT 104.105 189.545 104.665 189.715 ;
        RECT 105.110 189.575 106.185 189.745 ;
        RECT 106.355 189.845 107.035 190.175 ;
        RECT 107.250 189.845 107.500 190.175 ;
        RECT 107.670 189.885 107.920 190.345 ;
        RECT 104.495 189.405 104.665 189.545 ;
        RECT 103.340 189.365 104.305 189.375 ;
        RECT 103.000 189.195 103.170 189.285 ;
        RECT 103.630 189.205 104.305 189.365 ;
        RECT 101.040 189.005 101.780 189.035 ;
        RECT 101.040 188.705 101.955 189.005 ;
        RECT 101.630 188.530 101.955 188.705 ;
        RECT 100.660 187.975 100.915 188.505 ;
        RECT 101.085 187.795 101.390 188.255 ;
        RECT 101.635 188.175 101.955 188.530 ;
        RECT 102.125 188.745 102.665 189.115 ;
        RECT 103.000 189.025 103.405 189.195 ;
        RECT 102.125 188.345 102.365 188.745 ;
        RECT 102.845 188.575 103.065 188.855 ;
        RECT 102.535 188.405 103.065 188.575 ;
        RECT 102.535 188.175 102.705 188.405 ;
        RECT 103.235 188.245 103.405 189.025 ;
        RECT 103.575 188.415 103.925 189.035 ;
        RECT 104.095 188.415 104.305 189.205 ;
        RECT 104.495 189.235 105.995 189.405 ;
        RECT 104.495 188.545 104.665 189.235 ;
        RECT 106.355 189.065 106.525 189.845 ;
        RECT 107.330 189.715 107.500 189.845 ;
        RECT 104.835 188.895 106.525 189.065 ;
        RECT 106.695 189.285 107.160 189.675 ;
        RECT 107.330 189.545 107.725 189.715 ;
        RECT 104.835 188.715 105.005 188.895 ;
        RECT 101.635 188.005 102.705 188.175 ;
        RECT 102.875 187.795 103.065 188.235 ;
        RECT 103.235 187.965 104.185 188.245 ;
        RECT 104.495 188.155 104.755 188.545 ;
        RECT 105.175 188.475 105.965 188.725 ;
        RECT 104.405 187.985 104.755 188.155 ;
        RECT 104.965 187.795 105.295 188.255 ;
        RECT 106.170 188.185 106.340 188.895 ;
        RECT 106.695 188.695 106.865 189.285 ;
        RECT 106.510 188.475 106.865 188.695 ;
        RECT 107.035 188.475 107.385 189.095 ;
        RECT 107.555 188.185 107.725 189.545 ;
        RECT 108.090 189.375 108.415 190.160 ;
        RECT 107.895 188.325 108.355 189.375 ;
        RECT 106.170 188.015 107.025 188.185 ;
        RECT 107.230 188.015 107.725 188.185 ;
        RECT 107.895 187.795 108.225 188.155 ;
        RECT 108.585 188.055 108.755 190.175 ;
        RECT 108.925 189.845 109.255 190.345 ;
        RECT 109.425 189.675 109.680 190.175 ;
        RECT 108.930 189.505 109.680 189.675 ;
        RECT 108.930 188.515 109.160 189.505 ;
        RECT 109.330 188.685 109.680 189.335 ;
        RECT 109.855 189.270 110.125 190.175 ;
        RECT 110.295 189.585 110.625 190.345 ;
        RECT 110.805 189.415 110.975 190.175 ;
        RECT 108.930 188.345 109.680 188.515 ;
        RECT 108.925 187.795 109.255 188.175 ;
        RECT 109.425 188.055 109.680 188.345 ;
        RECT 109.855 188.470 110.025 189.270 ;
        RECT 110.310 189.245 110.975 189.415 ;
        RECT 112.155 189.255 113.365 190.345 ;
        RECT 110.310 189.100 110.480 189.245 ;
        RECT 110.195 188.770 110.480 189.100 ;
        RECT 110.310 188.515 110.480 188.770 ;
        RECT 110.715 188.695 111.045 189.065 ;
        RECT 112.155 188.715 112.675 189.255 ;
        RECT 112.845 188.545 113.365 189.085 ;
        RECT 109.855 187.965 110.115 188.470 ;
        RECT 110.310 188.345 110.975 188.515 ;
        RECT 110.295 187.795 110.625 188.175 ;
        RECT 110.805 187.965 110.975 188.345 ;
        RECT 112.155 187.795 113.365 188.545 ;
        RECT 26.970 187.625 113.450 187.795 ;
        RECT 27.055 186.875 28.265 187.625 ;
        RECT 28.900 186.915 29.155 187.445 ;
        RECT 29.325 187.165 29.630 187.625 ;
        RECT 29.875 187.245 30.945 187.415 ;
        RECT 27.055 186.335 27.575 186.875 ;
        RECT 27.745 186.165 28.265 186.705 ;
        RECT 27.055 185.075 28.265 186.165 ;
        RECT 28.900 186.265 29.110 186.915 ;
        RECT 29.875 186.890 30.195 187.245 ;
        RECT 29.870 186.715 30.195 186.890 ;
        RECT 29.280 186.415 30.195 186.715 ;
        RECT 30.365 186.675 30.605 187.075 ;
        RECT 30.775 187.015 30.945 187.245 ;
        RECT 31.115 187.185 31.305 187.625 ;
        RECT 31.475 187.175 32.425 187.455 ;
        RECT 32.645 187.265 32.995 187.435 ;
        RECT 30.775 186.845 31.305 187.015 ;
        RECT 29.280 186.385 30.020 186.415 ;
        RECT 28.900 185.385 29.155 186.265 ;
        RECT 29.325 185.075 29.630 186.215 ;
        RECT 29.850 185.795 30.020 186.385 ;
        RECT 30.365 186.305 30.905 186.675 ;
        RECT 31.085 186.565 31.305 186.845 ;
        RECT 31.475 186.395 31.645 187.175 ;
        RECT 31.240 186.225 31.645 186.395 ;
        RECT 31.815 186.385 32.165 187.005 ;
        RECT 31.240 186.135 31.410 186.225 ;
        RECT 32.335 186.215 32.545 187.005 ;
        RECT 30.190 185.965 31.410 186.135 ;
        RECT 31.870 186.055 32.545 186.215 ;
        RECT 29.850 185.625 30.650 185.795 ;
        RECT 29.970 185.075 30.300 185.455 ;
        RECT 30.480 185.335 30.650 185.625 ;
        RECT 31.240 185.585 31.410 185.965 ;
        RECT 31.580 186.045 32.545 186.055 ;
        RECT 32.735 186.875 32.995 187.265 ;
        RECT 33.205 187.165 33.535 187.625 ;
        RECT 34.410 187.235 35.265 187.405 ;
        RECT 35.470 187.235 35.965 187.405 ;
        RECT 36.135 187.265 36.465 187.625 ;
        RECT 32.735 186.185 32.905 186.875 ;
        RECT 33.075 186.525 33.245 186.705 ;
        RECT 33.415 186.695 34.205 186.945 ;
        RECT 34.410 186.525 34.580 187.235 ;
        RECT 34.750 186.725 35.105 186.945 ;
        RECT 33.075 186.355 34.765 186.525 ;
        RECT 31.580 185.755 32.040 186.045 ;
        RECT 32.735 186.015 34.235 186.185 ;
        RECT 32.735 185.875 32.905 186.015 ;
        RECT 32.345 185.705 32.905 185.875 ;
        RECT 30.820 185.075 31.070 185.535 ;
        RECT 31.240 185.245 32.110 185.585 ;
        RECT 32.345 185.245 32.515 185.705 ;
        RECT 33.350 185.675 34.425 185.845 ;
        RECT 32.685 185.075 33.055 185.535 ;
        RECT 33.350 185.335 33.520 185.675 ;
        RECT 33.690 185.075 34.020 185.505 ;
        RECT 34.255 185.335 34.425 185.675 ;
        RECT 34.595 185.575 34.765 186.355 ;
        RECT 34.935 186.135 35.105 186.725 ;
        RECT 35.275 186.325 35.625 186.945 ;
        RECT 34.935 185.745 35.400 186.135 ;
        RECT 35.795 185.875 35.965 187.235 ;
        RECT 36.135 186.045 36.595 187.095 ;
        RECT 35.570 185.705 35.965 185.875 ;
        RECT 35.570 185.575 35.740 185.705 ;
        RECT 34.595 185.245 35.275 185.575 ;
        RECT 35.490 185.245 35.740 185.575 ;
        RECT 35.910 185.075 36.160 185.535 ;
        RECT 36.330 185.260 36.655 186.045 ;
        RECT 36.825 185.245 36.995 187.365 ;
        RECT 37.165 187.245 37.495 187.625 ;
        RECT 37.665 187.075 37.920 187.365 ;
        RECT 37.170 186.905 37.920 187.075 ;
        RECT 38.100 186.915 38.355 187.445 ;
        RECT 38.525 187.165 38.830 187.625 ;
        RECT 39.075 187.245 40.145 187.415 ;
        RECT 37.170 185.915 37.400 186.905 ;
        RECT 37.570 186.085 37.920 186.735 ;
        RECT 38.100 186.265 38.310 186.915 ;
        RECT 39.075 186.890 39.395 187.245 ;
        RECT 39.070 186.715 39.395 186.890 ;
        RECT 38.480 186.415 39.395 186.715 ;
        RECT 39.565 186.675 39.805 187.075 ;
        RECT 39.975 187.015 40.145 187.245 ;
        RECT 40.315 187.185 40.505 187.625 ;
        RECT 40.675 187.175 41.625 187.455 ;
        RECT 41.845 187.265 42.195 187.435 ;
        RECT 39.975 186.845 40.505 187.015 ;
        RECT 38.480 186.385 39.220 186.415 ;
        RECT 37.170 185.745 37.920 185.915 ;
        RECT 37.165 185.075 37.495 185.575 ;
        RECT 37.665 185.245 37.920 185.745 ;
        RECT 38.100 185.385 38.355 186.265 ;
        RECT 38.525 185.075 38.830 186.215 ;
        RECT 39.050 185.795 39.220 186.385 ;
        RECT 39.565 186.305 40.105 186.675 ;
        RECT 40.285 186.565 40.505 186.845 ;
        RECT 40.675 186.395 40.845 187.175 ;
        RECT 40.440 186.225 40.845 186.395 ;
        RECT 41.015 186.385 41.365 187.005 ;
        RECT 40.440 186.135 40.610 186.225 ;
        RECT 41.535 186.215 41.745 187.005 ;
        RECT 39.390 185.965 40.610 186.135 ;
        RECT 41.070 186.055 41.745 186.215 ;
        RECT 39.050 185.625 39.850 185.795 ;
        RECT 39.170 185.075 39.500 185.455 ;
        RECT 39.680 185.335 39.850 185.625 ;
        RECT 40.440 185.585 40.610 185.965 ;
        RECT 40.780 186.045 41.745 186.055 ;
        RECT 41.935 186.875 42.195 187.265 ;
        RECT 42.405 187.165 42.735 187.625 ;
        RECT 43.610 187.235 44.465 187.405 ;
        RECT 44.670 187.235 45.165 187.405 ;
        RECT 45.335 187.265 45.665 187.625 ;
        RECT 41.935 186.185 42.105 186.875 ;
        RECT 42.275 186.525 42.445 186.705 ;
        RECT 42.615 186.695 43.405 186.945 ;
        RECT 43.610 186.525 43.780 187.235 ;
        RECT 43.950 186.725 44.305 186.945 ;
        RECT 42.275 186.355 43.965 186.525 ;
        RECT 40.780 185.755 41.240 186.045 ;
        RECT 41.935 186.015 43.435 186.185 ;
        RECT 41.935 185.875 42.105 186.015 ;
        RECT 41.545 185.705 42.105 185.875 ;
        RECT 40.020 185.075 40.270 185.535 ;
        RECT 40.440 185.245 41.310 185.585 ;
        RECT 41.545 185.245 41.715 185.705 ;
        RECT 42.550 185.675 43.625 185.845 ;
        RECT 41.885 185.075 42.255 185.535 ;
        RECT 42.550 185.335 42.720 185.675 ;
        RECT 42.890 185.075 43.220 185.505 ;
        RECT 43.455 185.335 43.625 185.675 ;
        RECT 43.795 185.575 43.965 186.355 ;
        RECT 44.135 186.135 44.305 186.725 ;
        RECT 44.475 186.325 44.825 186.945 ;
        RECT 44.135 185.745 44.600 186.135 ;
        RECT 44.995 185.875 45.165 187.235 ;
        RECT 45.335 186.045 45.795 187.095 ;
        RECT 44.770 185.705 45.165 185.875 ;
        RECT 44.770 185.575 44.940 185.705 ;
        RECT 43.795 185.245 44.475 185.575 ;
        RECT 44.690 185.245 44.940 185.575 ;
        RECT 45.110 185.075 45.360 185.535 ;
        RECT 45.530 185.260 45.855 186.045 ;
        RECT 46.025 185.245 46.195 187.365 ;
        RECT 46.365 187.245 46.695 187.625 ;
        RECT 46.865 187.075 47.120 187.365 ;
        RECT 46.370 186.905 47.120 187.075 ;
        RECT 47.385 187.075 47.555 187.455 ;
        RECT 47.735 187.245 48.065 187.625 ;
        RECT 47.385 186.905 48.050 187.075 ;
        RECT 48.245 186.950 48.505 187.455 ;
        RECT 46.370 185.915 46.600 186.905 ;
        RECT 46.770 186.085 47.120 186.735 ;
        RECT 47.315 186.355 47.645 186.725 ;
        RECT 47.880 186.650 48.050 186.905 ;
        RECT 47.880 186.320 48.165 186.650 ;
        RECT 47.880 186.175 48.050 186.320 ;
        RECT 47.385 186.005 48.050 186.175 ;
        RECT 48.335 186.150 48.505 186.950 ;
        RECT 48.675 186.900 48.965 187.625 ;
        RECT 49.600 186.885 49.855 187.455 ;
        RECT 50.025 187.225 50.355 187.625 ;
        RECT 50.780 187.090 51.310 187.455 ;
        RECT 51.500 187.285 51.775 187.455 ;
        RECT 51.495 187.115 51.775 187.285 ;
        RECT 50.780 187.055 50.955 187.090 ;
        RECT 50.025 186.885 50.955 187.055 ;
        RECT 46.370 185.745 47.120 185.915 ;
        RECT 46.365 185.075 46.695 185.575 ;
        RECT 46.865 185.245 47.120 185.745 ;
        RECT 47.385 185.245 47.555 186.005 ;
        RECT 47.735 185.075 48.065 185.835 ;
        RECT 48.235 185.245 48.505 186.150 ;
        RECT 48.675 185.075 48.965 186.240 ;
        RECT 49.600 186.215 49.770 186.885 ;
        RECT 50.025 186.715 50.195 186.885 ;
        RECT 49.940 186.385 50.195 186.715 ;
        RECT 50.420 186.385 50.615 186.715 ;
        RECT 49.600 185.245 49.935 186.215 ;
        RECT 50.105 185.075 50.275 186.215 ;
        RECT 50.445 185.415 50.615 186.385 ;
        RECT 50.785 185.755 50.955 186.885 ;
        RECT 51.125 186.095 51.295 186.895 ;
        RECT 51.500 186.295 51.775 187.115 ;
        RECT 51.945 186.095 52.135 187.455 ;
        RECT 52.315 187.090 52.825 187.625 ;
        RECT 53.045 186.815 53.290 187.420 ;
        RECT 53.825 187.075 53.995 187.455 ;
        RECT 54.175 187.245 54.505 187.625 ;
        RECT 53.825 186.905 54.490 187.075 ;
        RECT 54.685 186.950 54.945 187.455 ;
        RECT 52.335 186.645 53.565 186.815 ;
        RECT 51.125 185.925 52.135 186.095 ;
        RECT 52.305 186.080 53.055 186.270 ;
        RECT 50.785 185.585 51.910 185.755 ;
        RECT 52.305 185.415 52.475 186.080 ;
        RECT 53.225 185.835 53.565 186.645 ;
        RECT 53.755 186.355 54.085 186.725 ;
        RECT 54.320 186.650 54.490 186.905 ;
        RECT 54.320 186.320 54.605 186.650 ;
        RECT 54.320 186.175 54.490 186.320 ;
        RECT 50.445 185.245 52.475 185.415 ;
        RECT 52.645 185.075 52.815 185.835 ;
        RECT 53.050 185.425 53.565 185.835 ;
        RECT 53.825 186.005 54.490 186.175 ;
        RECT 54.775 186.150 54.945 186.950 ;
        RECT 53.825 185.245 53.995 186.005 ;
        RECT 54.175 185.075 54.505 185.835 ;
        RECT 54.675 185.245 54.945 186.150 ;
        RECT 55.115 186.885 55.500 187.455 ;
        RECT 55.670 187.165 55.995 187.625 ;
        RECT 56.515 186.995 56.795 187.455 ;
        RECT 55.115 186.215 55.395 186.885 ;
        RECT 55.670 186.825 56.795 186.995 ;
        RECT 55.670 186.715 56.120 186.825 ;
        RECT 55.565 186.385 56.120 186.715 ;
        RECT 56.985 186.655 57.385 187.455 ;
        RECT 57.785 187.165 58.055 187.625 ;
        RECT 58.225 186.995 58.510 187.455 ;
        RECT 55.115 185.245 55.500 186.215 ;
        RECT 55.670 185.925 56.120 186.385 ;
        RECT 56.290 186.095 57.385 186.655 ;
        RECT 55.670 185.705 56.795 185.925 ;
        RECT 55.670 185.075 55.995 185.535 ;
        RECT 56.515 185.245 56.795 185.705 ;
        RECT 56.985 185.245 57.385 186.095 ;
        RECT 57.555 186.825 58.510 186.995 ;
        RECT 58.800 186.885 59.055 187.455 ;
        RECT 59.225 187.225 59.555 187.625 ;
        RECT 59.980 187.090 60.510 187.455 ;
        RECT 59.980 187.055 60.155 187.090 ;
        RECT 59.225 186.885 60.155 187.055 ;
        RECT 57.555 185.925 57.765 186.825 ;
        RECT 57.935 186.095 58.625 186.655 ;
        RECT 58.800 186.215 58.970 186.885 ;
        RECT 59.225 186.715 59.395 186.885 ;
        RECT 59.140 186.385 59.395 186.715 ;
        RECT 59.620 186.385 59.815 186.715 ;
        RECT 57.555 185.705 58.510 185.925 ;
        RECT 57.785 185.075 58.055 185.535 ;
        RECT 58.225 185.245 58.510 185.705 ;
        RECT 58.800 185.245 59.135 186.215 ;
        RECT 59.305 185.075 59.475 186.215 ;
        RECT 59.645 185.415 59.815 186.385 ;
        RECT 59.985 185.755 60.155 186.885 ;
        RECT 60.325 186.095 60.495 186.895 ;
        RECT 60.700 186.605 60.975 187.455 ;
        RECT 60.695 186.435 60.975 186.605 ;
        RECT 60.700 186.295 60.975 186.435 ;
        RECT 61.145 186.095 61.335 187.455 ;
        RECT 61.515 187.090 62.025 187.625 ;
        RECT 62.245 186.815 62.490 187.420 ;
        RECT 61.535 186.645 62.765 186.815 ;
        RECT 63.860 186.785 64.120 187.625 ;
        RECT 64.295 186.880 64.550 187.455 ;
        RECT 64.720 187.245 65.050 187.625 ;
        RECT 65.265 187.075 65.435 187.455 ;
        RECT 64.720 186.905 65.435 187.075 ;
        RECT 66.000 187.055 66.170 187.305 ;
        RECT 60.325 185.925 61.335 186.095 ;
        RECT 61.505 186.080 62.255 186.270 ;
        RECT 59.985 185.585 61.110 185.755 ;
        RECT 61.505 185.415 61.675 186.080 ;
        RECT 62.425 185.835 62.765 186.645 ;
        RECT 59.645 185.245 61.675 185.415 ;
        RECT 61.845 185.075 62.015 185.835 ;
        RECT 62.250 185.425 62.765 185.835 ;
        RECT 63.860 185.075 64.120 186.225 ;
        RECT 64.295 186.150 64.465 186.880 ;
        RECT 64.720 186.715 64.890 186.905 ;
        RECT 65.695 186.885 66.170 187.055 ;
        RECT 66.405 186.885 66.735 187.625 ;
        RECT 66.905 187.055 67.105 187.400 ;
        RECT 67.275 187.225 67.605 187.625 ;
        RECT 67.775 187.055 67.975 187.410 ;
        RECT 68.145 187.230 68.475 187.625 ;
        RECT 66.905 186.885 68.745 187.055 ;
        RECT 64.635 186.385 64.890 186.715 ;
        RECT 64.720 186.175 64.890 186.385 ;
        RECT 65.170 186.355 65.525 186.725 ;
        RECT 64.295 185.245 64.550 186.150 ;
        RECT 64.720 186.005 65.435 186.175 ;
        RECT 64.720 185.075 65.050 185.835 ;
        RECT 65.265 185.245 65.435 186.005 ;
        RECT 65.695 185.915 65.865 186.885 ;
        RECT 66.035 186.095 66.385 186.715 ;
        RECT 66.555 186.095 66.875 186.715 ;
        RECT 67.045 186.095 67.375 186.715 ;
        RECT 67.545 186.095 67.845 186.715 ;
        RECT 68.085 185.915 68.305 186.715 ;
        RECT 65.695 185.705 68.305 185.915 ;
        RECT 66.405 185.075 66.735 185.525 ;
        RECT 68.485 185.260 68.745 186.885 ;
        RECT 68.915 185.245 69.175 187.455 ;
        RECT 69.345 187.245 69.675 187.625 ;
        RECT 69.885 186.715 70.080 187.290 ;
        RECT 70.350 186.715 70.535 187.295 ;
        RECT 69.345 185.795 69.515 186.715 ;
        RECT 69.825 186.385 70.080 186.715 ;
        RECT 70.305 186.385 70.535 186.715 ;
        RECT 70.785 187.285 72.265 187.455 ;
        RECT 70.785 186.385 70.955 187.285 ;
        RECT 71.125 186.785 71.675 187.115 ;
        RECT 71.865 186.955 72.265 187.285 ;
        RECT 72.445 187.245 72.775 187.625 ;
        RECT 73.085 187.125 73.345 187.455 ;
        RECT 69.885 186.075 70.080 186.385 ;
        RECT 70.350 186.075 70.535 186.385 ;
        RECT 71.125 185.795 71.295 186.785 ;
        RECT 71.865 186.475 72.035 186.955 ;
        RECT 72.615 186.765 72.825 186.945 ;
        RECT 72.205 186.595 72.825 186.765 ;
        RECT 69.345 185.625 71.295 185.795 ;
        RECT 71.465 186.305 72.035 186.475 ;
        RECT 73.175 186.425 73.345 187.125 ;
        RECT 74.435 186.900 74.725 187.625 ;
        RECT 74.895 186.975 75.155 187.455 ;
        RECT 75.325 187.085 75.575 187.625 ;
        RECT 71.465 185.795 71.635 186.305 ;
        RECT 72.215 186.255 73.345 186.425 ;
        RECT 72.215 186.135 72.385 186.255 ;
        RECT 71.805 185.965 72.385 186.135 ;
        RECT 71.465 185.625 72.205 185.795 ;
        RECT 72.655 185.755 73.005 186.085 ;
        RECT 69.345 185.075 69.675 185.455 ;
        RECT 70.100 185.245 70.270 185.625 ;
        RECT 70.530 185.075 70.860 185.455 ;
        RECT 71.055 185.245 71.225 185.625 ;
        RECT 71.435 185.075 71.765 185.455 ;
        RECT 72.015 185.245 72.205 185.625 ;
        RECT 73.175 185.575 73.345 186.255 ;
        RECT 72.445 185.075 72.775 185.455 ;
        RECT 73.085 185.245 73.345 185.575 ;
        RECT 74.435 185.075 74.725 186.240 ;
        RECT 74.895 185.945 75.065 186.975 ;
        RECT 75.745 186.945 75.965 187.405 ;
        RECT 75.715 186.920 75.965 186.945 ;
        RECT 75.235 186.325 75.465 186.720 ;
        RECT 75.635 186.495 75.965 186.920 ;
        RECT 76.135 187.245 77.025 187.415 ;
        RECT 76.135 186.520 76.305 187.245 ;
        RECT 76.475 186.690 77.025 187.075 ;
        RECT 77.195 186.825 77.535 187.455 ;
        RECT 77.705 186.825 77.955 187.625 ;
        RECT 78.145 186.975 78.475 187.455 ;
        RECT 78.645 187.165 78.870 187.625 ;
        RECT 79.040 186.975 79.370 187.455 ;
        RECT 76.135 186.450 77.025 186.520 ;
        RECT 76.130 186.425 77.025 186.450 ;
        RECT 76.120 186.410 77.025 186.425 ;
        RECT 76.115 186.395 77.025 186.410 ;
        RECT 76.105 186.390 77.025 186.395 ;
        RECT 76.100 186.380 77.025 186.390 ;
        RECT 76.095 186.370 77.025 186.380 ;
        RECT 76.085 186.365 77.025 186.370 ;
        RECT 76.075 186.355 77.025 186.365 ;
        RECT 76.065 186.350 77.025 186.355 ;
        RECT 76.065 186.345 76.400 186.350 ;
        RECT 76.050 186.340 76.400 186.345 ;
        RECT 76.035 186.330 76.400 186.340 ;
        RECT 76.010 186.325 76.400 186.330 ;
        RECT 75.235 186.320 76.400 186.325 ;
        RECT 75.235 186.285 76.370 186.320 ;
        RECT 75.235 186.260 76.335 186.285 ;
        RECT 75.235 186.230 76.305 186.260 ;
        RECT 75.235 186.200 76.285 186.230 ;
        RECT 75.235 186.170 76.265 186.200 ;
        RECT 75.235 186.160 76.195 186.170 ;
        RECT 75.235 186.150 76.170 186.160 ;
        RECT 75.235 186.135 76.150 186.150 ;
        RECT 75.235 186.120 76.130 186.135 ;
        RECT 75.340 186.110 76.125 186.120 ;
        RECT 75.340 186.075 76.110 186.110 ;
        RECT 74.895 185.245 75.170 185.945 ;
        RECT 75.340 185.825 76.095 186.075 ;
        RECT 76.265 185.755 76.595 186.000 ;
        RECT 76.765 185.900 77.025 186.350 ;
        RECT 77.195 186.215 77.370 186.825 ;
        RECT 78.145 186.805 79.370 186.975 ;
        RECT 80.000 186.845 80.500 187.455 ;
        RECT 80.880 186.915 81.135 187.445 ;
        RECT 81.305 187.165 81.610 187.625 ;
        RECT 81.855 187.245 82.925 187.415 ;
        RECT 77.540 186.465 78.235 186.635 ;
        RECT 78.065 186.215 78.235 186.465 ;
        RECT 78.410 186.435 78.830 186.635 ;
        RECT 79.000 186.435 79.330 186.635 ;
        RECT 79.500 186.435 79.830 186.635 ;
        RECT 80.000 186.215 80.170 186.845 ;
        RECT 80.355 186.385 80.705 186.635 ;
        RECT 80.880 186.265 81.090 186.915 ;
        RECT 81.855 186.890 82.175 187.245 ;
        RECT 81.850 186.715 82.175 186.890 ;
        RECT 81.260 186.415 82.175 186.715 ;
        RECT 82.345 186.675 82.585 187.075 ;
        RECT 82.755 187.015 82.925 187.245 ;
        RECT 83.095 187.185 83.285 187.625 ;
        RECT 83.455 187.175 84.405 187.455 ;
        RECT 84.625 187.265 84.975 187.435 ;
        RECT 82.755 186.845 83.285 187.015 ;
        RECT 81.260 186.385 82.000 186.415 ;
        RECT 76.410 185.730 76.595 185.755 ;
        RECT 76.410 185.630 77.025 185.730 ;
        RECT 75.340 185.075 75.595 185.620 ;
        RECT 75.765 185.245 76.245 185.585 ;
        RECT 76.420 185.075 77.025 185.630 ;
        RECT 77.195 185.245 77.535 186.215 ;
        RECT 77.705 185.075 77.875 186.215 ;
        RECT 78.065 186.045 80.500 186.215 ;
        RECT 78.145 185.075 78.395 185.875 ;
        RECT 79.040 185.245 79.370 186.045 ;
        RECT 79.670 185.075 80.000 185.875 ;
        RECT 80.170 185.245 80.500 186.045 ;
        RECT 80.880 185.385 81.135 186.265 ;
        RECT 81.305 185.075 81.610 186.215 ;
        RECT 81.830 185.795 82.000 186.385 ;
        RECT 82.345 186.305 82.885 186.675 ;
        RECT 83.065 186.565 83.285 186.845 ;
        RECT 83.455 186.395 83.625 187.175 ;
        RECT 83.220 186.225 83.625 186.395 ;
        RECT 83.795 186.385 84.145 187.005 ;
        RECT 83.220 186.135 83.390 186.225 ;
        RECT 84.315 186.215 84.525 187.005 ;
        RECT 82.170 185.965 83.390 186.135 ;
        RECT 83.850 186.055 84.525 186.215 ;
        RECT 81.830 185.625 82.630 185.795 ;
        RECT 81.950 185.075 82.280 185.455 ;
        RECT 82.460 185.335 82.630 185.625 ;
        RECT 83.220 185.585 83.390 185.965 ;
        RECT 83.560 186.045 84.525 186.055 ;
        RECT 84.715 186.875 84.975 187.265 ;
        RECT 85.185 187.165 85.515 187.625 ;
        RECT 86.390 187.235 87.245 187.405 ;
        RECT 87.450 187.235 87.945 187.405 ;
        RECT 88.115 187.265 88.445 187.625 ;
        RECT 84.715 186.185 84.885 186.875 ;
        RECT 85.055 186.525 85.225 186.705 ;
        RECT 85.395 186.695 86.185 186.945 ;
        RECT 86.390 186.525 86.560 187.235 ;
        RECT 86.730 186.725 87.085 186.945 ;
        RECT 85.055 186.355 86.745 186.525 ;
        RECT 83.560 185.755 84.020 186.045 ;
        RECT 84.715 186.015 86.215 186.185 ;
        RECT 84.715 185.875 84.885 186.015 ;
        RECT 84.325 185.705 84.885 185.875 ;
        RECT 82.800 185.075 83.050 185.535 ;
        RECT 83.220 185.245 84.090 185.585 ;
        RECT 84.325 185.245 84.495 185.705 ;
        RECT 85.330 185.675 86.405 185.845 ;
        RECT 84.665 185.075 85.035 185.535 ;
        RECT 85.330 185.335 85.500 185.675 ;
        RECT 85.670 185.075 86.000 185.505 ;
        RECT 86.235 185.335 86.405 185.675 ;
        RECT 86.575 185.575 86.745 186.355 ;
        RECT 86.915 186.135 87.085 186.725 ;
        RECT 87.255 186.325 87.605 186.945 ;
        RECT 86.915 185.745 87.380 186.135 ;
        RECT 87.775 185.875 87.945 187.235 ;
        RECT 88.115 186.045 88.575 187.095 ;
        RECT 87.550 185.705 87.945 185.875 ;
        RECT 87.550 185.575 87.720 185.705 ;
        RECT 86.575 185.245 87.255 185.575 ;
        RECT 87.470 185.245 87.720 185.575 ;
        RECT 87.890 185.075 88.140 185.535 ;
        RECT 88.310 185.260 88.635 186.045 ;
        RECT 88.805 185.245 88.975 187.365 ;
        RECT 89.145 187.245 89.475 187.625 ;
        RECT 89.645 187.075 89.900 187.365 ;
        RECT 89.150 186.905 89.900 187.075 ;
        RECT 90.190 186.995 90.475 187.455 ;
        RECT 90.645 187.165 90.915 187.625 ;
        RECT 89.150 185.915 89.380 186.905 ;
        RECT 90.190 186.825 91.145 186.995 ;
        RECT 89.550 186.085 89.900 186.735 ;
        RECT 90.075 186.095 90.765 186.655 ;
        RECT 90.935 185.925 91.145 186.825 ;
        RECT 89.150 185.745 89.900 185.915 ;
        RECT 89.145 185.075 89.475 185.575 ;
        RECT 89.645 185.245 89.900 185.745 ;
        RECT 90.190 185.705 91.145 185.925 ;
        RECT 91.315 186.655 91.715 187.455 ;
        RECT 91.905 186.995 92.185 187.455 ;
        RECT 92.705 187.165 93.030 187.625 ;
        RECT 91.905 186.825 93.030 186.995 ;
        RECT 93.200 186.885 93.585 187.455 ;
        RECT 92.580 186.715 93.030 186.825 ;
        RECT 91.315 186.095 92.410 186.655 ;
        RECT 92.580 186.385 93.135 186.715 ;
        RECT 90.190 185.245 90.475 185.705 ;
        RECT 90.645 185.075 90.915 185.535 ;
        RECT 91.315 185.245 91.715 186.095 ;
        RECT 92.580 185.925 93.030 186.385 ;
        RECT 93.305 186.215 93.585 186.885 ;
        RECT 91.905 185.705 93.030 185.925 ;
        RECT 91.905 185.245 92.185 185.705 ;
        RECT 92.705 185.075 93.030 185.535 ;
        RECT 93.200 185.245 93.585 186.215 ;
        RECT 93.755 186.825 94.095 187.455 ;
        RECT 94.265 186.825 94.515 187.625 ;
        RECT 94.705 186.975 95.035 187.455 ;
        RECT 95.205 187.165 95.430 187.625 ;
        RECT 95.600 186.975 95.930 187.455 ;
        RECT 93.755 186.215 93.930 186.825 ;
        RECT 94.705 186.805 95.930 186.975 ;
        RECT 96.560 186.845 97.060 187.455 ;
        RECT 97.525 186.975 97.695 187.455 ;
        RECT 97.875 187.145 98.115 187.625 ;
        RECT 98.365 186.975 98.535 187.455 ;
        RECT 98.705 187.145 99.035 187.625 ;
        RECT 99.205 186.975 99.375 187.455 ;
        RECT 94.100 186.465 94.795 186.635 ;
        RECT 94.625 186.215 94.795 186.465 ;
        RECT 94.970 186.435 95.390 186.635 ;
        RECT 95.560 186.435 95.890 186.635 ;
        RECT 96.060 186.435 96.390 186.635 ;
        RECT 96.560 186.215 96.730 186.845 ;
        RECT 97.525 186.805 98.160 186.975 ;
        RECT 98.365 186.805 99.375 186.975 ;
        RECT 99.545 186.825 99.875 187.625 ;
        RECT 100.195 186.900 100.485 187.625 ;
        RECT 100.930 186.815 101.175 187.420 ;
        RECT 101.395 187.090 101.905 187.625 ;
        RECT 97.990 186.635 98.160 186.805 ;
        RECT 96.915 186.385 97.265 186.635 ;
        RECT 97.440 186.395 97.820 186.635 ;
        RECT 97.990 186.465 98.490 186.635 ;
        RECT 97.990 186.225 98.160 186.465 ;
        RECT 98.880 186.265 99.375 186.805 ;
        RECT 93.755 185.245 94.095 186.215 ;
        RECT 94.265 185.075 94.435 186.215 ;
        RECT 94.625 186.045 97.060 186.215 ;
        RECT 94.705 185.075 94.955 185.875 ;
        RECT 95.600 185.245 95.930 186.045 ;
        RECT 96.230 185.075 96.560 185.875 ;
        RECT 96.730 185.245 97.060 186.045 ;
        RECT 97.445 186.055 98.160 186.225 ;
        RECT 98.365 186.095 99.375 186.265 ;
        RECT 100.655 186.645 101.885 186.815 ;
        RECT 97.445 185.245 97.775 186.055 ;
        RECT 97.945 185.075 98.185 185.875 ;
        RECT 98.365 185.245 98.535 186.095 ;
        RECT 98.705 185.075 99.035 185.875 ;
        RECT 99.205 185.245 99.375 186.095 ;
        RECT 99.545 185.075 99.875 186.225 ;
        RECT 100.195 185.075 100.485 186.240 ;
        RECT 100.655 185.835 100.995 186.645 ;
        RECT 101.165 186.080 101.915 186.270 ;
        RECT 100.655 185.425 101.170 185.835 ;
        RECT 101.405 185.075 101.575 185.835 ;
        RECT 101.745 185.415 101.915 186.080 ;
        RECT 102.085 186.095 102.275 187.455 ;
        RECT 102.445 186.945 102.720 187.455 ;
        RECT 102.910 187.090 103.440 187.455 ;
        RECT 103.865 187.225 104.195 187.625 ;
        RECT 103.265 187.055 103.440 187.090 ;
        RECT 102.445 186.775 102.725 186.945 ;
        RECT 102.445 186.295 102.720 186.775 ;
        RECT 102.925 186.095 103.095 186.895 ;
        RECT 102.085 185.925 103.095 186.095 ;
        RECT 103.265 186.885 104.195 187.055 ;
        RECT 104.365 186.885 104.620 187.455 ;
        RECT 103.265 185.755 103.435 186.885 ;
        RECT 104.025 186.715 104.195 186.885 ;
        RECT 102.310 185.585 103.435 185.755 ;
        RECT 103.605 186.385 103.800 186.715 ;
        RECT 104.025 186.385 104.280 186.715 ;
        RECT 103.605 185.415 103.775 186.385 ;
        RECT 104.450 186.215 104.620 186.885 ;
        RECT 101.745 185.245 103.775 185.415 ;
        RECT 103.945 185.075 104.115 186.215 ;
        RECT 104.285 185.245 104.620 186.215 ;
        RECT 104.795 186.885 105.180 187.455 ;
        RECT 105.350 187.165 105.675 187.625 ;
        RECT 106.195 186.995 106.475 187.455 ;
        RECT 104.795 186.215 105.075 186.885 ;
        RECT 105.350 186.825 106.475 186.995 ;
        RECT 105.350 186.715 105.800 186.825 ;
        RECT 105.245 186.385 105.800 186.715 ;
        RECT 106.665 186.655 107.065 187.455 ;
        RECT 107.465 187.165 107.735 187.625 ;
        RECT 107.905 186.995 108.190 187.455 ;
        RECT 104.795 185.245 105.180 186.215 ;
        RECT 105.350 185.925 105.800 186.385 ;
        RECT 105.970 186.095 107.065 186.655 ;
        RECT 105.350 185.705 106.475 185.925 ;
        RECT 105.350 185.075 105.675 185.535 ;
        RECT 106.195 185.245 106.475 185.705 ;
        RECT 106.665 185.245 107.065 186.095 ;
        RECT 107.235 186.825 108.190 186.995 ;
        RECT 108.680 186.845 109.180 187.455 ;
        RECT 107.235 185.925 107.445 186.825 ;
        RECT 107.615 186.095 108.305 186.655 ;
        RECT 108.475 186.385 108.825 186.635 ;
        RECT 109.010 186.215 109.180 186.845 ;
        RECT 109.810 186.975 110.140 187.455 ;
        RECT 110.310 187.165 110.535 187.625 ;
        RECT 110.705 186.975 111.035 187.455 ;
        RECT 109.810 186.805 111.035 186.975 ;
        RECT 111.225 186.825 111.475 187.625 ;
        RECT 111.645 186.825 111.985 187.455 ;
        RECT 112.155 186.875 113.365 187.625 ;
        RECT 109.350 186.435 109.680 186.635 ;
        RECT 109.850 186.435 110.180 186.635 ;
        RECT 110.350 186.435 110.770 186.635 ;
        RECT 110.945 186.465 111.640 186.635 ;
        RECT 110.945 186.215 111.115 186.465 ;
        RECT 111.810 186.265 111.985 186.825 ;
        RECT 111.755 186.215 111.985 186.265 ;
        RECT 108.680 186.045 111.115 186.215 ;
        RECT 107.235 185.705 108.190 185.925 ;
        RECT 107.465 185.075 107.735 185.535 ;
        RECT 107.905 185.245 108.190 185.705 ;
        RECT 108.680 185.245 109.010 186.045 ;
        RECT 109.180 185.075 109.510 185.875 ;
        RECT 109.810 185.245 110.140 186.045 ;
        RECT 110.785 185.075 111.035 185.875 ;
        RECT 111.305 185.075 111.475 186.215 ;
        RECT 111.645 185.245 111.985 186.215 ;
        RECT 112.155 186.165 112.675 186.705 ;
        RECT 112.845 186.335 113.365 186.875 ;
        RECT 112.155 185.075 113.365 186.165 ;
        RECT 26.970 184.905 113.450 185.075 ;
        RECT 27.055 183.815 28.265 184.905 ;
        RECT 27.055 183.105 27.575 183.645 ;
        RECT 27.745 183.275 28.265 183.815 ;
        RECT 28.955 183.765 29.165 184.905 ;
        RECT 29.335 183.755 29.665 184.735 ;
        RECT 29.835 183.765 30.065 184.905 ;
        RECT 30.315 183.765 30.545 184.905 ;
        RECT 30.715 183.755 31.045 184.735 ;
        RECT 31.215 183.765 31.425 184.905 ;
        RECT 31.660 183.765 31.995 184.735 ;
        RECT 32.165 183.765 32.335 184.905 ;
        RECT 32.505 184.565 34.535 184.735 ;
        RECT 27.055 182.355 28.265 183.105 ;
        RECT 28.955 182.355 29.165 183.175 ;
        RECT 29.335 183.155 29.585 183.755 ;
        RECT 29.755 183.345 30.085 183.595 ;
        RECT 30.295 183.345 30.625 183.595 ;
        RECT 29.335 182.525 29.665 183.155 ;
        RECT 29.835 182.355 30.065 183.175 ;
        RECT 30.315 182.355 30.545 183.175 ;
        RECT 30.795 183.155 31.045 183.755 ;
        RECT 30.715 182.525 31.045 183.155 ;
        RECT 31.215 182.355 31.425 183.175 ;
        RECT 31.660 183.095 31.830 183.765 ;
        RECT 32.505 183.595 32.675 184.565 ;
        RECT 32.000 183.265 32.255 183.595 ;
        RECT 32.480 183.265 32.675 183.595 ;
        RECT 32.845 184.225 33.970 184.395 ;
        RECT 32.085 183.095 32.255 183.265 ;
        RECT 32.845 183.095 33.015 184.225 ;
        RECT 31.660 182.525 31.915 183.095 ;
        RECT 32.085 182.925 33.015 183.095 ;
        RECT 33.185 183.885 34.195 184.055 ;
        RECT 33.185 183.085 33.355 183.885 ;
        RECT 33.560 183.545 33.835 183.685 ;
        RECT 33.555 183.375 33.835 183.545 ;
        RECT 32.840 182.890 33.015 182.925 ;
        RECT 32.085 182.355 32.415 182.755 ;
        RECT 32.840 182.525 33.370 182.890 ;
        RECT 33.560 182.525 33.835 183.375 ;
        RECT 34.005 182.525 34.195 183.885 ;
        RECT 34.365 183.900 34.535 184.565 ;
        RECT 34.705 184.145 34.875 184.905 ;
        RECT 35.110 184.145 35.625 184.555 ;
        RECT 34.365 183.710 35.115 183.900 ;
        RECT 35.285 183.335 35.625 184.145 ;
        RECT 35.795 183.740 36.085 184.905 ;
        RECT 36.720 183.765 37.055 184.735 ;
        RECT 37.225 183.765 37.395 184.905 ;
        RECT 37.565 184.565 39.595 184.735 ;
        RECT 34.395 183.165 35.625 183.335 ;
        RECT 34.375 182.355 34.885 182.890 ;
        RECT 35.105 182.560 35.350 183.165 ;
        RECT 36.720 183.095 36.890 183.765 ;
        RECT 37.565 183.595 37.735 184.565 ;
        RECT 37.060 183.265 37.315 183.595 ;
        RECT 37.540 183.265 37.735 183.595 ;
        RECT 37.905 184.225 39.030 184.395 ;
        RECT 37.145 183.095 37.315 183.265 ;
        RECT 37.905 183.095 38.075 184.225 ;
        RECT 35.795 182.355 36.085 183.080 ;
        RECT 36.720 182.525 36.975 183.095 ;
        RECT 37.145 182.925 38.075 183.095 ;
        RECT 38.245 183.885 39.255 184.055 ;
        RECT 38.245 183.085 38.415 183.885 ;
        RECT 38.620 183.205 38.895 183.685 ;
        RECT 38.615 183.035 38.895 183.205 ;
        RECT 37.900 182.890 38.075 182.925 ;
        RECT 37.145 182.355 37.475 182.755 ;
        RECT 37.900 182.525 38.430 182.890 ;
        RECT 38.620 182.525 38.895 183.035 ;
        RECT 39.065 182.525 39.255 183.885 ;
        RECT 39.425 183.900 39.595 184.565 ;
        RECT 39.765 184.145 39.935 184.905 ;
        RECT 40.170 184.145 40.685 184.555 ;
        RECT 39.425 183.710 40.175 183.900 ;
        RECT 40.345 183.335 40.685 184.145 ;
        RECT 39.455 183.165 40.685 183.335 ;
        RECT 41.320 183.765 41.655 184.735 ;
        RECT 41.825 183.765 41.995 184.905 ;
        RECT 42.165 184.565 44.195 184.735 ;
        RECT 39.435 182.355 39.945 182.890 ;
        RECT 40.165 182.560 40.410 183.165 ;
        RECT 41.320 183.095 41.490 183.765 ;
        RECT 42.165 183.595 42.335 184.565 ;
        RECT 41.660 183.265 41.915 183.595 ;
        RECT 42.140 183.265 42.335 183.595 ;
        RECT 42.505 184.225 43.630 184.395 ;
        RECT 41.745 183.095 41.915 183.265 ;
        RECT 42.505 183.095 42.675 184.225 ;
        RECT 41.320 182.525 41.575 183.095 ;
        RECT 41.745 182.925 42.675 183.095 ;
        RECT 42.845 183.885 43.855 184.055 ;
        RECT 42.845 183.085 43.015 183.885 ;
        RECT 43.220 183.545 43.495 183.685 ;
        RECT 43.215 183.375 43.495 183.545 ;
        RECT 42.500 182.890 42.675 182.925 ;
        RECT 41.745 182.355 42.075 182.755 ;
        RECT 42.500 182.525 43.030 182.890 ;
        RECT 43.220 182.525 43.495 183.375 ;
        RECT 43.665 182.525 43.855 183.885 ;
        RECT 44.025 183.900 44.195 184.565 ;
        RECT 44.365 184.145 44.535 184.905 ;
        RECT 44.770 184.145 45.285 184.555 ;
        RECT 44.025 183.710 44.775 183.900 ;
        RECT 44.945 183.335 45.285 184.145 ;
        RECT 44.055 183.165 45.285 183.335 ;
        RECT 45.460 183.715 45.715 184.595 ;
        RECT 45.885 183.765 46.190 184.905 ;
        RECT 46.530 184.525 46.860 184.905 ;
        RECT 47.040 184.355 47.210 184.645 ;
        RECT 47.380 184.445 47.630 184.905 ;
        RECT 46.410 184.185 47.210 184.355 ;
        RECT 47.800 184.395 48.670 184.735 ;
        RECT 44.035 182.355 44.545 182.890 ;
        RECT 44.765 182.560 45.010 183.165 ;
        RECT 45.460 183.065 45.670 183.715 ;
        RECT 46.410 183.595 46.580 184.185 ;
        RECT 47.800 184.015 47.970 184.395 ;
        RECT 48.905 184.275 49.075 184.735 ;
        RECT 49.245 184.445 49.615 184.905 ;
        RECT 49.910 184.305 50.080 184.645 ;
        RECT 50.250 184.475 50.580 184.905 ;
        RECT 50.815 184.305 50.985 184.645 ;
        RECT 46.750 183.845 47.970 184.015 ;
        RECT 48.140 183.935 48.600 184.225 ;
        RECT 48.905 184.105 49.465 184.275 ;
        RECT 49.910 184.135 50.985 184.305 ;
        RECT 51.155 184.405 51.835 184.735 ;
        RECT 52.050 184.405 52.300 184.735 ;
        RECT 52.470 184.445 52.720 184.905 ;
        RECT 49.295 183.965 49.465 184.105 ;
        RECT 48.140 183.925 49.105 183.935 ;
        RECT 47.800 183.755 47.970 183.845 ;
        RECT 48.430 183.765 49.105 183.925 ;
        RECT 45.840 183.565 46.580 183.595 ;
        RECT 45.840 183.265 46.755 183.565 ;
        RECT 46.430 183.090 46.755 183.265 ;
        RECT 45.460 182.535 45.715 183.065 ;
        RECT 45.885 182.355 46.190 182.815 ;
        RECT 46.435 182.735 46.755 183.090 ;
        RECT 46.925 183.305 47.465 183.675 ;
        RECT 47.800 183.585 48.205 183.755 ;
        RECT 46.925 182.905 47.165 183.305 ;
        RECT 47.645 183.135 47.865 183.415 ;
        RECT 47.335 182.965 47.865 183.135 ;
        RECT 47.335 182.735 47.505 182.965 ;
        RECT 48.035 182.805 48.205 183.585 ;
        RECT 48.375 182.975 48.725 183.595 ;
        RECT 48.895 182.975 49.105 183.765 ;
        RECT 49.295 183.795 50.795 183.965 ;
        RECT 49.295 183.105 49.465 183.795 ;
        RECT 51.155 183.625 51.325 184.405 ;
        RECT 52.130 184.275 52.300 184.405 ;
        RECT 49.635 183.455 51.325 183.625 ;
        RECT 51.495 183.845 51.960 184.235 ;
        RECT 52.130 184.105 52.525 184.275 ;
        RECT 49.635 183.275 49.805 183.455 ;
        RECT 46.435 182.565 47.505 182.735 ;
        RECT 47.675 182.355 47.865 182.795 ;
        RECT 48.035 182.525 48.985 182.805 ;
        RECT 49.295 182.715 49.555 183.105 ;
        RECT 49.975 183.035 50.765 183.285 ;
        RECT 49.205 182.545 49.555 182.715 ;
        RECT 49.765 182.355 50.095 182.815 ;
        RECT 50.970 182.745 51.140 183.455 ;
        RECT 51.495 183.255 51.665 183.845 ;
        RECT 51.310 183.035 51.665 183.255 ;
        RECT 51.835 183.035 52.185 183.655 ;
        RECT 52.355 182.745 52.525 184.105 ;
        RECT 52.890 183.935 53.215 184.720 ;
        RECT 52.695 182.885 53.155 183.935 ;
        RECT 50.970 182.575 51.825 182.745 ;
        RECT 52.030 182.575 52.525 182.745 ;
        RECT 52.695 182.355 53.025 182.715 ;
        RECT 53.385 182.615 53.555 184.735 ;
        RECT 53.725 184.405 54.055 184.905 ;
        RECT 54.225 184.235 54.480 184.735 ;
        RECT 53.730 184.065 54.480 184.235 ;
        RECT 53.730 183.075 53.960 184.065 ;
        RECT 54.710 184.035 54.995 184.905 ;
        RECT 55.165 184.275 55.425 184.735 ;
        RECT 55.600 184.445 55.855 184.905 ;
        RECT 56.025 184.275 56.285 184.735 ;
        RECT 55.165 184.105 56.285 184.275 ;
        RECT 56.455 184.105 56.765 184.905 ;
        RECT 54.130 183.245 54.480 183.895 ;
        RECT 55.165 183.855 55.425 184.105 ;
        RECT 56.935 183.935 57.245 184.735 ;
        RECT 54.670 183.685 55.425 183.855 ;
        RECT 56.215 183.765 57.245 183.935 ;
        RECT 54.670 183.175 55.075 183.685 ;
        RECT 56.215 183.515 56.385 183.765 ;
        RECT 55.245 183.345 56.385 183.515 ;
        RECT 53.730 182.905 54.480 183.075 ;
        RECT 54.670 183.005 56.320 183.175 ;
        RECT 56.555 183.025 56.905 183.595 ;
        RECT 53.725 182.355 54.055 182.735 ;
        RECT 54.225 182.615 54.480 182.905 ;
        RECT 54.715 182.355 54.995 182.835 ;
        RECT 55.165 182.615 55.425 183.005 ;
        RECT 55.600 182.355 55.855 182.835 ;
        RECT 56.025 182.615 56.320 183.005 ;
        RECT 57.075 182.855 57.245 183.765 ;
        RECT 57.415 184.145 57.930 184.555 ;
        RECT 58.165 184.145 58.335 184.905 ;
        RECT 58.505 184.565 60.535 184.735 ;
        RECT 57.415 183.335 57.755 184.145 ;
        RECT 58.505 183.900 58.675 184.565 ;
        RECT 59.070 184.225 60.195 184.395 ;
        RECT 57.925 183.710 58.675 183.900 ;
        RECT 58.845 183.885 59.855 184.055 ;
        RECT 57.415 183.165 58.645 183.335 ;
        RECT 56.500 182.355 56.775 182.835 ;
        RECT 56.945 182.525 57.245 182.855 ;
        RECT 57.690 182.560 57.935 183.165 ;
        RECT 58.155 182.355 58.665 182.890 ;
        RECT 58.845 182.525 59.035 183.885 ;
        RECT 59.205 183.205 59.480 183.685 ;
        RECT 59.205 183.035 59.485 183.205 ;
        RECT 59.685 183.085 59.855 183.885 ;
        RECT 60.025 183.095 60.195 184.225 ;
        RECT 60.365 183.595 60.535 184.565 ;
        RECT 60.705 183.765 60.875 184.905 ;
        RECT 61.045 183.765 61.380 184.735 ;
        RECT 60.365 183.265 60.560 183.595 ;
        RECT 60.785 183.265 61.040 183.595 ;
        RECT 60.785 183.095 60.955 183.265 ;
        RECT 61.210 183.095 61.380 183.765 ;
        RECT 61.555 183.740 61.845 184.905 ;
        RECT 62.015 183.765 62.400 184.735 ;
        RECT 62.570 184.445 62.895 184.905 ;
        RECT 63.415 184.275 63.695 184.735 ;
        RECT 62.570 184.055 63.695 184.275 ;
        RECT 59.205 182.525 59.480 183.035 ;
        RECT 60.025 182.925 60.955 183.095 ;
        RECT 60.025 182.890 60.200 182.925 ;
        RECT 59.670 182.525 60.200 182.890 ;
        RECT 60.625 182.355 60.955 182.755 ;
        RECT 61.125 182.525 61.380 183.095 ;
        RECT 62.015 183.095 62.295 183.765 ;
        RECT 62.570 183.595 63.020 184.055 ;
        RECT 63.885 183.885 64.285 184.735 ;
        RECT 64.685 184.445 64.955 184.905 ;
        RECT 65.125 184.275 65.410 184.735 ;
        RECT 62.465 183.265 63.020 183.595 ;
        RECT 63.190 183.325 64.285 183.885 ;
        RECT 62.570 183.155 63.020 183.265 ;
        RECT 61.555 182.355 61.845 183.080 ;
        RECT 62.015 182.525 62.400 183.095 ;
        RECT 62.570 182.985 63.695 183.155 ;
        RECT 62.570 182.355 62.895 182.815 ;
        RECT 63.415 182.525 63.695 182.985 ;
        RECT 63.885 182.525 64.285 183.325 ;
        RECT 64.455 184.055 65.410 184.275 ;
        RECT 64.455 183.155 64.665 184.055 ;
        RECT 64.835 183.325 65.525 183.885 ;
        RECT 65.695 183.765 66.080 184.735 ;
        RECT 66.250 184.445 66.575 184.905 ;
        RECT 67.095 184.275 67.375 184.735 ;
        RECT 66.250 184.055 67.375 184.275 ;
        RECT 64.455 182.985 65.410 183.155 ;
        RECT 64.685 182.355 64.955 182.815 ;
        RECT 65.125 182.525 65.410 182.985 ;
        RECT 65.695 183.095 65.975 183.765 ;
        RECT 66.250 183.595 66.700 184.055 ;
        RECT 67.565 183.885 67.965 184.735 ;
        RECT 68.365 184.445 68.635 184.905 ;
        RECT 68.805 184.275 69.090 184.735 ;
        RECT 66.145 183.265 66.700 183.595 ;
        RECT 66.870 183.325 67.965 183.885 ;
        RECT 66.250 183.155 66.700 183.265 ;
        RECT 65.695 182.525 66.080 183.095 ;
        RECT 66.250 182.985 67.375 183.155 ;
        RECT 66.250 182.355 66.575 182.815 ;
        RECT 67.095 182.525 67.375 182.985 ;
        RECT 67.565 182.525 67.965 183.325 ;
        RECT 68.135 184.055 69.090 184.275 ;
        RECT 68.135 183.155 68.345 184.055 ;
        RECT 70.500 183.935 70.830 184.735 ;
        RECT 71.000 184.105 71.330 184.905 ;
        RECT 71.630 183.935 71.960 184.735 ;
        RECT 72.605 184.105 72.855 184.905 ;
        RECT 68.515 183.325 69.205 183.885 ;
        RECT 70.500 183.765 72.935 183.935 ;
        RECT 73.125 183.765 73.295 184.905 ;
        RECT 73.465 183.765 73.805 184.735 ;
        RECT 70.295 183.345 70.645 183.595 ;
        RECT 68.135 182.985 69.090 183.155 ;
        RECT 70.830 183.135 71.000 183.765 ;
        RECT 71.170 183.345 71.500 183.545 ;
        RECT 71.670 183.345 72.000 183.545 ;
        RECT 72.170 183.345 72.590 183.545 ;
        RECT 72.765 183.515 72.935 183.765 ;
        RECT 73.575 183.715 73.805 183.765 ;
        RECT 72.765 183.345 73.460 183.515 ;
        RECT 68.365 182.355 68.635 182.815 ;
        RECT 68.805 182.525 69.090 182.985 ;
        RECT 70.500 182.525 71.000 183.135 ;
        RECT 71.630 183.005 72.855 183.175 ;
        RECT 73.630 183.155 73.805 183.715 ;
        RECT 71.630 182.525 71.960 183.005 ;
        RECT 72.130 182.355 72.355 182.815 ;
        RECT 72.525 182.525 72.855 183.005 ;
        RECT 73.045 182.355 73.295 183.155 ;
        RECT 73.465 182.525 73.805 183.155 ;
        RECT 73.975 183.765 74.315 184.735 ;
        RECT 74.485 183.765 74.655 184.905 ;
        RECT 74.925 184.105 75.175 184.905 ;
        RECT 75.820 183.935 76.150 184.735 ;
        RECT 76.450 184.105 76.780 184.905 ;
        RECT 76.950 183.935 77.280 184.735 ;
        RECT 74.845 183.765 77.280 183.935 ;
        RECT 77.655 183.765 77.995 184.735 ;
        RECT 78.165 183.765 78.335 184.905 ;
        RECT 78.605 184.105 78.855 184.905 ;
        RECT 79.500 183.935 79.830 184.735 ;
        RECT 80.130 184.105 80.460 184.905 ;
        RECT 80.630 183.935 80.960 184.735 ;
        RECT 81.850 184.105 82.150 184.905 ;
        RECT 82.320 183.935 82.650 184.735 ;
        RECT 82.820 184.105 82.990 184.905 ;
        RECT 83.160 183.935 83.490 184.735 ;
        RECT 83.660 184.105 83.830 184.905 ;
        RECT 84.000 183.935 84.330 184.735 ;
        RECT 84.500 184.105 84.670 184.905 ;
        RECT 84.840 183.935 85.170 184.735 ;
        RECT 85.340 184.105 85.595 184.905 ;
        RECT 78.525 183.765 80.960 183.935 ;
        RECT 81.795 183.765 85.765 183.935 ;
        RECT 85.975 183.765 86.205 184.905 ;
        RECT 73.975 183.155 74.150 183.765 ;
        RECT 74.845 183.515 75.015 183.765 ;
        RECT 74.320 183.345 75.015 183.515 ;
        RECT 75.190 183.345 75.610 183.545 ;
        RECT 75.780 183.345 76.110 183.545 ;
        RECT 76.280 183.345 76.610 183.545 ;
        RECT 73.975 182.525 74.315 183.155 ;
        RECT 74.485 182.355 74.735 183.155 ;
        RECT 74.925 183.005 76.150 183.175 ;
        RECT 74.925 182.525 75.255 183.005 ;
        RECT 75.425 182.355 75.650 182.815 ;
        RECT 75.820 182.525 76.150 183.005 ;
        RECT 76.780 183.135 76.950 183.765 ;
        RECT 77.135 183.345 77.485 183.595 ;
        RECT 77.655 183.155 77.830 183.765 ;
        RECT 78.525 183.515 78.695 183.765 ;
        RECT 78.000 183.345 78.695 183.515 ;
        RECT 78.870 183.345 79.290 183.545 ;
        RECT 79.460 183.345 79.790 183.545 ;
        RECT 79.960 183.345 80.290 183.545 ;
        RECT 76.780 182.525 77.280 183.135 ;
        RECT 77.655 182.525 77.995 183.155 ;
        RECT 78.165 182.355 78.415 183.155 ;
        RECT 78.605 183.005 79.830 183.175 ;
        RECT 78.605 182.525 78.935 183.005 ;
        RECT 79.105 182.355 79.330 182.815 ;
        RECT 79.500 182.525 79.830 183.005 ;
        RECT 80.460 183.135 80.630 183.765 ;
        RECT 80.815 183.345 81.165 183.595 ;
        RECT 81.795 183.175 82.115 183.765 ;
        RECT 82.315 183.545 85.170 183.595 ;
        RECT 82.315 183.375 85.245 183.545 ;
        RECT 82.315 183.345 85.170 183.375 ;
        RECT 85.420 183.175 85.765 183.765 ;
        RECT 86.375 183.755 86.705 184.735 ;
        RECT 86.875 183.765 87.085 184.905 ;
        RECT 85.955 183.345 86.285 183.595 ;
        RECT 80.460 182.525 80.960 183.135 ;
        RECT 81.795 182.985 85.765 183.175 ;
        RECT 81.845 182.355 82.150 182.815 ;
        RECT 82.320 182.525 82.650 182.985 ;
        RECT 82.820 182.355 82.990 182.815 ;
        RECT 83.160 182.525 83.490 182.985 ;
        RECT 83.660 182.355 83.830 182.815 ;
        RECT 84.000 182.525 84.330 182.985 ;
        RECT 84.500 182.355 84.670 182.815 ;
        RECT 84.840 182.525 85.170 182.985 ;
        RECT 85.340 182.355 85.595 182.815 ;
        RECT 85.975 182.355 86.205 183.175 ;
        RECT 86.455 183.155 86.705 183.755 ;
        RECT 87.315 183.740 87.605 184.905 ;
        RECT 88.900 183.935 89.230 184.735 ;
        RECT 89.400 184.105 89.730 184.905 ;
        RECT 90.030 183.935 90.360 184.735 ;
        RECT 91.005 184.105 91.255 184.905 ;
        RECT 88.900 183.765 91.335 183.935 ;
        RECT 91.525 183.765 91.695 184.905 ;
        RECT 91.865 183.765 92.205 184.735 ;
        RECT 92.490 184.275 92.775 184.735 ;
        RECT 92.945 184.445 93.215 184.905 ;
        RECT 92.490 184.055 93.445 184.275 ;
        RECT 88.695 183.345 89.045 183.595 ;
        RECT 86.375 182.525 86.705 183.155 ;
        RECT 86.875 182.355 87.085 183.175 ;
        RECT 89.230 183.135 89.400 183.765 ;
        RECT 89.570 183.345 89.900 183.545 ;
        RECT 90.070 183.345 90.400 183.545 ;
        RECT 90.570 183.345 90.990 183.545 ;
        RECT 91.165 183.515 91.335 183.765 ;
        RECT 91.165 183.345 91.860 183.515 ;
        RECT 87.315 182.355 87.605 183.080 ;
        RECT 88.900 182.525 89.400 183.135 ;
        RECT 90.030 183.005 91.255 183.175 ;
        RECT 92.030 183.155 92.205 183.765 ;
        RECT 92.375 183.325 93.065 183.885 ;
        RECT 93.235 183.155 93.445 184.055 ;
        RECT 90.030 182.525 90.360 183.005 ;
        RECT 90.530 182.355 90.755 182.815 ;
        RECT 90.925 182.525 91.255 183.005 ;
        RECT 91.445 182.355 91.695 183.155 ;
        RECT 91.865 182.525 92.205 183.155 ;
        RECT 92.490 182.985 93.445 183.155 ;
        RECT 93.615 183.885 94.015 184.735 ;
        RECT 94.205 184.275 94.485 184.735 ;
        RECT 95.005 184.445 95.330 184.905 ;
        RECT 94.205 184.055 95.330 184.275 ;
        RECT 93.615 183.325 94.710 183.885 ;
        RECT 94.880 183.595 95.330 184.055 ;
        RECT 95.500 183.765 95.885 184.735 ;
        RECT 96.115 183.765 96.325 184.905 ;
        RECT 92.490 182.525 92.775 182.985 ;
        RECT 92.945 182.355 93.215 182.815 ;
        RECT 93.615 182.525 94.015 183.325 ;
        RECT 94.880 183.265 95.435 183.595 ;
        RECT 94.880 183.155 95.330 183.265 ;
        RECT 94.205 182.985 95.330 183.155 ;
        RECT 95.605 183.095 95.885 183.765 ;
        RECT 96.495 183.755 96.825 184.735 ;
        RECT 96.995 183.765 97.225 184.905 ;
        RECT 97.495 183.765 97.705 184.905 ;
        RECT 97.875 183.755 98.205 184.735 ;
        RECT 98.375 183.765 98.605 184.905 ;
        RECT 99.390 184.275 99.675 184.735 ;
        RECT 99.845 184.445 100.115 184.905 ;
        RECT 99.390 184.055 100.345 184.275 ;
        RECT 94.205 182.525 94.485 182.985 ;
        RECT 95.005 182.355 95.330 182.815 ;
        RECT 95.500 182.525 95.885 183.095 ;
        RECT 96.115 182.355 96.325 183.175 ;
        RECT 96.495 183.155 96.745 183.755 ;
        RECT 96.915 183.345 97.245 183.595 ;
        RECT 96.495 182.525 96.825 183.155 ;
        RECT 96.995 182.355 97.225 183.175 ;
        RECT 97.495 182.355 97.705 183.175 ;
        RECT 97.875 183.155 98.125 183.755 ;
        RECT 98.295 183.345 98.625 183.595 ;
        RECT 99.275 183.325 99.965 183.885 ;
        RECT 97.875 182.525 98.205 183.155 ;
        RECT 98.375 182.355 98.605 183.175 ;
        RECT 100.135 183.155 100.345 184.055 ;
        RECT 99.390 182.985 100.345 183.155 ;
        RECT 100.515 183.885 100.915 184.735 ;
        RECT 101.105 184.275 101.385 184.735 ;
        RECT 101.905 184.445 102.230 184.905 ;
        RECT 101.105 184.055 102.230 184.275 ;
        RECT 100.515 183.325 101.610 183.885 ;
        RECT 101.780 183.595 102.230 184.055 ;
        RECT 102.400 183.765 102.785 184.735 ;
        RECT 103.070 184.275 103.355 184.735 ;
        RECT 103.525 184.445 103.795 184.905 ;
        RECT 103.070 184.055 104.025 184.275 ;
        RECT 99.390 182.525 99.675 182.985 ;
        RECT 99.845 182.355 100.115 182.815 ;
        RECT 100.515 182.525 100.915 183.325 ;
        RECT 101.780 183.265 102.335 183.595 ;
        RECT 101.780 183.155 102.230 183.265 ;
        RECT 101.105 182.985 102.230 183.155 ;
        RECT 102.505 183.095 102.785 183.765 ;
        RECT 102.955 183.325 103.645 183.885 ;
        RECT 103.815 183.155 104.025 184.055 ;
        RECT 101.105 182.525 101.385 182.985 ;
        RECT 101.905 182.355 102.230 182.815 ;
        RECT 102.400 182.525 102.785 183.095 ;
        RECT 103.070 182.985 104.025 183.155 ;
        RECT 104.195 183.885 104.595 184.735 ;
        RECT 104.785 184.275 105.065 184.735 ;
        RECT 105.585 184.445 105.910 184.905 ;
        RECT 104.785 184.055 105.910 184.275 ;
        RECT 104.195 183.325 105.290 183.885 ;
        RECT 105.460 183.595 105.910 184.055 ;
        RECT 106.080 183.765 106.465 184.735 ;
        RECT 106.750 184.275 107.035 184.735 ;
        RECT 107.205 184.445 107.475 184.905 ;
        RECT 106.750 184.055 107.705 184.275 ;
        RECT 103.070 182.525 103.355 182.985 ;
        RECT 103.525 182.355 103.795 182.815 ;
        RECT 104.195 182.525 104.595 183.325 ;
        RECT 105.460 183.265 106.015 183.595 ;
        RECT 105.460 183.155 105.910 183.265 ;
        RECT 104.785 182.985 105.910 183.155 ;
        RECT 106.185 183.095 106.465 183.765 ;
        RECT 106.635 183.325 107.325 183.885 ;
        RECT 107.495 183.155 107.705 184.055 ;
        RECT 104.785 182.525 105.065 182.985 ;
        RECT 105.585 182.355 105.910 182.815 ;
        RECT 106.080 182.525 106.465 183.095 ;
        RECT 106.750 182.985 107.705 183.155 ;
        RECT 107.875 183.885 108.275 184.735 ;
        RECT 108.465 184.275 108.745 184.735 ;
        RECT 109.265 184.445 109.590 184.905 ;
        RECT 108.465 184.055 109.590 184.275 ;
        RECT 107.875 183.325 108.970 183.885 ;
        RECT 109.140 183.595 109.590 184.055 ;
        RECT 109.760 183.765 110.145 184.735 ;
        RECT 106.750 182.525 107.035 182.985 ;
        RECT 107.205 182.355 107.475 182.815 ;
        RECT 107.875 182.525 108.275 183.325 ;
        RECT 109.140 183.265 109.695 183.595 ;
        RECT 109.140 183.155 109.590 183.265 ;
        RECT 108.465 182.985 109.590 183.155 ;
        RECT 109.865 183.095 110.145 183.765 ;
        RECT 108.465 182.525 108.745 182.985 ;
        RECT 109.265 182.355 109.590 182.815 ;
        RECT 109.760 182.525 110.145 183.095 ;
        RECT 110.775 183.830 111.045 184.735 ;
        RECT 111.215 184.145 111.545 184.905 ;
        RECT 111.725 183.975 111.895 184.735 ;
        RECT 110.775 183.030 110.945 183.830 ;
        RECT 111.230 183.805 111.895 183.975 ;
        RECT 112.155 183.815 113.365 184.905 ;
        RECT 111.230 183.660 111.400 183.805 ;
        RECT 111.115 183.330 111.400 183.660 ;
        RECT 111.230 183.075 111.400 183.330 ;
        RECT 111.635 183.255 111.965 183.625 ;
        RECT 112.155 183.275 112.675 183.815 ;
        RECT 112.845 183.105 113.365 183.645 ;
        RECT 110.775 182.525 111.035 183.030 ;
        RECT 111.230 182.905 111.895 183.075 ;
        RECT 111.215 182.355 111.545 182.735 ;
        RECT 111.725 182.525 111.895 182.905 ;
        RECT 112.155 182.355 113.365 183.105 ;
        RECT 26.970 182.185 113.450 182.355 ;
        RECT 27.055 181.435 28.265 182.185 ;
        RECT 27.055 180.895 27.575 181.435 ;
        RECT 29.415 181.365 29.625 182.185 ;
        RECT 29.795 181.385 30.125 182.015 ;
        RECT 27.745 180.725 28.265 181.265 ;
        RECT 29.795 180.785 30.045 181.385 ;
        RECT 30.295 181.365 30.525 182.185 ;
        RECT 30.740 181.475 30.995 182.005 ;
        RECT 31.165 181.725 31.470 182.185 ;
        RECT 31.715 181.805 32.785 181.975 ;
        RECT 30.215 180.945 30.545 181.195 ;
        RECT 30.740 180.825 30.950 181.475 ;
        RECT 31.715 181.450 32.035 181.805 ;
        RECT 31.710 181.275 32.035 181.450 ;
        RECT 31.120 180.975 32.035 181.275 ;
        RECT 32.205 181.235 32.445 181.635 ;
        RECT 32.615 181.575 32.785 181.805 ;
        RECT 32.955 181.745 33.145 182.185 ;
        RECT 33.315 181.735 34.265 182.015 ;
        RECT 34.485 181.825 34.835 181.995 ;
        RECT 32.615 181.405 33.145 181.575 ;
        RECT 31.120 180.945 31.860 180.975 ;
        RECT 27.055 179.635 28.265 180.725 ;
        RECT 29.415 179.635 29.625 180.775 ;
        RECT 29.795 179.805 30.125 180.785 ;
        RECT 30.295 179.635 30.525 180.775 ;
        RECT 30.740 179.945 30.995 180.825 ;
        RECT 31.165 179.635 31.470 180.775 ;
        RECT 31.690 180.355 31.860 180.945 ;
        RECT 32.205 180.865 32.745 181.235 ;
        RECT 32.925 181.125 33.145 181.405 ;
        RECT 33.315 180.955 33.485 181.735 ;
        RECT 33.080 180.785 33.485 180.955 ;
        RECT 33.655 180.945 34.005 181.565 ;
        RECT 33.080 180.695 33.250 180.785 ;
        RECT 34.175 180.775 34.385 181.565 ;
        RECT 32.030 180.525 33.250 180.695 ;
        RECT 33.710 180.615 34.385 180.775 ;
        RECT 31.690 180.185 32.490 180.355 ;
        RECT 31.810 179.635 32.140 180.015 ;
        RECT 32.320 179.895 32.490 180.185 ;
        RECT 33.080 180.145 33.250 180.525 ;
        RECT 33.420 180.605 34.385 180.615 ;
        RECT 34.575 181.435 34.835 181.825 ;
        RECT 35.045 181.725 35.375 182.185 ;
        RECT 36.250 181.795 37.105 181.965 ;
        RECT 37.310 181.795 37.805 181.965 ;
        RECT 37.975 181.825 38.305 182.185 ;
        RECT 34.575 180.745 34.745 181.435 ;
        RECT 34.915 181.085 35.085 181.265 ;
        RECT 35.255 181.255 36.045 181.505 ;
        RECT 36.250 181.085 36.420 181.795 ;
        RECT 36.590 181.285 36.945 181.505 ;
        RECT 34.915 180.915 36.605 181.085 ;
        RECT 33.420 180.315 33.880 180.605 ;
        RECT 34.575 180.575 36.075 180.745 ;
        RECT 34.575 180.435 34.745 180.575 ;
        RECT 34.185 180.265 34.745 180.435 ;
        RECT 32.660 179.635 32.910 180.095 ;
        RECT 33.080 179.805 33.950 180.145 ;
        RECT 34.185 179.805 34.355 180.265 ;
        RECT 35.190 180.235 36.265 180.405 ;
        RECT 34.525 179.635 34.895 180.095 ;
        RECT 35.190 179.895 35.360 180.235 ;
        RECT 35.530 179.635 35.860 180.065 ;
        RECT 36.095 179.895 36.265 180.235 ;
        RECT 36.435 180.135 36.605 180.915 ;
        RECT 36.775 180.695 36.945 181.285 ;
        RECT 37.115 180.885 37.465 181.505 ;
        RECT 36.775 180.305 37.240 180.695 ;
        RECT 37.635 180.435 37.805 181.795 ;
        RECT 37.975 180.605 38.435 181.655 ;
        RECT 37.410 180.265 37.805 180.435 ;
        RECT 37.410 180.135 37.580 180.265 ;
        RECT 36.435 179.805 37.115 180.135 ;
        RECT 37.330 179.805 37.580 180.135 ;
        RECT 37.750 179.635 38.000 180.095 ;
        RECT 38.170 179.820 38.495 180.605 ;
        RECT 38.665 179.805 38.835 181.925 ;
        RECT 39.005 181.805 39.335 182.185 ;
        RECT 39.505 181.635 39.760 181.925 ;
        RECT 39.010 181.465 39.760 181.635 ;
        RECT 39.010 180.475 39.240 181.465 ;
        RECT 39.975 181.365 40.205 182.185 ;
        RECT 40.375 181.385 40.705 182.015 ;
        RECT 39.410 180.645 39.760 181.295 ;
        RECT 39.955 180.945 40.285 181.195 ;
        RECT 40.455 180.785 40.705 181.385 ;
        RECT 40.875 181.365 41.085 182.185 ;
        RECT 41.430 181.555 41.715 182.015 ;
        RECT 41.885 181.725 42.155 182.185 ;
        RECT 41.430 181.385 42.385 181.555 ;
        RECT 39.010 180.305 39.760 180.475 ;
        RECT 39.005 179.635 39.335 180.135 ;
        RECT 39.505 179.805 39.760 180.305 ;
        RECT 39.975 179.635 40.205 180.775 ;
        RECT 40.375 179.805 40.705 180.785 ;
        RECT 40.875 179.635 41.085 180.775 ;
        RECT 41.315 180.655 42.005 181.215 ;
        RECT 42.175 180.485 42.385 181.385 ;
        RECT 41.430 180.265 42.385 180.485 ;
        RECT 42.555 181.215 42.955 182.015 ;
        RECT 43.145 181.555 43.425 182.015 ;
        RECT 43.945 181.725 44.270 182.185 ;
        RECT 43.145 181.385 44.270 181.555 ;
        RECT 44.440 181.445 44.825 182.015 ;
        RECT 43.820 181.275 44.270 181.385 ;
        RECT 42.555 180.655 43.650 181.215 ;
        RECT 43.820 180.945 44.375 181.275 ;
        RECT 41.430 179.805 41.715 180.265 ;
        RECT 41.885 179.635 42.155 180.095 ;
        RECT 42.555 179.805 42.955 180.655 ;
        RECT 43.820 180.485 44.270 180.945 ;
        RECT 44.545 180.775 44.825 181.445 ;
        RECT 43.145 180.265 44.270 180.485 ;
        RECT 43.145 179.805 43.425 180.265 ;
        RECT 43.945 179.635 44.270 180.095 ;
        RECT 44.440 179.805 44.825 180.775 ;
        RECT 44.995 181.385 45.335 182.015 ;
        RECT 45.505 181.385 45.755 182.185 ;
        RECT 45.945 181.535 46.275 182.015 ;
        RECT 46.445 181.725 46.670 182.185 ;
        RECT 46.840 181.535 47.170 182.015 ;
        RECT 44.995 180.825 45.170 181.385 ;
        RECT 45.945 181.365 47.170 181.535 ;
        RECT 47.800 181.405 48.300 182.015 ;
        RECT 48.675 181.460 48.965 182.185 ;
        RECT 49.135 181.675 49.440 182.185 ;
        RECT 45.340 181.025 46.035 181.195 ;
        RECT 44.995 180.775 45.225 180.825 ;
        RECT 45.865 180.775 46.035 181.025 ;
        RECT 46.210 180.995 46.630 181.195 ;
        RECT 46.800 180.995 47.130 181.195 ;
        RECT 47.300 180.995 47.630 181.195 ;
        RECT 47.800 180.775 47.970 181.405 ;
        RECT 48.155 180.945 48.505 181.195 ;
        RECT 49.135 180.945 49.450 181.505 ;
        RECT 49.620 181.195 49.870 182.005 ;
        RECT 50.040 181.660 50.300 182.185 ;
        RECT 50.480 181.195 50.730 182.005 ;
        RECT 50.900 181.625 51.160 182.185 ;
        RECT 51.330 181.535 51.590 181.990 ;
        RECT 51.760 181.705 52.020 182.185 ;
        RECT 52.190 181.535 52.450 181.990 ;
        RECT 52.620 181.705 52.880 182.185 ;
        RECT 53.050 181.535 53.310 181.990 ;
        RECT 53.480 181.705 53.725 182.185 ;
        RECT 53.895 181.535 54.170 181.990 ;
        RECT 54.340 181.705 54.585 182.185 ;
        RECT 54.755 181.535 55.015 181.990 ;
        RECT 55.195 181.705 55.445 182.185 ;
        RECT 55.615 181.535 55.875 181.990 ;
        RECT 56.055 181.705 56.305 182.185 ;
        RECT 56.475 181.535 56.735 181.990 ;
        RECT 56.915 181.705 57.175 182.185 ;
        RECT 57.345 181.535 57.605 181.990 ;
        RECT 57.775 181.705 58.075 182.185 ;
        RECT 51.330 181.365 58.075 181.535 ;
        RECT 49.620 180.945 56.740 181.195 ;
        RECT 44.995 179.805 45.335 180.775 ;
        RECT 45.505 179.635 45.675 180.775 ;
        RECT 45.865 180.605 48.300 180.775 ;
        RECT 45.945 179.635 46.195 180.435 ;
        RECT 46.840 179.805 47.170 180.605 ;
        RECT 47.470 179.635 47.800 180.435 ;
        RECT 47.970 179.805 48.300 180.605 ;
        RECT 48.675 179.635 48.965 180.800 ;
        RECT 49.145 179.635 49.440 180.445 ;
        RECT 49.620 179.805 49.865 180.945 ;
        RECT 50.040 179.635 50.300 180.445 ;
        RECT 50.480 179.810 50.730 180.945 ;
        RECT 56.910 180.775 58.075 181.365 ;
        RECT 51.330 180.550 58.075 180.775 ;
        RECT 58.340 181.475 58.595 182.005 ;
        RECT 58.765 181.725 59.070 182.185 ;
        RECT 59.315 181.805 60.385 181.975 ;
        RECT 58.340 180.825 58.550 181.475 ;
        RECT 59.315 181.450 59.635 181.805 ;
        RECT 59.310 181.275 59.635 181.450 ;
        RECT 58.720 180.975 59.635 181.275 ;
        RECT 59.805 181.235 60.045 181.635 ;
        RECT 60.215 181.575 60.385 181.805 ;
        RECT 60.555 181.745 60.745 182.185 ;
        RECT 60.915 181.735 61.865 182.015 ;
        RECT 62.085 181.825 62.435 181.995 ;
        RECT 60.215 181.405 60.745 181.575 ;
        RECT 58.720 180.945 59.460 180.975 ;
        RECT 51.330 180.535 56.735 180.550 ;
        RECT 50.900 179.640 51.160 180.435 ;
        RECT 51.330 179.810 51.590 180.535 ;
        RECT 51.760 179.640 52.020 180.365 ;
        RECT 52.190 179.810 52.450 180.535 ;
        RECT 52.620 179.640 52.880 180.365 ;
        RECT 53.050 179.810 53.310 180.535 ;
        RECT 53.480 179.640 53.740 180.365 ;
        RECT 53.910 179.810 54.170 180.535 ;
        RECT 54.340 179.640 54.585 180.365 ;
        RECT 54.755 179.810 55.015 180.535 ;
        RECT 55.200 179.640 55.445 180.365 ;
        RECT 55.615 179.810 55.875 180.535 ;
        RECT 56.060 179.640 56.305 180.365 ;
        RECT 56.475 179.810 56.735 180.535 ;
        RECT 56.920 179.640 57.175 180.365 ;
        RECT 57.345 179.810 57.635 180.550 ;
        RECT 50.900 179.635 57.175 179.640 ;
        RECT 57.805 179.635 58.075 180.380 ;
        RECT 58.340 179.945 58.595 180.825 ;
        RECT 58.765 179.635 59.070 180.775 ;
        RECT 59.290 180.355 59.460 180.945 ;
        RECT 59.805 180.865 60.345 181.235 ;
        RECT 60.525 181.125 60.745 181.405 ;
        RECT 60.915 180.955 61.085 181.735 ;
        RECT 60.680 180.785 61.085 180.955 ;
        RECT 61.255 180.945 61.605 181.565 ;
        RECT 60.680 180.695 60.850 180.785 ;
        RECT 61.775 180.775 61.985 181.565 ;
        RECT 59.630 180.525 60.850 180.695 ;
        RECT 61.310 180.615 61.985 180.775 ;
        RECT 59.290 180.185 60.090 180.355 ;
        RECT 59.410 179.635 59.740 180.015 ;
        RECT 59.920 179.895 60.090 180.185 ;
        RECT 60.680 180.145 60.850 180.525 ;
        RECT 61.020 180.605 61.985 180.615 ;
        RECT 62.175 181.435 62.435 181.825 ;
        RECT 62.645 181.725 62.975 182.185 ;
        RECT 63.850 181.795 64.705 181.965 ;
        RECT 64.910 181.795 65.405 181.965 ;
        RECT 65.575 181.825 65.905 182.185 ;
        RECT 62.175 180.745 62.345 181.435 ;
        RECT 62.515 181.085 62.685 181.265 ;
        RECT 62.855 181.255 63.645 181.505 ;
        RECT 63.850 181.085 64.020 181.795 ;
        RECT 64.190 181.285 64.545 181.505 ;
        RECT 62.515 180.915 64.205 181.085 ;
        RECT 61.020 180.315 61.480 180.605 ;
        RECT 62.175 180.575 63.675 180.745 ;
        RECT 62.175 180.435 62.345 180.575 ;
        RECT 61.785 180.265 62.345 180.435 ;
        RECT 60.260 179.635 60.510 180.095 ;
        RECT 60.680 179.805 61.550 180.145 ;
        RECT 61.785 179.805 61.955 180.265 ;
        RECT 62.790 180.235 63.865 180.405 ;
        RECT 62.125 179.635 62.495 180.095 ;
        RECT 62.790 179.895 62.960 180.235 ;
        RECT 63.130 179.635 63.460 180.065 ;
        RECT 63.695 179.895 63.865 180.235 ;
        RECT 64.035 180.135 64.205 180.915 ;
        RECT 64.375 180.695 64.545 181.285 ;
        RECT 64.715 180.885 65.065 181.505 ;
        RECT 64.375 180.305 64.840 180.695 ;
        RECT 65.235 180.435 65.405 181.795 ;
        RECT 65.575 180.605 66.035 181.655 ;
        RECT 65.010 180.265 65.405 180.435 ;
        RECT 65.010 180.135 65.180 180.265 ;
        RECT 64.035 179.805 64.715 180.135 ;
        RECT 64.930 179.805 65.180 180.135 ;
        RECT 65.350 179.635 65.600 180.095 ;
        RECT 65.770 179.820 66.095 180.605 ;
        RECT 66.265 179.805 66.435 181.925 ;
        RECT 66.605 181.805 66.935 182.185 ;
        RECT 67.105 181.635 67.360 181.925 ;
        RECT 66.610 181.465 67.360 181.635 ;
        RECT 68.005 181.655 68.335 182.015 ;
        RECT 68.505 181.825 68.835 182.185 ;
        RECT 69.035 181.655 69.365 182.015 ;
        RECT 66.610 180.475 66.840 181.465 ;
        RECT 68.005 181.445 69.365 181.655 ;
        RECT 69.875 181.425 70.585 182.015 ;
        RECT 71.025 181.790 71.355 182.185 ;
        RECT 71.525 181.615 71.725 181.970 ;
        RECT 71.895 181.785 72.225 182.185 ;
        RECT 72.395 181.615 72.595 181.960 ;
        RECT 67.010 180.645 67.360 181.295 ;
        RECT 67.995 180.945 68.305 181.275 ;
        RECT 68.515 180.945 68.890 181.275 ;
        RECT 69.210 180.945 69.705 181.275 ;
        RECT 66.610 180.305 67.360 180.475 ;
        RECT 66.605 179.635 66.935 180.135 ;
        RECT 67.105 179.805 67.360 180.305 ;
        RECT 68.005 179.635 68.335 180.695 ;
        RECT 68.515 180.020 68.685 180.945 ;
        RECT 68.855 180.455 69.185 180.675 ;
        RECT 69.380 180.655 69.705 180.945 ;
        RECT 69.880 180.655 70.210 181.195 ;
        RECT 70.380 180.455 70.585 181.425 ;
        RECT 68.855 180.225 70.585 180.455 ;
        RECT 68.855 179.825 69.185 180.225 ;
        RECT 69.355 179.635 69.685 179.995 ;
        RECT 69.885 179.805 70.585 180.225 ;
        RECT 70.755 181.445 72.595 181.615 ;
        RECT 72.765 181.445 73.095 182.185 ;
        RECT 73.330 181.615 73.500 181.865 ;
        RECT 73.330 181.445 73.805 181.615 ;
        RECT 74.435 181.460 74.725 182.185 ;
        RECT 74.985 181.635 75.155 182.015 ;
        RECT 75.370 181.805 75.700 182.185 ;
        RECT 74.985 181.465 75.700 181.635 ;
        RECT 70.755 179.820 71.015 181.445 ;
        RECT 71.195 180.475 71.415 181.275 ;
        RECT 71.655 180.655 71.955 181.275 ;
        RECT 72.125 180.655 72.455 181.275 ;
        RECT 72.625 180.655 72.945 181.275 ;
        RECT 73.115 180.655 73.465 181.275 ;
        RECT 73.635 180.475 73.805 181.445 ;
        RECT 74.895 180.915 75.250 181.285 ;
        RECT 75.530 181.275 75.700 181.465 ;
        RECT 75.870 181.440 76.125 182.015 ;
        RECT 75.530 180.945 75.785 181.275 ;
        RECT 71.195 180.265 73.805 180.475 ;
        RECT 72.765 179.635 73.095 180.085 ;
        RECT 74.435 179.635 74.725 180.800 ;
        RECT 75.530 180.735 75.700 180.945 ;
        RECT 74.985 180.565 75.700 180.735 ;
        RECT 75.955 180.710 76.125 181.440 ;
        RECT 76.300 181.345 76.560 182.185 ;
        RECT 77.470 181.375 77.715 181.980 ;
        RECT 77.935 181.650 78.445 182.185 ;
        RECT 77.195 181.205 78.425 181.375 ;
        RECT 74.985 179.805 75.155 180.565 ;
        RECT 75.370 179.635 75.700 180.395 ;
        RECT 75.870 179.805 76.125 180.710 ;
        RECT 76.300 179.635 76.560 180.785 ;
        RECT 77.195 180.395 77.535 181.205 ;
        RECT 77.705 180.640 78.455 180.830 ;
        RECT 77.195 179.985 77.710 180.395 ;
        RECT 77.945 179.635 78.115 180.395 ;
        RECT 78.285 179.975 78.455 180.640 ;
        RECT 78.625 180.655 78.815 182.015 ;
        RECT 78.985 181.165 79.260 182.015 ;
        RECT 79.450 181.650 79.980 182.015 ;
        RECT 80.405 181.785 80.735 182.185 ;
        RECT 79.805 181.615 79.980 181.650 ;
        RECT 78.985 180.995 79.265 181.165 ;
        RECT 78.985 180.855 79.260 180.995 ;
        RECT 79.465 180.655 79.635 181.455 ;
        RECT 78.625 180.485 79.635 180.655 ;
        RECT 79.805 181.445 80.735 181.615 ;
        RECT 80.905 181.445 81.160 182.015 ;
        RECT 79.805 180.315 79.975 181.445 ;
        RECT 80.565 181.275 80.735 181.445 ;
        RECT 78.850 180.145 79.975 180.315 ;
        RECT 80.145 180.945 80.340 181.275 ;
        RECT 80.565 180.945 80.820 181.275 ;
        RECT 80.145 179.975 80.315 180.945 ;
        RECT 80.990 180.775 81.160 181.445 ;
        RECT 78.285 179.805 80.315 179.975 ;
        RECT 80.485 179.635 80.655 180.775 ;
        RECT 80.825 179.805 81.160 180.775 ;
        RECT 81.335 181.385 81.675 182.015 ;
        RECT 81.845 181.385 82.095 182.185 ;
        RECT 82.285 181.535 82.615 182.015 ;
        RECT 82.785 181.725 83.010 182.185 ;
        RECT 83.180 181.535 83.510 182.015 ;
        RECT 81.335 180.825 81.510 181.385 ;
        RECT 82.285 181.365 83.510 181.535 ;
        RECT 84.140 181.405 84.640 182.015 ;
        RECT 85.020 181.635 85.275 181.925 ;
        RECT 85.445 181.805 85.775 182.185 ;
        RECT 85.020 181.465 85.770 181.635 ;
        RECT 81.680 181.025 82.375 181.195 ;
        RECT 81.335 180.775 81.565 180.825 ;
        RECT 82.205 180.775 82.375 181.025 ;
        RECT 82.550 180.995 82.970 181.195 ;
        RECT 83.140 180.995 83.470 181.195 ;
        RECT 83.640 180.995 83.970 181.195 ;
        RECT 84.140 180.775 84.310 181.405 ;
        RECT 84.495 180.945 84.845 181.195 ;
        RECT 81.335 179.805 81.675 180.775 ;
        RECT 81.845 179.635 82.015 180.775 ;
        RECT 82.205 180.605 84.640 180.775 ;
        RECT 85.020 180.645 85.370 181.295 ;
        RECT 82.285 179.635 82.535 180.435 ;
        RECT 83.180 179.805 83.510 180.605 ;
        RECT 83.810 179.635 84.140 180.435 ;
        RECT 84.310 179.805 84.640 180.605 ;
        RECT 85.540 180.475 85.770 181.465 ;
        RECT 85.020 180.305 85.770 180.475 ;
        RECT 85.020 179.805 85.275 180.305 ;
        RECT 85.445 179.635 85.775 180.135 ;
        RECT 85.945 179.805 86.115 181.925 ;
        RECT 86.475 181.825 86.805 182.185 ;
        RECT 86.975 181.795 87.470 181.965 ;
        RECT 87.675 181.795 88.530 181.965 ;
        RECT 86.345 180.605 86.805 181.655 ;
        RECT 86.285 179.820 86.610 180.605 ;
        RECT 86.975 180.435 87.145 181.795 ;
        RECT 87.315 180.885 87.665 181.505 ;
        RECT 87.835 181.285 88.190 181.505 ;
        RECT 87.835 180.695 88.005 181.285 ;
        RECT 88.360 181.085 88.530 181.795 ;
        RECT 89.405 181.725 89.735 182.185 ;
        RECT 89.945 181.825 90.295 181.995 ;
        RECT 88.735 181.255 89.525 181.505 ;
        RECT 89.945 181.435 90.205 181.825 ;
        RECT 90.515 181.735 91.465 182.015 ;
        RECT 91.635 181.745 91.825 182.185 ;
        RECT 91.995 181.805 93.065 181.975 ;
        RECT 89.695 181.085 89.865 181.265 ;
        RECT 86.975 180.265 87.370 180.435 ;
        RECT 87.540 180.305 88.005 180.695 ;
        RECT 88.175 180.915 89.865 181.085 ;
        RECT 87.200 180.135 87.370 180.265 ;
        RECT 88.175 180.135 88.345 180.915 ;
        RECT 90.035 180.745 90.205 181.435 ;
        RECT 88.705 180.575 90.205 180.745 ;
        RECT 90.395 180.775 90.605 181.565 ;
        RECT 90.775 180.945 91.125 181.565 ;
        RECT 91.295 180.955 91.465 181.735 ;
        RECT 91.995 181.575 92.165 181.805 ;
        RECT 91.635 181.405 92.165 181.575 ;
        RECT 91.635 181.125 91.855 181.405 ;
        RECT 92.335 181.235 92.575 181.635 ;
        RECT 91.295 180.785 91.700 180.955 ;
        RECT 92.035 180.865 92.575 181.235 ;
        RECT 92.745 181.450 93.065 181.805 ;
        RECT 93.310 181.725 93.615 182.185 ;
        RECT 93.785 181.475 94.040 182.005 ;
        RECT 92.745 181.275 93.070 181.450 ;
        RECT 92.745 180.975 93.660 181.275 ;
        RECT 92.920 180.945 93.660 180.975 ;
        RECT 90.395 180.615 91.070 180.775 ;
        RECT 91.530 180.695 91.700 180.785 ;
        RECT 90.395 180.605 91.360 180.615 ;
        RECT 90.035 180.435 90.205 180.575 ;
        RECT 86.780 179.635 87.030 180.095 ;
        RECT 87.200 179.805 87.450 180.135 ;
        RECT 87.665 179.805 88.345 180.135 ;
        RECT 88.515 180.235 89.590 180.405 ;
        RECT 90.035 180.265 90.595 180.435 ;
        RECT 90.900 180.315 91.360 180.605 ;
        RECT 91.530 180.525 92.750 180.695 ;
        RECT 88.515 179.895 88.685 180.235 ;
        RECT 88.920 179.635 89.250 180.065 ;
        RECT 89.420 179.895 89.590 180.235 ;
        RECT 89.885 179.635 90.255 180.095 ;
        RECT 90.425 179.805 90.595 180.265 ;
        RECT 91.530 180.145 91.700 180.525 ;
        RECT 92.920 180.355 93.090 180.945 ;
        RECT 93.830 180.825 94.040 181.475 ;
        RECT 94.220 181.345 94.480 182.185 ;
        RECT 94.655 181.440 94.910 182.015 ;
        RECT 95.080 181.805 95.410 182.185 ;
        RECT 95.625 181.635 95.795 182.015 ;
        RECT 95.080 181.465 95.795 181.635 ;
        RECT 90.830 179.805 91.700 180.145 ;
        RECT 92.290 180.185 93.090 180.355 ;
        RECT 91.870 179.635 92.120 180.095 ;
        RECT 92.290 179.895 92.460 180.185 ;
        RECT 92.640 179.635 92.970 180.015 ;
        RECT 93.310 179.635 93.615 180.775 ;
        RECT 93.785 179.945 94.040 180.825 ;
        RECT 94.220 179.635 94.480 180.785 ;
        RECT 94.655 180.710 94.825 181.440 ;
        RECT 95.080 181.275 95.250 181.465 ;
        RECT 96.060 181.445 96.315 182.015 ;
        RECT 96.485 181.785 96.815 182.185 ;
        RECT 97.240 181.650 97.770 182.015 ;
        RECT 97.240 181.615 97.415 181.650 ;
        RECT 96.485 181.445 97.415 181.615 ;
        RECT 94.995 180.945 95.250 181.275 ;
        RECT 95.080 180.735 95.250 180.945 ;
        RECT 95.530 180.915 95.885 181.285 ;
        RECT 96.060 180.775 96.230 181.445 ;
        RECT 96.485 181.275 96.655 181.445 ;
        RECT 96.400 180.945 96.655 181.275 ;
        RECT 96.880 180.945 97.075 181.275 ;
        RECT 94.655 179.805 94.910 180.710 ;
        RECT 95.080 180.565 95.795 180.735 ;
        RECT 95.080 179.635 95.410 180.395 ;
        RECT 95.625 179.805 95.795 180.565 ;
        RECT 96.060 179.805 96.395 180.775 ;
        RECT 96.565 179.635 96.735 180.775 ;
        RECT 96.905 179.975 97.075 180.945 ;
        RECT 97.245 180.315 97.415 181.445 ;
        RECT 97.585 180.655 97.755 181.455 ;
        RECT 97.960 181.165 98.235 182.015 ;
        RECT 97.955 180.995 98.235 181.165 ;
        RECT 97.960 180.855 98.235 180.995 ;
        RECT 98.405 180.655 98.595 182.015 ;
        RECT 98.775 181.650 99.285 182.185 ;
        RECT 99.505 181.375 99.750 181.980 ;
        RECT 100.195 181.460 100.485 182.185 ;
        RECT 100.660 181.785 100.995 182.185 ;
        RECT 101.165 181.615 101.370 182.015 ;
        RECT 101.580 181.705 101.855 182.185 ;
        RECT 102.065 181.685 102.325 182.015 ;
        RECT 100.685 181.445 101.370 181.615 ;
        RECT 98.795 181.205 100.025 181.375 ;
        RECT 97.585 180.485 98.595 180.655 ;
        RECT 98.765 180.640 99.515 180.830 ;
        RECT 97.245 180.145 98.370 180.315 ;
        RECT 98.765 179.975 98.935 180.640 ;
        RECT 99.685 180.395 100.025 181.205 ;
        RECT 96.905 179.805 98.935 179.975 ;
        RECT 99.105 179.635 99.275 180.395 ;
        RECT 99.510 179.985 100.025 180.395 ;
        RECT 100.195 179.635 100.485 180.800 ;
        RECT 100.685 180.415 101.025 181.445 ;
        RECT 101.195 180.775 101.445 181.275 ;
        RECT 101.625 180.945 101.985 181.525 ;
        RECT 102.155 180.775 102.325 181.685 ;
        RECT 102.500 181.635 102.755 181.925 ;
        RECT 102.925 181.805 103.255 182.185 ;
        RECT 102.500 181.465 103.250 181.635 ;
        RECT 101.195 180.605 102.325 180.775 ;
        RECT 102.500 180.645 102.850 181.295 ;
        RECT 100.685 180.240 101.350 180.415 ;
        RECT 100.660 179.635 100.995 180.060 ;
        RECT 101.165 179.835 101.350 180.240 ;
        RECT 101.555 179.635 101.885 180.415 ;
        RECT 102.055 179.835 102.325 180.605 ;
        RECT 103.020 180.475 103.250 181.465 ;
        RECT 102.500 180.305 103.250 180.475 ;
        RECT 102.500 179.805 102.755 180.305 ;
        RECT 102.925 179.635 103.255 180.135 ;
        RECT 103.425 179.805 103.595 181.925 ;
        RECT 103.955 181.825 104.285 182.185 ;
        RECT 104.455 181.795 104.950 181.965 ;
        RECT 105.155 181.795 106.010 181.965 ;
        RECT 103.825 180.605 104.285 181.655 ;
        RECT 103.765 179.820 104.090 180.605 ;
        RECT 104.455 180.435 104.625 181.795 ;
        RECT 104.795 180.885 105.145 181.505 ;
        RECT 105.315 181.285 105.670 181.505 ;
        RECT 105.315 180.695 105.485 181.285 ;
        RECT 105.840 181.085 106.010 181.795 ;
        RECT 106.885 181.725 107.215 182.185 ;
        RECT 107.425 181.825 107.775 181.995 ;
        RECT 106.215 181.255 107.005 181.505 ;
        RECT 107.425 181.435 107.685 181.825 ;
        RECT 107.995 181.735 108.945 182.015 ;
        RECT 109.115 181.745 109.305 182.185 ;
        RECT 109.475 181.805 110.545 181.975 ;
        RECT 107.175 181.085 107.345 181.265 ;
        RECT 104.455 180.265 104.850 180.435 ;
        RECT 105.020 180.305 105.485 180.695 ;
        RECT 105.655 180.915 107.345 181.085 ;
        RECT 104.680 180.135 104.850 180.265 ;
        RECT 105.655 180.135 105.825 180.915 ;
        RECT 107.515 180.745 107.685 181.435 ;
        RECT 106.185 180.575 107.685 180.745 ;
        RECT 107.875 180.775 108.085 181.565 ;
        RECT 108.255 180.945 108.605 181.565 ;
        RECT 108.775 180.955 108.945 181.735 ;
        RECT 109.475 181.575 109.645 181.805 ;
        RECT 109.115 181.405 109.645 181.575 ;
        RECT 109.115 181.125 109.335 181.405 ;
        RECT 109.815 181.235 110.055 181.635 ;
        RECT 108.775 180.785 109.180 180.955 ;
        RECT 109.515 180.865 110.055 181.235 ;
        RECT 110.225 181.450 110.545 181.805 ;
        RECT 110.790 181.725 111.095 182.185 ;
        RECT 111.265 181.475 111.520 182.005 ;
        RECT 110.225 181.275 110.550 181.450 ;
        RECT 110.225 180.975 111.140 181.275 ;
        RECT 110.400 180.945 111.140 180.975 ;
        RECT 107.875 180.615 108.550 180.775 ;
        RECT 109.010 180.695 109.180 180.785 ;
        RECT 107.875 180.605 108.840 180.615 ;
        RECT 107.515 180.435 107.685 180.575 ;
        RECT 104.260 179.635 104.510 180.095 ;
        RECT 104.680 179.805 104.930 180.135 ;
        RECT 105.145 179.805 105.825 180.135 ;
        RECT 105.995 180.235 107.070 180.405 ;
        RECT 107.515 180.265 108.075 180.435 ;
        RECT 108.380 180.315 108.840 180.605 ;
        RECT 109.010 180.525 110.230 180.695 ;
        RECT 105.995 179.895 106.165 180.235 ;
        RECT 106.400 179.635 106.730 180.065 ;
        RECT 106.900 179.895 107.070 180.235 ;
        RECT 107.365 179.635 107.735 180.095 ;
        RECT 107.905 179.805 108.075 180.265 ;
        RECT 109.010 180.145 109.180 180.525 ;
        RECT 110.400 180.355 110.570 180.945 ;
        RECT 111.310 180.825 111.520 181.475 ;
        RECT 112.155 181.435 113.365 182.185 ;
        RECT 108.310 179.805 109.180 180.145 ;
        RECT 109.770 180.185 110.570 180.355 ;
        RECT 109.350 179.635 109.600 180.095 ;
        RECT 109.770 179.895 109.940 180.185 ;
        RECT 110.120 179.635 110.450 180.015 ;
        RECT 110.790 179.635 111.095 180.775 ;
        RECT 111.265 179.945 111.520 180.825 ;
        RECT 112.155 180.725 112.675 181.265 ;
        RECT 112.845 180.895 113.365 181.435 ;
        RECT 112.155 179.635 113.365 180.725 ;
        RECT 26.970 179.465 113.450 179.635 ;
        RECT 27.055 178.375 28.265 179.465 ;
        RECT 27.055 177.665 27.575 178.205 ;
        RECT 27.745 177.835 28.265 178.375 ;
        RECT 28.985 178.535 29.155 179.295 ;
        RECT 29.335 178.705 29.665 179.465 ;
        RECT 28.985 178.365 29.650 178.535 ;
        RECT 29.835 178.390 30.105 179.295 ;
        RECT 29.480 178.220 29.650 178.365 ;
        RECT 28.915 177.815 29.245 178.185 ;
        RECT 29.480 177.890 29.765 178.220 ;
        RECT 27.055 176.915 28.265 177.665 ;
        RECT 29.480 177.635 29.650 177.890 ;
        RECT 28.985 177.465 29.650 177.635 ;
        RECT 29.935 177.590 30.105 178.390 ;
        RECT 30.315 178.325 30.545 179.465 ;
        RECT 30.715 178.315 31.045 179.295 ;
        RECT 31.215 178.325 31.425 179.465 ;
        RECT 31.660 178.325 31.995 179.295 ;
        RECT 32.165 178.325 32.335 179.465 ;
        RECT 32.505 179.125 34.535 179.295 ;
        RECT 30.295 177.905 30.625 178.155 ;
        RECT 28.985 177.085 29.155 177.465 ;
        RECT 29.335 176.915 29.665 177.295 ;
        RECT 29.845 177.085 30.105 177.590 ;
        RECT 30.315 176.915 30.545 177.735 ;
        RECT 30.795 177.715 31.045 178.315 ;
        RECT 30.715 177.085 31.045 177.715 ;
        RECT 31.215 176.915 31.425 177.735 ;
        RECT 31.660 177.655 31.830 178.325 ;
        RECT 32.505 178.155 32.675 179.125 ;
        RECT 32.000 177.825 32.255 178.155 ;
        RECT 32.480 177.825 32.675 178.155 ;
        RECT 32.845 178.785 33.970 178.955 ;
        RECT 32.085 177.655 32.255 177.825 ;
        RECT 32.845 177.655 33.015 178.785 ;
        RECT 31.660 177.085 31.915 177.655 ;
        RECT 32.085 177.485 33.015 177.655 ;
        RECT 33.185 178.445 34.195 178.615 ;
        RECT 33.185 177.645 33.355 178.445 ;
        RECT 32.840 177.450 33.015 177.485 ;
        RECT 32.085 176.915 32.415 177.315 ;
        RECT 32.840 177.085 33.370 177.450 ;
        RECT 33.560 177.425 33.835 178.245 ;
        RECT 33.555 177.255 33.835 177.425 ;
        RECT 33.560 177.085 33.835 177.255 ;
        RECT 34.005 177.085 34.195 178.445 ;
        RECT 34.365 178.460 34.535 179.125 ;
        RECT 34.705 178.705 34.875 179.465 ;
        RECT 35.110 178.705 35.625 179.115 ;
        RECT 34.365 178.270 35.115 178.460 ;
        RECT 35.285 177.895 35.625 178.705 ;
        RECT 35.795 178.300 36.085 179.465 ;
        RECT 36.805 178.535 36.975 179.295 ;
        RECT 37.155 178.705 37.485 179.465 ;
        RECT 36.805 178.365 37.470 178.535 ;
        RECT 37.655 178.390 37.925 179.295 ;
        RECT 37.300 178.220 37.470 178.365 ;
        RECT 34.395 177.725 35.625 177.895 ;
        RECT 36.735 177.815 37.065 178.185 ;
        RECT 37.300 177.890 37.585 178.220 ;
        RECT 34.375 176.915 34.885 177.450 ;
        RECT 35.105 177.120 35.350 177.725 ;
        RECT 35.795 176.915 36.085 177.640 ;
        RECT 37.300 177.635 37.470 177.890 ;
        RECT 36.805 177.465 37.470 177.635 ;
        RECT 37.755 177.590 37.925 178.390 ;
        RECT 38.135 178.325 38.365 179.465 ;
        RECT 38.535 178.315 38.865 179.295 ;
        RECT 39.035 178.325 39.245 179.465 ;
        RECT 39.680 178.495 40.010 179.295 ;
        RECT 40.180 178.665 40.510 179.465 ;
        RECT 40.810 178.495 41.140 179.295 ;
        RECT 41.785 178.665 42.035 179.465 ;
        RECT 39.680 178.325 42.115 178.495 ;
        RECT 42.305 178.325 42.475 179.465 ;
        RECT 42.645 178.325 42.985 179.295 ;
        RECT 43.360 178.495 43.690 179.295 ;
        RECT 43.860 178.665 44.190 179.465 ;
        RECT 44.490 178.495 44.820 179.295 ;
        RECT 45.465 178.665 45.715 179.465 ;
        RECT 43.360 178.325 45.795 178.495 ;
        RECT 45.985 178.325 46.155 179.465 ;
        RECT 46.325 178.325 46.665 179.295 ;
        RECT 38.115 177.905 38.445 178.155 ;
        RECT 36.805 177.085 36.975 177.465 ;
        RECT 37.155 176.915 37.485 177.295 ;
        RECT 37.665 177.085 37.925 177.590 ;
        RECT 38.135 176.915 38.365 177.735 ;
        RECT 38.615 177.715 38.865 178.315 ;
        RECT 39.475 177.905 39.825 178.155 ;
        RECT 38.535 177.085 38.865 177.715 ;
        RECT 39.035 176.915 39.245 177.735 ;
        RECT 40.010 177.695 40.180 178.325 ;
        RECT 40.350 177.905 40.680 178.105 ;
        RECT 40.850 177.905 41.180 178.105 ;
        RECT 41.350 177.905 41.770 178.105 ;
        RECT 41.945 178.075 42.115 178.325 ;
        RECT 41.945 177.905 42.640 178.075 ;
        RECT 39.680 177.085 40.180 177.695 ;
        RECT 40.810 177.565 42.035 177.735 ;
        RECT 42.810 177.715 42.985 178.325 ;
        RECT 43.155 177.905 43.505 178.155 ;
        RECT 40.810 177.085 41.140 177.565 ;
        RECT 41.310 176.915 41.535 177.375 ;
        RECT 41.705 177.085 42.035 177.565 ;
        RECT 42.225 176.915 42.475 177.715 ;
        RECT 42.645 177.085 42.985 177.715 ;
        RECT 43.690 177.695 43.860 178.325 ;
        RECT 44.030 177.905 44.360 178.105 ;
        RECT 44.530 177.905 44.860 178.105 ;
        RECT 45.030 177.905 45.450 178.105 ;
        RECT 45.625 178.075 45.795 178.325 ;
        RECT 45.625 177.905 46.320 178.075 ;
        RECT 43.360 177.085 43.860 177.695 ;
        RECT 44.490 177.565 45.715 177.735 ;
        RECT 46.490 177.715 46.665 178.325 ;
        RECT 44.490 177.085 44.820 177.565 ;
        RECT 44.990 176.915 45.215 177.375 ;
        RECT 45.385 177.085 45.715 177.565 ;
        RECT 45.905 176.915 46.155 177.715 ;
        RECT 46.325 177.085 46.665 177.715 ;
        RECT 46.835 178.325 47.220 179.295 ;
        RECT 47.390 179.005 47.715 179.465 ;
        RECT 48.235 178.835 48.515 179.295 ;
        RECT 47.390 178.615 48.515 178.835 ;
        RECT 46.835 177.655 47.115 178.325 ;
        RECT 47.390 178.155 47.840 178.615 ;
        RECT 48.705 178.445 49.105 179.295 ;
        RECT 49.505 179.005 49.775 179.465 ;
        RECT 49.945 178.835 50.230 179.295 ;
        RECT 47.285 177.825 47.840 178.155 ;
        RECT 48.010 177.885 49.105 178.445 ;
        RECT 47.390 177.715 47.840 177.825 ;
        RECT 46.835 177.085 47.220 177.655 ;
        RECT 47.390 177.545 48.515 177.715 ;
        RECT 47.390 176.915 47.715 177.375 ;
        RECT 48.235 177.085 48.515 177.545 ;
        RECT 48.705 177.085 49.105 177.885 ;
        RECT 49.275 178.615 50.230 178.835 ;
        RECT 49.275 177.715 49.485 178.615 ;
        RECT 49.655 177.885 50.345 178.445 ;
        RECT 51.440 178.315 51.700 179.465 ;
        RECT 51.875 178.390 52.130 179.295 ;
        RECT 52.300 178.705 52.630 179.465 ;
        RECT 52.845 178.535 53.015 179.295 ;
        RECT 53.330 178.665 53.630 179.465 ;
        RECT 49.275 177.545 50.230 177.715 ;
        RECT 49.505 176.915 49.775 177.375 ;
        RECT 49.945 177.085 50.230 177.545 ;
        RECT 51.440 176.915 51.700 177.755 ;
        RECT 51.875 177.660 52.045 178.390 ;
        RECT 52.300 178.365 53.015 178.535 ;
        RECT 53.800 178.495 54.130 179.295 ;
        RECT 54.300 178.665 54.470 179.465 ;
        RECT 54.640 178.495 54.970 179.295 ;
        RECT 55.140 178.665 55.310 179.465 ;
        RECT 55.480 178.495 55.810 179.295 ;
        RECT 55.980 178.665 56.150 179.465 ;
        RECT 56.320 178.495 56.650 179.295 ;
        RECT 56.820 178.665 57.075 179.465 ;
        RECT 52.300 178.155 52.470 178.365 ;
        RECT 53.275 178.325 57.245 178.495 ;
        RECT 52.215 177.825 52.470 178.155 ;
        RECT 51.875 177.085 52.130 177.660 ;
        RECT 52.300 177.635 52.470 177.825 ;
        RECT 52.750 177.815 53.105 178.185 ;
        RECT 53.275 177.735 53.595 178.325 ;
        RECT 53.795 177.905 56.650 178.155 ;
        RECT 56.900 177.735 57.245 178.325 ;
        RECT 52.300 177.465 53.015 177.635 ;
        RECT 53.275 177.545 57.245 177.735 ;
        RECT 57.875 178.325 58.215 179.295 ;
        RECT 58.385 178.325 58.555 179.465 ;
        RECT 58.825 178.665 59.075 179.465 ;
        RECT 59.720 178.495 60.050 179.295 ;
        RECT 60.350 178.665 60.680 179.465 ;
        RECT 60.850 178.495 61.180 179.295 ;
        RECT 58.745 178.325 61.180 178.495 ;
        RECT 57.875 177.715 58.050 178.325 ;
        RECT 58.745 178.075 58.915 178.325 ;
        RECT 58.220 177.905 58.915 178.075 ;
        RECT 59.090 177.905 59.510 178.105 ;
        RECT 59.680 177.905 60.010 178.105 ;
        RECT 60.180 177.905 60.510 178.105 ;
        RECT 52.300 176.915 52.630 177.295 ;
        RECT 52.845 177.085 53.015 177.465 ;
        RECT 53.325 176.915 53.630 177.375 ;
        RECT 53.800 177.085 54.130 177.545 ;
        RECT 54.300 176.915 54.470 177.375 ;
        RECT 54.640 177.085 54.970 177.545 ;
        RECT 55.140 176.915 55.310 177.375 ;
        RECT 55.480 177.085 55.810 177.545 ;
        RECT 55.980 176.915 56.150 177.375 ;
        RECT 56.320 177.085 56.650 177.545 ;
        RECT 56.820 176.915 57.075 177.375 ;
        RECT 57.875 177.085 58.215 177.715 ;
        RECT 58.385 176.915 58.635 177.715 ;
        RECT 58.825 177.565 60.050 177.735 ;
        RECT 58.825 177.085 59.155 177.565 ;
        RECT 59.325 176.915 59.550 177.375 ;
        RECT 59.720 177.085 60.050 177.565 ;
        RECT 60.680 177.695 60.850 178.325 ;
        RECT 61.555 178.300 61.845 179.465 ;
        RECT 62.015 178.325 62.355 179.295 ;
        RECT 62.525 178.325 62.695 179.465 ;
        RECT 62.965 178.665 63.215 179.465 ;
        RECT 63.860 178.495 64.190 179.295 ;
        RECT 64.490 178.665 64.820 179.465 ;
        RECT 64.990 178.495 65.320 179.295 ;
        RECT 62.885 178.325 65.320 178.495 ;
        RECT 65.695 178.325 66.035 179.295 ;
        RECT 66.205 178.325 66.375 179.465 ;
        RECT 66.645 178.665 66.895 179.465 ;
        RECT 67.540 178.495 67.870 179.295 ;
        RECT 68.170 178.665 68.500 179.465 ;
        RECT 68.670 178.495 69.000 179.295 ;
        RECT 66.565 178.325 69.000 178.495 ;
        RECT 61.035 177.905 61.385 178.155 ;
        RECT 62.015 177.715 62.190 178.325 ;
        RECT 62.885 178.075 63.055 178.325 ;
        RECT 62.360 177.905 63.055 178.075 ;
        RECT 63.230 177.905 63.650 178.105 ;
        RECT 63.820 177.905 64.150 178.105 ;
        RECT 64.320 177.905 64.650 178.105 ;
        RECT 60.680 177.085 61.180 177.695 ;
        RECT 61.555 176.915 61.845 177.640 ;
        RECT 62.015 177.085 62.355 177.715 ;
        RECT 62.525 176.915 62.775 177.715 ;
        RECT 62.965 177.565 64.190 177.735 ;
        RECT 62.965 177.085 63.295 177.565 ;
        RECT 63.465 176.915 63.690 177.375 ;
        RECT 63.860 177.085 64.190 177.565 ;
        RECT 64.820 177.695 64.990 178.325 ;
        RECT 65.175 177.905 65.525 178.155 ;
        RECT 65.695 177.715 65.870 178.325 ;
        RECT 66.565 178.075 66.735 178.325 ;
        RECT 66.040 177.905 66.735 178.075 ;
        RECT 66.910 177.905 67.330 178.105 ;
        RECT 67.500 177.905 67.830 178.105 ;
        RECT 68.000 177.905 68.330 178.105 ;
        RECT 64.820 177.085 65.320 177.695 ;
        RECT 65.695 177.085 66.035 177.715 ;
        RECT 66.205 176.915 66.455 177.715 ;
        RECT 66.645 177.565 67.870 177.735 ;
        RECT 66.645 177.085 66.975 177.565 ;
        RECT 67.145 176.915 67.370 177.375 ;
        RECT 67.540 177.085 67.870 177.565 ;
        RECT 68.500 177.695 68.670 178.325 ;
        RECT 69.380 178.315 69.640 179.465 ;
        RECT 69.815 178.390 70.070 179.295 ;
        RECT 70.240 178.705 70.570 179.465 ;
        RECT 70.785 178.535 70.955 179.295 ;
        RECT 68.855 177.905 69.205 178.155 ;
        RECT 68.500 177.085 69.000 177.695 ;
        RECT 69.380 176.915 69.640 177.755 ;
        RECT 69.815 177.660 69.985 178.390 ;
        RECT 70.240 178.365 70.955 178.535 ;
        RECT 71.215 178.495 71.525 179.295 ;
        RECT 71.695 178.665 72.005 179.465 ;
        RECT 72.175 178.835 72.435 179.295 ;
        RECT 72.605 179.005 72.860 179.465 ;
        RECT 73.035 178.835 73.295 179.295 ;
        RECT 72.175 178.665 73.295 178.835 ;
        RECT 70.240 178.155 70.410 178.365 ;
        RECT 71.215 178.325 72.245 178.495 ;
        RECT 70.155 177.825 70.410 178.155 ;
        RECT 69.815 177.085 70.070 177.660 ;
        RECT 70.240 177.635 70.410 177.825 ;
        RECT 70.690 177.815 71.045 178.185 ;
        RECT 70.240 177.465 70.955 177.635 ;
        RECT 70.240 176.915 70.570 177.295 ;
        RECT 70.785 177.085 70.955 177.465 ;
        RECT 71.215 177.415 71.385 178.325 ;
        RECT 71.555 177.585 71.905 178.155 ;
        RECT 72.075 178.075 72.245 178.325 ;
        RECT 73.035 178.415 73.295 178.665 ;
        RECT 73.465 178.595 73.750 179.465 ;
        RECT 73.035 178.245 73.790 178.415 ;
        RECT 73.980 178.315 74.240 179.465 ;
        RECT 74.415 178.390 74.670 179.295 ;
        RECT 74.840 178.705 75.170 179.465 ;
        RECT 75.385 178.535 75.555 179.295 ;
        RECT 76.825 178.720 77.095 179.465 ;
        RECT 77.725 179.460 84.000 179.465 ;
        RECT 77.265 178.550 77.555 179.290 ;
        RECT 77.725 178.735 77.980 179.460 ;
        RECT 78.165 178.565 78.425 179.290 ;
        RECT 78.595 178.735 78.840 179.460 ;
        RECT 79.025 178.565 79.285 179.290 ;
        RECT 79.455 178.735 79.700 179.460 ;
        RECT 79.885 178.565 80.145 179.290 ;
        RECT 80.315 178.735 80.560 179.460 ;
        RECT 80.730 178.565 80.990 179.290 ;
        RECT 81.160 178.735 81.420 179.460 ;
        RECT 81.590 178.565 81.850 179.290 ;
        RECT 82.020 178.735 82.280 179.460 ;
        RECT 82.450 178.565 82.710 179.290 ;
        RECT 82.880 178.735 83.140 179.460 ;
        RECT 83.310 178.565 83.570 179.290 ;
        RECT 83.740 178.665 84.000 179.460 ;
        RECT 78.165 178.550 83.570 178.565 ;
        RECT 72.075 177.905 73.215 178.075 ;
        RECT 73.385 177.735 73.790 178.245 ;
        RECT 72.140 177.565 73.790 177.735 ;
        RECT 71.215 177.085 71.515 177.415 ;
        RECT 71.685 176.915 71.960 177.395 ;
        RECT 72.140 177.175 72.435 177.565 ;
        RECT 72.605 176.915 72.860 177.395 ;
        RECT 73.035 177.175 73.295 177.565 ;
        RECT 73.465 176.915 73.745 177.395 ;
        RECT 73.980 176.915 74.240 177.755 ;
        RECT 74.415 177.660 74.585 178.390 ;
        RECT 74.840 178.365 75.555 178.535 ;
        RECT 74.840 178.155 75.010 178.365 ;
        RECT 76.825 178.325 83.570 178.550 ;
        RECT 74.755 177.825 75.010 178.155 ;
        RECT 74.415 177.085 74.670 177.660 ;
        RECT 74.840 177.635 75.010 177.825 ;
        RECT 75.290 177.815 75.645 178.185 ;
        RECT 76.825 177.735 77.990 178.325 ;
        RECT 84.170 178.155 84.420 179.290 ;
        RECT 84.600 178.655 84.860 179.465 ;
        RECT 85.035 178.155 85.280 179.295 ;
        RECT 85.460 178.655 85.755 179.465 ;
        RECT 85.995 178.325 86.205 179.465 ;
        RECT 86.375 178.315 86.705 179.295 ;
        RECT 86.875 178.325 87.105 179.465 ;
        RECT 78.160 177.905 85.280 178.155 ;
        RECT 74.840 177.465 75.555 177.635 ;
        RECT 76.825 177.565 83.570 177.735 ;
        RECT 74.840 176.915 75.170 177.295 ;
        RECT 75.385 177.085 75.555 177.465 ;
        RECT 76.825 176.915 77.125 177.395 ;
        RECT 77.295 177.110 77.555 177.565 ;
        RECT 77.725 176.915 77.985 177.395 ;
        RECT 78.165 177.110 78.425 177.565 ;
        RECT 78.595 176.915 78.845 177.395 ;
        RECT 79.025 177.110 79.285 177.565 ;
        RECT 79.455 176.915 79.705 177.395 ;
        RECT 79.885 177.110 80.145 177.565 ;
        RECT 80.315 176.915 80.560 177.395 ;
        RECT 80.730 177.110 81.005 177.565 ;
        RECT 81.175 176.915 81.420 177.395 ;
        RECT 81.590 177.110 81.850 177.565 ;
        RECT 82.020 176.915 82.280 177.395 ;
        RECT 82.450 177.110 82.710 177.565 ;
        RECT 82.880 176.915 83.140 177.395 ;
        RECT 83.310 177.110 83.570 177.565 ;
        RECT 83.740 176.915 84.000 177.475 ;
        RECT 84.170 177.095 84.420 177.905 ;
        RECT 84.600 176.915 84.860 177.440 ;
        RECT 85.030 177.095 85.280 177.905 ;
        RECT 85.450 177.595 85.765 178.155 ;
        RECT 85.460 176.915 85.765 177.425 ;
        RECT 85.995 176.915 86.205 177.735 ;
        RECT 86.375 177.715 86.625 178.315 ;
        RECT 87.315 178.300 87.605 179.465 ;
        RECT 87.775 178.630 88.160 179.465 ;
        RECT 88.330 178.460 88.590 179.265 ;
        RECT 88.760 178.630 89.020 179.465 ;
        RECT 89.190 178.460 89.445 179.265 ;
        RECT 89.620 178.630 89.880 179.465 ;
        RECT 90.050 178.460 90.305 179.265 ;
        RECT 90.480 178.630 90.825 179.465 ;
        RECT 91.000 178.795 91.255 179.295 ;
        RECT 91.425 178.965 91.755 179.465 ;
        RECT 91.000 178.625 91.750 178.795 ;
        RECT 87.775 178.290 90.805 178.460 ;
        RECT 86.795 177.905 87.125 178.155 ;
        RECT 86.375 177.085 86.705 177.715 ;
        RECT 86.875 176.915 87.105 177.735 ;
        RECT 87.775 177.725 88.075 178.290 ;
        RECT 88.250 177.895 90.465 178.120 ;
        RECT 90.635 177.725 90.805 178.290 ;
        RECT 91.000 177.805 91.350 178.455 ;
        RECT 87.315 176.915 87.605 177.640 ;
        RECT 87.775 177.555 90.805 177.725 ;
        RECT 91.520 177.635 91.750 178.625 ;
        RECT 88.295 176.915 88.595 177.385 ;
        RECT 88.765 177.110 89.020 177.555 ;
        RECT 89.190 176.915 89.450 177.385 ;
        RECT 89.620 177.110 89.880 177.555 ;
        RECT 91.000 177.465 91.750 177.635 ;
        RECT 90.050 176.915 90.345 177.385 ;
        RECT 91.000 177.175 91.255 177.465 ;
        RECT 91.425 176.915 91.755 177.295 ;
        RECT 91.925 177.175 92.095 179.295 ;
        RECT 92.265 178.495 92.590 179.280 ;
        RECT 92.760 179.005 93.010 179.465 ;
        RECT 93.180 178.965 93.430 179.295 ;
        RECT 93.645 178.965 94.325 179.295 ;
        RECT 93.180 178.835 93.350 178.965 ;
        RECT 92.955 178.665 93.350 178.835 ;
        RECT 92.325 177.445 92.785 178.495 ;
        RECT 92.955 177.305 93.125 178.665 ;
        RECT 93.520 178.405 93.985 178.795 ;
        RECT 93.295 177.595 93.645 178.215 ;
        RECT 93.815 177.815 93.985 178.405 ;
        RECT 94.155 178.185 94.325 178.965 ;
        RECT 94.495 178.865 94.665 179.205 ;
        RECT 94.900 179.035 95.230 179.465 ;
        RECT 95.400 178.865 95.570 179.205 ;
        RECT 95.865 179.005 96.235 179.465 ;
        RECT 94.495 178.695 95.570 178.865 ;
        RECT 96.405 178.835 96.575 179.295 ;
        RECT 96.810 178.955 97.680 179.295 ;
        RECT 97.850 179.005 98.100 179.465 ;
        RECT 96.015 178.665 96.575 178.835 ;
        RECT 96.015 178.525 96.185 178.665 ;
        RECT 94.685 178.355 96.185 178.525 ;
        RECT 96.880 178.495 97.340 178.785 ;
        RECT 94.155 178.015 95.845 178.185 ;
        RECT 93.815 177.595 94.170 177.815 ;
        RECT 94.340 177.305 94.510 178.015 ;
        RECT 94.715 177.595 95.505 177.845 ;
        RECT 95.675 177.835 95.845 178.015 ;
        RECT 96.015 177.665 96.185 178.355 ;
        RECT 92.455 176.915 92.785 177.275 ;
        RECT 92.955 177.135 93.450 177.305 ;
        RECT 93.655 177.135 94.510 177.305 ;
        RECT 95.385 176.915 95.715 177.375 ;
        RECT 95.925 177.275 96.185 177.665 ;
        RECT 96.375 178.485 97.340 178.495 ;
        RECT 97.510 178.575 97.680 178.955 ;
        RECT 98.270 178.915 98.440 179.205 ;
        RECT 98.620 179.085 98.950 179.465 ;
        RECT 98.270 178.745 99.070 178.915 ;
        RECT 96.375 178.325 97.050 178.485 ;
        RECT 97.510 178.405 98.730 178.575 ;
        RECT 96.375 177.535 96.585 178.325 ;
        RECT 97.510 178.315 97.680 178.405 ;
        RECT 96.755 177.535 97.105 178.155 ;
        RECT 97.275 178.145 97.680 178.315 ;
        RECT 97.275 177.365 97.445 178.145 ;
        RECT 97.615 177.695 97.835 177.975 ;
        RECT 98.015 177.865 98.555 178.235 ;
        RECT 98.900 178.155 99.070 178.745 ;
        RECT 99.290 178.325 99.595 179.465 ;
        RECT 99.765 178.275 100.020 179.155 ;
        RECT 100.285 178.535 100.455 179.295 ;
        RECT 100.670 178.705 101.000 179.465 ;
        RECT 100.285 178.365 101.000 178.535 ;
        RECT 101.170 178.390 101.425 179.295 ;
        RECT 98.900 178.125 99.640 178.155 ;
        RECT 97.615 177.525 98.145 177.695 ;
        RECT 95.925 177.105 96.275 177.275 ;
        RECT 96.495 177.085 97.445 177.365 ;
        RECT 97.615 176.915 97.805 177.355 ;
        RECT 97.975 177.295 98.145 177.525 ;
        RECT 98.315 177.465 98.555 177.865 ;
        RECT 98.725 177.825 99.640 178.125 ;
        RECT 98.725 177.650 99.050 177.825 ;
        RECT 98.725 177.295 99.045 177.650 ;
        RECT 99.810 177.625 100.020 178.275 ;
        RECT 100.195 177.815 100.550 178.185 ;
        RECT 100.830 178.155 101.000 178.365 ;
        RECT 100.830 177.825 101.085 178.155 ;
        RECT 100.830 177.635 101.000 177.825 ;
        RECT 101.255 177.660 101.425 178.390 ;
        RECT 101.600 178.315 101.860 179.465 ;
        RECT 102.500 178.275 102.755 179.155 ;
        RECT 102.925 178.325 103.230 179.465 ;
        RECT 103.570 179.085 103.900 179.465 ;
        RECT 104.080 178.915 104.250 179.205 ;
        RECT 104.420 179.005 104.670 179.465 ;
        RECT 103.450 178.745 104.250 178.915 ;
        RECT 104.840 178.955 105.710 179.295 ;
        RECT 97.975 177.125 99.045 177.295 ;
        RECT 99.290 176.915 99.595 177.375 ;
        RECT 99.765 177.095 100.020 177.625 ;
        RECT 100.285 177.465 101.000 177.635 ;
        RECT 100.285 177.085 100.455 177.465 ;
        RECT 100.670 176.915 101.000 177.295 ;
        RECT 101.170 177.085 101.425 177.660 ;
        RECT 101.600 176.915 101.860 177.755 ;
        RECT 102.500 177.625 102.710 178.275 ;
        RECT 103.450 178.155 103.620 178.745 ;
        RECT 104.840 178.575 105.010 178.955 ;
        RECT 105.945 178.835 106.115 179.295 ;
        RECT 106.285 179.005 106.655 179.465 ;
        RECT 106.950 178.865 107.120 179.205 ;
        RECT 107.290 179.035 107.620 179.465 ;
        RECT 107.855 178.865 108.025 179.205 ;
        RECT 103.790 178.405 105.010 178.575 ;
        RECT 105.180 178.495 105.640 178.785 ;
        RECT 105.945 178.665 106.505 178.835 ;
        RECT 106.950 178.695 108.025 178.865 ;
        RECT 108.195 178.965 108.875 179.295 ;
        RECT 109.090 178.965 109.340 179.295 ;
        RECT 109.510 179.005 109.760 179.465 ;
        RECT 106.335 178.525 106.505 178.665 ;
        RECT 105.180 178.485 106.145 178.495 ;
        RECT 104.840 178.315 105.010 178.405 ;
        RECT 105.470 178.325 106.145 178.485 ;
        RECT 102.880 178.125 103.620 178.155 ;
        RECT 102.880 177.825 103.795 178.125 ;
        RECT 103.470 177.650 103.795 177.825 ;
        RECT 102.500 177.095 102.755 177.625 ;
        RECT 102.925 176.915 103.230 177.375 ;
        RECT 103.475 177.295 103.795 177.650 ;
        RECT 103.965 177.865 104.505 178.235 ;
        RECT 104.840 178.145 105.245 178.315 ;
        RECT 103.965 177.465 104.205 177.865 ;
        RECT 104.685 177.695 104.905 177.975 ;
        RECT 104.375 177.525 104.905 177.695 ;
        RECT 104.375 177.295 104.545 177.525 ;
        RECT 105.075 177.365 105.245 178.145 ;
        RECT 105.415 177.535 105.765 178.155 ;
        RECT 105.935 177.535 106.145 178.325 ;
        RECT 106.335 178.355 107.835 178.525 ;
        RECT 106.335 177.665 106.505 178.355 ;
        RECT 108.195 178.185 108.365 178.965 ;
        RECT 109.170 178.835 109.340 178.965 ;
        RECT 106.675 178.015 108.365 178.185 ;
        RECT 108.535 178.405 109.000 178.795 ;
        RECT 109.170 178.665 109.565 178.835 ;
        RECT 106.675 177.835 106.845 178.015 ;
        RECT 103.475 177.125 104.545 177.295 ;
        RECT 104.715 176.915 104.905 177.355 ;
        RECT 105.075 177.085 106.025 177.365 ;
        RECT 106.335 177.275 106.595 177.665 ;
        RECT 107.015 177.595 107.805 177.845 ;
        RECT 106.245 177.105 106.595 177.275 ;
        RECT 106.805 176.915 107.135 177.375 ;
        RECT 108.010 177.305 108.180 178.015 ;
        RECT 108.535 177.815 108.705 178.405 ;
        RECT 108.350 177.595 108.705 177.815 ;
        RECT 108.875 177.595 109.225 178.215 ;
        RECT 109.395 177.305 109.565 178.665 ;
        RECT 109.930 178.495 110.255 179.280 ;
        RECT 109.735 177.445 110.195 178.495 ;
        RECT 108.010 177.135 108.865 177.305 ;
        RECT 109.070 177.135 109.565 177.305 ;
        RECT 109.735 176.915 110.065 177.275 ;
        RECT 110.425 177.175 110.595 179.295 ;
        RECT 110.765 178.965 111.095 179.465 ;
        RECT 111.265 178.795 111.520 179.295 ;
        RECT 110.770 178.625 111.520 178.795 ;
        RECT 110.770 177.635 111.000 178.625 ;
        RECT 111.170 177.805 111.520 178.455 ;
        RECT 112.155 178.375 113.365 179.465 ;
        RECT 112.155 177.835 112.675 178.375 ;
        RECT 112.845 177.665 113.365 178.205 ;
        RECT 110.770 177.465 111.520 177.635 ;
        RECT 110.765 176.915 111.095 177.295 ;
        RECT 111.265 177.175 111.520 177.465 ;
        RECT 112.155 176.915 113.365 177.665 ;
        RECT 26.970 176.745 113.450 176.915 ;
        RECT 27.055 175.995 28.265 176.745 ;
        RECT 28.525 176.195 28.695 176.485 ;
        RECT 28.865 176.365 29.195 176.745 ;
        RECT 28.525 176.025 29.190 176.195 ;
        RECT 27.055 175.455 27.575 175.995 ;
        RECT 27.745 175.285 28.265 175.825 ;
        RECT 27.055 174.195 28.265 175.285 ;
        RECT 28.440 175.205 28.790 175.855 ;
        RECT 28.960 175.035 29.190 176.025 ;
        RECT 28.525 174.865 29.190 175.035 ;
        RECT 28.525 174.365 28.695 174.865 ;
        RECT 28.865 174.195 29.195 174.695 ;
        RECT 29.365 174.365 29.590 176.485 ;
        RECT 29.805 176.365 30.135 176.745 ;
        RECT 30.305 176.195 30.475 176.525 ;
        RECT 30.775 176.365 31.790 176.565 ;
        RECT 29.780 176.005 30.475 176.195 ;
        RECT 29.780 175.035 29.950 176.005 ;
        RECT 30.120 175.205 30.530 175.825 ;
        RECT 30.700 175.255 30.920 176.125 ;
        RECT 31.100 175.815 31.450 176.185 ;
        RECT 31.620 175.635 31.790 176.365 ;
        RECT 31.960 176.305 32.370 176.745 ;
        RECT 32.660 176.105 32.910 176.535 ;
        RECT 33.110 176.285 33.430 176.745 ;
        RECT 33.990 176.355 34.840 176.525 ;
        RECT 31.960 175.765 32.370 176.095 ;
        RECT 32.660 175.765 33.080 176.105 ;
        RECT 31.370 175.595 31.790 175.635 ;
        RECT 31.370 175.425 32.720 175.595 ;
        RECT 29.780 174.865 30.475 175.035 ;
        RECT 30.700 174.875 31.200 175.255 ;
        RECT 29.805 174.195 30.135 174.695 ;
        RECT 30.305 174.365 30.475 174.865 ;
        RECT 31.370 174.580 31.540 175.425 ;
        RECT 32.470 175.265 32.720 175.425 ;
        RECT 31.710 174.995 31.960 175.255 ;
        RECT 32.890 174.995 33.080 175.765 ;
        RECT 31.710 174.745 33.080 174.995 ;
        RECT 33.250 175.935 34.500 176.105 ;
        RECT 33.250 175.175 33.420 175.935 ;
        RECT 34.170 175.815 34.500 175.935 ;
        RECT 33.590 175.355 33.770 175.765 ;
        RECT 34.670 175.595 34.840 176.355 ;
        RECT 35.040 176.265 35.700 176.745 ;
        RECT 35.880 176.150 36.200 176.480 ;
        RECT 35.030 175.825 35.690 176.095 ;
        RECT 35.030 175.765 35.360 175.825 ;
        RECT 35.510 175.595 35.840 175.655 ;
        RECT 33.940 175.425 35.840 175.595 ;
        RECT 33.250 174.865 33.770 175.175 ;
        RECT 33.940 174.915 34.110 175.425 ;
        RECT 36.010 175.255 36.200 176.150 ;
        RECT 34.280 175.085 36.200 175.255 ;
        RECT 35.880 175.065 36.200 175.085 ;
        RECT 36.400 175.835 36.650 176.485 ;
        RECT 36.830 176.285 37.115 176.745 ;
        RECT 37.295 176.035 37.550 176.565 ;
        RECT 36.400 175.505 37.200 175.835 ;
        RECT 33.940 174.745 35.150 174.915 ;
        RECT 30.710 174.410 31.540 174.580 ;
        RECT 31.780 174.195 32.160 174.575 ;
        RECT 32.340 174.455 32.510 174.745 ;
        RECT 33.940 174.665 34.110 174.745 ;
        RECT 32.680 174.195 33.010 174.575 ;
        RECT 33.480 174.415 34.110 174.665 ;
        RECT 34.290 174.195 34.710 174.575 ;
        RECT 34.910 174.455 35.150 174.745 ;
        RECT 35.380 174.195 35.710 174.885 ;
        RECT 35.880 174.455 36.050 175.065 ;
        RECT 36.400 174.915 36.650 175.505 ;
        RECT 37.370 175.175 37.550 176.035 ;
        RECT 38.100 176.195 38.355 176.485 ;
        RECT 38.525 176.365 38.855 176.745 ;
        RECT 38.100 176.025 38.850 176.195 ;
        RECT 38.100 175.205 38.450 175.855 ;
        RECT 36.320 174.405 36.650 174.915 ;
        RECT 36.830 174.195 37.115 174.995 ;
        RECT 37.295 174.705 37.550 175.175 ;
        RECT 38.620 175.035 38.850 176.025 ;
        RECT 38.100 174.865 38.850 175.035 ;
        RECT 37.295 174.535 37.635 174.705 ;
        RECT 37.295 174.505 37.550 174.535 ;
        RECT 38.100 174.365 38.355 174.865 ;
        RECT 38.525 174.195 38.855 174.695 ;
        RECT 39.025 174.365 39.195 176.485 ;
        RECT 39.555 176.385 39.885 176.745 ;
        RECT 40.055 176.355 40.550 176.525 ;
        RECT 40.755 176.355 41.610 176.525 ;
        RECT 39.425 175.165 39.885 176.215 ;
        RECT 39.365 174.380 39.690 175.165 ;
        RECT 40.055 174.995 40.225 176.355 ;
        RECT 40.395 175.445 40.745 176.065 ;
        RECT 40.915 175.845 41.270 176.065 ;
        RECT 40.915 175.255 41.085 175.845 ;
        RECT 41.440 175.645 41.610 176.355 ;
        RECT 42.485 176.285 42.815 176.745 ;
        RECT 43.025 176.385 43.375 176.555 ;
        RECT 41.815 175.815 42.605 176.065 ;
        RECT 43.025 175.995 43.285 176.385 ;
        RECT 43.595 176.295 44.545 176.575 ;
        RECT 44.715 176.305 44.905 176.745 ;
        RECT 45.075 176.365 46.145 176.535 ;
        RECT 42.775 175.645 42.945 175.825 ;
        RECT 40.055 174.825 40.450 174.995 ;
        RECT 40.620 174.865 41.085 175.255 ;
        RECT 41.255 175.475 42.945 175.645 ;
        RECT 40.280 174.695 40.450 174.825 ;
        RECT 41.255 174.695 41.425 175.475 ;
        RECT 43.115 175.305 43.285 175.995 ;
        RECT 41.785 175.135 43.285 175.305 ;
        RECT 43.475 175.335 43.685 176.125 ;
        RECT 43.855 175.505 44.205 176.125 ;
        RECT 44.375 175.515 44.545 176.295 ;
        RECT 45.075 176.135 45.245 176.365 ;
        RECT 44.715 175.965 45.245 176.135 ;
        RECT 44.715 175.685 44.935 175.965 ;
        RECT 45.415 175.795 45.655 176.195 ;
        RECT 44.375 175.345 44.780 175.515 ;
        RECT 45.115 175.425 45.655 175.795 ;
        RECT 45.825 176.010 46.145 176.365 ;
        RECT 46.390 176.285 46.695 176.745 ;
        RECT 46.865 176.035 47.120 176.565 ;
        RECT 45.825 175.835 46.150 176.010 ;
        RECT 45.825 175.535 46.740 175.835 ;
        RECT 46.000 175.505 46.740 175.535 ;
        RECT 43.475 175.175 44.150 175.335 ;
        RECT 44.610 175.255 44.780 175.345 ;
        RECT 43.475 175.165 44.440 175.175 ;
        RECT 43.115 174.995 43.285 175.135 ;
        RECT 39.860 174.195 40.110 174.655 ;
        RECT 40.280 174.365 40.530 174.695 ;
        RECT 40.745 174.365 41.425 174.695 ;
        RECT 41.595 174.795 42.670 174.965 ;
        RECT 43.115 174.825 43.675 174.995 ;
        RECT 43.980 174.875 44.440 175.165 ;
        RECT 44.610 175.085 45.830 175.255 ;
        RECT 41.595 174.455 41.765 174.795 ;
        RECT 42.000 174.195 42.330 174.625 ;
        RECT 42.500 174.455 42.670 174.795 ;
        RECT 42.965 174.195 43.335 174.655 ;
        RECT 43.505 174.365 43.675 174.825 ;
        RECT 44.610 174.705 44.780 175.085 ;
        RECT 46.000 174.915 46.170 175.505 ;
        RECT 46.910 175.385 47.120 176.035 ;
        RECT 47.335 175.925 47.565 176.745 ;
        RECT 47.735 175.945 48.065 176.575 ;
        RECT 47.315 175.505 47.645 175.755 ;
        RECT 43.910 174.365 44.780 174.705 ;
        RECT 45.370 174.745 46.170 174.915 ;
        RECT 44.950 174.195 45.200 174.655 ;
        RECT 45.370 174.455 45.540 174.745 ;
        RECT 45.720 174.195 46.050 174.575 ;
        RECT 46.390 174.195 46.695 175.335 ;
        RECT 46.865 174.505 47.120 175.385 ;
        RECT 47.815 175.345 48.065 175.945 ;
        RECT 48.235 175.925 48.445 176.745 ;
        RECT 48.675 176.020 48.965 176.745 ;
        RECT 49.250 176.115 49.535 176.575 ;
        RECT 49.705 176.285 49.975 176.745 ;
        RECT 49.250 175.945 50.205 176.115 ;
        RECT 47.335 174.195 47.565 175.335 ;
        RECT 47.735 174.365 48.065 175.345 ;
        RECT 48.235 174.195 48.445 175.335 ;
        RECT 48.675 174.195 48.965 175.360 ;
        RECT 49.135 175.215 49.825 175.775 ;
        RECT 49.995 175.045 50.205 175.945 ;
        RECT 49.250 174.825 50.205 175.045 ;
        RECT 50.375 175.775 50.775 176.575 ;
        RECT 50.965 176.115 51.245 176.575 ;
        RECT 51.765 176.285 52.090 176.745 ;
        RECT 50.965 175.945 52.090 176.115 ;
        RECT 52.260 176.005 52.645 176.575 ;
        RECT 51.640 175.835 52.090 175.945 ;
        RECT 50.375 175.215 51.470 175.775 ;
        RECT 51.640 175.505 52.195 175.835 ;
        RECT 49.250 174.365 49.535 174.825 ;
        RECT 49.705 174.195 49.975 174.655 ;
        RECT 50.375 174.365 50.775 175.215 ;
        RECT 51.640 175.045 52.090 175.505 ;
        RECT 52.365 175.335 52.645 176.005 ;
        RECT 52.930 176.115 53.215 176.575 ;
        RECT 53.385 176.285 53.655 176.745 ;
        RECT 52.930 175.945 53.885 176.115 ;
        RECT 50.965 174.825 52.090 175.045 ;
        RECT 50.965 174.365 51.245 174.825 ;
        RECT 51.765 174.195 52.090 174.655 ;
        RECT 52.260 174.365 52.645 175.335 ;
        RECT 52.815 175.215 53.505 175.775 ;
        RECT 53.675 175.045 53.885 175.945 ;
        RECT 52.930 174.825 53.885 175.045 ;
        RECT 54.055 175.775 54.455 176.575 ;
        RECT 54.645 176.115 54.925 176.575 ;
        RECT 55.445 176.285 55.770 176.745 ;
        RECT 54.645 175.945 55.770 176.115 ;
        RECT 55.940 176.005 56.325 176.575 ;
        RECT 55.320 175.835 55.770 175.945 ;
        RECT 54.055 175.215 55.150 175.775 ;
        RECT 55.320 175.505 55.875 175.835 ;
        RECT 52.930 174.365 53.215 174.825 ;
        RECT 53.385 174.195 53.655 174.655 ;
        RECT 54.055 174.365 54.455 175.215 ;
        RECT 55.320 175.045 55.770 175.505 ;
        RECT 56.045 175.335 56.325 176.005 ;
        RECT 54.645 174.825 55.770 175.045 ;
        RECT 54.645 174.365 54.925 174.825 ;
        RECT 55.445 174.195 55.770 174.655 ;
        RECT 55.940 174.365 56.325 175.335 ;
        RECT 56.960 176.035 57.215 176.565 ;
        RECT 57.385 176.285 57.690 176.745 ;
        RECT 57.935 176.365 59.005 176.535 ;
        RECT 56.960 175.385 57.170 176.035 ;
        RECT 57.935 176.010 58.255 176.365 ;
        RECT 57.930 175.835 58.255 176.010 ;
        RECT 57.340 175.535 58.255 175.835 ;
        RECT 58.425 175.795 58.665 176.195 ;
        RECT 58.835 176.135 59.005 176.365 ;
        RECT 59.175 176.305 59.365 176.745 ;
        RECT 59.535 176.295 60.485 176.575 ;
        RECT 60.705 176.385 61.055 176.555 ;
        RECT 58.835 175.965 59.365 176.135 ;
        RECT 57.340 175.505 58.080 175.535 ;
        RECT 56.960 174.505 57.215 175.385 ;
        RECT 57.385 174.195 57.690 175.335 ;
        RECT 57.910 174.915 58.080 175.505 ;
        RECT 58.425 175.425 58.965 175.795 ;
        RECT 59.145 175.685 59.365 175.965 ;
        RECT 59.535 175.515 59.705 176.295 ;
        RECT 59.300 175.345 59.705 175.515 ;
        RECT 59.875 175.505 60.225 176.125 ;
        RECT 59.300 175.255 59.470 175.345 ;
        RECT 60.395 175.335 60.605 176.125 ;
        RECT 58.250 175.085 59.470 175.255 ;
        RECT 59.930 175.175 60.605 175.335 ;
        RECT 57.910 174.745 58.710 174.915 ;
        RECT 58.030 174.195 58.360 174.575 ;
        RECT 58.540 174.455 58.710 174.745 ;
        RECT 59.300 174.705 59.470 175.085 ;
        RECT 59.640 175.165 60.605 175.175 ;
        RECT 60.795 175.995 61.055 176.385 ;
        RECT 61.265 176.285 61.595 176.745 ;
        RECT 62.470 176.355 63.325 176.525 ;
        RECT 63.530 176.355 64.025 176.525 ;
        RECT 64.195 176.385 64.525 176.745 ;
        RECT 60.795 175.305 60.965 175.995 ;
        RECT 61.135 175.645 61.305 175.825 ;
        RECT 61.475 175.815 62.265 176.065 ;
        RECT 62.470 175.645 62.640 176.355 ;
        RECT 62.810 175.845 63.165 176.065 ;
        RECT 61.135 175.475 62.825 175.645 ;
        RECT 59.640 174.875 60.100 175.165 ;
        RECT 60.795 175.135 62.295 175.305 ;
        RECT 60.795 174.995 60.965 175.135 ;
        RECT 60.405 174.825 60.965 174.995 ;
        RECT 58.880 174.195 59.130 174.655 ;
        RECT 59.300 174.365 60.170 174.705 ;
        RECT 60.405 174.365 60.575 174.825 ;
        RECT 61.410 174.795 62.485 174.965 ;
        RECT 60.745 174.195 61.115 174.655 ;
        RECT 61.410 174.455 61.580 174.795 ;
        RECT 61.750 174.195 62.080 174.625 ;
        RECT 62.315 174.455 62.485 174.795 ;
        RECT 62.655 174.695 62.825 175.475 ;
        RECT 62.995 175.255 63.165 175.845 ;
        RECT 63.335 175.445 63.685 176.065 ;
        RECT 62.995 174.865 63.460 175.255 ;
        RECT 63.855 174.995 64.025 176.355 ;
        RECT 64.195 175.165 64.655 176.215 ;
        RECT 63.630 174.825 64.025 174.995 ;
        RECT 63.630 174.695 63.800 174.825 ;
        RECT 62.655 174.365 63.335 174.695 ;
        RECT 63.550 174.365 63.800 174.695 ;
        RECT 63.970 174.195 64.220 174.655 ;
        RECT 64.390 174.380 64.715 175.165 ;
        RECT 64.885 174.365 65.055 176.485 ;
        RECT 65.225 176.365 65.555 176.745 ;
        RECT 65.725 176.195 65.980 176.485 ;
        RECT 66.215 176.265 66.495 176.745 ;
        RECT 65.230 176.025 65.980 176.195 ;
        RECT 66.665 176.095 66.925 176.485 ;
        RECT 67.100 176.265 67.355 176.745 ;
        RECT 67.525 176.095 67.820 176.485 ;
        RECT 68.000 176.265 68.275 176.745 ;
        RECT 68.445 176.245 68.745 176.575 ;
        RECT 65.230 175.035 65.460 176.025 ;
        RECT 66.170 175.925 67.820 176.095 ;
        RECT 65.630 175.205 65.980 175.855 ;
        RECT 66.170 175.415 66.575 175.925 ;
        RECT 66.745 175.585 67.885 175.755 ;
        RECT 66.170 175.245 66.925 175.415 ;
        RECT 65.230 174.865 65.980 175.035 ;
        RECT 65.225 174.195 65.555 174.695 ;
        RECT 65.725 174.365 65.980 174.865 ;
        RECT 66.210 174.195 66.495 175.065 ;
        RECT 66.665 174.995 66.925 175.245 ;
        RECT 67.715 175.335 67.885 175.585 ;
        RECT 68.055 175.505 68.405 176.075 ;
        RECT 68.575 175.335 68.745 176.245 ;
        RECT 69.005 176.195 69.175 176.575 ;
        RECT 69.390 176.365 69.720 176.745 ;
        RECT 69.005 176.025 69.720 176.195 ;
        RECT 68.915 175.475 69.270 175.845 ;
        RECT 69.550 175.835 69.720 176.025 ;
        RECT 69.890 176.000 70.145 176.575 ;
        RECT 69.550 175.505 69.805 175.835 ;
        RECT 67.715 175.165 68.745 175.335 ;
        RECT 69.550 175.295 69.720 175.505 ;
        RECT 66.665 174.825 67.785 174.995 ;
        RECT 66.665 174.365 66.925 174.825 ;
        RECT 67.100 174.195 67.355 174.655 ;
        RECT 67.525 174.365 67.785 174.825 ;
        RECT 67.955 174.195 68.265 174.995 ;
        RECT 68.435 174.365 68.745 175.165 ;
        RECT 69.005 175.125 69.720 175.295 ;
        RECT 69.975 175.270 70.145 176.000 ;
        RECT 70.320 175.905 70.580 176.745 ;
        RECT 70.755 175.985 71.465 176.575 ;
        RECT 71.975 176.215 72.305 176.575 ;
        RECT 72.505 176.385 72.835 176.745 ;
        RECT 73.005 176.215 73.335 176.575 ;
        RECT 71.975 176.005 73.335 176.215 ;
        RECT 74.435 176.020 74.725 176.745 ;
        RECT 70.755 175.895 70.985 175.985 ;
        RECT 74.935 175.925 75.165 176.745 ;
        RECT 75.335 175.945 75.665 176.575 ;
        RECT 69.005 174.365 69.175 175.125 ;
        RECT 69.390 174.195 69.720 174.955 ;
        RECT 69.890 174.365 70.145 175.270 ;
        RECT 70.320 174.195 70.580 175.345 ;
        RECT 70.755 175.015 70.960 175.895 ;
        RECT 71.130 175.215 71.460 175.755 ;
        RECT 71.635 175.505 72.130 175.835 ;
        RECT 72.450 175.505 72.825 175.835 ;
        RECT 73.035 175.505 73.345 175.835 ;
        RECT 74.915 175.505 75.245 175.755 ;
        RECT 71.635 175.215 71.960 175.505 ;
        RECT 72.155 175.015 72.485 175.235 ;
        RECT 70.755 174.785 72.485 175.015 ;
        RECT 70.755 174.365 71.455 174.785 ;
        RECT 71.655 174.195 71.985 174.555 ;
        RECT 72.155 174.385 72.485 174.785 ;
        RECT 72.655 174.580 72.825 175.505 ;
        RECT 73.005 174.195 73.335 175.255 ;
        RECT 74.435 174.195 74.725 175.360 ;
        RECT 75.415 175.345 75.665 175.945 ;
        RECT 75.835 175.925 76.045 176.745 ;
        RECT 76.650 176.035 76.905 176.565 ;
        RECT 77.085 176.285 77.370 176.745 ;
        RECT 76.650 175.385 76.830 176.035 ;
        RECT 77.550 175.835 77.800 176.485 ;
        RECT 77.000 175.505 77.800 175.835 ;
        RECT 74.935 174.195 75.165 175.335 ;
        RECT 75.335 174.365 75.665 175.345 ;
        RECT 75.835 174.195 76.045 175.335 ;
        RECT 76.565 175.215 76.830 175.385 ;
        RECT 76.650 175.175 76.830 175.215 ;
        RECT 76.650 174.505 76.905 175.175 ;
        RECT 77.085 174.195 77.370 174.995 ;
        RECT 77.550 174.915 77.800 175.505 ;
        RECT 78.000 176.150 78.320 176.480 ;
        RECT 78.500 176.265 79.160 176.745 ;
        RECT 79.360 176.355 80.210 176.525 ;
        RECT 78.000 175.255 78.190 176.150 ;
        RECT 78.510 175.825 79.170 176.095 ;
        RECT 78.840 175.765 79.170 175.825 ;
        RECT 78.360 175.595 78.690 175.655 ;
        RECT 79.360 175.595 79.530 176.355 ;
        RECT 80.770 176.285 81.090 176.745 ;
        RECT 81.290 176.105 81.540 176.535 ;
        RECT 81.830 176.305 82.240 176.745 ;
        RECT 82.410 176.365 83.425 176.565 ;
        RECT 79.700 175.935 80.950 176.105 ;
        RECT 79.700 175.815 80.030 175.935 ;
        RECT 78.360 175.425 80.260 175.595 ;
        RECT 78.000 175.085 79.920 175.255 ;
        RECT 78.000 175.065 78.320 175.085 ;
        RECT 77.550 174.405 77.880 174.915 ;
        RECT 78.150 174.455 78.320 175.065 ;
        RECT 80.090 174.915 80.260 175.425 ;
        RECT 80.430 175.355 80.610 175.765 ;
        RECT 80.780 175.175 80.950 175.935 ;
        RECT 78.490 174.195 78.820 174.885 ;
        RECT 79.050 174.745 80.260 174.915 ;
        RECT 80.430 174.865 80.950 175.175 ;
        RECT 81.120 175.765 81.540 176.105 ;
        RECT 81.830 175.765 82.240 176.095 ;
        RECT 81.120 174.995 81.310 175.765 ;
        RECT 82.410 175.635 82.580 176.365 ;
        RECT 83.725 176.195 83.895 176.525 ;
        RECT 84.065 176.365 84.395 176.745 ;
        RECT 82.750 175.815 83.100 176.185 ;
        RECT 82.410 175.595 82.830 175.635 ;
        RECT 81.480 175.425 82.830 175.595 ;
        RECT 81.480 175.265 81.730 175.425 ;
        RECT 82.240 174.995 82.490 175.255 ;
        RECT 81.120 174.745 82.490 174.995 ;
        RECT 79.050 174.455 79.290 174.745 ;
        RECT 80.090 174.665 80.260 174.745 ;
        RECT 79.490 174.195 79.910 174.575 ;
        RECT 80.090 174.415 80.720 174.665 ;
        RECT 81.190 174.195 81.520 174.575 ;
        RECT 81.690 174.455 81.860 174.745 ;
        RECT 82.660 174.580 82.830 175.425 ;
        RECT 83.280 175.255 83.500 176.125 ;
        RECT 83.725 176.005 84.420 176.195 ;
        RECT 83.000 174.875 83.500 175.255 ;
        RECT 83.670 175.205 84.080 175.825 ;
        RECT 84.250 175.035 84.420 176.005 ;
        RECT 83.725 174.865 84.420 175.035 ;
        RECT 82.040 174.195 82.420 174.575 ;
        RECT 82.660 174.410 83.490 174.580 ;
        RECT 83.725 174.365 83.895 174.865 ;
        RECT 84.065 174.195 84.395 174.695 ;
        RECT 84.610 174.365 84.835 176.485 ;
        RECT 85.005 176.365 85.335 176.745 ;
        RECT 85.505 176.195 85.675 176.485 ;
        RECT 85.935 176.235 86.240 176.745 ;
        RECT 85.010 176.025 85.675 176.195 ;
        RECT 85.010 175.035 85.240 176.025 ;
        RECT 85.410 175.205 85.760 175.855 ;
        RECT 85.935 175.505 86.250 176.065 ;
        RECT 86.420 175.755 86.670 176.565 ;
        RECT 86.840 176.220 87.100 176.745 ;
        RECT 87.280 175.755 87.530 176.565 ;
        RECT 87.700 176.185 87.960 176.745 ;
        RECT 88.130 176.095 88.390 176.550 ;
        RECT 88.560 176.265 88.820 176.745 ;
        RECT 88.990 176.095 89.250 176.550 ;
        RECT 89.420 176.265 89.680 176.745 ;
        RECT 89.850 176.095 90.110 176.550 ;
        RECT 90.280 176.265 90.525 176.745 ;
        RECT 90.695 176.095 90.970 176.550 ;
        RECT 91.140 176.265 91.385 176.745 ;
        RECT 91.555 176.095 91.815 176.550 ;
        RECT 91.995 176.265 92.245 176.745 ;
        RECT 92.415 176.095 92.675 176.550 ;
        RECT 92.855 176.265 93.105 176.745 ;
        RECT 93.275 176.095 93.535 176.550 ;
        RECT 93.715 176.265 93.975 176.745 ;
        RECT 94.145 176.095 94.405 176.550 ;
        RECT 94.575 176.265 94.875 176.745 ;
        RECT 88.130 176.065 94.875 176.095 ;
        RECT 88.130 175.925 94.905 176.065 ;
        RECT 95.410 175.935 95.655 176.540 ;
        RECT 95.875 176.210 96.385 176.745 ;
        RECT 93.710 175.895 94.905 175.925 ;
        RECT 86.420 175.505 93.540 175.755 ;
        RECT 85.010 174.865 85.675 175.035 ;
        RECT 85.005 174.195 85.335 174.695 ;
        RECT 85.505 174.365 85.675 174.865 ;
        RECT 85.945 174.195 86.240 175.005 ;
        RECT 86.420 174.365 86.665 175.505 ;
        RECT 86.840 174.195 87.100 175.005 ;
        RECT 87.280 174.370 87.530 175.505 ;
        RECT 93.710 175.335 94.875 175.895 ;
        RECT 88.130 175.110 94.875 175.335 ;
        RECT 95.135 175.765 96.365 175.935 ;
        RECT 88.130 175.095 93.535 175.110 ;
        RECT 87.700 174.200 87.960 174.995 ;
        RECT 88.130 174.370 88.390 175.095 ;
        RECT 88.560 174.200 88.820 174.925 ;
        RECT 88.990 174.370 89.250 175.095 ;
        RECT 89.420 174.200 89.680 174.925 ;
        RECT 89.850 174.370 90.110 175.095 ;
        RECT 90.280 174.200 90.540 174.925 ;
        RECT 90.710 174.370 90.970 175.095 ;
        RECT 91.140 174.200 91.385 174.925 ;
        RECT 91.555 174.370 91.815 175.095 ;
        RECT 92.000 174.200 92.245 174.925 ;
        RECT 92.415 174.370 92.675 175.095 ;
        RECT 92.860 174.200 93.105 174.925 ;
        RECT 93.275 174.370 93.535 175.095 ;
        RECT 93.720 174.200 93.975 174.925 ;
        RECT 94.145 174.370 94.435 175.110 ;
        RECT 95.135 174.955 95.475 175.765 ;
        RECT 95.645 175.200 96.395 175.390 ;
        RECT 87.700 174.195 93.975 174.200 ;
        RECT 94.605 174.195 94.875 174.940 ;
        RECT 95.135 174.545 95.650 174.955 ;
        RECT 95.885 174.195 96.055 174.955 ;
        RECT 96.225 174.535 96.395 175.200 ;
        RECT 96.565 175.215 96.755 176.575 ;
        RECT 96.925 176.065 97.200 176.575 ;
        RECT 97.390 176.210 97.920 176.575 ;
        RECT 98.345 176.345 98.675 176.745 ;
        RECT 97.745 176.175 97.920 176.210 ;
        RECT 96.925 175.895 97.205 176.065 ;
        RECT 96.925 175.415 97.200 175.895 ;
        RECT 97.405 175.215 97.575 176.015 ;
        RECT 96.565 175.045 97.575 175.215 ;
        RECT 97.745 176.005 98.675 176.175 ;
        RECT 98.845 176.005 99.100 176.575 ;
        RECT 100.195 176.020 100.485 176.745 ;
        RECT 97.745 174.875 97.915 176.005 ;
        RECT 98.505 175.835 98.675 176.005 ;
        RECT 96.790 174.705 97.915 174.875 ;
        RECT 98.085 175.505 98.280 175.835 ;
        RECT 98.505 175.505 98.760 175.835 ;
        RECT 98.085 174.535 98.255 175.505 ;
        RECT 98.930 175.335 99.100 176.005 ;
        RECT 101.390 175.935 101.635 176.540 ;
        RECT 101.855 176.210 102.365 176.745 ;
        RECT 101.115 175.765 102.345 175.935 ;
        RECT 96.225 174.365 98.255 174.535 ;
        RECT 98.425 174.195 98.595 175.335 ;
        RECT 98.765 174.365 99.100 175.335 ;
        RECT 100.195 174.195 100.485 175.360 ;
        RECT 101.115 174.955 101.455 175.765 ;
        RECT 101.625 175.200 102.375 175.390 ;
        RECT 101.115 174.545 101.630 174.955 ;
        RECT 101.865 174.195 102.035 174.955 ;
        RECT 102.205 174.535 102.375 175.200 ;
        RECT 102.545 175.215 102.735 176.575 ;
        RECT 102.905 175.725 103.180 176.575 ;
        RECT 103.370 176.210 103.900 176.575 ;
        RECT 104.325 176.345 104.655 176.745 ;
        RECT 103.725 176.175 103.900 176.210 ;
        RECT 102.905 175.555 103.185 175.725 ;
        RECT 102.905 175.415 103.180 175.555 ;
        RECT 103.385 175.215 103.555 176.015 ;
        RECT 102.545 175.045 103.555 175.215 ;
        RECT 103.725 176.005 104.655 176.175 ;
        RECT 104.825 176.005 105.080 176.575 ;
        RECT 103.725 174.875 103.895 176.005 ;
        RECT 104.485 175.835 104.655 176.005 ;
        RECT 102.770 174.705 103.895 174.875 ;
        RECT 104.065 175.505 104.260 175.835 ;
        RECT 104.485 175.505 104.740 175.835 ;
        RECT 104.065 174.535 104.235 175.505 ;
        RECT 104.910 175.335 105.080 176.005 ;
        RECT 105.530 175.935 105.775 176.540 ;
        RECT 105.995 176.210 106.505 176.745 ;
        RECT 102.205 174.365 104.235 174.535 ;
        RECT 104.405 174.195 104.575 175.335 ;
        RECT 104.745 174.365 105.080 175.335 ;
        RECT 105.255 175.765 106.485 175.935 ;
        RECT 105.255 174.955 105.595 175.765 ;
        RECT 105.765 175.200 106.515 175.390 ;
        RECT 105.255 174.545 105.770 174.955 ;
        RECT 106.005 174.195 106.175 174.955 ;
        RECT 106.345 174.535 106.515 175.200 ;
        RECT 106.685 175.215 106.875 176.575 ;
        RECT 107.045 176.405 107.320 176.575 ;
        RECT 107.045 176.235 107.325 176.405 ;
        RECT 107.045 175.415 107.320 176.235 ;
        RECT 107.510 176.210 108.040 176.575 ;
        RECT 108.465 176.345 108.795 176.745 ;
        RECT 107.865 176.175 108.040 176.210 ;
        RECT 107.525 175.215 107.695 176.015 ;
        RECT 106.685 175.045 107.695 175.215 ;
        RECT 107.865 176.005 108.795 176.175 ;
        RECT 108.965 176.005 109.220 176.575 ;
        RECT 107.865 174.875 108.035 176.005 ;
        RECT 108.625 175.835 108.795 176.005 ;
        RECT 106.910 174.705 108.035 174.875 ;
        RECT 108.205 175.505 108.400 175.835 ;
        RECT 108.625 175.505 108.880 175.835 ;
        RECT 108.205 174.535 108.375 175.505 ;
        RECT 109.050 175.335 109.220 176.005 ;
        RECT 109.485 176.095 109.655 176.575 ;
        RECT 109.835 176.265 110.075 176.745 ;
        RECT 110.325 176.095 110.495 176.575 ;
        RECT 110.665 176.265 110.995 176.745 ;
        RECT 111.165 176.095 111.335 176.575 ;
        RECT 109.485 175.925 110.120 176.095 ;
        RECT 110.325 175.925 111.335 176.095 ;
        RECT 111.505 175.945 111.835 176.745 ;
        RECT 112.155 175.995 113.365 176.745 ;
        RECT 109.950 175.755 110.120 175.925 ;
        RECT 109.400 175.515 109.780 175.755 ;
        RECT 109.950 175.585 110.450 175.755 ;
        RECT 109.950 175.345 110.120 175.585 ;
        RECT 110.840 175.385 111.335 175.925 ;
        RECT 106.345 174.365 108.375 174.535 ;
        RECT 108.545 174.195 108.715 175.335 ;
        RECT 108.885 174.365 109.220 175.335 ;
        RECT 109.405 175.175 110.120 175.345 ;
        RECT 110.325 175.215 111.335 175.385 ;
        RECT 109.405 174.365 109.735 175.175 ;
        RECT 109.905 174.195 110.145 174.995 ;
        RECT 110.325 174.365 110.495 175.215 ;
        RECT 110.665 174.195 110.995 174.995 ;
        RECT 111.165 174.365 111.335 175.215 ;
        RECT 111.505 174.195 111.835 175.345 ;
        RECT 112.155 175.285 112.675 175.825 ;
        RECT 112.845 175.455 113.365 175.995 ;
        RECT 112.155 174.195 113.365 175.285 ;
        RECT 26.970 174.025 113.450 174.195 ;
        RECT 27.055 172.935 28.265 174.025 ;
        RECT 28.635 173.355 28.915 174.025 ;
        RECT 29.085 173.135 29.385 173.685 ;
        RECT 29.585 173.305 29.915 174.025 ;
        RECT 30.105 173.305 30.565 173.855 ;
        RECT 27.055 172.225 27.575 172.765 ;
        RECT 27.745 172.395 28.265 172.935 ;
        RECT 28.450 172.715 28.715 173.075 ;
        RECT 29.085 172.965 30.025 173.135 ;
        RECT 29.855 172.715 30.025 172.965 ;
        RECT 28.450 172.465 29.125 172.715 ;
        RECT 29.345 172.465 29.685 172.715 ;
        RECT 29.855 172.385 30.145 172.715 ;
        RECT 29.855 172.295 30.025 172.385 ;
        RECT 27.055 171.475 28.265 172.225 ;
        RECT 28.635 172.105 30.025 172.295 ;
        RECT 28.635 171.745 28.965 172.105 ;
        RECT 30.315 171.935 30.565 173.305 ;
        RECT 29.585 171.475 29.835 171.935 ;
        RECT 30.005 171.645 30.565 171.935 ;
        RECT 31.660 172.885 31.995 173.855 ;
        RECT 32.165 172.885 32.335 174.025 ;
        RECT 32.505 173.685 34.535 173.855 ;
        RECT 31.660 172.215 31.830 172.885 ;
        RECT 32.505 172.715 32.675 173.685 ;
        RECT 32.000 172.385 32.255 172.715 ;
        RECT 32.480 172.385 32.675 172.715 ;
        RECT 32.845 173.345 33.970 173.515 ;
        RECT 32.085 172.215 32.255 172.385 ;
        RECT 32.845 172.215 33.015 173.345 ;
        RECT 31.660 171.645 31.915 172.215 ;
        RECT 32.085 172.045 33.015 172.215 ;
        RECT 33.185 173.005 34.195 173.175 ;
        RECT 33.185 172.205 33.355 173.005 ;
        RECT 32.840 172.010 33.015 172.045 ;
        RECT 32.085 171.475 32.415 171.875 ;
        RECT 32.840 171.645 33.370 172.010 ;
        RECT 33.560 171.985 33.835 172.805 ;
        RECT 33.555 171.815 33.835 171.985 ;
        RECT 33.560 171.645 33.835 171.815 ;
        RECT 34.005 171.645 34.195 173.005 ;
        RECT 34.365 173.020 34.535 173.685 ;
        RECT 34.705 173.265 34.875 174.025 ;
        RECT 35.110 173.265 35.625 173.675 ;
        RECT 34.365 172.830 35.115 173.020 ;
        RECT 35.285 172.455 35.625 173.265 ;
        RECT 35.795 172.860 36.085 174.025 ;
        RECT 36.310 173.225 36.610 174.025 ;
        RECT 36.780 173.055 37.110 173.855 ;
        RECT 37.280 173.225 37.450 174.025 ;
        RECT 37.620 173.055 37.950 173.855 ;
        RECT 38.120 173.225 38.290 174.025 ;
        RECT 38.460 173.055 38.790 173.855 ;
        RECT 38.960 173.225 39.130 174.025 ;
        RECT 39.300 173.055 39.630 173.855 ;
        RECT 39.800 173.225 40.055 174.025 ;
        RECT 40.400 173.355 40.655 173.855 ;
        RECT 40.825 173.525 41.155 174.025 ;
        RECT 40.400 173.185 41.150 173.355 ;
        RECT 36.255 172.885 40.225 173.055 ;
        RECT 34.395 172.285 35.625 172.455 ;
        RECT 36.255 172.295 36.575 172.885 ;
        RECT 36.775 172.665 39.630 172.715 ;
        RECT 36.775 172.495 39.705 172.665 ;
        RECT 36.775 172.465 39.630 172.495 ;
        RECT 39.880 172.295 40.225 172.885 ;
        RECT 40.400 172.365 40.750 173.015 ;
        RECT 34.375 171.475 34.885 172.010 ;
        RECT 35.105 171.680 35.350 172.285 ;
        RECT 35.795 171.475 36.085 172.200 ;
        RECT 36.255 172.105 40.225 172.295 ;
        RECT 40.920 172.195 41.150 173.185 ;
        RECT 36.305 171.475 36.610 171.935 ;
        RECT 36.780 171.645 37.110 172.105 ;
        RECT 37.280 171.475 37.450 171.935 ;
        RECT 37.620 171.645 37.950 172.105 ;
        RECT 38.120 171.475 38.290 171.935 ;
        RECT 38.460 171.645 38.790 172.105 ;
        RECT 38.960 171.475 39.130 171.935 ;
        RECT 39.300 171.645 39.630 172.105 ;
        RECT 40.400 172.025 41.150 172.195 ;
        RECT 39.800 171.475 40.055 171.935 ;
        RECT 40.400 171.735 40.655 172.025 ;
        RECT 40.825 171.475 41.155 171.855 ;
        RECT 41.325 171.735 41.495 173.855 ;
        RECT 41.665 173.055 41.990 173.840 ;
        RECT 42.160 173.565 42.410 174.025 ;
        RECT 42.580 173.525 42.830 173.855 ;
        RECT 43.045 173.525 43.725 173.855 ;
        RECT 42.580 173.395 42.750 173.525 ;
        RECT 42.355 173.225 42.750 173.395 ;
        RECT 41.725 172.005 42.185 173.055 ;
        RECT 42.355 171.865 42.525 173.225 ;
        RECT 42.920 172.965 43.385 173.355 ;
        RECT 42.695 172.155 43.045 172.775 ;
        RECT 43.215 172.375 43.385 172.965 ;
        RECT 43.555 172.745 43.725 173.525 ;
        RECT 43.895 173.425 44.065 173.765 ;
        RECT 44.300 173.595 44.630 174.025 ;
        RECT 44.800 173.425 44.970 173.765 ;
        RECT 45.265 173.565 45.635 174.025 ;
        RECT 43.895 173.255 44.970 173.425 ;
        RECT 45.805 173.395 45.975 173.855 ;
        RECT 46.210 173.515 47.080 173.855 ;
        RECT 47.250 173.565 47.500 174.025 ;
        RECT 45.415 173.225 45.975 173.395 ;
        RECT 45.415 173.085 45.585 173.225 ;
        RECT 44.085 172.915 45.585 173.085 ;
        RECT 46.280 173.055 46.740 173.345 ;
        RECT 43.555 172.575 45.245 172.745 ;
        RECT 43.215 172.155 43.570 172.375 ;
        RECT 43.740 171.865 43.910 172.575 ;
        RECT 44.115 172.155 44.905 172.405 ;
        RECT 45.075 172.395 45.245 172.575 ;
        RECT 45.415 172.225 45.585 172.915 ;
        RECT 41.855 171.475 42.185 171.835 ;
        RECT 42.355 171.695 42.850 171.865 ;
        RECT 43.055 171.695 43.910 171.865 ;
        RECT 44.785 171.475 45.115 171.935 ;
        RECT 45.325 171.835 45.585 172.225 ;
        RECT 45.775 173.045 46.740 173.055 ;
        RECT 46.910 173.135 47.080 173.515 ;
        RECT 47.670 173.475 47.840 173.765 ;
        RECT 48.020 173.645 48.350 174.025 ;
        RECT 47.670 173.305 48.470 173.475 ;
        RECT 45.775 172.885 46.450 173.045 ;
        RECT 46.910 172.965 48.130 173.135 ;
        RECT 45.775 172.095 45.985 172.885 ;
        RECT 46.910 172.875 47.080 172.965 ;
        RECT 46.155 172.095 46.505 172.715 ;
        RECT 46.675 172.705 47.080 172.875 ;
        RECT 46.675 171.925 46.845 172.705 ;
        RECT 47.015 172.255 47.235 172.535 ;
        RECT 47.415 172.425 47.955 172.795 ;
        RECT 48.300 172.715 48.470 173.305 ;
        RECT 48.690 172.885 48.995 174.025 ;
        RECT 49.165 172.835 49.420 173.715 ;
        RECT 49.600 173.355 49.855 173.855 ;
        RECT 50.025 173.525 50.355 174.025 ;
        RECT 49.600 173.185 50.350 173.355 ;
        RECT 48.300 172.685 49.040 172.715 ;
        RECT 47.015 172.085 47.545 172.255 ;
        RECT 45.325 171.665 45.675 171.835 ;
        RECT 45.895 171.645 46.845 171.925 ;
        RECT 47.015 171.475 47.205 171.915 ;
        RECT 47.375 171.855 47.545 172.085 ;
        RECT 47.715 172.025 47.955 172.425 ;
        RECT 48.125 172.385 49.040 172.685 ;
        RECT 48.125 172.210 48.450 172.385 ;
        RECT 48.125 171.855 48.445 172.210 ;
        RECT 49.210 172.185 49.420 172.835 ;
        RECT 49.600 172.365 49.950 173.015 ;
        RECT 50.120 172.195 50.350 173.185 ;
        RECT 47.375 171.685 48.445 171.855 ;
        RECT 48.690 171.475 48.995 171.935 ;
        RECT 49.165 171.655 49.420 172.185 ;
        RECT 49.600 172.025 50.350 172.195 ;
        RECT 49.600 171.735 49.855 172.025 ;
        RECT 50.025 171.475 50.355 171.855 ;
        RECT 50.525 171.735 50.695 173.855 ;
        RECT 50.865 173.055 51.190 173.840 ;
        RECT 51.360 173.565 51.610 174.025 ;
        RECT 51.780 173.525 52.030 173.855 ;
        RECT 52.245 173.525 52.925 173.855 ;
        RECT 51.780 173.395 51.950 173.525 ;
        RECT 51.555 173.225 51.950 173.395 ;
        RECT 50.925 172.005 51.385 173.055 ;
        RECT 51.555 171.865 51.725 173.225 ;
        RECT 52.120 172.965 52.585 173.355 ;
        RECT 51.895 172.155 52.245 172.775 ;
        RECT 52.415 172.375 52.585 172.965 ;
        RECT 52.755 172.745 52.925 173.525 ;
        RECT 53.095 173.425 53.265 173.765 ;
        RECT 53.500 173.595 53.830 174.025 ;
        RECT 54.000 173.425 54.170 173.765 ;
        RECT 54.465 173.565 54.835 174.025 ;
        RECT 53.095 173.255 54.170 173.425 ;
        RECT 55.005 173.395 55.175 173.855 ;
        RECT 55.410 173.515 56.280 173.855 ;
        RECT 56.450 173.565 56.700 174.025 ;
        RECT 54.615 173.225 55.175 173.395 ;
        RECT 54.615 173.085 54.785 173.225 ;
        RECT 53.285 172.915 54.785 173.085 ;
        RECT 55.480 173.055 55.940 173.345 ;
        RECT 52.755 172.575 54.445 172.745 ;
        RECT 52.415 172.155 52.770 172.375 ;
        RECT 52.940 171.865 53.110 172.575 ;
        RECT 53.315 172.155 54.105 172.405 ;
        RECT 54.275 172.395 54.445 172.575 ;
        RECT 54.615 172.225 54.785 172.915 ;
        RECT 51.055 171.475 51.385 171.835 ;
        RECT 51.555 171.695 52.050 171.865 ;
        RECT 52.255 171.695 53.110 171.865 ;
        RECT 53.985 171.475 54.315 171.935 ;
        RECT 54.525 171.835 54.785 172.225 ;
        RECT 54.975 173.045 55.940 173.055 ;
        RECT 56.110 173.135 56.280 173.515 ;
        RECT 56.870 173.475 57.040 173.765 ;
        RECT 57.220 173.645 57.550 174.025 ;
        RECT 56.870 173.305 57.670 173.475 ;
        RECT 54.975 172.885 55.650 173.045 ;
        RECT 56.110 172.965 57.330 173.135 ;
        RECT 54.975 172.095 55.185 172.885 ;
        RECT 56.110 172.875 56.280 172.965 ;
        RECT 55.355 172.095 55.705 172.715 ;
        RECT 55.875 172.705 56.280 172.875 ;
        RECT 55.875 171.925 56.045 172.705 ;
        RECT 56.215 172.255 56.435 172.535 ;
        RECT 56.615 172.425 57.155 172.795 ;
        RECT 57.500 172.715 57.670 173.305 ;
        RECT 57.890 172.885 58.195 174.025 ;
        RECT 58.365 172.835 58.620 173.715 ;
        RECT 58.945 172.875 59.275 174.025 ;
        RECT 59.445 173.005 59.615 173.855 ;
        RECT 59.785 173.225 60.115 174.025 ;
        RECT 60.285 173.005 60.455 173.855 ;
        RECT 60.635 173.225 60.875 174.025 ;
        RECT 61.045 173.045 61.375 173.855 ;
        RECT 57.500 172.685 58.240 172.715 ;
        RECT 56.215 172.085 56.745 172.255 ;
        RECT 54.525 171.665 54.875 171.835 ;
        RECT 55.095 171.645 56.045 171.925 ;
        RECT 56.215 171.475 56.405 171.915 ;
        RECT 56.575 171.855 56.745 172.085 ;
        RECT 56.915 172.025 57.155 172.425 ;
        RECT 57.325 172.385 58.240 172.685 ;
        RECT 57.325 172.210 57.650 172.385 ;
        RECT 57.325 171.855 57.645 172.210 ;
        RECT 58.410 172.185 58.620 172.835 ;
        RECT 59.445 172.835 60.455 173.005 ;
        RECT 60.660 172.875 61.375 173.045 ;
        RECT 59.445 172.295 59.940 172.835 ;
        RECT 60.660 172.635 60.830 172.875 ;
        RECT 61.555 172.860 61.845 174.025 ;
        RECT 62.020 172.835 62.275 173.715 ;
        RECT 62.445 172.885 62.750 174.025 ;
        RECT 63.090 173.645 63.420 174.025 ;
        RECT 63.600 173.475 63.770 173.765 ;
        RECT 63.940 173.565 64.190 174.025 ;
        RECT 62.970 173.305 63.770 173.475 ;
        RECT 64.360 173.515 65.230 173.855 ;
        RECT 60.330 172.465 60.830 172.635 ;
        RECT 61.000 172.465 61.380 172.705 ;
        RECT 60.660 172.295 60.830 172.465 ;
        RECT 56.575 171.685 57.645 171.855 ;
        RECT 57.890 171.475 58.195 171.935 ;
        RECT 58.365 171.655 58.620 172.185 ;
        RECT 58.945 171.475 59.275 172.275 ;
        RECT 59.445 172.125 60.455 172.295 ;
        RECT 60.660 172.125 61.295 172.295 ;
        RECT 59.445 171.645 59.615 172.125 ;
        RECT 59.785 171.475 60.115 171.955 ;
        RECT 60.285 171.645 60.455 172.125 ;
        RECT 60.705 171.475 60.945 171.955 ;
        RECT 61.125 171.645 61.295 172.125 ;
        RECT 61.555 171.475 61.845 172.200 ;
        RECT 62.020 172.185 62.230 172.835 ;
        RECT 62.970 172.715 63.140 173.305 ;
        RECT 64.360 173.135 64.530 173.515 ;
        RECT 65.465 173.395 65.635 173.855 ;
        RECT 65.805 173.565 66.175 174.025 ;
        RECT 66.470 173.425 66.640 173.765 ;
        RECT 66.810 173.595 67.140 174.025 ;
        RECT 67.375 173.425 67.545 173.765 ;
        RECT 63.310 172.965 64.530 173.135 ;
        RECT 64.700 173.055 65.160 173.345 ;
        RECT 65.465 173.225 66.025 173.395 ;
        RECT 66.470 173.255 67.545 173.425 ;
        RECT 67.715 173.525 68.395 173.855 ;
        RECT 68.610 173.525 68.860 173.855 ;
        RECT 69.030 173.565 69.280 174.025 ;
        RECT 65.855 173.085 66.025 173.225 ;
        RECT 64.700 173.045 65.665 173.055 ;
        RECT 64.360 172.875 64.530 172.965 ;
        RECT 64.990 172.885 65.665 173.045 ;
        RECT 62.400 172.685 63.140 172.715 ;
        RECT 62.400 172.385 63.315 172.685 ;
        RECT 62.990 172.210 63.315 172.385 ;
        RECT 62.020 171.655 62.275 172.185 ;
        RECT 62.445 171.475 62.750 171.935 ;
        RECT 62.995 171.855 63.315 172.210 ;
        RECT 63.485 172.425 64.025 172.795 ;
        RECT 64.360 172.705 64.765 172.875 ;
        RECT 63.485 172.025 63.725 172.425 ;
        RECT 64.205 172.255 64.425 172.535 ;
        RECT 63.895 172.085 64.425 172.255 ;
        RECT 63.895 171.855 64.065 172.085 ;
        RECT 64.595 171.925 64.765 172.705 ;
        RECT 64.935 172.095 65.285 172.715 ;
        RECT 65.455 172.095 65.665 172.885 ;
        RECT 65.855 172.915 67.355 173.085 ;
        RECT 65.855 172.225 66.025 172.915 ;
        RECT 67.715 172.745 67.885 173.525 ;
        RECT 68.690 173.395 68.860 173.525 ;
        RECT 66.195 172.575 67.885 172.745 ;
        RECT 68.055 172.965 68.520 173.355 ;
        RECT 68.690 173.225 69.085 173.395 ;
        RECT 66.195 172.395 66.365 172.575 ;
        RECT 62.995 171.685 64.065 171.855 ;
        RECT 64.235 171.475 64.425 171.915 ;
        RECT 64.595 171.645 65.545 171.925 ;
        RECT 65.855 171.835 66.115 172.225 ;
        RECT 66.535 172.155 67.325 172.405 ;
        RECT 65.765 171.665 66.115 171.835 ;
        RECT 66.325 171.475 66.655 171.935 ;
        RECT 67.530 171.865 67.700 172.575 ;
        RECT 68.055 172.375 68.225 172.965 ;
        RECT 67.870 172.155 68.225 172.375 ;
        RECT 68.395 172.155 68.745 172.775 ;
        RECT 68.915 171.865 69.085 173.225 ;
        RECT 69.450 173.055 69.775 173.840 ;
        RECT 69.255 172.005 69.715 173.055 ;
        RECT 67.530 171.695 68.385 171.865 ;
        RECT 68.590 171.695 69.085 171.865 ;
        RECT 69.255 171.475 69.585 171.835 ;
        RECT 69.945 171.735 70.115 173.855 ;
        RECT 70.285 173.525 70.615 174.025 ;
        RECT 70.785 173.355 71.040 173.855 ;
        RECT 70.290 173.185 71.040 173.355 ;
        RECT 70.290 172.195 70.520 173.185 ;
        RECT 71.270 173.155 71.555 174.025 ;
        RECT 71.725 173.395 71.985 173.855 ;
        RECT 72.160 173.565 72.415 174.025 ;
        RECT 72.585 173.395 72.845 173.855 ;
        RECT 71.725 173.225 72.845 173.395 ;
        RECT 73.015 173.225 73.325 174.025 ;
        RECT 70.690 172.365 71.040 173.015 ;
        RECT 71.725 172.975 71.985 173.225 ;
        RECT 73.495 173.055 73.805 173.855 ;
        RECT 75.270 173.345 75.525 173.715 ;
        RECT 75.185 173.175 75.525 173.345 ;
        RECT 75.705 173.225 75.990 174.025 ;
        RECT 76.170 173.305 76.500 173.815 ;
        RECT 71.230 172.805 71.985 172.975 ;
        RECT 72.775 172.885 73.805 173.055 ;
        RECT 71.230 172.295 71.635 172.805 ;
        RECT 72.775 172.635 72.945 172.885 ;
        RECT 71.805 172.465 72.945 172.635 ;
        RECT 70.290 172.025 71.040 172.195 ;
        RECT 71.230 172.125 72.880 172.295 ;
        RECT 73.115 172.145 73.465 172.715 ;
        RECT 70.285 171.475 70.615 171.855 ;
        RECT 70.785 171.735 71.040 172.025 ;
        RECT 71.275 171.475 71.555 171.955 ;
        RECT 71.725 171.735 71.985 172.125 ;
        RECT 72.160 171.475 72.415 171.955 ;
        RECT 72.585 171.735 72.880 172.125 ;
        RECT 73.635 171.975 73.805 172.885 ;
        RECT 73.060 171.475 73.335 171.955 ;
        RECT 73.505 171.645 73.805 171.975 ;
        RECT 75.270 173.045 75.525 173.175 ;
        RECT 75.270 172.185 75.450 173.045 ;
        RECT 76.170 172.715 76.420 173.305 ;
        RECT 76.770 173.155 76.940 173.765 ;
        RECT 77.110 173.335 77.440 174.025 ;
        RECT 77.670 173.475 77.910 173.765 ;
        RECT 78.110 173.645 78.530 174.025 ;
        RECT 78.710 173.555 79.340 173.805 ;
        RECT 79.810 173.645 80.140 174.025 ;
        RECT 78.710 173.475 78.880 173.555 ;
        RECT 80.310 173.475 80.480 173.765 ;
        RECT 80.660 173.645 81.040 174.025 ;
        RECT 81.280 173.640 82.110 173.810 ;
        RECT 77.670 173.305 78.880 173.475 ;
        RECT 75.620 172.385 76.420 172.715 ;
        RECT 75.270 171.655 75.525 172.185 ;
        RECT 75.705 171.475 75.990 171.935 ;
        RECT 76.170 171.735 76.420 172.385 ;
        RECT 76.620 173.135 76.940 173.155 ;
        RECT 76.620 172.965 78.540 173.135 ;
        RECT 76.620 172.070 76.810 172.965 ;
        RECT 78.710 172.795 78.880 173.305 ;
        RECT 79.050 173.045 79.570 173.355 ;
        RECT 76.980 172.625 78.880 172.795 ;
        RECT 76.980 172.565 77.310 172.625 ;
        RECT 77.460 172.395 77.790 172.455 ;
        RECT 77.130 172.125 77.790 172.395 ;
        RECT 76.620 171.740 76.940 172.070 ;
        RECT 77.120 171.475 77.780 171.955 ;
        RECT 77.980 171.865 78.150 172.625 ;
        RECT 79.050 172.455 79.230 172.865 ;
        RECT 78.320 172.285 78.650 172.405 ;
        RECT 79.400 172.285 79.570 173.045 ;
        RECT 78.320 172.115 79.570 172.285 ;
        RECT 79.740 173.225 81.110 173.475 ;
        RECT 79.740 172.455 79.930 173.225 ;
        RECT 80.860 172.965 81.110 173.225 ;
        RECT 80.100 172.795 80.350 172.955 ;
        RECT 81.280 172.795 81.450 173.640 ;
        RECT 82.345 173.355 82.515 173.855 ;
        RECT 82.685 173.525 83.015 174.025 ;
        RECT 81.620 172.965 82.120 173.345 ;
        RECT 82.345 173.185 83.040 173.355 ;
        RECT 80.100 172.625 81.450 172.795 ;
        RECT 81.030 172.585 81.450 172.625 ;
        RECT 79.740 172.115 80.160 172.455 ;
        RECT 80.450 172.125 80.860 172.455 ;
        RECT 77.980 171.695 78.830 171.865 ;
        RECT 79.390 171.475 79.710 171.935 ;
        RECT 79.910 171.685 80.160 172.115 ;
        RECT 80.450 171.475 80.860 171.915 ;
        RECT 81.030 171.855 81.200 172.585 ;
        RECT 81.370 172.035 81.720 172.405 ;
        RECT 81.900 172.095 82.120 172.965 ;
        RECT 82.290 172.395 82.700 173.015 ;
        RECT 82.870 172.215 83.040 173.185 ;
        RECT 82.345 172.025 83.040 172.215 ;
        RECT 81.030 171.655 82.045 171.855 ;
        RECT 82.345 171.695 82.515 172.025 ;
        RECT 82.685 171.475 83.015 171.855 ;
        RECT 83.230 171.735 83.455 173.855 ;
        RECT 83.625 173.525 83.955 174.025 ;
        RECT 84.125 173.355 84.295 173.855 ;
        RECT 83.630 173.185 84.295 173.355 ;
        RECT 83.630 172.195 83.860 173.185 ;
        RECT 84.645 173.095 84.815 173.855 ;
        RECT 85.030 173.265 85.360 174.025 ;
        RECT 84.030 172.365 84.380 173.015 ;
        RECT 84.645 172.925 85.360 173.095 ;
        RECT 85.530 172.950 85.785 173.855 ;
        RECT 84.555 172.375 84.910 172.745 ;
        RECT 85.190 172.715 85.360 172.925 ;
        RECT 85.190 172.385 85.445 172.715 ;
        RECT 85.190 172.195 85.360 172.385 ;
        RECT 85.615 172.220 85.785 172.950 ;
        RECT 85.960 172.875 86.220 174.025 ;
        RECT 87.315 172.860 87.605 174.025 ;
        RECT 88.150 173.045 88.405 173.715 ;
        RECT 88.585 173.225 88.870 174.025 ;
        RECT 89.050 173.305 89.380 173.815 ;
        RECT 83.630 172.025 84.295 172.195 ;
        RECT 83.625 171.475 83.955 171.855 ;
        RECT 84.125 171.735 84.295 172.025 ;
        RECT 84.645 172.025 85.360 172.195 ;
        RECT 84.645 171.645 84.815 172.025 ;
        RECT 85.030 171.475 85.360 171.855 ;
        RECT 85.530 171.645 85.785 172.220 ;
        RECT 85.960 171.475 86.220 172.315 ;
        RECT 87.315 171.475 87.605 172.200 ;
        RECT 88.150 172.185 88.330 173.045 ;
        RECT 89.050 172.715 89.300 173.305 ;
        RECT 89.650 173.155 89.820 173.765 ;
        RECT 89.990 173.335 90.320 174.025 ;
        RECT 90.550 173.475 90.790 173.765 ;
        RECT 90.990 173.645 91.410 174.025 ;
        RECT 91.590 173.555 92.220 173.805 ;
        RECT 92.690 173.645 93.020 174.025 ;
        RECT 91.590 173.475 91.760 173.555 ;
        RECT 93.190 173.475 93.360 173.765 ;
        RECT 93.540 173.645 93.920 174.025 ;
        RECT 94.160 173.640 94.990 173.810 ;
        RECT 90.550 173.305 91.760 173.475 ;
        RECT 88.500 172.385 89.300 172.715 ;
        RECT 88.150 171.985 88.405 172.185 ;
        RECT 88.065 171.815 88.405 171.985 ;
        RECT 88.150 171.655 88.405 171.815 ;
        RECT 88.585 171.475 88.870 171.935 ;
        RECT 89.050 171.735 89.300 172.385 ;
        RECT 89.500 173.135 89.820 173.155 ;
        RECT 89.500 172.965 91.420 173.135 ;
        RECT 89.500 172.070 89.690 172.965 ;
        RECT 91.590 172.795 91.760 173.305 ;
        RECT 91.930 173.045 92.450 173.355 ;
        RECT 89.860 172.625 91.760 172.795 ;
        RECT 89.860 172.565 90.190 172.625 ;
        RECT 90.340 172.395 90.670 172.455 ;
        RECT 90.010 172.125 90.670 172.395 ;
        RECT 89.500 171.740 89.820 172.070 ;
        RECT 90.000 171.475 90.660 171.955 ;
        RECT 90.860 171.865 91.030 172.625 ;
        RECT 91.930 172.455 92.110 172.865 ;
        RECT 91.200 172.285 91.530 172.405 ;
        RECT 92.280 172.285 92.450 173.045 ;
        RECT 91.200 172.115 92.450 172.285 ;
        RECT 92.620 173.225 93.990 173.475 ;
        RECT 92.620 172.455 92.810 173.225 ;
        RECT 93.740 172.965 93.990 173.225 ;
        RECT 92.980 172.795 93.230 172.955 ;
        RECT 94.160 172.795 94.330 173.640 ;
        RECT 95.225 173.355 95.395 173.855 ;
        RECT 95.565 173.525 95.895 174.025 ;
        RECT 94.500 172.965 95.000 173.345 ;
        RECT 95.225 173.185 95.920 173.355 ;
        RECT 92.980 172.625 94.330 172.795 ;
        RECT 93.910 172.585 94.330 172.625 ;
        RECT 92.620 172.115 93.040 172.455 ;
        RECT 93.330 172.125 93.740 172.455 ;
        RECT 90.860 171.695 91.710 171.865 ;
        RECT 92.270 171.475 92.590 171.935 ;
        RECT 92.790 171.685 93.040 172.115 ;
        RECT 93.330 171.475 93.740 171.915 ;
        RECT 93.910 171.855 94.080 172.585 ;
        RECT 94.250 172.035 94.600 172.405 ;
        RECT 94.780 172.095 95.000 172.965 ;
        RECT 95.170 172.395 95.580 173.015 ;
        RECT 95.750 172.215 95.920 173.185 ;
        RECT 95.225 172.025 95.920 172.215 ;
        RECT 93.910 171.655 94.925 171.855 ;
        RECT 95.225 171.695 95.395 172.025 ;
        RECT 95.565 171.475 95.895 171.855 ;
        RECT 96.110 171.735 96.335 173.855 ;
        RECT 96.505 173.525 96.835 174.025 ;
        RECT 97.005 173.355 97.175 173.855 ;
        RECT 96.510 173.185 97.175 173.355 ;
        RECT 97.435 173.265 97.950 173.675 ;
        RECT 98.185 173.265 98.355 174.025 ;
        RECT 98.525 173.685 100.555 173.855 ;
        RECT 96.510 172.195 96.740 173.185 ;
        RECT 96.910 172.365 97.260 173.015 ;
        RECT 97.435 172.455 97.775 173.265 ;
        RECT 98.525 173.020 98.695 173.685 ;
        RECT 99.090 173.345 100.215 173.515 ;
        RECT 97.945 172.830 98.695 173.020 ;
        RECT 98.865 173.005 99.875 173.175 ;
        RECT 97.435 172.285 98.665 172.455 ;
        RECT 96.510 172.025 97.175 172.195 ;
        RECT 96.505 171.475 96.835 171.855 ;
        RECT 97.005 171.735 97.175 172.025 ;
        RECT 97.710 171.680 97.955 172.285 ;
        RECT 98.175 171.475 98.685 172.010 ;
        RECT 98.865 171.645 99.055 173.005 ;
        RECT 99.225 171.985 99.500 172.805 ;
        RECT 99.705 172.205 99.875 173.005 ;
        RECT 100.045 172.215 100.215 173.345 ;
        RECT 100.385 172.715 100.555 173.685 ;
        RECT 100.725 172.885 100.895 174.025 ;
        RECT 101.065 172.885 101.400 173.855 ;
        RECT 100.385 172.385 100.580 172.715 ;
        RECT 100.805 172.385 101.060 172.715 ;
        RECT 100.805 172.215 100.975 172.385 ;
        RECT 101.230 172.215 101.400 172.885 ;
        RECT 100.045 172.045 100.975 172.215 ;
        RECT 100.045 172.010 100.220 172.045 ;
        RECT 99.225 171.815 99.505 171.985 ;
        RECT 99.225 171.645 99.500 171.815 ;
        RECT 99.690 171.645 100.220 172.010 ;
        RECT 100.645 171.475 100.975 171.875 ;
        RECT 101.145 171.645 101.400 172.215 ;
        RECT 101.580 172.835 101.835 173.715 ;
        RECT 102.005 172.885 102.310 174.025 ;
        RECT 102.650 173.645 102.980 174.025 ;
        RECT 103.160 173.475 103.330 173.765 ;
        RECT 103.500 173.565 103.750 174.025 ;
        RECT 102.530 173.305 103.330 173.475 ;
        RECT 103.920 173.515 104.790 173.855 ;
        RECT 101.580 172.185 101.790 172.835 ;
        RECT 102.530 172.715 102.700 173.305 ;
        RECT 103.920 173.135 104.090 173.515 ;
        RECT 105.025 173.395 105.195 173.855 ;
        RECT 105.365 173.565 105.735 174.025 ;
        RECT 106.030 173.425 106.200 173.765 ;
        RECT 106.370 173.595 106.700 174.025 ;
        RECT 106.935 173.425 107.105 173.765 ;
        RECT 102.870 172.965 104.090 173.135 ;
        RECT 104.260 173.055 104.720 173.345 ;
        RECT 105.025 173.225 105.585 173.395 ;
        RECT 106.030 173.255 107.105 173.425 ;
        RECT 107.275 173.525 107.955 173.855 ;
        RECT 108.170 173.525 108.420 173.855 ;
        RECT 108.590 173.565 108.840 174.025 ;
        RECT 105.415 173.085 105.585 173.225 ;
        RECT 104.260 173.045 105.225 173.055 ;
        RECT 103.920 172.875 104.090 172.965 ;
        RECT 104.550 172.885 105.225 173.045 ;
        RECT 101.960 172.685 102.700 172.715 ;
        RECT 101.960 172.385 102.875 172.685 ;
        RECT 102.550 172.210 102.875 172.385 ;
        RECT 101.580 171.655 101.835 172.185 ;
        RECT 102.005 171.475 102.310 171.935 ;
        RECT 102.555 171.855 102.875 172.210 ;
        RECT 103.045 172.425 103.585 172.795 ;
        RECT 103.920 172.705 104.325 172.875 ;
        RECT 103.045 172.025 103.285 172.425 ;
        RECT 103.765 172.255 103.985 172.535 ;
        RECT 103.455 172.085 103.985 172.255 ;
        RECT 103.455 171.855 103.625 172.085 ;
        RECT 104.155 171.925 104.325 172.705 ;
        RECT 104.495 172.095 104.845 172.715 ;
        RECT 105.015 172.095 105.225 172.885 ;
        RECT 105.415 172.915 106.915 173.085 ;
        RECT 105.415 172.225 105.585 172.915 ;
        RECT 107.275 172.745 107.445 173.525 ;
        RECT 108.250 173.395 108.420 173.525 ;
        RECT 105.755 172.575 107.445 172.745 ;
        RECT 107.615 172.965 108.080 173.355 ;
        RECT 108.250 173.225 108.645 173.395 ;
        RECT 105.755 172.395 105.925 172.575 ;
        RECT 102.555 171.685 103.625 171.855 ;
        RECT 103.795 171.475 103.985 171.915 ;
        RECT 104.155 171.645 105.105 171.925 ;
        RECT 105.415 171.835 105.675 172.225 ;
        RECT 106.095 172.155 106.885 172.405 ;
        RECT 105.325 171.665 105.675 171.835 ;
        RECT 105.885 171.475 106.215 171.935 ;
        RECT 107.090 171.865 107.260 172.575 ;
        RECT 107.615 172.375 107.785 172.965 ;
        RECT 107.430 172.155 107.785 172.375 ;
        RECT 107.955 172.155 108.305 172.775 ;
        RECT 108.475 171.865 108.645 173.225 ;
        RECT 109.010 173.055 109.335 173.840 ;
        RECT 108.815 172.005 109.275 173.055 ;
        RECT 107.090 171.695 107.945 171.865 ;
        RECT 108.150 171.695 108.645 171.865 ;
        RECT 108.815 171.475 109.145 171.835 ;
        RECT 109.505 171.735 109.675 173.855 ;
        RECT 109.845 173.525 110.175 174.025 ;
        RECT 110.345 173.355 110.600 173.855 ;
        RECT 109.850 173.185 110.600 173.355 ;
        RECT 109.850 172.195 110.080 173.185 ;
        RECT 110.250 172.365 110.600 173.015 ;
        RECT 110.835 172.885 111.045 174.025 ;
        RECT 111.215 172.875 111.545 173.855 ;
        RECT 111.715 172.885 111.945 174.025 ;
        RECT 112.155 172.935 113.365 174.025 ;
        RECT 109.850 172.025 110.600 172.195 ;
        RECT 109.845 171.475 110.175 171.855 ;
        RECT 110.345 171.735 110.600 172.025 ;
        RECT 110.835 171.475 111.045 172.295 ;
        RECT 111.215 172.275 111.465 172.875 ;
        RECT 111.635 172.465 111.965 172.715 ;
        RECT 112.155 172.395 112.675 172.935 ;
        RECT 111.215 171.645 111.545 172.275 ;
        RECT 111.715 171.475 111.945 172.295 ;
        RECT 112.845 172.225 113.365 172.765 ;
        RECT 112.155 171.475 113.365 172.225 ;
        RECT 26.970 171.305 113.450 171.475 ;
        RECT 27.055 170.555 28.265 171.305 ;
        RECT 28.525 170.755 28.695 171.045 ;
        RECT 28.865 170.925 29.195 171.305 ;
        RECT 28.525 170.585 29.190 170.755 ;
        RECT 27.055 170.015 27.575 170.555 ;
        RECT 27.745 169.845 28.265 170.385 ;
        RECT 27.055 168.755 28.265 169.845 ;
        RECT 28.440 169.765 28.790 170.415 ;
        RECT 28.960 169.595 29.190 170.585 ;
        RECT 28.525 169.425 29.190 169.595 ;
        RECT 28.525 168.925 28.695 169.425 ;
        RECT 28.865 168.755 29.195 169.255 ;
        RECT 29.365 168.925 29.590 171.045 ;
        RECT 29.805 170.925 30.135 171.305 ;
        RECT 30.305 170.755 30.475 171.085 ;
        RECT 30.775 170.925 31.790 171.125 ;
        RECT 29.780 170.565 30.475 170.755 ;
        RECT 29.780 169.595 29.950 170.565 ;
        RECT 30.120 169.765 30.530 170.385 ;
        RECT 30.700 169.815 30.920 170.685 ;
        RECT 31.100 170.375 31.450 170.745 ;
        RECT 31.620 170.195 31.790 170.925 ;
        RECT 31.960 170.865 32.370 171.305 ;
        RECT 32.660 170.665 32.910 171.095 ;
        RECT 33.110 170.845 33.430 171.305 ;
        RECT 33.990 170.915 34.840 171.085 ;
        RECT 31.960 170.325 32.370 170.655 ;
        RECT 32.660 170.325 33.080 170.665 ;
        RECT 31.370 170.155 31.790 170.195 ;
        RECT 31.370 169.985 32.720 170.155 ;
        RECT 29.780 169.425 30.475 169.595 ;
        RECT 30.700 169.435 31.200 169.815 ;
        RECT 29.805 168.755 30.135 169.255 ;
        RECT 30.305 168.925 30.475 169.425 ;
        RECT 31.370 169.140 31.540 169.985 ;
        RECT 32.470 169.825 32.720 169.985 ;
        RECT 31.710 169.555 31.960 169.815 ;
        RECT 32.890 169.555 33.080 170.325 ;
        RECT 31.710 169.305 33.080 169.555 ;
        RECT 33.250 170.495 34.500 170.665 ;
        RECT 33.250 169.735 33.420 170.495 ;
        RECT 34.170 170.375 34.500 170.495 ;
        RECT 33.590 169.915 33.770 170.325 ;
        RECT 34.670 170.155 34.840 170.915 ;
        RECT 35.040 170.825 35.700 171.305 ;
        RECT 35.880 170.710 36.200 171.040 ;
        RECT 35.030 170.385 35.690 170.655 ;
        RECT 35.030 170.325 35.360 170.385 ;
        RECT 35.510 170.155 35.840 170.215 ;
        RECT 33.940 169.985 35.840 170.155 ;
        RECT 33.250 169.425 33.770 169.735 ;
        RECT 33.940 169.475 34.110 169.985 ;
        RECT 36.010 169.815 36.200 170.710 ;
        RECT 34.280 169.645 36.200 169.815 ;
        RECT 35.880 169.625 36.200 169.645 ;
        RECT 36.400 170.395 36.650 171.045 ;
        RECT 36.830 170.845 37.115 171.305 ;
        RECT 37.295 170.965 37.550 171.125 ;
        RECT 37.295 170.795 37.635 170.965 ;
        RECT 38.185 170.825 38.485 171.305 ;
        RECT 37.295 170.595 37.550 170.795 ;
        RECT 38.655 170.655 38.915 171.110 ;
        RECT 39.085 170.825 39.345 171.305 ;
        RECT 39.525 170.655 39.785 171.110 ;
        RECT 39.955 170.825 40.205 171.305 ;
        RECT 40.385 170.655 40.645 171.110 ;
        RECT 40.815 170.825 41.065 171.305 ;
        RECT 41.245 170.655 41.505 171.110 ;
        RECT 41.675 170.825 41.920 171.305 ;
        RECT 42.090 170.655 42.365 171.110 ;
        RECT 42.535 170.825 42.780 171.305 ;
        RECT 42.950 170.655 43.210 171.110 ;
        RECT 43.380 170.825 43.640 171.305 ;
        RECT 43.810 170.655 44.070 171.110 ;
        RECT 44.240 170.825 44.500 171.305 ;
        RECT 44.670 170.655 44.930 171.110 ;
        RECT 45.100 170.745 45.360 171.305 ;
        RECT 36.400 170.065 37.200 170.395 ;
        RECT 33.940 169.305 35.150 169.475 ;
        RECT 30.710 168.970 31.540 169.140 ;
        RECT 31.780 168.755 32.160 169.135 ;
        RECT 32.340 169.015 32.510 169.305 ;
        RECT 33.940 169.225 34.110 169.305 ;
        RECT 32.680 168.755 33.010 169.135 ;
        RECT 33.480 168.975 34.110 169.225 ;
        RECT 34.290 168.755 34.710 169.135 ;
        RECT 34.910 169.015 35.150 169.305 ;
        RECT 35.380 168.755 35.710 169.445 ;
        RECT 35.880 169.015 36.050 169.625 ;
        RECT 36.400 169.475 36.650 170.065 ;
        RECT 37.370 169.735 37.550 170.595 ;
        RECT 36.320 168.965 36.650 169.475 ;
        RECT 36.830 168.755 37.115 169.555 ;
        RECT 37.295 169.065 37.550 169.735 ;
        RECT 38.185 170.485 44.930 170.655 ;
        RECT 38.185 169.895 39.350 170.485 ;
        RECT 45.530 170.315 45.780 171.125 ;
        RECT 45.960 170.780 46.220 171.305 ;
        RECT 46.390 170.315 46.640 171.125 ;
        RECT 46.820 170.795 47.125 171.305 ;
        RECT 47.385 170.755 47.555 171.135 ;
        RECT 47.735 170.925 48.065 171.305 ;
        RECT 39.520 170.065 46.640 170.315 ;
        RECT 46.810 170.065 47.125 170.625 ;
        RECT 47.385 170.585 48.050 170.755 ;
        RECT 48.245 170.630 48.505 171.135 ;
        RECT 38.185 169.670 44.930 169.895 ;
        RECT 38.185 168.755 38.455 169.500 ;
        RECT 38.625 168.930 38.915 169.670 ;
        RECT 39.525 169.655 44.930 169.670 ;
        RECT 39.085 168.760 39.340 169.485 ;
        RECT 39.525 168.930 39.785 169.655 ;
        RECT 39.955 168.760 40.200 169.485 ;
        RECT 40.385 168.930 40.645 169.655 ;
        RECT 40.815 168.760 41.060 169.485 ;
        RECT 41.245 168.930 41.505 169.655 ;
        RECT 41.675 168.760 41.920 169.485 ;
        RECT 42.090 168.930 42.350 169.655 ;
        RECT 42.520 168.760 42.780 169.485 ;
        RECT 42.950 168.930 43.210 169.655 ;
        RECT 43.380 168.760 43.640 169.485 ;
        RECT 43.810 168.930 44.070 169.655 ;
        RECT 44.240 168.760 44.500 169.485 ;
        RECT 44.670 168.930 44.930 169.655 ;
        RECT 45.100 168.760 45.360 169.555 ;
        RECT 45.530 168.930 45.780 170.065 ;
        RECT 39.085 168.755 45.360 168.760 ;
        RECT 45.960 168.755 46.220 169.565 ;
        RECT 46.395 168.925 46.640 170.065 ;
        RECT 47.315 170.035 47.645 170.405 ;
        RECT 47.880 170.330 48.050 170.585 ;
        RECT 47.880 170.000 48.165 170.330 ;
        RECT 47.880 169.855 48.050 170.000 ;
        RECT 47.385 169.685 48.050 169.855 ;
        RECT 48.335 169.830 48.505 170.630 ;
        RECT 48.675 170.580 48.965 171.305 ;
        RECT 49.140 170.565 49.395 171.135 ;
        RECT 49.565 170.905 49.895 171.305 ;
        RECT 50.320 170.770 50.850 171.135 ;
        RECT 50.320 170.735 50.495 170.770 ;
        RECT 49.565 170.565 50.495 170.735 ;
        RECT 51.040 170.625 51.315 171.135 ;
        RECT 46.820 168.755 47.115 169.565 ;
        RECT 47.385 168.925 47.555 169.685 ;
        RECT 47.735 168.755 48.065 169.515 ;
        RECT 48.235 168.925 48.505 169.830 ;
        RECT 48.675 168.755 48.965 169.920 ;
        RECT 49.140 169.895 49.310 170.565 ;
        RECT 49.565 170.395 49.735 170.565 ;
        RECT 49.480 170.065 49.735 170.395 ;
        RECT 49.960 170.065 50.155 170.395 ;
        RECT 49.140 168.925 49.475 169.895 ;
        RECT 49.645 168.755 49.815 169.895 ;
        RECT 49.985 169.095 50.155 170.065 ;
        RECT 50.325 169.435 50.495 170.565 ;
        RECT 50.665 169.775 50.835 170.575 ;
        RECT 51.035 170.455 51.315 170.625 ;
        RECT 51.040 169.975 51.315 170.455 ;
        RECT 51.485 169.775 51.675 171.135 ;
        RECT 51.855 170.770 52.365 171.305 ;
        RECT 52.585 170.495 52.830 171.100 ;
        RECT 53.280 170.565 53.535 171.135 ;
        RECT 53.705 170.905 54.035 171.305 ;
        RECT 54.460 170.770 54.990 171.135 ;
        RECT 55.180 170.965 55.455 171.135 ;
        RECT 55.175 170.795 55.455 170.965 ;
        RECT 54.460 170.735 54.635 170.770 ;
        RECT 53.705 170.565 54.635 170.735 ;
        RECT 51.875 170.325 53.105 170.495 ;
        RECT 50.665 169.605 51.675 169.775 ;
        RECT 51.845 169.760 52.595 169.950 ;
        RECT 50.325 169.265 51.450 169.435 ;
        RECT 51.845 169.095 52.015 169.760 ;
        RECT 52.765 169.515 53.105 170.325 ;
        RECT 49.985 168.925 52.015 169.095 ;
        RECT 52.185 168.755 52.355 169.515 ;
        RECT 52.590 169.105 53.105 169.515 ;
        RECT 53.280 169.895 53.450 170.565 ;
        RECT 53.705 170.395 53.875 170.565 ;
        RECT 53.620 170.065 53.875 170.395 ;
        RECT 54.100 170.065 54.295 170.395 ;
        RECT 53.280 168.925 53.615 169.895 ;
        RECT 53.785 168.755 53.955 169.895 ;
        RECT 54.125 169.095 54.295 170.065 ;
        RECT 54.465 169.435 54.635 170.565 ;
        RECT 54.805 169.775 54.975 170.575 ;
        RECT 55.180 169.975 55.455 170.795 ;
        RECT 55.625 169.775 55.815 171.135 ;
        RECT 55.995 170.770 56.505 171.305 ;
        RECT 56.725 170.495 56.970 171.100 ;
        RECT 57.420 170.565 57.675 171.135 ;
        RECT 57.845 170.905 58.175 171.305 ;
        RECT 58.600 170.770 59.130 171.135 ;
        RECT 58.600 170.735 58.775 170.770 ;
        RECT 57.845 170.565 58.775 170.735 ;
        RECT 59.320 170.625 59.595 171.135 ;
        RECT 56.015 170.325 57.245 170.495 ;
        RECT 54.805 169.605 55.815 169.775 ;
        RECT 55.985 169.760 56.735 169.950 ;
        RECT 54.465 169.265 55.590 169.435 ;
        RECT 55.985 169.095 56.155 169.760 ;
        RECT 56.905 169.515 57.245 170.325 ;
        RECT 54.125 168.925 56.155 169.095 ;
        RECT 56.325 168.755 56.495 169.515 ;
        RECT 56.730 169.105 57.245 169.515 ;
        RECT 57.420 169.895 57.590 170.565 ;
        RECT 57.845 170.395 58.015 170.565 ;
        RECT 57.760 170.065 58.015 170.395 ;
        RECT 58.240 170.065 58.435 170.395 ;
        RECT 57.420 168.925 57.755 169.895 ;
        RECT 57.925 168.755 58.095 169.895 ;
        RECT 58.265 169.095 58.435 170.065 ;
        RECT 58.605 169.435 58.775 170.565 ;
        RECT 58.945 169.775 59.115 170.575 ;
        RECT 59.315 170.455 59.595 170.625 ;
        RECT 59.320 169.975 59.595 170.455 ;
        RECT 59.765 169.775 59.955 171.135 ;
        RECT 60.135 170.770 60.645 171.305 ;
        RECT 60.865 170.495 61.110 171.100 ;
        RECT 61.830 170.495 62.075 171.100 ;
        RECT 62.295 170.770 62.805 171.305 ;
        RECT 60.155 170.325 61.385 170.495 ;
        RECT 58.945 169.605 59.955 169.775 ;
        RECT 60.125 169.760 60.875 169.950 ;
        RECT 58.605 169.265 59.730 169.435 ;
        RECT 60.125 169.095 60.295 169.760 ;
        RECT 61.045 169.515 61.385 170.325 ;
        RECT 58.265 168.925 60.295 169.095 ;
        RECT 60.465 168.755 60.635 169.515 ;
        RECT 60.870 169.105 61.385 169.515 ;
        RECT 61.555 170.325 62.785 170.495 ;
        RECT 61.555 169.515 61.895 170.325 ;
        RECT 62.065 169.760 62.815 169.950 ;
        RECT 61.555 169.105 62.070 169.515 ;
        RECT 62.305 168.755 62.475 169.515 ;
        RECT 62.645 169.095 62.815 169.760 ;
        RECT 62.985 169.775 63.175 171.135 ;
        RECT 63.345 170.965 63.620 171.135 ;
        RECT 63.345 170.795 63.625 170.965 ;
        RECT 63.345 169.975 63.620 170.795 ;
        RECT 63.810 170.770 64.340 171.135 ;
        RECT 64.765 170.905 65.095 171.305 ;
        RECT 64.165 170.735 64.340 170.770 ;
        RECT 63.825 169.775 63.995 170.575 ;
        RECT 62.985 169.605 63.995 169.775 ;
        RECT 64.165 170.565 65.095 170.735 ;
        RECT 65.265 170.565 65.520 171.135 ;
        RECT 64.165 169.435 64.335 170.565 ;
        RECT 64.925 170.395 65.095 170.565 ;
        RECT 63.210 169.265 64.335 169.435 ;
        RECT 64.505 170.065 64.700 170.395 ;
        RECT 64.925 170.065 65.180 170.395 ;
        RECT 64.505 169.095 64.675 170.065 ;
        RECT 65.350 169.895 65.520 170.565 ;
        RECT 62.645 168.925 64.675 169.095 ;
        RECT 64.845 168.755 65.015 169.895 ;
        RECT 65.185 168.925 65.520 169.895 ;
        RECT 65.695 170.565 66.080 171.135 ;
        RECT 66.250 170.845 66.575 171.305 ;
        RECT 67.095 170.675 67.375 171.135 ;
        RECT 65.695 169.895 65.975 170.565 ;
        RECT 66.250 170.505 67.375 170.675 ;
        RECT 66.250 170.395 66.700 170.505 ;
        RECT 66.145 170.065 66.700 170.395 ;
        RECT 67.565 170.335 67.965 171.135 ;
        RECT 68.365 170.845 68.635 171.305 ;
        RECT 68.805 170.675 69.090 171.135 ;
        RECT 65.695 168.925 66.080 169.895 ;
        RECT 66.250 169.605 66.700 170.065 ;
        RECT 66.870 169.775 67.965 170.335 ;
        RECT 66.250 169.385 67.375 169.605 ;
        RECT 66.250 168.755 66.575 169.215 ;
        RECT 67.095 168.925 67.375 169.385 ;
        RECT 67.565 168.925 67.965 169.775 ;
        RECT 68.135 170.505 69.090 170.675 ;
        RECT 69.525 170.505 69.855 171.305 ;
        RECT 70.025 170.655 70.195 171.135 ;
        RECT 70.365 170.825 70.695 171.305 ;
        RECT 70.865 170.655 71.035 171.135 ;
        RECT 71.285 170.825 71.525 171.305 ;
        RECT 71.705 170.655 71.875 171.135 ;
        RECT 68.135 169.605 68.345 170.505 ;
        RECT 70.025 170.485 71.035 170.655 ;
        RECT 71.240 170.485 71.875 170.655 ;
        RECT 68.515 169.775 69.205 170.335 ;
        RECT 70.025 170.285 70.520 170.485 ;
        RECT 71.240 170.315 71.410 170.485 ;
        RECT 72.140 170.465 72.400 171.305 ;
        RECT 72.575 170.560 72.830 171.135 ;
        RECT 73.000 170.925 73.330 171.305 ;
        RECT 73.545 170.755 73.715 171.135 ;
        RECT 73.000 170.585 73.715 170.755 ;
        RECT 70.025 170.115 70.525 170.285 ;
        RECT 70.910 170.145 71.410 170.315 ;
        RECT 70.025 169.945 70.520 170.115 ;
        RECT 68.135 169.385 69.090 169.605 ;
        RECT 68.365 168.755 68.635 169.215 ;
        RECT 68.805 168.925 69.090 169.385 ;
        RECT 69.525 168.755 69.855 169.905 ;
        RECT 70.025 169.775 71.035 169.945 ;
        RECT 70.025 168.925 70.195 169.775 ;
        RECT 70.365 168.755 70.695 169.555 ;
        RECT 70.865 168.925 71.035 169.775 ;
        RECT 71.240 169.905 71.410 170.145 ;
        RECT 71.580 170.075 71.960 170.315 ;
        RECT 71.240 169.735 71.955 169.905 ;
        RECT 71.215 168.755 71.455 169.555 ;
        RECT 71.625 168.925 71.955 169.735 ;
        RECT 72.140 168.755 72.400 169.905 ;
        RECT 72.575 169.830 72.745 170.560 ;
        RECT 73.000 170.395 73.170 170.585 ;
        RECT 74.435 170.580 74.725 171.305 ;
        RECT 74.895 170.630 75.155 171.135 ;
        RECT 75.335 170.925 75.665 171.305 ;
        RECT 75.845 170.755 76.015 171.135 ;
        RECT 72.915 170.065 73.170 170.395 ;
        RECT 73.000 169.855 73.170 170.065 ;
        RECT 73.450 170.035 73.805 170.405 ;
        RECT 72.575 168.925 72.830 169.830 ;
        RECT 73.000 169.685 73.715 169.855 ;
        RECT 73.000 168.755 73.330 169.515 ;
        RECT 73.545 168.925 73.715 169.685 ;
        RECT 74.435 168.755 74.725 169.920 ;
        RECT 74.895 169.830 75.065 170.630 ;
        RECT 75.350 170.585 76.015 170.755 ;
        RECT 75.350 170.330 75.520 170.585 ;
        RECT 76.550 170.495 76.795 171.100 ;
        RECT 77.015 170.770 77.525 171.305 ;
        RECT 75.235 170.000 75.520 170.330 ;
        RECT 75.755 170.035 76.085 170.405 ;
        RECT 76.275 170.325 77.505 170.495 ;
        RECT 75.350 169.855 75.520 170.000 ;
        RECT 74.895 168.925 75.165 169.830 ;
        RECT 75.350 169.685 76.015 169.855 ;
        RECT 75.335 168.755 75.665 169.515 ;
        RECT 75.845 168.925 76.015 169.685 ;
        RECT 76.275 169.515 76.615 170.325 ;
        RECT 76.785 169.760 77.535 169.950 ;
        RECT 76.275 169.105 76.790 169.515 ;
        RECT 77.025 168.755 77.195 169.515 ;
        RECT 77.365 169.095 77.535 169.760 ;
        RECT 77.705 169.775 77.895 171.135 ;
        RECT 78.065 170.285 78.340 171.135 ;
        RECT 78.530 170.770 79.060 171.135 ;
        RECT 79.485 170.905 79.815 171.305 ;
        RECT 78.885 170.735 79.060 170.770 ;
        RECT 78.065 170.115 78.345 170.285 ;
        RECT 78.065 169.975 78.340 170.115 ;
        RECT 78.545 169.775 78.715 170.575 ;
        RECT 77.705 169.605 78.715 169.775 ;
        RECT 78.885 170.565 79.815 170.735 ;
        RECT 79.985 170.565 80.240 171.135 ;
        RECT 78.885 169.435 79.055 170.565 ;
        RECT 79.645 170.395 79.815 170.565 ;
        RECT 77.930 169.265 79.055 169.435 ;
        RECT 79.225 170.065 79.420 170.395 ;
        RECT 79.645 170.065 79.900 170.395 ;
        RECT 79.225 169.095 79.395 170.065 ;
        RECT 80.070 169.895 80.240 170.565 ;
        RECT 80.475 170.485 80.685 171.305 ;
        RECT 80.855 170.505 81.185 171.135 ;
        RECT 80.855 169.905 81.105 170.505 ;
        RECT 81.355 170.485 81.585 171.305 ;
        RECT 82.170 170.595 82.425 171.125 ;
        RECT 82.605 170.845 82.890 171.305 ;
        RECT 81.275 170.065 81.605 170.315 ;
        RECT 77.365 168.925 79.395 169.095 ;
        RECT 79.565 168.755 79.735 169.895 ;
        RECT 79.905 168.925 80.240 169.895 ;
        RECT 80.475 168.755 80.685 169.895 ;
        RECT 80.855 168.925 81.185 169.905 ;
        RECT 81.355 168.755 81.585 169.895 ;
        RECT 82.170 169.735 82.350 170.595 ;
        RECT 83.070 170.395 83.320 171.045 ;
        RECT 82.520 170.065 83.320 170.395 ;
        RECT 82.170 169.605 82.425 169.735 ;
        RECT 82.085 169.435 82.425 169.605 ;
        RECT 82.170 169.065 82.425 169.435 ;
        RECT 82.605 168.755 82.890 169.555 ;
        RECT 83.070 169.475 83.320 170.065 ;
        RECT 83.520 170.710 83.840 171.040 ;
        RECT 84.020 170.825 84.680 171.305 ;
        RECT 84.880 170.915 85.730 171.085 ;
        RECT 83.520 169.815 83.710 170.710 ;
        RECT 84.030 170.385 84.690 170.655 ;
        RECT 84.360 170.325 84.690 170.385 ;
        RECT 83.880 170.155 84.210 170.215 ;
        RECT 84.880 170.155 85.050 170.915 ;
        RECT 86.290 170.845 86.610 171.305 ;
        RECT 86.810 170.665 87.060 171.095 ;
        RECT 87.350 170.865 87.760 171.305 ;
        RECT 87.930 170.925 88.945 171.125 ;
        RECT 85.220 170.495 86.470 170.665 ;
        RECT 85.220 170.375 85.550 170.495 ;
        RECT 83.880 169.985 85.780 170.155 ;
        RECT 83.520 169.645 85.440 169.815 ;
        RECT 83.520 169.625 83.840 169.645 ;
        RECT 83.070 168.965 83.400 169.475 ;
        RECT 83.670 169.015 83.840 169.625 ;
        RECT 85.610 169.475 85.780 169.985 ;
        RECT 85.950 169.915 86.130 170.325 ;
        RECT 86.300 169.735 86.470 170.495 ;
        RECT 84.010 168.755 84.340 169.445 ;
        RECT 84.570 169.305 85.780 169.475 ;
        RECT 85.950 169.425 86.470 169.735 ;
        RECT 86.640 170.325 87.060 170.665 ;
        RECT 87.350 170.325 87.760 170.655 ;
        RECT 86.640 169.555 86.830 170.325 ;
        RECT 87.930 170.195 88.100 170.925 ;
        RECT 89.245 170.755 89.415 171.085 ;
        RECT 89.585 170.925 89.915 171.305 ;
        RECT 88.270 170.375 88.620 170.745 ;
        RECT 87.930 170.155 88.350 170.195 ;
        RECT 87.000 169.985 88.350 170.155 ;
        RECT 87.000 169.825 87.250 169.985 ;
        RECT 87.760 169.555 88.010 169.815 ;
        RECT 86.640 169.305 88.010 169.555 ;
        RECT 84.570 169.015 84.810 169.305 ;
        RECT 85.610 169.225 85.780 169.305 ;
        RECT 85.010 168.755 85.430 169.135 ;
        RECT 85.610 168.975 86.240 169.225 ;
        RECT 86.710 168.755 87.040 169.135 ;
        RECT 87.210 169.015 87.380 169.305 ;
        RECT 88.180 169.140 88.350 169.985 ;
        RECT 88.800 169.815 89.020 170.685 ;
        RECT 89.245 170.565 89.940 170.755 ;
        RECT 88.520 169.435 89.020 169.815 ;
        RECT 89.190 169.765 89.600 170.385 ;
        RECT 89.770 169.595 89.940 170.565 ;
        RECT 89.245 169.425 89.940 169.595 ;
        RECT 87.560 168.755 87.940 169.135 ;
        RECT 88.180 168.970 89.010 169.140 ;
        RECT 89.245 168.925 89.415 169.425 ;
        RECT 89.585 168.755 89.915 169.255 ;
        RECT 90.130 168.925 90.355 171.045 ;
        RECT 90.525 170.925 90.855 171.305 ;
        RECT 91.025 170.755 91.195 171.045 ;
        RECT 90.530 170.585 91.195 170.755 ;
        RECT 90.530 169.595 90.760 170.585 ;
        RECT 91.730 170.495 91.975 171.100 ;
        RECT 92.195 170.770 92.705 171.305 ;
        RECT 90.930 169.765 91.280 170.415 ;
        RECT 91.455 170.325 92.685 170.495 ;
        RECT 90.530 169.425 91.195 169.595 ;
        RECT 90.525 168.755 90.855 169.255 ;
        RECT 91.025 168.925 91.195 169.425 ;
        RECT 91.455 169.515 91.795 170.325 ;
        RECT 91.965 169.760 92.715 169.950 ;
        RECT 91.455 169.105 91.970 169.515 ;
        RECT 92.205 168.755 92.375 169.515 ;
        RECT 92.545 169.095 92.715 169.760 ;
        RECT 92.885 169.775 93.075 171.135 ;
        RECT 93.245 170.625 93.520 171.135 ;
        RECT 93.710 170.770 94.240 171.135 ;
        RECT 94.665 170.905 94.995 171.305 ;
        RECT 94.065 170.735 94.240 170.770 ;
        RECT 93.245 170.455 93.525 170.625 ;
        RECT 93.245 169.975 93.520 170.455 ;
        RECT 93.725 169.775 93.895 170.575 ;
        RECT 92.885 169.605 93.895 169.775 ;
        RECT 94.065 170.565 94.995 170.735 ;
        RECT 95.165 170.565 95.420 171.135 ;
        RECT 94.065 169.435 94.235 170.565 ;
        RECT 94.825 170.395 94.995 170.565 ;
        RECT 93.110 169.265 94.235 169.435 ;
        RECT 94.405 170.065 94.600 170.395 ;
        RECT 94.825 170.065 95.080 170.395 ;
        RECT 94.405 169.095 94.575 170.065 ;
        RECT 95.250 169.895 95.420 170.565 ;
        RECT 92.545 168.925 94.575 169.095 ;
        RECT 94.745 168.755 94.915 169.895 ;
        RECT 95.085 168.925 95.420 169.895 ;
        RECT 96.515 170.505 96.855 171.135 ;
        RECT 97.025 170.505 97.275 171.305 ;
        RECT 97.465 170.655 97.795 171.135 ;
        RECT 97.965 170.845 98.190 171.305 ;
        RECT 98.360 170.655 98.690 171.135 ;
        RECT 96.515 169.895 96.690 170.505 ;
        RECT 97.465 170.485 98.690 170.655 ;
        RECT 99.320 170.525 99.820 171.135 ;
        RECT 100.195 170.580 100.485 171.305 ;
        RECT 96.860 170.145 97.555 170.315 ;
        RECT 97.385 169.895 97.555 170.145 ;
        RECT 97.730 170.115 98.150 170.315 ;
        RECT 98.320 170.115 98.650 170.315 ;
        RECT 98.820 170.115 99.150 170.315 ;
        RECT 99.320 169.895 99.490 170.525 ;
        RECT 100.655 170.505 100.995 171.135 ;
        RECT 101.165 170.505 101.415 171.305 ;
        RECT 101.605 170.655 101.935 171.135 ;
        RECT 102.105 170.845 102.330 171.305 ;
        RECT 102.500 170.655 102.830 171.135 ;
        RECT 99.675 170.065 100.025 170.315 ;
        RECT 96.515 168.925 96.855 169.895 ;
        RECT 97.025 168.755 97.195 169.895 ;
        RECT 97.385 169.725 99.820 169.895 ;
        RECT 97.465 168.755 97.715 169.555 ;
        RECT 98.360 168.925 98.690 169.725 ;
        RECT 98.990 168.755 99.320 169.555 ;
        RECT 99.490 168.925 99.820 169.725 ;
        RECT 100.195 168.755 100.485 169.920 ;
        RECT 100.655 169.895 100.830 170.505 ;
        RECT 101.605 170.485 102.830 170.655 ;
        RECT 103.460 170.525 103.960 171.135 ;
        RECT 104.335 170.565 104.720 171.135 ;
        RECT 104.890 170.845 105.215 171.305 ;
        RECT 105.735 170.675 106.015 171.135 ;
        RECT 101.000 170.145 101.695 170.315 ;
        RECT 101.525 169.895 101.695 170.145 ;
        RECT 101.870 170.115 102.290 170.315 ;
        RECT 102.460 170.115 102.790 170.315 ;
        RECT 102.960 170.115 103.290 170.315 ;
        RECT 103.460 169.895 103.630 170.525 ;
        RECT 103.815 170.065 104.165 170.315 ;
        RECT 104.335 169.895 104.615 170.565 ;
        RECT 104.890 170.505 106.015 170.675 ;
        RECT 104.890 170.395 105.340 170.505 ;
        RECT 104.785 170.065 105.340 170.395 ;
        RECT 106.205 170.335 106.605 171.135 ;
        RECT 107.005 170.845 107.275 171.305 ;
        RECT 107.445 170.675 107.730 171.135 ;
        RECT 100.655 168.925 100.995 169.895 ;
        RECT 101.165 168.755 101.335 169.895 ;
        RECT 101.525 169.725 103.960 169.895 ;
        RECT 101.605 168.755 101.855 169.555 ;
        RECT 102.500 168.925 102.830 169.725 ;
        RECT 103.130 168.755 103.460 169.555 ;
        RECT 103.630 168.925 103.960 169.725 ;
        RECT 104.335 168.925 104.720 169.895 ;
        RECT 104.890 169.605 105.340 170.065 ;
        RECT 105.510 169.775 106.605 170.335 ;
        RECT 104.890 169.385 106.015 169.605 ;
        RECT 104.890 168.755 105.215 169.215 ;
        RECT 105.735 168.925 106.015 169.385 ;
        RECT 106.205 168.925 106.605 169.775 ;
        RECT 106.775 170.505 107.730 170.675 ;
        RECT 108.220 170.525 108.720 171.135 ;
        RECT 106.775 169.605 106.985 170.505 ;
        RECT 107.155 169.775 107.845 170.335 ;
        RECT 108.015 170.065 108.365 170.315 ;
        RECT 108.550 169.895 108.720 170.525 ;
        RECT 109.350 170.655 109.680 171.135 ;
        RECT 109.850 170.845 110.075 171.305 ;
        RECT 110.245 170.655 110.575 171.135 ;
        RECT 109.350 170.485 110.575 170.655 ;
        RECT 110.765 170.505 111.015 171.305 ;
        RECT 111.185 170.505 111.525 171.135 ;
        RECT 112.155 170.555 113.365 171.305 ;
        RECT 108.890 170.115 109.220 170.315 ;
        RECT 109.390 170.115 109.720 170.315 ;
        RECT 109.890 170.115 110.310 170.315 ;
        RECT 110.485 170.145 111.180 170.315 ;
        RECT 110.485 169.895 110.655 170.145 ;
        RECT 111.350 169.895 111.525 170.505 ;
        RECT 108.220 169.725 110.655 169.895 ;
        RECT 106.775 169.385 107.730 169.605 ;
        RECT 107.005 168.755 107.275 169.215 ;
        RECT 107.445 168.925 107.730 169.385 ;
        RECT 108.220 168.925 108.550 169.725 ;
        RECT 108.720 168.755 109.050 169.555 ;
        RECT 109.350 168.925 109.680 169.725 ;
        RECT 110.325 168.755 110.575 169.555 ;
        RECT 110.845 168.755 111.015 169.895 ;
        RECT 111.185 168.925 111.525 169.895 ;
        RECT 112.155 169.845 112.675 170.385 ;
        RECT 112.845 170.015 113.365 170.555 ;
        RECT 112.155 168.755 113.365 169.845 ;
        RECT 26.970 168.585 113.450 168.755 ;
        RECT 27.055 167.495 28.265 168.585 ;
        RECT 29.555 167.915 29.835 168.585 ;
        RECT 30.005 167.695 30.305 168.245 ;
        RECT 30.505 167.865 30.835 168.585 ;
        RECT 31.025 167.865 31.485 168.415 ;
        RECT 27.055 166.785 27.575 167.325 ;
        RECT 27.745 166.955 28.265 167.495 ;
        RECT 29.370 167.275 29.635 167.635 ;
        RECT 30.005 167.525 30.945 167.695 ;
        RECT 30.775 167.275 30.945 167.525 ;
        RECT 29.370 167.025 30.045 167.275 ;
        RECT 30.265 167.025 30.605 167.275 ;
        RECT 30.775 166.945 31.065 167.275 ;
        RECT 30.775 166.855 30.945 166.945 ;
        RECT 27.055 166.035 28.265 166.785 ;
        RECT 29.555 166.665 30.945 166.855 ;
        RECT 29.555 166.305 29.885 166.665 ;
        RECT 31.235 166.495 31.485 167.865 ;
        RECT 30.505 166.035 30.755 166.495 ;
        RECT 30.925 166.205 31.485 166.495 ;
        RECT 31.660 167.445 31.995 168.415 ;
        RECT 32.165 167.445 32.335 168.585 ;
        RECT 32.505 168.245 34.535 168.415 ;
        RECT 31.660 166.775 31.830 167.445 ;
        RECT 32.505 167.275 32.675 168.245 ;
        RECT 32.000 166.945 32.255 167.275 ;
        RECT 32.480 166.945 32.675 167.275 ;
        RECT 32.845 167.905 33.970 168.075 ;
        RECT 32.085 166.775 32.255 166.945 ;
        RECT 32.845 166.775 33.015 167.905 ;
        RECT 31.660 166.205 31.915 166.775 ;
        RECT 32.085 166.605 33.015 166.775 ;
        RECT 33.185 167.565 34.195 167.735 ;
        RECT 33.185 166.765 33.355 167.565 ;
        RECT 32.840 166.570 33.015 166.605 ;
        RECT 32.085 166.035 32.415 166.435 ;
        RECT 32.840 166.205 33.370 166.570 ;
        RECT 33.560 166.545 33.835 167.365 ;
        RECT 33.555 166.375 33.835 166.545 ;
        RECT 33.560 166.205 33.835 166.375 ;
        RECT 34.005 166.205 34.195 167.565 ;
        RECT 34.365 167.580 34.535 168.245 ;
        RECT 34.705 167.825 34.875 168.585 ;
        RECT 35.110 167.825 35.625 168.235 ;
        RECT 34.365 167.390 35.115 167.580 ;
        RECT 35.285 167.015 35.625 167.825 ;
        RECT 35.795 167.420 36.085 168.585 ;
        RECT 36.805 167.655 36.975 168.415 ;
        RECT 37.155 167.825 37.485 168.585 ;
        RECT 36.805 167.485 37.470 167.655 ;
        RECT 37.655 167.510 37.925 168.415 ;
        RECT 37.300 167.340 37.470 167.485 ;
        RECT 34.395 166.845 35.625 167.015 ;
        RECT 36.735 166.935 37.065 167.305 ;
        RECT 37.300 167.010 37.585 167.340 ;
        RECT 34.375 166.035 34.885 166.570 ;
        RECT 35.105 166.240 35.350 166.845 ;
        RECT 35.795 166.035 36.085 166.760 ;
        RECT 37.300 166.755 37.470 167.010 ;
        RECT 36.805 166.585 37.470 166.755 ;
        RECT 37.755 166.710 37.925 167.510 ;
        RECT 38.300 167.615 38.630 168.415 ;
        RECT 38.800 167.785 39.130 168.585 ;
        RECT 39.430 167.615 39.760 168.415 ;
        RECT 40.405 167.785 40.655 168.585 ;
        RECT 38.300 167.445 40.735 167.615 ;
        RECT 40.925 167.445 41.095 168.585 ;
        RECT 41.265 167.445 41.605 168.415 ;
        RECT 38.095 167.025 38.445 167.275 ;
        RECT 38.630 166.815 38.800 167.445 ;
        RECT 38.970 167.025 39.300 167.225 ;
        RECT 39.470 167.025 39.800 167.225 ;
        RECT 39.970 167.025 40.390 167.225 ;
        RECT 40.565 167.195 40.735 167.445 ;
        RECT 41.375 167.395 41.605 167.445 ;
        RECT 40.565 167.025 41.260 167.195 ;
        RECT 36.805 166.205 36.975 166.585 ;
        RECT 37.155 166.035 37.485 166.415 ;
        RECT 37.665 166.205 37.925 166.710 ;
        RECT 38.300 166.205 38.800 166.815 ;
        RECT 39.430 166.685 40.655 166.855 ;
        RECT 41.430 166.835 41.605 167.395 ;
        RECT 39.430 166.205 39.760 166.685 ;
        RECT 39.930 166.035 40.155 166.495 ;
        RECT 40.325 166.205 40.655 166.685 ;
        RECT 40.845 166.035 41.095 166.835 ;
        RECT 41.265 166.205 41.605 166.835 ;
        RECT 42.150 167.605 42.405 168.275 ;
        RECT 42.585 167.785 42.870 168.585 ;
        RECT 43.050 167.865 43.380 168.375 ;
        RECT 42.150 166.745 42.330 167.605 ;
        RECT 43.050 167.275 43.300 167.865 ;
        RECT 43.650 167.715 43.820 168.325 ;
        RECT 43.990 167.895 44.320 168.585 ;
        RECT 44.550 168.035 44.790 168.325 ;
        RECT 44.990 168.205 45.410 168.585 ;
        RECT 45.590 168.115 46.220 168.365 ;
        RECT 46.690 168.205 47.020 168.585 ;
        RECT 45.590 168.035 45.760 168.115 ;
        RECT 47.190 168.035 47.360 168.325 ;
        RECT 47.540 168.205 47.920 168.585 ;
        RECT 48.160 168.200 48.990 168.370 ;
        RECT 44.550 167.865 45.760 168.035 ;
        RECT 42.500 166.945 43.300 167.275 ;
        RECT 42.150 166.545 42.405 166.745 ;
        RECT 42.065 166.375 42.405 166.545 ;
        RECT 42.150 166.215 42.405 166.375 ;
        RECT 42.585 166.035 42.870 166.495 ;
        RECT 43.050 166.295 43.300 166.945 ;
        RECT 43.500 167.695 43.820 167.715 ;
        RECT 43.500 167.525 45.420 167.695 ;
        RECT 43.500 166.630 43.690 167.525 ;
        RECT 45.590 167.355 45.760 167.865 ;
        RECT 45.930 167.605 46.450 167.915 ;
        RECT 43.860 167.185 45.760 167.355 ;
        RECT 43.860 167.125 44.190 167.185 ;
        RECT 44.340 166.955 44.670 167.015 ;
        RECT 44.010 166.685 44.670 166.955 ;
        RECT 43.500 166.300 43.820 166.630 ;
        RECT 44.000 166.035 44.660 166.515 ;
        RECT 44.860 166.425 45.030 167.185 ;
        RECT 45.930 167.015 46.110 167.425 ;
        RECT 45.200 166.845 45.530 166.965 ;
        RECT 46.280 166.845 46.450 167.605 ;
        RECT 45.200 166.675 46.450 166.845 ;
        RECT 46.620 167.785 47.990 168.035 ;
        RECT 46.620 167.015 46.810 167.785 ;
        RECT 47.740 167.525 47.990 167.785 ;
        RECT 46.980 167.355 47.230 167.515 ;
        RECT 48.160 167.355 48.330 168.200 ;
        RECT 49.225 167.915 49.395 168.415 ;
        RECT 49.565 168.085 49.895 168.585 ;
        RECT 48.500 167.525 49.000 167.905 ;
        RECT 49.225 167.745 49.920 167.915 ;
        RECT 46.980 167.185 48.330 167.355 ;
        RECT 47.910 167.145 48.330 167.185 ;
        RECT 46.620 166.675 47.040 167.015 ;
        RECT 47.330 166.685 47.740 167.015 ;
        RECT 44.860 166.255 45.710 166.425 ;
        RECT 46.270 166.035 46.590 166.495 ;
        RECT 46.790 166.245 47.040 166.675 ;
        RECT 47.330 166.035 47.740 166.475 ;
        RECT 47.910 166.415 48.080 167.145 ;
        RECT 48.250 166.595 48.600 166.965 ;
        RECT 48.780 166.655 49.000 167.525 ;
        RECT 49.170 166.955 49.580 167.575 ;
        RECT 49.750 166.775 49.920 167.745 ;
        RECT 49.225 166.585 49.920 166.775 ;
        RECT 47.910 166.215 48.925 166.415 ;
        RECT 49.225 166.255 49.395 166.585 ;
        RECT 49.565 166.035 49.895 166.415 ;
        RECT 50.110 166.295 50.335 168.415 ;
        RECT 50.505 168.085 50.835 168.585 ;
        RECT 51.005 167.915 51.175 168.415 ;
        RECT 50.510 167.745 51.175 167.915 ;
        RECT 50.510 166.755 50.740 167.745 ;
        RECT 50.910 166.925 51.260 167.575 ;
        RECT 51.440 167.445 51.775 168.415 ;
        RECT 51.945 167.445 52.115 168.585 ;
        RECT 52.285 168.245 54.315 168.415 ;
        RECT 51.440 166.775 51.610 167.445 ;
        RECT 52.285 167.275 52.455 168.245 ;
        RECT 51.780 166.945 52.035 167.275 ;
        RECT 52.260 166.945 52.455 167.275 ;
        RECT 52.625 167.905 53.750 168.075 ;
        RECT 51.865 166.775 52.035 166.945 ;
        RECT 52.625 166.775 52.795 167.905 ;
        RECT 50.510 166.585 51.175 166.755 ;
        RECT 50.505 166.035 50.835 166.415 ;
        RECT 51.005 166.295 51.175 166.585 ;
        RECT 51.440 166.205 51.695 166.775 ;
        RECT 51.865 166.605 52.795 166.775 ;
        RECT 52.965 167.565 53.975 167.735 ;
        RECT 52.965 166.765 53.135 167.565 ;
        RECT 53.340 166.885 53.615 167.365 ;
        RECT 53.335 166.715 53.615 166.885 ;
        RECT 52.620 166.570 52.795 166.605 ;
        RECT 51.865 166.035 52.195 166.435 ;
        RECT 52.620 166.205 53.150 166.570 ;
        RECT 53.340 166.205 53.615 166.715 ;
        RECT 53.785 166.205 53.975 167.565 ;
        RECT 54.145 167.580 54.315 168.245 ;
        RECT 54.485 167.825 54.655 168.585 ;
        RECT 54.890 167.825 55.405 168.235 ;
        RECT 54.145 167.390 54.895 167.580 ;
        RECT 55.065 167.015 55.405 167.825 ;
        RECT 56.585 167.655 56.755 168.415 ;
        RECT 56.935 167.825 57.265 168.585 ;
        RECT 56.585 167.485 57.250 167.655 ;
        RECT 57.435 167.510 57.705 168.415 ;
        RECT 57.080 167.340 57.250 167.485 ;
        RECT 54.175 166.845 55.405 167.015 ;
        RECT 56.515 166.935 56.845 167.305 ;
        RECT 57.080 167.010 57.365 167.340 ;
        RECT 54.155 166.035 54.665 166.570 ;
        RECT 54.885 166.240 55.130 166.845 ;
        RECT 57.080 166.755 57.250 167.010 ;
        RECT 56.585 166.585 57.250 166.755 ;
        RECT 57.535 166.710 57.705 167.510 ;
        RECT 56.585 166.205 56.755 166.585 ;
        RECT 56.935 166.035 57.265 166.415 ;
        RECT 57.445 166.205 57.705 166.710 ;
        RECT 57.875 167.445 58.215 168.415 ;
        RECT 58.385 167.445 58.555 168.585 ;
        RECT 58.825 167.785 59.075 168.585 ;
        RECT 59.720 167.615 60.050 168.415 ;
        RECT 60.350 167.785 60.680 168.585 ;
        RECT 60.850 167.615 61.180 168.415 ;
        RECT 58.745 167.445 61.180 167.615 ;
        RECT 57.875 166.885 58.050 167.445 ;
        RECT 58.745 167.195 58.915 167.445 ;
        RECT 58.220 167.025 58.915 167.195 ;
        RECT 59.090 167.025 59.510 167.225 ;
        RECT 59.680 167.025 60.010 167.225 ;
        RECT 60.180 167.025 60.510 167.225 ;
        RECT 57.875 166.835 58.105 166.885 ;
        RECT 57.875 166.205 58.215 166.835 ;
        RECT 58.385 166.035 58.635 166.835 ;
        RECT 58.825 166.685 60.050 166.855 ;
        RECT 58.825 166.205 59.155 166.685 ;
        RECT 59.325 166.035 59.550 166.495 ;
        RECT 59.720 166.205 60.050 166.685 ;
        RECT 60.680 166.815 60.850 167.445 ;
        RECT 61.555 167.420 61.845 168.585 ;
        RECT 62.015 167.445 62.355 168.415 ;
        RECT 62.525 167.445 62.695 168.585 ;
        RECT 62.965 167.785 63.215 168.585 ;
        RECT 63.860 167.615 64.190 168.415 ;
        RECT 64.490 167.785 64.820 168.585 ;
        RECT 64.990 167.615 65.320 168.415 ;
        RECT 62.885 167.445 65.320 167.615 ;
        RECT 66.165 167.605 66.495 168.415 ;
        RECT 66.665 167.785 66.905 168.585 ;
        RECT 61.035 167.025 61.385 167.275 ;
        RECT 62.015 166.835 62.190 167.445 ;
        RECT 62.885 167.195 63.055 167.445 ;
        RECT 62.360 167.025 63.055 167.195 ;
        RECT 63.225 167.055 63.650 167.225 ;
        RECT 63.230 167.025 63.650 167.055 ;
        RECT 63.820 167.025 64.150 167.225 ;
        RECT 64.320 167.025 64.650 167.225 ;
        RECT 60.680 166.205 61.180 166.815 ;
        RECT 61.555 166.035 61.845 166.760 ;
        RECT 62.015 166.205 62.355 166.835 ;
        RECT 62.525 166.035 62.775 166.835 ;
        RECT 62.965 166.685 64.190 166.855 ;
        RECT 62.965 166.205 63.295 166.685 ;
        RECT 63.465 166.035 63.690 166.495 ;
        RECT 63.860 166.205 64.190 166.685 ;
        RECT 64.820 166.815 64.990 167.445 ;
        RECT 66.165 167.435 66.880 167.605 ;
        RECT 65.175 167.025 65.525 167.275 ;
        RECT 66.160 167.025 66.540 167.265 ;
        RECT 66.710 167.195 66.880 167.435 ;
        RECT 67.085 167.565 67.255 168.415 ;
        RECT 67.425 167.785 67.755 168.585 ;
        RECT 67.925 167.565 68.095 168.415 ;
        RECT 67.085 167.395 68.095 167.565 ;
        RECT 68.265 167.435 68.595 168.585 ;
        RECT 69.120 167.615 69.450 168.415 ;
        RECT 69.620 167.785 69.950 168.585 ;
        RECT 70.250 167.615 70.580 168.415 ;
        RECT 71.225 167.785 71.475 168.585 ;
        RECT 69.120 167.445 71.555 167.615 ;
        RECT 71.745 167.445 71.915 168.585 ;
        RECT 72.085 167.445 72.425 168.415 ;
        RECT 66.710 167.025 67.210 167.195 ;
        RECT 66.710 166.855 66.880 167.025 ;
        RECT 67.600 166.855 68.095 167.395 ;
        RECT 68.915 167.025 69.265 167.275 ;
        RECT 64.820 166.205 65.320 166.815 ;
        RECT 66.245 166.685 66.880 166.855 ;
        RECT 67.085 166.685 68.095 166.855 ;
        RECT 66.245 166.205 66.415 166.685 ;
        RECT 66.595 166.035 66.835 166.515 ;
        RECT 67.085 166.205 67.255 166.685 ;
        RECT 67.425 166.035 67.755 166.515 ;
        RECT 67.925 166.205 68.095 166.685 ;
        RECT 68.265 166.035 68.595 166.835 ;
        RECT 69.450 166.815 69.620 167.445 ;
        RECT 69.790 167.025 70.120 167.225 ;
        RECT 70.290 167.025 70.620 167.225 ;
        RECT 70.790 167.025 71.210 167.225 ;
        RECT 71.385 167.195 71.555 167.445 ;
        RECT 72.195 167.395 72.425 167.445 ;
        RECT 71.385 167.025 72.080 167.195 ;
        RECT 69.120 166.205 69.620 166.815 ;
        RECT 70.250 166.685 71.475 166.855 ;
        RECT 72.250 166.835 72.425 167.395 ;
        RECT 70.250 166.205 70.580 166.685 ;
        RECT 70.750 166.035 70.975 166.495 ;
        RECT 71.145 166.205 71.475 166.685 ;
        RECT 71.665 166.035 71.915 166.835 ;
        RECT 72.085 166.205 72.425 166.835 ;
        RECT 72.595 167.445 72.935 168.415 ;
        RECT 73.105 167.445 73.275 168.585 ;
        RECT 73.545 167.785 73.795 168.585 ;
        RECT 74.440 167.615 74.770 168.415 ;
        RECT 75.070 167.785 75.400 168.585 ;
        RECT 75.570 167.615 75.900 168.415 ;
        RECT 73.465 167.445 75.900 167.615 ;
        RECT 76.650 167.605 76.905 168.275 ;
        RECT 77.085 167.785 77.370 168.585 ;
        RECT 77.550 167.865 77.880 168.375 ;
        RECT 72.595 166.885 72.770 167.445 ;
        RECT 73.465 167.195 73.635 167.445 ;
        RECT 72.940 167.025 73.635 167.195 ;
        RECT 73.810 167.025 74.230 167.225 ;
        RECT 74.400 167.025 74.730 167.225 ;
        RECT 74.900 167.025 75.230 167.225 ;
        RECT 72.595 166.835 72.825 166.885 ;
        RECT 72.595 166.205 72.935 166.835 ;
        RECT 73.105 166.035 73.355 166.835 ;
        RECT 73.545 166.685 74.770 166.855 ;
        RECT 73.545 166.205 73.875 166.685 ;
        RECT 74.045 166.035 74.270 166.495 ;
        RECT 74.440 166.205 74.770 166.685 ;
        RECT 75.400 166.815 75.570 167.445 ;
        RECT 75.755 167.025 76.105 167.275 ;
        RECT 75.400 166.205 75.900 166.815 ;
        RECT 76.650 166.745 76.830 167.605 ;
        RECT 77.550 167.275 77.800 167.865 ;
        RECT 78.150 167.715 78.320 168.325 ;
        RECT 78.490 167.895 78.820 168.585 ;
        RECT 79.050 168.035 79.290 168.325 ;
        RECT 79.490 168.205 79.910 168.585 ;
        RECT 80.090 168.115 80.720 168.365 ;
        RECT 81.190 168.205 81.520 168.585 ;
        RECT 80.090 168.035 80.260 168.115 ;
        RECT 81.690 168.035 81.860 168.325 ;
        RECT 82.040 168.205 82.420 168.585 ;
        RECT 82.660 168.200 83.490 168.370 ;
        RECT 79.050 167.865 80.260 168.035 ;
        RECT 77.000 166.945 77.800 167.275 ;
        RECT 76.650 166.545 76.905 166.745 ;
        RECT 76.565 166.375 76.905 166.545 ;
        RECT 76.650 166.215 76.905 166.375 ;
        RECT 77.085 166.035 77.370 166.495 ;
        RECT 77.550 166.295 77.800 166.945 ;
        RECT 78.000 167.695 78.320 167.715 ;
        RECT 78.000 167.525 79.920 167.695 ;
        RECT 78.000 166.630 78.190 167.525 ;
        RECT 80.090 167.355 80.260 167.865 ;
        RECT 80.430 167.605 80.950 167.915 ;
        RECT 78.360 167.185 80.260 167.355 ;
        RECT 78.360 167.125 78.690 167.185 ;
        RECT 78.840 166.955 79.170 167.015 ;
        RECT 78.510 166.685 79.170 166.955 ;
        RECT 78.000 166.300 78.320 166.630 ;
        RECT 78.500 166.035 79.160 166.515 ;
        RECT 79.360 166.425 79.530 167.185 ;
        RECT 80.430 167.015 80.610 167.425 ;
        RECT 79.700 166.845 80.030 166.965 ;
        RECT 80.780 166.845 80.950 167.605 ;
        RECT 79.700 166.675 80.950 166.845 ;
        RECT 81.120 167.785 82.490 168.035 ;
        RECT 81.120 167.015 81.310 167.785 ;
        RECT 82.240 167.525 82.490 167.785 ;
        RECT 81.480 167.355 81.730 167.515 ;
        RECT 82.660 167.355 82.830 168.200 ;
        RECT 83.725 167.915 83.895 168.415 ;
        RECT 84.065 168.085 84.395 168.585 ;
        RECT 83.000 167.525 83.500 167.905 ;
        RECT 83.725 167.745 84.420 167.915 ;
        RECT 81.480 167.185 82.830 167.355 ;
        RECT 82.410 167.145 82.830 167.185 ;
        RECT 81.120 166.675 81.540 167.015 ;
        RECT 81.830 166.685 82.240 167.015 ;
        RECT 79.360 166.255 80.210 166.425 ;
        RECT 80.770 166.035 81.090 166.495 ;
        RECT 81.290 166.245 81.540 166.675 ;
        RECT 81.830 166.035 82.240 166.475 ;
        RECT 82.410 166.415 82.580 167.145 ;
        RECT 82.750 166.595 83.100 166.965 ;
        RECT 83.280 166.655 83.500 167.525 ;
        RECT 83.670 166.955 84.080 167.575 ;
        RECT 84.250 166.775 84.420 167.745 ;
        RECT 83.725 166.585 84.420 166.775 ;
        RECT 82.410 166.215 83.425 166.415 ;
        RECT 83.725 166.255 83.895 166.585 ;
        RECT 84.065 166.035 84.395 166.415 ;
        RECT 84.610 166.295 84.835 168.415 ;
        RECT 85.005 168.085 85.335 168.585 ;
        RECT 85.505 167.915 85.675 168.415 ;
        RECT 85.010 167.745 85.675 167.915 ;
        RECT 85.010 166.755 85.240 167.745 ;
        RECT 85.410 166.925 85.760 167.575 ;
        RECT 85.935 167.510 86.205 168.415 ;
        RECT 86.375 167.825 86.705 168.585 ;
        RECT 86.885 167.655 87.055 168.415 ;
        RECT 85.010 166.585 85.675 166.755 ;
        RECT 85.005 166.035 85.335 166.415 ;
        RECT 85.505 166.295 85.675 166.585 ;
        RECT 85.935 166.710 86.105 167.510 ;
        RECT 86.390 167.485 87.055 167.655 ;
        RECT 86.390 167.340 86.560 167.485 ;
        RECT 87.315 167.420 87.605 168.585 ;
        RECT 87.775 167.825 88.290 168.235 ;
        RECT 88.525 167.825 88.695 168.585 ;
        RECT 88.865 168.245 90.895 168.415 ;
        RECT 86.275 167.010 86.560 167.340 ;
        RECT 86.390 166.755 86.560 167.010 ;
        RECT 86.795 166.935 87.125 167.305 ;
        RECT 87.775 167.015 88.115 167.825 ;
        RECT 88.865 167.580 89.035 168.245 ;
        RECT 89.430 167.905 90.555 168.075 ;
        RECT 88.285 167.390 89.035 167.580 ;
        RECT 89.205 167.565 90.215 167.735 ;
        RECT 87.775 166.845 89.005 167.015 ;
        RECT 85.935 166.205 86.195 166.710 ;
        RECT 86.390 166.585 87.055 166.755 ;
        RECT 86.375 166.035 86.705 166.415 ;
        RECT 86.885 166.205 87.055 166.585 ;
        RECT 87.315 166.035 87.605 166.760 ;
        RECT 88.050 166.240 88.295 166.845 ;
        RECT 88.515 166.035 89.025 166.570 ;
        RECT 89.205 166.205 89.395 167.565 ;
        RECT 89.565 167.225 89.840 167.365 ;
        RECT 89.565 167.055 89.845 167.225 ;
        RECT 89.565 166.205 89.840 167.055 ;
        RECT 90.045 166.765 90.215 167.565 ;
        RECT 90.385 166.775 90.555 167.905 ;
        RECT 90.725 167.275 90.895 168.245 ;
        RECT 91.065 167.445 91.235 168.585 ;
        RECT 91.405 167.445 91.740 168.415 ;
        RECT 90.725 166.945 90.920 167.275 ;
        RECT 91.145 166.945 91.400 167.275 ;
        RECT 91.145 166.775 91.315 166.945 ;
        RECT 91.570 166.775 91.740 167.445 ;
        RECT 90.385 166.605 91.315 166.775 ;
        RECT 90.385 166.570 90.560 166.605 ;
        RECT 90.030 166.205 90.560 166.570 ;
        RECT 90.985 166.035 91.315 166.435 ;
        RECT 91.485 166.205 91.740 166.775 ;
        RECT 91.915 167.445 92.300 168.415 ;
        RECT 92.470 168.125 92.795 168.585 ;
        RECT 93.315 167.955 93.595 168.415 ;
        RECT 92.470 167.735 93.595 167.955 ;
        RECT 91.915 166.775 92.195 167.445 ;
        RECT 92.470 167.275 92.920 167.735 ;
        RECT 93.785 167.565 94.185 168.415 ;
        RECT 94.585 168.125 94.855 168.585 ;
        RECT 95.025 167.955 95.310 168.415 ;
        RECT 92.365 166.945 92.920 167.275 ;
        RECT 93.090 167.005 94.185 167.565 ;
        RECT 92.470 166.835 92.920 166.945 ;
        RECT 91.915 166.205 92.300 166.775 ;
        RECT 92.470 166.665 93.595 166.835 ;
        RECT 92.470 166.035 92.795 166.495 ;
        RECT 93.315 166.205 93.595 166.665 ;
        RECT 93.785 166.205 94.185 167.005 ;
        RECT 94.355 167.735 95.310 167.955 ;
        RECT 94.355 166.835 94.565 167.735 ;
        RECT 94.735 167.005 95.425 167.565 ;
        RECT 95.595 167.445 95.935 168.415 ;
        RECT 96.105 167.445 96.275 168.585 ;
        RECT 96.545 167.785 96.795 168.585 ;
        RECT 97.440 167.615 97.770 168.415 ;
        RECT 98.070 167.785 98.400 168.585 ;
        RECT 98.570 167.615 98.900 168.415 ;
        RECT 96.465 167.445 98.900 167.615 ;
        RECT 99.745 167.605 100.075 168.415 ;
        RECT 100.245 167.785 100.485 168.585 ;
        RECT 95.595 166.835 95.770 167.445 ;
        RECT 96.465 167.195 96.635 167.445 ;
        RECT 95.940 167.025 96.635 167.195 ;
        RECT 96.810 167.025 97.230 167.225 ;
        RECT 97.400 167.025 97.730 167.225 ;
        RECT 97.900 167.025 98.230 167.225 ;
        RECT 94.355 166.665 95.310 166.835 ;
        RECT 94.585 166.035 94.855 166.495 ;
        RECT 95.025 166.205 95.310 166.665 ;
        RECT 95.595 166.205 95.935 166.835 ;
        RECT 96.105 166.035 96.355 166.835 ;
        RECT 96.545 166.685 97.770 166.855 ;
        RECT 96.545 166.205 96.875 166.685 ;
        RECT 97.045 166.035 97.270 166.495 ;
        RECT 97.440 166.205 97.770 166.685 ;
        RECT 98.400 166.815 98.570 167.445 ;
        RECT 99.745 167.435 100.460 167.605 ;
        RECT 98.755 167.025 99.105 167.275 ;
        RECT 99.740 167.025 100.120 167.265 ;
        RECT 100.290 167.195 100.460 167.435 ;
        RECT 100.665 167.565 100.835 168.415 ;
        RECT 101.005 167.785 101.335 168.585 ;
        RECT 101.505 167.565 101.675 168.415 ;
        RECT 100.665 167.395 101.675 167.565 ;
        RECT 101.845 167.435 102.175 168.585 ;
        RECT 101.180 167.225 101.675 167.395 ;
        RECT 100.290 167.025 100.790 167.195 ;
        RECT 101.175 167.055 101.675 167.225 ;
        RECT 100.290 166.855 100.460 167.025 ;
        RECT 101.180 166.855 101.675 167.055 ;
        RECT 98.400 166.205 98.900 166.815 ;
        RECT 99.825 166.685 100.460 166.855 ;
        RECT 100.665 166.685 101.675 166.855 ;
        RECT 102.500 167.395 102.755 168.275 ;
        RECT 102.925 167.445 103.230 168.585 ;
        RECT 103.570 168.205 103.900 168.585 ;
        RECT 104.080 168.035 104.250 168.325 ;
        RECT 104.420 168.125 104.670 168.585 ;
        RECT 103.450 167.865 104.250 168.035 ;
        RECT 104.840 168.075 105.710 168.415 ;
        RECT 99.825 166.205 99.995 166.685 ;
        RECT 100.175 166.035 100.415 166.515 ;
        RECT 100.665 166.205 100.835 166.685 ;
        RECT 101.005 166.035 101.335 166.515 ;
        RECT 101.505 166.205 101.675 166.685 ;
        RECT 101.845 166.035 102.175 166.835 ;
        RECT 102.500 166.745 102.710 167.395 ;
        RECT 103.450 167.275 103.620 167.865 ;
        RECT 104.840 167.695 105.010 168.075 ;
        RECT 105.945 167.955 106.115 168.415 ;
        RECT 106.285 168.125 106.655 168.585 ;
        RECT 106.950 167.985 107.120 168.325 ;
        RECT 107.290 168.155 107.620 168.585 ;
        RECT 107.855 167.985 108.025 168.325 ;
        RECT 103.790 167.525 105.010 167.695 ;
        RECT 105.180 167.615 105.640 167.905 ;
        RECT 105.945 167.785 106.505 167.955 ;
        RECT 106.950 167.815 108.025 167.985 ;
        RECT 108.195 168.085 108.875 168.415 ;
        RECT 109.090 168.085 109.340 168.415 ;
        RECT 109.510 168.125 109.760 168.585 ;
        RECT 106.335 167.645 106.505 167.785 ;
        RECT 105.180 167.605 106.145 167.615 ;
        RECT 104.840 167.435 105.010 167.525 ;
        RECT 105.470 167.445 106.145 167.605 ;
        RECT 102.880 167.245 103.620 167.275 ;
        RECT 102.880 166.945 103.795 167.245 ;
        RECT 103.470 166.770 103.795 166.945 ;
        RECT 102.500 166.215 102.755 166.745 ;
        RECT 102.925 166.035 103.230 166.495 ;
        RECT 103.475 166.415 103.795 166.770 ;
        RECT 103.965 166.985 104.505 167.355 ;
        RECT 104.840 167.265 105.245 167.435 ;
        RECT 103.965 166.585 104.205 166.985 ;
        RECT 104.685 166.815 104.905 167.095 ;
        RECT 104.375 166.645 104.905 166.815 ;
        RECT 104.375 166.415 104.545 166.645 ;
        RECT 105.075 166.485 105.245 167.265 ;
        RECT 105.415 166.655 105.765 167.275 ;
        RECT 105.935 166.655 106.145 167.445 ;
        RECT 106.335 167.475 107.835 167.645 ;
        RECT 106.335 166.785 106.505 167.475 ;
        RECT 108.195 167.305 108.365 168.085 ;
        RECT 109.170 167.955 109.340 168.085 ;
        RECT 106.675 167.135 108.365 167.305 ;
        RECT 108.535 167.525 109.000 167.915 ;
        RECT 109.170 167.785 109.565 167.955 ;
        RECT 106.675 166.955 106.845 167.135 ;
        RECT 103.475 166.245 104.545 166.415 ;
        RECT 104.715 166.035 104.905 166.475 ;
        RECT 105.075 166.205 106.025 166.485 ;
        RECT 106.335 166.395 106.595 166.785 ;
        RECT 107.015 166.715 107.805 166.965 ;
        RECT 106.245 166.225 106.595 166.395 ;
        RECT 106.805 166.035 107.135 166.495 ;
        RECT 108.010 166.425 108.180 167.135 ;
        RECT 108.535 166.935 108.705 167.525 ;
        RECT 108.350 166.715 108.705 166.935 ;
        RECT 108.875 166.715 109.225 167.335 ;
        RECT 109.395 166.425 109.565 167.785 ;
        RECT 109.930 167.615 110.255 168.400 ;
        RECT 109.735 166.565 110.195 167.615 ;
        RECT 108.010 166.255 108.865 166.425 ;
        RECT 109.070 166.255 109.565 166.425 ;
        RECT 109.735 166.035 110.065 166.395 ;
        RECT 110.425 166.295 110.595 168.415 ;
        RECT 110.765 168.085 111.095 168.585 ;
        RECT 111.265 167.915 111.520 168.415 ;
        RECT 110.770 167.745 111.520 167.915 ;
        RECT 110.770 166.755 111.000 167.745 ;
        RECT 111.170 166.925 111.520 167.575 ;
        RECT 112.155 167.495 113.365 168.585 ;
        RECT 112.155 166.955 112.675 167.495 ;
        RECT 112.845 166.785 113.365 167.325 ;
        RECT 110.770 166.585 111.520 166.755 ;
        RECT 110.765 166.035 111.095 166.415 ;
        RECT 111.265 166.295 111.520 166.585 ;
        RECT 112.155 166.035 113.365 166.785 ;
        RECT 26.970 165.865 113.450 166.035 ;
        RECT 27.055 165.115 28.265 165.865 ;
        RECT 28.810 165.155 29.065 165.685 ;
        RECT 29.245 165.405 29.530 165.865 ;
        RECT 27.055 164.575 27.575 165.115 ;
        RECT 27.745 164.405 28.265 164.945 ;
        RECT 27.055 163.315 28.265 164.405 ;
        RECT 28.810 164.295 28.990 165.155 ;
        RECT 29.710 164.955 29.960 165.605 ;
        RECT 29.160 164.625 29.960 164.955 ;
        RECT 28.810 163.825 29.065 164.295 ;
        RECT 28.725 163.655 29.065 163.825 ;
        RECT 28.810 163.625 29.065 163.655 ;
        RECT 29.245 163.315 29.530 164.115 ;
        RECT 29.710 164.035 29.960 164.625 ;
        RECT 30.160 165.270 30.480 165.600 ;
        RECT 30.660 165.385 31.320 165.865 ;
        RECT 31.520 165.475 32.370 165.645 ;
        RECT 30.160 164.375 30.350 165.270 ;
        RECT 30.670 164.945 31.330 165.215 ;
        RECT 31.000 164.885 31.330 164.945 ;
        RECT 30.520 164.715 30.850 164.775 ;
        RECT 31.520 164.715 31.690 165.475 ;
        RECT 32.930 165.405 33.250 165.865 ;
        RECT 33.450 165.225 33.700 165.655 ;
        RECT 33.990 165.425 34.400 165.865 ;
        RECT 34.570 165.485 35.585 165.685 ;
        RECT 31.860 165.055 33.110 165.225 ;
        RECT 31.860 164.935 32.190 165.055 ;
        RECT 30.520 164.545 32.420 164.715 ;
        RECT 30.160 164.205 32.080 164.375 ;
        RECT 30.160 164.185 30.480 164.205 ;
        RECT 29.710 163.525 30.040 164.035 ;
        RECT 30.310 163.575 30.480 164.185 ;
        RECT 32.250 164.035 32.420 164.545 ;
        RECT 32.590 164.475 32.770 164.885 ;
        RECT 32.940 164.295 33.110 165.055 ;
        RECT 30.650 163.315 30.980 164.005 ;
        RECT 31.210 163.865 32.420 164.035 ;
        RECT 32.590 163.985 33.110 164.295 ;
        RECT 33.280 164.885 33.700 165.225 ;
        RECT 33.990 164.885 34.400 165.215 ;
        RECT 33.280 164.115 33.470 164.885 ;
        RECT 34.570 164.755 34.740 165.485 ;
        RECT 35.885 165.315 36.055 165.645 ;
        RECT 36.225 165.485 36.555 165.865 ;
        RECT 34.910 164.935 35.260 165.305 ;
        RECT 34.570 164.715 34.990 164.755 ;
        RECT 33.640 164.545 34.990 164.715 ;
        RECT 33.640 164.385 33.890 164.545 ;
        RECT 34.400 164.115 34.650 164.375 ;
        RECT 33.280 163.865 34.650 164.115 ;
        RECT 31.210 163.575 31.450 163.865 ;
        RECT 32.250 163.785 32.420 163.865 ;
        RECT 31.650 163.315 32.070 163.695 ;
        RECT 32.250 163.535 32.880 163.785 ;
        RECT 33.350 163.315 33.680 163.695 ;
        RECT 33.850 163.575 34.020 163.865 ;
        RECT 34.820 163.700 34.990 164.545 ;
        RECT 35.440 164.375 35.660 165.245 ;
        RECT 35.885 165.125 36.580 165.315 ;
        RECT 35.160 163.995 35.660 164.375 ;
        RECT 35.830 164.325 36.240 164.945 ;
        RECT 36.410 164.155 36.580 165.125 ;
        RECT 35.885 163.985 36.580 164.155 ;
        RECT 34.200 163.315 34.580 163.695 ;
        RECT 34.820 163.530 35.650 163.700 ;
        RECT 35.885 163.485 36.055 163.985 ;
        RECT 36.225 163.315 36.555 163.815 ;
        RECT 36.770 163.485 36.995 165.605 ;
        RECT 37.165 165.485 37.495 165.865 ;
        RECT 37.665 165.315 37.835 165.605 ;
        RECT 37.170 165.145 37.835 165.315 ;
        RECT 38.095 165.190 38.355 165.695 ;
        RECT 38.535 165.485 38.865 165.865 ;
        RECT 39.045 165.315 39.215 165.695 ;
        RECT 37.170 164.155 37.400 165.145 ;
        RECT 37.570 164.325 37.920 164.975 ;
        RECT 38.095 164.390 38.265 165.190 ;
        RECT 38.550 165.145 39.215 165.315 ;
        RECT 38.550 164.890 38.720 165.145 ;
        RECT 40.400 165.125 40.655 165.695 ;
        RECT 40.825 165.465 41.155 165.865 ;
        RECT 41.580 165.330 42.110 165.695 ;
        RECT 42.300 165.525 42.575 165.695 ;
        RECT 42.295 165.355 42.575 165.525 ;
        RECT 41.580 165.295 41.755 165.330 ;
        RECT 40.825 165.125 41.755 165.295 ;
        RECT 38.435 164.560 38.720 164.890 ;
        RECT 38.955 164.595 39.285 164.965 ;
        RECT 38.550 164.415 38.720 164.560 ;
        RECT 40.400 164.455 40.570 165.125 ;
        RECT 40.825 164.955 40.995 165.125 ;
        RECT 40.740 164.625 40.995 164.955 ;
        RECT 41.220 164.625 41.415 164.955 ;
        RECT 37.170 163.985 37.835 164.155 ;
        RECT 37.165 163.315 37.495 163.815 ;
        RECT 37.665 163.485 37.835 163.985 ;
        RECT 38.095 163.485 38.365 164.390 ;
        RECT 38.550 164.245 39.215 164.415 ;
        RECT 38.535 163.315 38.865 164.075 ;
        RECT 39.045 163.485 39.215 164.245 ;
        RECT 40.400 163.485 40.735 164.455 ;
        RECT 40.905 163.315 41.075 164.455 ;
        RECT 41.245 163.655 41.415 164.625 ;
        RECT 41.585 163.995 41.755 165.125 ;
        RECT 41.925 164.335 42.095 165.135 ;
        RECT 42.300 164.535 42.575 165.355 ;
        RECT 42.745 164.335 42.935 165.695 ;
        RECT 43.115 165.330 43.625 165.865 ;
        RECT 43.845 165.055 44.090 165.660 ;
        RECT 45.110 165.235 45.395 165.695 ;
        RECT 45.565 165.405 45.835 165.865 ;
        RECT 45.110 165.065 46.065 165.235 ;
        RECT 43.135 164.885 44.365 165.055 ;
        RECT 41.925 164.165 42.935 164.335 ;
        RECT 43.105 164.320 43.855 164.510 ;
        RECT 41.585 163.825 42.710 163.995 ;
        RECT 43.105 163.655 43.275 164.320 ;
        RECT 44.025 164.075 44.365 164.885 ;
        RECT 44.995 164.335 45.685 164.895 ;
        RECT 45.855 164.165 46.065 165.065 ;
        RECT 41.245 163.485 43.275 163.655 ;
        RECT 43.445 163.315 43.615 164.075 ;
        RECT 43.850 163.665 44.365 164.075 ;
        RECT 45.110 163.945 46.065 164.165 ;
        RECT 46.235 164.895 46.635 165.695 ;
        RECT 46.825 165.235 47.105 165.695 ;
        RECT 47.625 165.405 47.950 165.865 ;
        RECT 46.825 165.065 47.950 165.235 ;
        RECT 48.120 165.125 48.505 165.695 ;
        RECT 48.675 165.140 48.965 165.865 ;
        RECT 49.335 165.235 49.665 165.595 ;
        RECT 50.285 165.405 50.535 165.865 ;
        RECT 50.705 165.405 51.265 165.695 ;
        RECT 47.500 164.955 47.950 165.065 ;
        RECT 46.235 164.335 47.330 164.895 ;
        RECT 47.500 164.625 48.055 164.955 ;
        RECT 45.110 163.485 45.395 163.945 ;
        RECT 45.565 163.315 45.835 163.775 ;
        RECT 46.235 163.485 46.635 164.335 ;
        RECT 47.500 164.165 47.950 164.625 ;
        RECT 48.225 164.455 48.505 165.125 ;
        RECT 49.335 165.045 50.725 165.235 ;
        RECT 50.555 164.955 50.725 165.045 ;
        RECT 49.150 164.625 49.825 164.875 ;
        RECT 50.045 164.625 50.385 164.875 ;
        RECT 50.555 164.625 50.845 164.955 ;
        RECT 46.825 163.945 47.950 164.165 ;
        RECT 46.825 163.485 47.105 163.945 ;
        RECT 47.625 163.315 47.950 163.775 ;
        RECT 48.120 163.485 48.505 164.455 ;
        RECT 48.675 163.315 48.965 164.480 ;
        RECT 49.150 164.265 49.415 164.625 ;
        RECT 50.555 164.375 50.725 164.625 ;
        RECT 49.785 164.205 50.725 164.375 ;
        RECT 49.335 163.315 49.615 163.985 ;
        RECT 49.785 163.655 50.085 164.205 ;
        RECT 51.015 164.035 51.265 165.405 ;
        RECT 50.285 163.315 50.615 164.035 ;
        RECT 50.805 163.485 51.265 164.035 ;
        RECT 51.435 165.065 51.775 165.695 ;
        RECT 51.945 165.065 52.195 165.865 ;
        RECT 52.385 165.215 52.715 165.695 ;
        RECT 52.885 165.405 53.110 165.865 ;
        RECT 53.280 165.215 53.610 165.695 ;
        RECT 51.435 164.455 51.610 165.065 ;
        RECT 52.385 165.045 53.610 165.215 ;
        RECT 54.240 165.085 54.740 165.695 ;
        RECT 55.320 165.085 55.820 165.695 ;
        RECT 51.780 164.705 52.475 164.875 ;
        RECT 52.305 164.455 52.475 164.705 ;
        RECT 52.650 164.675 53.070 164.875 ;
        RECT 53.240 164.675 53.570 164.875 ;
        RECT 53.740 164.675 54.070 164.875 ;
        RECT 54.240 164.455 54.410 165.085 ;
        RECT 54.595 164.625 54.945 164.875 ;
        RECT 55.115 164.625 55.465 164.875 ;
        RECT 55.650 164.455 55.820 165.085 ;
        RECT 56.450 165.215 56.780 165.695 ;
        RECT 56.950 165.405 57.175 165.865 ;
        RECT 57.345 165.215 57.675 165.695 ;
        RECT 56.450 165.045 57.675 165.215 ;
        RECT 57.865 165.065 58.115 165.865 ;
        RECT 58.285 165.065 58.625 165.695 ;
        RECT 55.990 164.675 56.320 164.875 ;
        RECT 56.490 164.675 56.820 164.875 ;
        RECT 56.990 164.675 57.410 164.875 ;
        RECT 57.585 164.705 58.280 164.875 ;
        RECT 57.585 164.455 57.755 164.705 ;
        RECT 58.450 164.455 58.625 165.065 ;
        RECT 51.435 163.485 51.775 164.455 ;
        RECT 51.945 163.315 52.115 164.455 ;
        RECT 52.305 164.285 54.740 164.455 ;
        RECT 52.385 163.315 52.635 164.115 ;
        RECT 53.280 163.485 53.610 164.285 ;
        RECT 53.910 163.315 54.240 164.115 ;
        RECT 54.410 163.485 54.740 164.285 ;
        RECT 55.320 164.285 57.755 164.455 ;
        RECT 55.320 163.485 55.650 164.285 ;
        RECT 55.820 163.315 56.150 164.115 ;
        RECT 56.450 163.485 56.780 164.285 ;
        RECT 57.425 163.315 57.675 164.115 ;
        RECT 57.945 163.315 58.115 164.455 ;
        RECT 58.285 163.485 58.625 164.455 ;
        RECT 59.630 165.155 59.885 165.685 ;
        RECT 60.065 165.405 60.350 165.865 ;
        RECT 59.630 164.295 59.810 165.155 ;
        RECT 60.530 164.955 60.780 165.605 ;
        RECT 59.980 164.625 60.780 164.955 ;
        RECT 59.630 163.825 59.885 164.295 ;
        RECT 59.545 163.655 59.885 163.825 ;
        RECT 59.630 163.625 59.885 163.655 ;
        RECT 60.065 163.315 60.350 164.115 ;
        RECT 60.530 164.035 60.780 164.625 ;
        RECT 60.980 165.270 61.300 165.600 ;
        RECT 61.480 165.385 62.140 165.865 ;
        RECT 62.340 165.475 63.190 165.645 ;
        RECT 60.980 164.375 61.170 165.270 ;
        RECT 61.490 164.945 62.150 165.215 ;
        RECT 61.820 164.885 62.150 164.945 ;
        RECT 61.340 164.715 61.670 164.775 ;
        RECT 62.340 164.715 62.510 165.475 ;
        RECT 63.750 165.405 64.070 165.865 ;
        RECT 64.270 165.225 64.520 165.655 ;
        RECT 64.810 165.425 65.220 165.865 ;
        RECT 65.390 165.485 66.405 165.685 ;
        RECT 62.680 165.055 63.930 165.225 ;
        RECT 62.680 164.935 63.010 165.055 ;
        RECT 61.340 164.545 63.240 164.715 ;
        RECT 60.980 164.205 62.900 164.375 ;
        RECT 60.980 164.185 61.300 164.205 ;
        RECT 60.530 163.525 60.860 164.035 ;
        RECT 61.130 163.575 61.300 164.185 ;
        RECT 63.070 164.035 63.240 164.545 ;
        RECT 63.410 164.475 63.590 164.885 ;
        RECT 63.760 164.295 63.930 165.055 ;
        RECT 61.470 163.315 61.800 164.005 ;
        RECT 62.030 163.865 63.240 164.035 ;
        RECT 63.410 163.985 63.930 164.295 ;
        RECT 64.100 164.885 64.520 165.225 ;
        RECT 64.810 164.885 65.220 165.215 ;
        RECT 64.100 164.115 64.290 164.885 ;
        RECT 65.390 164.755 65.560 165.485 ;
        RECT 66.705 165.315 66.875 165.645 ;
        RECT 67.045 165.485 67.375 165.865 ;
        RECT 65.730 164.935 66.080 165.305 ;
        RECT 65.390 164.715 65.810 164.755 ;
        RECT 64.460 164.545 65.810 164.715 ;
        RECT 64.460 164.385 64.710 164.545 ;
        RECT 65.220 164.115 65.470 164.375 ;
        RECT 64.100 163.865 65.470 164.115 ;
        RECT 62.030 163.575 62.270 163.865 ;
        RECT 63.070 163.785 63.240 163.865 ;
        RECT 62.470 163.315 62.890 163.695 ;
        RECT 63.070 163.535 63.700 163.785 ;
        RECT 64.170 163.315 64.500 163.695 ;
        RECT 64.670 163.575 64.840 163.865 ;
        RECT 65.640 163.700 65.810 164.545 ;
        RECT 66.260 164.375 66.480 165.245 ;
        RECT 66.705 165.125 67.400 165.315 ;
        RECT 65.980 163.995 66.480 164.375 ;
        RECT 66.650 164.325 67.060 164.945 ;
        RECT 67.230 164.155 67.400 165.125 ;
        RECT 66.705 163.985 67.400 164.155 ;
        RECT 65.020 163.315 65.400 163.695 ;
        RECT 65.640 163.530 66.470 163.700 ;
        RECT 66.705 163.485 66.875 163.985 ;
        RECT 67.045 163.315 67.375 163.815 ;
        RECT 67.590 163.485 67.815 165.605 ;
        RECT 67.985 165.485 68.315 165.865 ;
        RECT 68.485 165.315 68.655 165.605 ;
        RECT 67.990 165.145 68.655 165.315 ;
        RECT 67.990 164.155 68.220 165.145 ;
        RECT 68.920 165.025 69.180 165.865 ;
        RECT 69.355 165.120 69.610 165.695 ;
        RECT 69.780 165.485 70.110 165.865 ;
        RECT 70.325 165.315 70.495 165.695 ;
        RECT 69.780 165.145 70.495 165.315 ;
        RECT 68.390 164.325 68.740 164.975 ;
        RECT 67.990 163.985 68.655 164.155 ;
        RECT 67.985 163.315 68.315 163.815 ;
        RECT 68.485 163.485 68.655 163.985 ;
        RECT 68.920 163.315 69.180 164.465 ;
        RECT 69.355 164.390 69.525 165.120 ;
        RECT 69.780 164.955 69.950 165.145 ;
        RECT 70.755 165.065 71.095 165.695 ;
        RECT 71.265 165.065 71.515 165.865 ;
        RECT 71.705 165.215 72.035 165.695 ;
        RECT 72.205 165.405 72.430 165.865 ;
        RECT 72.600 165.215 72.930 165.695 ;
        RECT 70.755 165.015 70.985 165.065 ;
        RECT 71.705 165.045 72.930 165.215 ;
        RECT 73.560 165.085 74.060 165.695 ;
        RECT 74.435 165.140 74.725 165.865 ;
        RECT 69.695 164.625 69.950 164.955 ;
        RECT 69.780 164.415 69.950 164.625 ;
        RECT 70.230 164.595 70.585 164.965 ;
        RECT 70.755 164.455 70.930 165.015 ;
        RECT 71.100 164.705 71.795 164.875 ;
        RECT 71.625 164.455 71.795 164.705 ;
        RECT 71.970 164.675 72.390 164.875 ;
        RECT 72.560 164.675 72.890 164.875 ;
        RECT 73.060 164.675 73.390 164.875 ;
        RECT 73.560 164.455 73.730 165.085 ;
        RECT 74.900 165.025 75.160 165.865 ;
        RECT 75.335 165.120 75.590 165.695 ;
        RECT 75.760 165.485 76.090 165.865 ;
        RECT 76.305 165.315 76.475 165.695 ;
        RECT 75.760 165.145 76.475 165.315 ;
        RECT 73.915 164.625 74.265 164.875 ;
        RECT 69.355 163.485 69.610 164.390 ;
        RECT 69.780 164.245 70.495 164.415 ;
        RECT 69.780 163.315 70.110 164.075 ;
        RECT 70.325 163.485 70.495 164.245 ;
        RECT 70.755 163.485 71.095 164.455 ;
        RECT 71.265 163.315 71.435 164.455 ;
        RECT 71.625 164.285 74.060 164.455 ;
        RECT 71.705 163.315 71.955 164.115 ;
        RECT 72.600 163.485 72.930 164.285 ;
        RECT 73.230 163.315 73.560 164.115 ;
        RECT 73.730 163.485 74.060 164.285 ;
        RECT 74.435 163.315 74.725 164.480 ;
        RECT 74.900 163.315 75.160 164.465 ;
        RECT 75.335 164.390 75.505 165.120 ;
        RECT 75.760 164.955 75.930 165.145 ;
        RECT 76.795 165.045 77.005 165.865 ;
        RECT 77.175 165.065 77.505 165.695 ;
        RECT 75.675 164.625 75.930 164.955 ;
        RECT 75.760 164.415 75.930 164.625 ;
        RECT 76.210 164.595 76.565 164.965 ;
        RECT 77.175 164.465 77.425 165.065 ;
        RECT 77.675 165.045 77.905 165.865 ;
        RECT 78.390 165.055 78.635 165.660 ;
        RECT 78.855 165.330 79.365 165.865 ;
        RECT 78.115 164.885 79.345 165.055 ;
        RECT 77.595 164.625 77.925 164.875 ;
        RECT 75.335 163.485 75.590 164.390 ;
        RECT 75.760 164.245 76.475 164.415 ;
        RECT 75.760 163.315 76.090 164.075 ;
        RECT 76.305 163.485 76.475 164.245 ;
        RECT 76.795 163.315 77.005 164.455 ;
        RECT 77.175 163.485 77.505 164.465 ;
        RECT 77.675 163.315 77.905 164.455 ;
        RECT 78.115 164.075 78.455 164.885 ;
        RECT 78.625 164.320 79.375 164.510 ;
        RECT 78.115 163.665 78.630 164.075 ;
        RECT 78.865 163.315 79.035 164.075 ;
        RECT 79.205 163.655 79.375 164.320 ;
        RECT 79.545 164.335 79.735 165.695 ;
        RECT 79.905 164.845 80.180 165.695 ;
        RECT 80.370 165.330 80.900 165.695 ;
        RECT 81.325 165.465 81.655 165.865 ;
        RECT 80.725 165.295 80.900 165.330 ;
        RECT 79.905 164.675 80.185 164.845 ;
        RECT 79.905 164.535 80.180 164.675 ;
        RECT 80.385 164.335 80.555 165.135 ;
        RECT 79.545 164.165 80.555 164.335 ;
        RECT 80.725 165.125 81.655 165.295 ;
        RECT 81.825 165.125 82.080 165.695 ;
        RECT 82.345 165.315 82.515 165.695 ;
        RECT 82.695 165.485 83.025 165.865 ;
        RECT 82.345 165.145 83.010 165.315 ;
        RECT 83.205 165.190 83.465 165.695 ;
        RECT 80.725 163.995 80.895 165.125 ;
        RECT 81.485 164.955 81.655 165.125 ;
        RECT 79.770 163.825 80.895 163.995 ;
        RECT 81.065 164.625 81.260 164.955 ;
        RECT 81.485 164.625 81.740 164.955 ;
        RECT 81.065 163.655 81.235 164.625 ;
        RECT 81.910 164.455 82.080 165.125 ;
        RECT 82.275 164.595 82.605 164.965 ;
        RECT 82.840 164.890 83.010 165.145 ;
        RECT 79.205 163.485 81.235 163.655 ;
        RECT 81.405 163.315 81.575 164.455 ;
        RECT 81.745 163.485 82.080 164.455 ;
        RECT 82.840 164.560 83.125 164.890 ;
        RECT 82.840 164.415 83.010 164.560 ;
        RECT 82.345 164.245 83.010 164.415 ;
        RECT 83.295 164.390 83.465 165.190 ;
        RECT 84.595 165.045 84.825 165.865 ;
        RECT 84.995 165.065 85.325 165.695 ;
        RECT 84.575 164.625 84.905 164.875 ;
        RECT 85.075 164.465 85.325 165.065 ;
        RECT 85.495 165.045 85.705 165.865 ;
        RECT 86.025 165.315 86.195 165.695 ;
        RECT 86.375 165.485 86.705 165.865 ;
        RECT 86.025 165.145 86.690 165.315 ;
        RECT 86.885 165.190 87.145 165.695 ;
        RECT 85.955 164.595 86.285 164.965 ;
        RECT 86.520 164.890 86.690 165.145 ;
        RECT 82.345 163.485 82.515 164.245 ;
        RECT 82.695 163.315 83.025 164.075 ;
        RECT 83.195 163.485 83.465 164.390 ;
        RECT 84.595 163.315 84.825 164.455 ;
        RECT 84.995 163.485 85.325 164.465 ;
        RECT 86.520 164.560 86.805 164.890 ;
        RECT 85.495 163.315 85.705 164.455 ;
        RECT 86.520 164.415 86.690 164.560 ;
        RECT 86.025 164.245 86.690 164.415 ;
        RECT 86.975 164.390 87.145 165.190 ;
        RECT 86.025 163.485 86.195 164.245 ;
        RECT 86.375 163.315 86.705 164.075 ;
        RECT 86.875 163.485 87.145 164.390 ;
        RECT 87.315 165.190 87.585 165.535 ;
        RECT 87.775 165.465 88.155 165.865 ;
        RECT 88.325 165.295 88.495 165.645 ;
        RECT 88.665 165.465 88.995 165.865 ;
        RECT 89.195 165.295 89.365 165.645 ;
        RECT 89.565 165.365 89.895 165.865 ;
        RECT 87.315 164.455 87.485 165.190 ;
        RECT 87.755 165.125 89.365 165.295 ;
        RECT 87.755 164.955 87.925 165.125 ;
        RECT 87.655 164.625 87.925 164.955 ;
        RECT 88.095 164.625 88.500 164.955 ;
        RECT 87.755 164.455 87.925 164.625 ;
        RECT 88.670 164.505 89.380 164.955 ;
        RECT 89.550 164.625 89.900 165.195 ;
        RECT 90.075 165.065 90.415 165.695 ;
        RECT 90.585 165.065 90.835 165.865 ;
        RECT 91.025 165.215 91.355 165.695 ;
        RECT 91.525 165.405 91.750 165.865 ;
        RECT 91.920 165.215 92.250 165.695 ;
        RECT 87.315 163.485 87.585 164.455 ;
        RECT 87.755 164.285 88.480 164.455 ;
        RECT 88.670 164.335 89.385 164.505 ;
        RECT 90.075 164.455 90.250 165.065 ;
        RECT 91.025 165.045 92.250 165.215 ;
        RECT 92.880 165.085 93.380 165.695 ;
        RECT 90.420 164.705 91.115 164.875 ;
        RECT 90.945 164.455 91.115 164.705 ;
        RECT 91.290 164.675 91.710 164.875 ;
        RECT 91.880 164.675 92.210 164.875 ;
        RECT 92.380 164.675 92.710 164.875 ;
        RECT 92.880 164.455 93.050 165.085 ;
        RECT 93.755 165.065 94.095 165.695 ;
        RECT 94.265 165.065 94.515 165.865 ;
        RECT 94.705 165.215 95.035 165.695 ;
        RECT 95.205 165.405 95.430 165.865 ;
        RECT 95.600 165.215 95.930 165.695 ;
        RECT 93.235 164.625 93.585 164.875 ;
        RECT 93.755 164.455 93.930 165.065 ;
        RECT 94.705 165.045 95.930 165.215 ;
        RECT 96.560 165.085 97.060 165.695 ;
        RECT 97.435 165.190 97.705 165.535 ;
        RECT 97.895 165.465 98.275 165.865 ;
        RECT 98.445 165.295 98.615 165.645 ;
        RECT 98.785 165.465 99.115 165.865 ;
        RECT 99.315 165.295 99.485 165.645 ;
        RECT 99.685 165.365 100.015 165.865 ;
        RECT 94.100 164.705 94.795 164.875 ;
        RECT 94.625 164.455 94.795 164.705 ;
        RECT 94.970 164.675 95.390 164.875 ;
        RECT 95.560 164.675 95.890 164.875 ;
        RECT 96.060 164.675 96.390 164.875 ;
        RECT 96.560 164.455 96.730 165.085 ;
        RECT 96.915 164.625 97.265 164.875 ;
        RECT 97.435 164.455 97.605 165.190 ;
        RECT 97.875 165.125 99.485 165.295 ;
        RECT 97.875 164.955 98.045 165.125 ;
        RECT 97.775 164.625 98.045 164.955 ;
        RECT 98.215 164.625 98.620 164.955 ;
        RECT 97.875 164.455 98.045 164.625 ;
        RECT 98.790 164.505 99.500 164.955 ;
        RECT 99.670 164.625 100.020 165.195 ;
        RECT 100.195 165.140 100.485 165.865 ;
        RECT 100.655 165.190 100.915 165.695 ;
        RECT 101.095 165.485 101.425 165.865 ;
        RECT 101.605 165.315 101.775 165.695 ;
        RECT 88.310 164.165 88.480 164.285 ;
        RECT 89.580 164.165 89.900 164.455 ;
        RECT 87.795 163.315 88.075 164.115 ;
        RECT 88.310 163.995 89.900 164.165 ;
        RECT 88.245 163.535 89.900 163.825 ;
        RECT 90.075 163.485 90.415 164.455 ;
        RECT 90.585 163.315 90.755 164.455 ;
        RECT 90.945 164.285 93.380 164.455 ;
        RECT 91.025 163.315 91.275 164.115 ;
        RECT 91.920 163.485 92.250 164.285 ;
        RECT 92.550 163.315 92.880 164.115 ;
        RECT 93.050 163.485 93.380 164.285 ;
        RECT 93.755 163.485 94.095 164.455 ;
        RECT 94.265 163.315 94.435 164.455 ;
        RECT 94.625 164.285 97.060 164.455 ;
        RECT 94.705 163.315 94.955 164.115 ;
        RECT 95.600 163.485 95.930 164.285 ;
        RECT 96.230 163.315 96.560 164.115 ;
        RECT 96.730 163.485 97.060 164.285 ;
        RECT 97.435 163.485 97.705 164.455 ;
        RECT 97.875 164.285 98.600 164.455 ;
        RECT 98.790 164.335 99.505 164.505 ;
        RECT 98.430 164.165 98.600 164.285 ;
        RECT 99.700 164.165 100.020 164.455 ;
        RECT 97.915 163.315 98.195 164.115 ;
        RECT 98.430 163.995 100.020 164.165 ;
        RECT 98.365 163.535 100.020 163.825 ;
        RECT 100.195 163.315 100.485 164.480 ;
        RECT 100.655 164.390 100.825 165.190 ;
        RECT 101.110 165.145 101.775 165.315 ;
        RECT 102.870 165.155 103.125 165.685 ;
        RECT 103.305 165.405 103.590 165.865 ;
        RECT 101.110 164.890 101.280 165.145 ;
        RECT 100.995 164.560 101.280 164.890 ;
        RECT 101.515 164.595 101.845 164.965 ;
        RECT 101.110 164.415 101.280 164.560 ;
        RECT 100.655 163.485 100.925 164.390 ;
        RECT 101.110 164.245 101.775 164.415 ;
        RECT 101.095 163.315 101.425 164.075 ;
        RECT 101.605 163.485 101.775 164.245 ;
        RECT 102.870 164.295 103.050 165.155 ;
        RECT 103.770 164.955 104.020 165.605 ;
        RECT 103.220 164.625 104.020 164.955 ;
        RECT 102.870 163.825 103.125 164.295 ;
        RECT 102.785 163.655 103.125 163.825 ;
        RECT 102.870 163.625 103.125 163.655 ;
        RECT 103.305 163.315 103.590 164.115 ;
        RECT 103.770 164.035 104.020 164.625 ;
        RECT 104.220 165.270 104.540 165.600 ;
        RECT 104.720 165.385 105.380 165.865 ;
        RECT 105.580 165.475 106.430 165.645 ;
        RECT 104.220 164.375 104.410 165.270 ;
        RECT 104.730 164.945 105.390 165.215 ;
        RECT 105.060 164.885 105.390 164.945 ;
        RECT 104.580 164.715 104.910 164.775 ;
        RECT 105.580 164.715 105.750 165.475 ;
        RECT 106.990 165.405 107.310 165.865 ;
        RECT 107.510 165.225 107.760 165.655 ;
        RECT 108.050 165.425 108.460 165.865 ;
        RECT 108.630 165.485 109.645 165.685 ;
        RECT 105.920 165.055 107.170 165.225 ;
        RECT 105.920 164.935 106.250 165.055 ;
        RECT 104.580 164.545 106.480 164.715 ;
        RECT 104.220 164.205 106.140 164.375 ;
        RECT 104.220 164.185 104.540 164.205 ;
        RECT 103.770 163.525 104.100 164.035 ;
        RECT 104.370 163.575 104.540 164.185 ;
        RECT 106.310 164.035 106.480 164.545 ;
        RECT 106.650 164.475 106.830 164.885 ;
        RECT 107.000 164.295 107.170 165.055 ;
        RECT 104.710 163.315 105.040 164.005 ;
        RECT 105.270 163.865 106.480 164.035 ;
        RECT 106.650 163.985 107.170 164.295 ;
        RECT 107.340 164.885 107.760 165.225 ;
        RECT 108.050 164.885 108.460 165.215 ;
        RECT 107.340 164.115 107.530 164.885 ;
        RECT 108.630 164.755 108.800 165.485 ;
        RECT 109.945 165.315 110.115 165.645 ;
        RECT 110.285 165.485 110.615 165.865 ;
        RECT 108.970 164.935 109.320 165.305 ;
        RECT 108.630 164.715 109.050 164.755 ;
        RECT 107.700 164.545 109.050 164.715 ;
        RECT 107.700 164.385 107.950 164.545 ;
        RECT 108.460 164.115 108.710 164.375 ;
        RECT 107.340 163.865 108.710 164.115 ;
        RECT 105.270 163.575 105.510 163.865 ;
        RECT 106.310 163.785 106.480 163.865 ;
        RECT 105.710 163.315 106.130 163.695 ;
        RECT 106.310 163.535 106.940 163.785 ;
        RECT 107.410 163.315 107.740 163.695 ;
        RECT 107.910 163.575 108.080 163.865 ;
        RECT 108.880 163.700 109.050 164.545 ;
        RECT 109.500 164.375 109.720 165.245 ;
        RECT 109.945 165.125 110.640 165.315 ;
        RECT 109.220 163.995 109.720 164.375 ;
        RECT 109.890 164.325 110.300 164.945 ;
        RECT 110.470 164.155 110.640 165.125 ;
        RECT 109.945 163.985 110.640 164.155 ;
        RECT 108.260 163.315 108.640 163.695 ;
        RECT 108.880 163.530 109.710 163.700 ;
        RECT 109.945 163.485 110.115 163.985 ;
        RECT 110.285 163.315 110.615 163.815 ;
        RECT 110.830 163.485 111.055 165.605 ;
        RECT 111.225 165.485 111.555 165.865 ;
        RECT 111.725 165.315 111.895 165.605 ;
        RECT 111.230 165.145 111.895 165.315 ;
        RECT 111.230 164.155 111.460 165.145 ;
        RECT 112.155 165.115 113.365 165.865 ;
        RECT 111.630 164.325 111.980 164.975 ;
        RECT 112.155 164.405 112.675 164.945 ;
        RECT 112.845 164.575 113.365 165.115 ;
        RECT 111.230 163.985 111.895 164.155 ;
        RECT 111.225 163.315 111.555 163.815 ;
        RECT 111.725 163.485 111.895 163.985 ;
        RECT 112.155 163.315 113.365 164.405 ;
        RECT 26.970 163.145 113.450 163.315 ;
        RECT 27.055 162.055 28.265 163.145 ;
        RECT 29.555 162.475 29.835 163.145 ;
        RECT 30.005 162.255 30.305 162.805 ;
        RECT 30.505 162.425 30.835 163.145 ;
        RECT 31.025 162.425 31.485 162.975 ;
        RECT 27.055 161.345 27.575 161.885 ;
        RECT 27.745 161.515 28.265 162.055 ;
        RECT 29.370 161.835 29.635 162.195 ;
        RECT 30.005 162.085 30.945 162.255 ;
        RECT 30.775 161.835 30.945 162.085 ;
        RECT 29.370 161.585 30.045 161.835 ;
        RECT 30.265 161.585 30.605 161.835 ;
        RECT 30.775 161.505 31.065 161.835 ;
        RECT 30.775 161.415 30.945 161.505 ;
        RECT 27.055 160.595 28.265 161.345 ;
        RECT 29.555 161.225 30.945 161.415 ;
        RECT 29.555 160.865 29.885 161.225 ;
        RECT 31.235 161.055 31.485 162.425 ;
        RECT 31.655 162.385 32.170 162.795 ;
        RECT 32.405 162.385 32.575 163.145 ;
        RECT 32.745 162.805 34.775 162.975 ;
        RECT 31.655 161.575 31.995 162.385 ;
        RECT 32.745 162.140 32.915 162.805 ;
        RECT 33.310 162.465 34.435 162.635 ;
        RECT 32.165 161.950 32.915 162.140 ;
        RECT 33.085 162.125 34.095 162.295 ;
        RECT 31.655 161.405 32.885 161.575 ;
        RECT 30.505 160.595 30.755 161.055 ;
        RECT 30.925 160.765 31.485 161.055 ;
        RECT 31.930 160.800 32.175 161.405 ;
        RECT 32.395 160.595 32.905 161.130 ;
        RECT 33.085 160.765 33.275 162.125 ;
        RECT 33.445 161.105 33.720 161.925 ;
        RECT 33.925 161.325 34.095 162.125 ;
        RECT 34.265 161.335 34.435 162.465 ;
        RECT 34.605 161.835 34.775 162.805 ;
        RECT 34.945 162.005 35.115 163.145 ;
        RECT 35.285 162.005 35.620 162.975 ;
        RECT 34.605 161.505 34.800 161.835 ;
        RECT 35.025 161.505 35.280 161.835 ;
        RECT 35.025 161.335 35.195 161.505 ;
        RECT 35.450 161.335 35.620 162.005 ;
        RECT 35.795 161.980 36.085 163.145 ;
        RECT 36.345 162.475 36.515 162.975 ;
        RECT 36.685 162.645 37.015 163.145 ;
        RECT 36.345 162.305 37.010 162.475 ;
        RECT 36.260 161.485 36.610 162.135 ;
        RECT 34.265 161.165 35.195 161.335 ;
        RECT 34.265 161.130 34.440 161.165 ;
        RECT 33.445 160.935 33.725 161.105 ;
        RECT 33.445 160.765 33.720 160.935 ;
        RECT 33.910 160.765 34.440 161.130 ;
        RECT 34.865 160.595 35.195 160.995 ;
        RECT 35.365 160.765 35.620 161.335 ;
        RECT 35.795 160.595 36.085 161.320 ;
        RECT 36.780 161.315 37.010 162.305 ;
        RECT 36.345 161.145 37.010 161.315 ;
        RECT 36.345 160.855 36.515 161.145 ;
        RECT 36.685 160.595 37.015 160.975 ;
        RECT 37.185 160.855 37.410 162.975 ;
        RECT 37.625 162.645 37.955 163.145 ;
        RECT 38.125 162.475 38.295 162.975 ;
        RECT 38.530 162.760 39.360 162.930 ;
        RECT 39.600 162.765 39.980 163.145 ;
        RECT 37.600 162.305 38.295 162.475 ;
        RECT 37.600 161.335 37.770 162.305 ;
        RECT 37.940 161.515 38.350 162.135 ;
        RECT 38.520 162.085 39.020 162.465 ;
        RECT 37.600 161.145 38.295 161.335 ;
        RECT 38.520 161.215 38.740 162.085 ;
        RECT 39.190 161.915 39.360 162.760 ;
        RECT 40.160 162.595 40.330 162.885 ;
        RECT 40.500 162.765 40.830 163.145 ;
        RECT 41.300 162.675 41.930 162.925 ;
        RECT 42.110 162.765 42.530 163.145 ;
        RECT 41.760 162.595 41.930 162.675 ;
        RECT 42.730 162.595 42.970 162.885 ;
        RECT 39.530 162.345 40.900 162.595 ;
        RECT 39.530 162.085 39.780 162.345 ;
        RECT 40.290 161.915 40.540 162.075 ;
        RECT 39.190 161.745 40.540 161.915 ;
        RECT 39.190 161.705 39.610 161.745 ;
        RECT 38.920 161.155 39.270 161.525 ;
        RECT 37.625 160.595 37.955 160.975 ;
        RECT 38.125 160.815 38.295 161.145 ;
        RECT 39.440 160.975 39.610 161.705 ;
        RECT 40.710 161.575 40.900 162.345 ;
        RECT 39.780 161.245 40.190 161.575 ;
        RECT 40.480 161.235 40.900 161.575 ;
        RECT 41.070 162.165 41.590 162.475 ;
        RECT 41.760 162.425 42.970 162.595 ;
        RECT 43.200 162.455 43.530 163.145 ;
        RECT 41.070 161.405 41.240 162.165 ;
        RECT 41.410 161.575 41.590 161.985 ;
        RECT 41.760 161.915 41.930 162.425 ;
        RECT 43.700 162.275 43.870 162.885 ;
        RECT 44.140 162.425 44.470 162.935 ;
        RECT 43.700 162.255 44.020 162.275 ;
        RECT 42.100 162.085 44.020 162.255 ;
        RECT 41.760 161.745 43.660 161.915 ;
        RECT 41.990 161.405 42.320 161.525 ;
        RECT 41.070 161.235 42.320 161.405 ;
        RECT 38.595 160.775 39.610 160.975 ;
        RECT 39.780 160.595 40.190 161.035 ;
        RECT 40.480 160.805 40.730 161.235 ;
        RECT 40.930 160.595 41.250 161.055 ;
        RECT 42.490 160.985 42.660 161.745 ;
        RECT 43.330 161.685 43.660 161.745 ;
        RECT 42.850 161.515 43.180 161.575 ;
        RECT 42.850 161.245 43.510 161.515 ;
        RECT 43.830 161.190 44.020 162.085 ;
        RECT 41.810 160.815 42.660 160.985 ;
        RECT 42.860 160.595 43.520 161.075 ;
        RECT 43.700 160.860 44.020 161.190 ;
        RECT 44.220 161.835 44.470 162.425 ;
        RECT 44.650 162.345 44.935 163.145 ;
        RECT 45.115 162.165 45.370 162.835 ;
        RECT 44.220 161.505 45.020 161.835 ;
        RECT 44.220 160.855 44.470 161.505 ;
        RECT 45.190 161.305 45.370 162.165 ;
        RECT 45.115 161.105 45.370 161.305 ;
        RECT 45.915 162.005 46.255 162.975 ;
        RECT 46.425 162.005 46.595 163.145 ;
        RECT 46.865 162.345 47.115 163.145 ;
        RECT 47.760 162.175 48.090 162.975 ;
        RECT 48.390 162.345 48.720 163.145 ;
        RECT 48.890 162.175 49.220 162.975 ;
        RECT 46.785 162.005 49.220 162.175 ;
        RECT 50.055 162.005 50.395 162.975 ;
        RECT 50.565 162.005 50.735 163.145 ;
        RECT 51.005 162.345 51.255 163.145 ;
        RECT 51.900 162.175 52.230 162.975 ;
        RECT 52.530 162.345 52.860 163.145 ;
        RECT 53.030 162.175 53.360 162.975 ;
        RECT 50.925 162.005 53.360 162.175 ;
        RECT 53.775 162.005 54.005 163.145 ;
        RECT 45.915 161.955 46.145 162.005 ;
        RECT 45.915 161.395 46.090 161.955 ;
        RECT 46.785 161.755 46.955 162.005 ;
        RECT 46.260 161.585 46.955 161.755 ;
        RECT 47.130 161.585 47.550 161.785 ;
        RECT 47.720 161.585 48.050 161.785 ;
        RECT 48.220 161.585 48.550 161.785 ;
        RECT 44.650 160.595 44.935 161.055 ;
        RECT 45.115 160.935 45.455 161.105 ;
        RECT 45.115 160.775 45.370 160.935 ;
        RECT 45.915 160.765 46.255 161.395 ;
        RECT 46.425 160.595 46.675 161.395 ;
        RECT 46.865 161.245 48.090 161.415 ;
        RECT 46.865 160.765 47.195 161.245 ;
        RECT 47.365 160.595 47.590 161.055 ;
        RECT 47.760 160.765 48.090 161.245 ;
        RECT 48.720 161.375 48.890 162.005 ;
        RECT 49.075 161.585 49.425 161.835 ;
        RECT 50.055 161.395 50.230 162.005 ;
        RECT 50.925 161.755 51.095 162.005 ;
        RECT 50.400 161.585 51.095 161.755 ;
        RECT 51.270 161.585 51.690 161.785 ;
        RECT 51.860 161.585 52.190 161.785 ;
        RECT 52.360 161.585 52.690 161.785 ;
        RECT 48.720 160.765 49.220 161.375 ;
        RECT 50.055 160.765 50.395 161.395 ;
        RECT 50.565 160.595 50.815 161.395 ;
        RECT 51.005 161.245 52.230 161.415 ;
        RECT 51.005 160.765 51.335 161.245 ;
        RECT 51.505 160.595 51.730 161.055 ;
        RECT 51.900 160.765 52.230 161.245 ;
        RECT 52.860 161.375 53.030 162.005 ;
        RECT 54.175 161.995 54.505 162.975 ;
        RECT 54.675 162.005 54.885 163.145 ;
        RECT 56.075 162.005 56.305 163.145 ;
        RECT 56.475 161.995 56.805 162.975 ;
        RECT 56.975 162.005 57.185 163.145 ;
        RECT 57.415 162.005 57.755 162.975 ;
        RECT 57.925 162.005 58.095 163.145 ;
        RECT 58.365 162.345 58.615 163.145 ;
        RECT 59.260 162.175 59.590 162.975 ;
        RECT 59.890 162.345 60.220 163.145 ;
        RECT 60.390 162.175 60.720 162.975 ;
        RECT 58.285 162.005 60.720 162.175 ;
        RECT 53.215 161.585 53.565 161.835 ;
        RECT 53.755 161.585 54.085 161.835 ;
        RECT 52.860 160.765 53.360 161.375 ;
        RECT 53.775 160.595 54.005 161.415 ;
        RECT 54.255 161.395 54.505 161.995 ;
        RECT 56.055 161.585 56.385 161.835 ;
        RECT 54.175 160.765 54.505 161.395 ;
        RECT 54.675 160.595 54.885 161.415 ;
        RECT 56.075 160.595 56.305 161.415 ;
        RECT 56.555 161.395 56.805 161.995 ;
        RECT 56.475 160.765 56.805 161.395 ;
        RECT 56.975 160.595 57.185 161.415 ;
        RECT 57.415 161.395 57.590 162.005 ;
        RECT 58.285 161.755 58.455 162.005 ;
        RECT 57.760 161.585 58.455 161.755 ;
        RECT 58.630 161.585 59.050 161.785 ;
        RECT 59.220 161.585 59.550 161.785 ;
        RECT 59.720 161.585 60.050 161.785 ;
        RECT 57.415 160.765 57.755 161.395 ;
        RECT 57.925 160.595 58.175 161.395 ;
        RECT 58.365 161.245 59.590 161.415 ;
        RECT 58.365 160.765 58.695 161.245 ;
        RECT 58.865 160.595 59.090 161.055 ;
        RECT 59.260 160.765 59.590 161.245 ;
        RECT 60.220 161.375 60.390 162.005 ;
        RECT 61.555 161.980 61.845 163.145 ;
        RECT 62.105 162.400 62.375 163.145 ;
        RECT 63.005 163.140 69.280 163.145 ;
        RECT 62.545 162.230 62.835 162.970 ;
        RECT 63.005 162.415 63.260 163.140 ;
        RECT 63.445 162.245 63.705 162.970 ;
        RECT 63.875 162.415 64.120 163.140 ;
        RECT 64.305 162.245 64.565 162.970 ;
        RECT 64.735 162.415 64.980 163.140 ;
        RECT 65.165 162.245 65.425 162.970 ;
        RECT 65.595 162.415 65.840 163.140 ;
        RECT 66.010 162.245 66.270 162.970 ;
        RECT 66.440 162.415 66.700 163.140 ;
        RECT 66.870 162.245 67.130 162.970 ;
        RECT 67.300 162.415 67.560 163.140 ;
        RECT 67.730 162.245 67.990 162.970 ;
        RECT 68.160 162.415 68.420 163.140 ;
        RECT 68.590 162.245 68.850 162.970 ;
        RECT 69.020 162.345 69.280 163.140 ;
        RECT 63.445 162.230 68.850 162.245 ;
        RECT 62.105 162.005 68.850 162.230 ;
        RECT 60.575 161.585 60.925 161.835 ;
        RECT 62.105 161.415 63.270 162.005 ;
        RECT 69.450 161.835 69.700 162.970 ;
        RECT 69.880 162.335 70.140 163.145 ;
        RECT 70.315 161.835 70.560 162.975 ;
        RECT 70.740 162.335 71.035 163.145 ;
        RECT 72.145 162.085 72.475 163.145 ;
        RECT 72.655 161.835 72.825 162.805 ;
        RECT 72.995 162.555 73.325 162.955 ;
        RECT 73.495 162.785 73.825 163.145 ;
        RECT 74.025 162.555 74.725 162.975 ;
        RECT 72.995 162.325 74.725 162.555 ;
        RECT 72.995 162.105 73.325 162.325 ;
        RECT 73.520 161.835 73.845 162.125 ;
        RECT 63.440 161.585 70.560 161.835 ;
        RECT 60.220 160.765 60.720 161.375 ;
        RECT 61.555 160.595 61.845 161.320 ;
        RECT 62.105 161.245 68.850 161.415 ;
        RECT 62.105 160.595 62.405 161.075 ;
        RECT 62.575 160.790 62.835 161.245 ;
        RECT 63.005 160.595 63.265 161.075 ;
        RECT 63.445 160.790 63.705 161.245 ;
        RECT 63.875 160.595 64.125 161.075 ;
        RECT 64.305 160.790 64.565 161.245 ;
        RECT 64.735 160.595 64.985 161.075 ;
        RECT 65.165 160.790 65.425 161.245 ;
        RECT 65.595 160.595 65.840 161.075 ;
        RECT 66.010 160.790 66.285 161.245 ;
        RECT 66.455 160.595 66.700 161.075 ;
        RECT 66.870 160.790 67.130 161.245 ;
        RECT 67.300 160.595 67.560 161.075 ;
        RECT 67.730 160.790 67.990 161.245 ;
        RECT 68.160 160.595 68.420 161.075 ;
        RECT 68.590 160.790 68.850 161.245 ;
        RECT 69.020 160.595 69.280 161.155 ;
        RECT 69.450 160.775 69.700 161.585 ;
        RECT 69.880 160.595 70.140 161.120 ;
        RECT 70.310 160.775 70.560 161.585 ;
        RECT 70.730 161.275 71.045 161.835 ;
        RECT 72.135 161.505 72.445 161.835 ;
        RECT 72.655 161.505 73.030 161.835 ;
        RECT 73.350 161.505 73.845 161.835 ;
        RECT 74.020 161.585 74.350 162.125 ;
        RECT 74.520 161.355 74.725 162.325 ;
        RECT 72.145 161.125 73.505 161.335 ;
        RECT 70.740 160.595 71.045 161.105 ;
        RECT 72.145 160.765 72.475 161.125 ;
        RECT 72.645 160.595 72.975 160.955 ;
        RECT 73.175 160.765 73.505 161.125 ;
        RECT 74.015 160.765 74.725 161.355 ;
        RECT 74.895 162.005 75.235 162.975 ;
        RECT 75.405 162.005 75.575 163.145 ;
        RECT 75.845 162.345 76.095 163.145 ;
        RECT 76.740 162.175 77.070 162.975 ;
        RECT 77.370 162.345 77.700 163.145 ;
        RECT 77.870 162.175 78.200 162.975 ;
        RECT 75.765 162.005 78.200 162.175 ;
        RECT 79.075 162.005 79.305 163.145 ;
        RECT 74.895 161.395 75.070 162.005 ;
        RECT 75.765 161.755 75.935 162.005 ;
        RECT 75.240 161.585 75.935 161.755 ;
        RECT 76.110 161.585 76.530 161.785 ;
        RECT 76.700 161.585 77.030 161.785 ;
        RECT 77.200 161.585 77.530 161.785 ;
        RECT 74.895 160.765 75.235 161.395 ;
        RECT 75.405 160.595 75.655 161.395 ;
        RECT 75.845 161.245 77.070 161.415 ;
        RECT 75.845 160.765 76.175 161.245 ;
        RECT 76.345 160.595 76.570 161.055 ;
        RECT 76.740 160.765 77.070 161.245 ;
        RECT 77.700 161.375 77.870 162.005 ;
        RECT 79.475 161.995 79.805 162.975 ;
        RECT 79.975 162.005 80.185 163.145 ;
        RECT 80.475 162.005 80.685 163.145 ;
        RECT 78.055 161.585 78.405 161.835 ;
        RECT 79.055 161.585 79.385 161.835 ;
        RECT 77.700 160.765 78.200 161.375 ;
        RECT 79.075 160.595 79.305 161.415 ;
        RECT 79.555 161.395 79.805 161.995 ;
        RECT 80.855 161.995 81.185 162.975 ;
        RECT 81.355 162.005 81.585 163.145 ;
        RECT 81.835 162.005 82.065 163.145 ;
        RECT 82.235 161.995 82.565 162.975 ;
        RECT 82.735 162.005 82.945 163.145 ;
        RECT 83.175 162.385 83.690 162.795 ;
        RECT 83.925 162.385 84.095 163.145 ;
        RECT 84.265 162.805 86.295 162.975 ;
        RECT 79.475 160.765 79.805 161.395 ;
        RECT 79.975 160.595 80.185 161.415 ;
        RECT 80.475 160.595 80.685 161.415 ;
        RECT 80.855 161.395 81.105 161.995 ;
        RECT 81.275 161.585 81.605 161.835 ;
        RECT 81.815 161.585 82.145 161.835 ;
        RECT 80.855 160.765 81.185 161.395 ;
        RECT 81.355 160.595 81.585 161.415 ;
        RECT 81.835 160.595 82.065 161.415 ;
        RECT 82.315 161.395 82.565 161.995 ;
        RECT 83.175 161.575 83.515 162.385 ;
        RECT 84.265 162.140 84.435 162.805 ;
        RECT 84.830 162.465 85.955 162.635 ;
        RECT 83.685 161.950 84.435 162.140 ;
        RECT 84.605 162.125 85.615 162.295 ;
        RECT 82.235 160.765 82.565 161.395 ;
        RECT 82.735 160.595 82.945 161.415 ;
        RECT 83.175 161.405 84.405 161.575 ;
        RECT 83.450 160.800 83.695 161.405 ;
        RECT 83.915 160.595 84.425 161.130 ;
        RECT 84.605 160.765 84.795 162.125 ;
        RECT 84.965 161.445 85.240 161.925 ;
        RECT 84.965 161.275 85.245 161.445 ;
        RECT 85.445 161.325 85.615 162.125 ;
        RECT 85.785 161.335 85.955 162.465 ;
        RECT 86.125 161.835 86.295 162.805 ;
        RECT 86.465 162.005 86.635 163.145 ;
        RECT 86.805 162.005 87.140 162.975 ;
        RECT 86.125 161.505 86.320 161.835 ;
        RECT 86.545 161.505 86.800 161.835 ;
        RECT 86.545 161.335 86.715 161.505 ;
        RECT 86.970 161.335 87.140 162.005 ;
        RECT 87.315 161.980 87.605 163.145 ;
        RECT 87.815 162.005 88.045 163.145 ;
        RECT 88.215 161.995 88.545 162.975 ;
        RECT 88.715 162.005 88.925 163.145 ;
        RECT 90.190 162.515 90.475 162.975 ;
        RECT 90.645 162.685 90.915 163.145 ;
        RECT 90.190 162.295 91.145 162.515 ;
        RECT 87.795 161.585 88.125 161.835 ;
        RECT 84.965 160.765 85.240 161.275 ;
        RECT 85.785 161.165 86.715 161.335 ;
        RECT 85.785 161.130 85.960 161.165 ;
        RECT 85.430 160.765 85.960 161.130 ;
        RECT 86.385 160.595 86.715 160.995 ;
        RECT 86.885 160.765 87.140 161.335 ;
        RECT 87.315 160.595 87.605 161.320 ;
        RECT 87.815 160.595 88.045 161.415 ;
        RECT 88.295 161.395 88.545 161.995 ;
        RECT 90.075 161.565 90.765 162.125 ;
        RECT 88.215 160.765 88.545 161.395 ;
        RECT 88.715 160.595 88.925 161.415 ;
        RECT 90.935 161.395 91.145 162.295 ;
        RECT 90.190 161.225 91.145 161.395 ;
        RECT 91.315 162.125 91.715 162.975 ;
        RECT 91.905 162.515 92.185 162.975 ;
        RECT 92.705 162.685 93.030 163.145 ;
        RECT 91.905 162.295 93.030 162.515 ;
        RECT 91.315 161.565 92.410 162.125 ;
        RECT 92.580 161.835 93.030 162.295 ;
        RECT 93.200 162.005 93.585 162.975 ;
        RECT 90.190 160.765 90.475 161.225 ;
        RECT 90.645 160.595 90.915 161.055 ;
        RECT 91.315 160.765 91.715 161.565 ;
        RECT 92.580 161.505 93.135 161.835 ;
        RECT 92.580 161.395 93.030 161.505 ;
        RECT 91.905 161.225 93.030 161.395 ;
        RECT 93.305 161.335 93.585 162.005 ;
        RECT 91.905 160.765 92.185 161.225 ;
        RECT 92.705 160.595 93.030 161.055 ;
        RECT 93.200 160.765 93.585 161.335 ;
        RECT 93.755 162.005 94.095 162.975 ;
        RECT 94.265 162.005 94.435 163.145 ;
        RECT 94.705 162.345 94.955 163.145 ;
        RECT 95.600 162.175 95.930 162.975 ;
        RECT 96.230 162.345 96.560 163.145 ;
        RECT 96.730 162.175 97.060 162.975 ;
        RECT 94.625 162.005 97.060 162.175 ;
        RECT 98.100 162.175 98.430 162.975 ;
        RECT 98.600 162.345 98.930 163.145 ;
        RECT 99.230 162.175 99.560 162.975 ;
        RECT 100.205 162.345 100.455 163.145 ;
        RECT 98.100 162.005 100.535 162.175 ;
        RECT 100.725 162.005 100.895 163.145 ;
        RECT 101.065 162.005 101.405 162.975 ;
        RECT 93.755 161.395 93.930 162.005 ;
        RECT 94.625 161.755 94.795 162.005 ;
        RECT 94.100 161.585 94.795 161.755 ;
        RECT 94.970 161.585 95.390 161.785 ;
        RECT 95.560 161.585 95.890 161.785 ;
        RECT 96.060 161.585 96.390 161.785 ;
        RECT 93.755 160.765 94.095 161.395 ;
        RECT 94.265 160.595 94.515 161.395 ;
        RECT 94.705 161.245 95.930 161.415 ;
        RECT 94.705 160.765 95.035 161.245 ;
        RECT 95.205 160.595 95.430 161.055 ;
        RECT 95.600 160.765 95.930 161.245 ;
        RECT 96.560 161.375 96.730 162.005 ;
        RECT 96.915 161.585 97.265 161.835 ;
        RECT 97.895 161.585 98.245 161.835 ;
        RECT 98.430 161.375 98.600 162.005 ;
        RECT 98.770 161.585 99.100 161.785 ;
        RECT 99.270 161.585 99.600 161.785 ;
        RECT 99.770 161.585 100.190 161.785 ;
        RECT 100.365 161.755 100.535 162.005 ;
        RECT 100.365 161.585 101.060 161.755 ;
        RECT 96.560 160.765 97.060 161.375 ;
        RECT 98.100 160.765 98.600 161.375 ;
        RECT 99.230 161.245 100.455 161.415 ;
        RECT 101.230 161.395 101.405 162.005 ;
        RECT 101.575 162.385 102.090 162.795 ;
        RECT 102.325 162.385 102.495 163.145 ;
        RECT 102.665 162.805 104.695 162.975 ;
        RECT 101.575 161.575 101.915 162.385 ;
        RECT 102.665 162.140 102.835 162.805 ;
        RECT 103.230 162.465 104.355 162.635 ;
        RECT 102.085 161.950 102.835 162.140 ;
        RECT 103.005 162.125 104.015 162.295 ;
        RECT 101.575 161.405 102.805 161.575 ;
        RECT 99.230 160.765 99.560 161.245 ;
        RECT 99.730 160.595 99.955 161.055 ;
        RECT 100.125 160.765 100.455 161.245 ;
        RECT 100.645 160.595 100.895 161.395 ;
        RECT 101.065 160.765 101.405 161.395 ;
        RECT 101.850 160.800 102.095 161.405 ;
        RECT 102.315 160.595 102.825 161.130 ;
        RECT 103.005 160.765 103.195 162.125 ;
        RECT 103.365 161.105 103.640 161.925 ;
        RECT 103.845 161.325 104.015 162.125 ;
        RECT 104.185 161.335 104.355 162.465 ;
        RECT 104.525 161.835 104.695 162.805 ;
        RECT 104.865 162.005 105.035 163.145 ;
        RECT 105.205 162.005 105.540 162.975 ;
        RECT 104.525 161.505 104.720 161.835 ;
        RECT 104.945 161.505 105.200 161.835 ;
        RECT 104.945 161.335 105.115 161.505 ;
        RECT 105.370 161.335 105.540 162.005 ;
        RECT 105.715 162.385 106.230 162.795 ;
        RECT 106.465 162.385 106.635 163.145 ;
        RECT 106.805 162.805 108.835 162.975 ;
        RECT 105.715 161.575 106.055 162.385 ;
        RECT 106.805 162.140 106.975 162.805 ;
        RECT 107.370 162.465 108.495 162.635 ;
        RECT 106.225 161.950 106.975 162.140 ;
        RECT 107.145 162.125 108.155 162.295 ;
        RECT 105.715 161.405 106.945 161.575 ;
        RECT 104.185 161.165 105.115 161.335 ;
        RECT 104.185 161.130 104.360 161.165 ;
        RECT 103.365 160.935 103.645 161.105 ;
        RECT 103.365 160.765 103.640 160.935 ;
        RECT 103.830 160.765 104.360 161.130 ;
        RECT 104.785 160.595 105.115 160.995 ;
        RECT 105.285 160.765 105.540 161.335 ;
        RECT 105.990 160.800 106.235 161.405 ;
        RECT 106.455 160.595 106.965 161.130 ;
        RECT 107.145 160.765 107.335 162.125 ;
        RECT 107.505 161.445 107.780 161.925 ;
        RECT 107.505 161.275 107.785 161.445 ;
        RECT 107.985 161.325 108.155 162.125 ;
        RECT 108.325 161.335 108.495 162.465 ;
        RECT 108.665 161.835 108.835 162.805 ;
        RECT 109.005 162.005 109.175 163.145 ;
        RECT 109.345 162.005 109.680 162.975 ;
        RECT 109.945 162.215 110.115 162.975 ;
        RECT 110.295 162.385 110.625 163.145 ;
        RECT 109.945 162.045 110.610 162.215 ;
        RECT 110.795 162.070 111.065 162.975 ;
        RECT 108.665 161.505 108.860 161.835 ;
        RECT 109.085 161.505 109.340 161.835 ;
        RECT 109.085 161.335 109.255 161.505 ;
        RECT 109.510 161.335 109.680 162.005 ;
        RECT 110.440 161.900 110.610 162.045 ;
        RECT 109.875 161.495 110.205 161.865 ;
        RECT 110.440 161.570 110.725 161.900 ;
        RECT 107.505 160.765 107.780 161.275 ;
        RECT 108.325 161.165 109.255 161.335 ;
        RECT 108.325 161.130 108.500 161.165 ;
        RECT 107.970 160.765 108.500 161.130 ;
        RECT 108.925 160.595 109.255 160.995 ;
        RECT 109.425 160.765 109.680 161.335 ;
        RECT 110.440 161.315 110.610 161.570 ;
        RECT 109.945 161.145 110.610 161.315 ;
        RECT 110.895 161.270 111.065 162.070 ;
        RECT 112.155 162.055 113.365 163.145 ;
        RECT 112.155 161.515 112.675 162.055 ;
        RECT 112.845 161.345 113.365 161.885 ;
        RECT 109.945 160.765 110.115 161.145 ;
        RECT 110.295 160.595 110.625 160.975 ;
        RECT 110.805 160.765 111.065 161.270 ;
        RECT 112.155 160.595 113.365 161.345 ;
        RECT 26.970 160.425 113.450 160.595 ;
        RECT 27.055 159.675 28.265 160.425 ;
        RECT 28.435 159.750 28.705 160.095 ;
        RECT 28.895 160.025 29.275 160.425 ;
        RECT 29.445 159.855 29.615 160.205 ;
        RECT 29.785 160.025 30.115 160.425 ;
        RECT 30.315 159.855 30.485 160.205 ;
        RECT 30.685 159.925 31.015 160.425 ;
        RECT 27.055 159.135 27.575 159.675 ;
        RECT 27.745 158.965 28.265 159.505 ;
        RECT 27.055 157.875 28.265 158.965 ;
        RECT 28.435 159.015 28.605 159.750 ;
        RECT 28.875 159.685 30.485 159.855 ;
        RECT 28.875 159.515 29.045 159.685 ;
        RECT 28.775 159.185 29.045 159.515 ;
        RECT 29.215 159.185 29.620 159.515 ;
        RECT 28.875 159.015 29.045 159.185 ;
        RECT 29.790 159.065 30.500 159.515 ;
        RECT 30.670 159.185 31.020 159.755 ;
        RECT 31.195 159.750 31.465 160.095 ;
        RECT 31.655 160.025 32.035 160.425 ;
        RECT 32.205 159.855 32.375 160.205 ;
        RECT 32.545 160.025 32.875 160.425 ;
        RECT 33.075 159.855 33.245 160.205 ;
        RECT 33.445 159.925 33.775 160.425 ;
        RECT 28.435 158.045 28.705 159.015 ;
        RECT 28.875 158.845 29.600 159.015 ;
        RECT 29.790 158.895 30.505 159.065 ;
        RECT 31.195 159.015 31.365 159.750 ;
        RECT 31.635 159.685 33.245 159.855 ;
        RECT 31.635 159.515 31.805 159.685 ;
        RECT 31.535 159.185 31.805 159.515 ;
        RECT 31.975 159.185 32.380 159.515 ;
        RECT 31.635 159.015 31.805 159.185 ;
        RECT 32.550 159.065 33.260 159.515 ;
        RECT 33.430 159.185 33.780 159.755 ;
        RECT 33.955 159.685 34.340 160.255 ;
        RECT 34.510 159.965 34.835 160.425 ;
        RECT 35.355 159.795 35.635 160.255 ;
        RECT 29.430 158.725 29.600 158.845 ;
        RECT 30.700 158.725 31.020 159.015 ;
        RECT 28.915 157.875 29.195 158.675 ;
        RECT 29.430 158.555 31.020 158.725 ;
        RECT 29.365 158.095 31.020 158.385 ;
        RECT 31.195 158.045 31.465 159.015 ;
        RECT 31.635 158.845 32.360 159.015 ;
        RECT 32.550 158.895 33.265 159.065 ;
        RECT 33.955 159.015 34.235 159.685 ;
        RECT 34.510 159.625 35.635 159.795 ;
        RECT 34.510 159.515 34.960 159.625 ;
        RECT 34.405 159.185 34.960 159.515 ;
        RECT 35.825 159.455 36.225 160.255 ;
        RECT 36.625 159.965 36.895 160.425 ;
        RECT 37.065 159.795 37.350 160.255 ;
        RECT 32.190 158.725 32.360 158.845 ;
        RECT 33.460 158.725 33.780 159.015 ;
        RECT 31.675 157.875 31.955 158.675 ;
        RECT 32.190 158.555 33.780 158.725 ;
        RECT 32.125 158.095 33.780 158.385 ;
        RECT 33.955 158.045 34.340 159.015 ;
        RECT 34.510 158.725 34.960 159.185 ;
        RECT 35.130 158.895 36.225 159.455 ;
        RECT 34.510 158.505 35.635 158.725 ;
        RECT 34.510 157.875 34.835 158.335 ;
        RECT 35.355 158.045 35.635 158.505 ;
        RECT 35.825 158.045 36.225 158.895 ;
        RECT 36.395 159.625 37.350 159.795 ;
        RECT 37.635 159.625 37.975 160.255 ;
        RECT 38.145 159.625 38.395 160.425 ;
        RECT 38.585 159.775 38.915 160.255 ;
        RECT 39.085 159.965 39.310 160.425 ;
        RECT 39.480 159.775 39.810 160.255 ;
        RECT 36.395 158.725 36.605 159.625 ;
        RECT 37.635 159.575 37.865 159.625 ;
        RECT 38.585 159.605 39.810 159.775 ;
        RECT 40.440 159.645 40.940 160.255 ;
        RECT 36.775 158.895 37.465 159.455 ;
        RECT 37.635 159.015 37.810 159.575 ;
        RECT 37.980 159.265 38.675 159.435 ;
        RECT 38.505 159.015 38.675 159.265 ;
        RECT 38.850 159.235 39.270 159.435 ;
        RECT 39.440 159.235 39.770 159.435 ;
        RECT 39.940 159.235 40.270 159.435 ;
        RECT 40.440 159.015 40.610 159.645 ;
        RECT 41.315 159.625 41.655 160.255 ;
        RECT 41.825 159.625 42.075 160.425 ;
        RECT 42.265 159.775 42.595 160.255 ;
        RECT 42.765 159.965 42.990 160.425 ;
        RECT 43.160 159.775 43.490 160.255 ;
        RECT 40.795 159.185 41.145 159.435 ;
        RECT 41.315 159.015 41.490 159.625 ;
        RECT 42.265 159.605 43.490 159.775 ;
        RECT 44.120 159.645 44.620 160.255 ;
        RECT 41.660 159.265 42.355 159.435 ;
        RECT 42.185 159.015 42.355 159.265 ;
        RECT 42.530 159.235 42.950 159.435 ;
        RECT 43.120 159.235 43.450 159.435 ;
        RECT 43.620 159.235 43.950 159.435 ;
        RECT 44.120 159.015 44.290 159.645 ;
        RECT 44.995 159.625 45.335 160.255 ;
        RECT 45.505 159.625 45.755 160.425 ;
        RECT 45.945 159.775 46.275 160.255 ;
        RECT 46.445 159.965 46.670 160.425 ;
        RECT 46.840 159.775 47.170 160.255 ;
        RECT 44.475 159.185 44.825 159.435 ;
        RECT 44.995 159.015 45.170 159.625 ;
        RECT 45.945 159.605 47.170 159.775 ;
        RECT 47.800 159.645 48.300 160.255 ;
        RECT 48.675 159.700 48.965 160.425 ;
        RECT 49.225 159.875 49.395 160.165 ;
        RECT 49.565 160.045 49.895 160.425 ;
        RECT 49.225 159.705 49.890 159.875 ;
        RECT 45.340 159.265 46.035 159.435 ;
        RECT 45.865 159.015 46.035 159.265 ;
        RECT 46.210 159.235 46.630 159.435 ;
        RECT 46.800 159.235 47.130 159.435 ;
        RECT 47.300 159.235 47.630 159.435 ;
        RECT 47.800 159.015 47.970 159.645 ;
        RECT 48.155 159.185 48.505 159.435 ;
        RECT 36.395 158.505 37.350 158.725 ;
        RECT 36.625 157.875 36.895 158.335 ;
        RECT 37.065 158.045 37.350 158.505 ;
        RECT 37.635 158.045 37.975 159.015 ;
        RECT 38.145 157.875 38.315 159.015 ;
        RECT 38.505 158.845 40.940 159.015 ;
        RECT 38.585 157.875 38.835 158.675 ;
        RECT 39.480 158.045 39.810 158.845 ;
        RECT 40.110 157.875 40.440 158.675 ;
        RECT 40.610 158.045 40.940 158.845 ;
        RECT 41.315 158.045 41.655 159.015 ;
        RECT 41.825 157.875 41.995 159.015 ;
        RECT 42.185 158.845 44.620 159.015 ;
        RECT 42.265 157.875 42.515 158.675 ;
        RECT 43.160 158.045 43.490 158.845 ;
        RECT 43.790 157.875 44.120 158.675 ;
        RECT 44.290 158.045 44.620 158.845 ;
        RECT 44.995 158.045 45.335 159.015 ;
        RECT 45.505 157.875 45.675 159.015 ;
        RECT 45.865 158.845 48.300 159.015 ;
        RECT 45.945 157.875 46.195 158.675 ;
        RECT 46.840 158.045 47.170 158.845 ;
        RECT 47.470 157.875 47.800 158.675 ;
        RECT 47.970 158.045 48.300 158.845 ;
        RECT 48.675 157.875 48.965 159.040 ;
        RECT 49.140 158.885 49.490 159.535 ;
        RECT 49.660 158.715 49.890 159.705 ;
        RECT 49.225 158.545 49.890 158.715 ;
        RECT 49.225 158.045 49.395 158.545 ;
        RECT 49.565 157.875 49.895 158.375 ;
        RECT 50.065 158.045 50.290 160.165 ;
        RECT 50.505 160.045 50.835 160.425 ;
        RECT 51.005 159.875 51.175 160.205 ;
        RECT 51.475 160.045 52.490 160.245 ;
        RECT 50.480 159.685 51.175 159.875 ;
        RECT 50.480 158.715 50.650 159.685 ;
        RECT 50.820 158.885 51.230 159.505 ;
        RECT 51.400 158.935 51.620 159.805 ;
        RECT 51.800 159.495 52.150 159.865 ;
        RECT 52.320 159.315 52.490 160.045 ;
        RECT 52.660 159.985 53.070 160.425 ;
        RECT 53.360 159.785 53.610 160.215 ;
        RECT 53.810 159.965 54.130 160.425 ;
        RECT 54.690 160.035 55.540 160.205 ;
        RECT 52.660 159.445 53.070 159.775 ;
        RECT 53.360 159.445 53.780 159.785 ;
        RECT 52.070 159.275 52.490 159.315 ;
        RECT 52.070 159.105 53.420 159.275 ;
        RECT 50.480 158.545 51.175 158.715 ;
        RECT 51.400 158.555 51.900 158.935 ;
        RECT 50.505 157.875 50.835 158.375 ;
        RECT 51.005 158.045 51.175 158.545 ;
        RECT 52.070 158.260 52.240 159.105 ;
        RECT 53.170 158.945 53.420 159.105 ;
        RECT 52.410 158.675 52.660 158.935 ;
        RECT 53.590 158.675 53.780 159.445 ;
        RECT 52.410 158.425 53.780 158.675 ;
        RECT 53.950 159.615 55.200 159.785 ;
        RECT 53.950 158.855 54.120 159.615 ;
        RECT 54.870 159.495 55.200 159.615 ;
        RECT 54.290 159.035 54.470 159.445 ;
        RECT 55.370 159.275 55.540 160.035 ;
        RECT 55.740 159.945 56.400 160.425 ;
        RECT 56.580 159.830 56.900 160.160 ;
        RECT 55.730 159.505 56.390 159.775 ;
        RECT 55.730 159.445 56.060 159.505 ;
        RECT 56.210 159.275 56.540 159.335 ;
        RECT 54.640 159.105 56.540 159.275 ;
        RECT 53.950 158.545 54.470 158.855 ;
        RECT 54.640 158.595 54.810 159.105 ;
        RECT 56.710 158.935 56.900 159.830 ;
        RECT 54.980 158.765 56.900 158.935 ;
        RECT 56.580 158.745 56.900 158.765 ;
        RECT 57.100 159.515 57.350 160.165 ;
        RECT 57.530 159.965 57.815 160.425 ;
        RECT 57.995 159.715 58.250 160.245 ;
        RECT 57.100 159.185 57.900 159.515 ;
        RECT 54.640 158.425 55.850 158.595 ;
        RECT 51.410 158.090 52.240 158.260 ;
        RECT 52.480 157.875 52.860 158.255 ;
        RECT 53.040 158.135 53.210 158.425 ;
        RECT 54.640 158.345 54.810 158.425 ;
        RECT 53.380 157.875 53.710 158.255 ;
        RECT 54.180 158.095 54.810 158.345 ;
        RECT 54.990 157.875 55.410 158.255 ;
        RECT 55.610 158.135 55.850 158.425 ;
        RECT 56.080 157.875 56.410 158.565 ;
        RECT 56.580 158.135 56.750 158.745 ;
        RECT 57.100 158.595 57.350 159.185 ;
        RECT 58.070 159.065 58.250 159.715 ;
        RECT 59.070 159.615 59.315 160.220 ;
        RECT 59.535 159.890 60.045 160.425 ;
        RECT 58.795 159.445 60.025 159.615 ;
        RECT 58.070 158.895 58.335 159.065 ;
        RECT 58.070 158.855 58.250 158.895 ;
        RECT 57.020 158.085 57.350 158.595 ;
        RECT 57.530 157.875 57.815 158.675 ;
        RECT 57.995 158.185 58.250 158.855 ;
        RECT 58.795 158.635 59.135 159.445 ;
        RECT 59.305 158.880 60.055 159.070 ;
        RECT 58.795 158.225 59.310 158.635 ;
        RECT 59.545 157.875 59.715 158.635 ;
        RECT 59.885 158.215 60.055 158.880 ;
        RECT 60.225 158.895 60.415 160.255 ;
        RECT 60.585 159.405 60.860 160.255 ;
        RECT 61.050 159.890 61.580 160.255 ;
        RECT 62.005 160.025 62.335 160.425 ;
        RECT 61.405 159.855 61.580 159.890 ;
        RECT 60.585 159.235 60.865 159.405 ;
        RECT 60.585 159.095 60.860 159.235 ;
        RECT 61.065 158.895 61.235 159.695 ;
        RECT 60.225 158.725 61.235 158.895 ;
        RECT 61.405 159.685 62.335 159.855 ;
        RECT 62.505 159.685 62.760 160.255 ;
        RECT 63.945 159.875 64.115 160.255 ;
        RECT 64.295 160.045 64.625 160.425 ;
        RECT 63.945 159.705 64.610 159.875 ;
        RECT 64.805 159.750 65.065 160.255 ;
        RECT 61.405 158.555 61.575 159.685 ;
        RECT 62.165 159.515 62.335 159.685 ;
        RECT 60.450 158.385 61.575 158.555 ;
        RECT 61.745 159.185 61.940 159.515 ;
        RECT 62.165 159.185 62.420 159.515 ;
        RECT 61.745 158.215 61.915 159.185 ;
        RECT 62.590 159.015 62.760 159.685 ;
        RECT 63.875 159.155 64.205 159.525 ;
        RECT 64.440 159.450 64.610 159.705 ;
        RECT 59.885 158.045 61.915 158.215 ;
        RECT 62.085 157.875 62.255 159.015 ;
        RECT 62.425 158.045 62.760 159.015 ;
        RECT 64.440 159.120 64.725 159.450 ;
        RECT 64.440 158.975 64.610 159.120 ;
        RECT 63.945 158.805 64.610 158.975 ;
        RECT 64.895 158.950 65.065 159.750 ;
        RECT 65.240 159.585 65.500 160.425 ;
        RECT 65.675 159.680 65.930 160.255 ;
        RECT 66.100 160.045 66.430 160.425 ;
        RECT 66.645 159.875 66.815 160.255 ;
        RECT 67.135 159.945 67.415 160.425 ;
        RECT 66.100 159.705 66.815 159.875 ;
        RECT 67.585 159.775 67.845 160.165 ;
        RECT 68.020 159.945 68.275 160.425 ;
        RECT 68.445 159.775 68.740 160.165 ;
        RECT 68.920 159.945 69.195 160.425 ;
        RECT 69.365 159.925 69.665 160.255 ;
        RECT 63.945 158.045 64.115 158.805 ;
        RECT 64.295 157.875 64.625 158.635 ;
        RECT 64.795 158.045 65.065 158.950 ;
        RECT 65.240 157.875 65.500 159.025 ;
        RECT 65.675 158.950 65.845 159.680 ;
        RECT 66.100 159.515 66.270 159.705 ;
        RECT 67.090 159.605 68.740 159.775 ;
        RECT 66.015 159.185 66.270 159.515 ;
        RECT 66.100 158.975 66.270 159.185 ;
        RECT 66.550 159.155 66.905 159.525 ;
        RECT 67.090 159.095 67.495 159.605 ;
        RECT 67.665 159.265 68.805 159.435 ;
        RECT 65.675 158.045 65.930 158.950 ;
        RECT 66.100 158.805 66.815 158.975 ;
        RECT 67.090 158.925 67.845 159.095 ;
        RECT 66.100 157.875 66.430 158.635 ;
        RECT 66.645 158.045 66.815 158.805 ;
        RECT 67.130 157.875 67.415 158.745 ;
        RECT 67.585 158.675 67.845 158.925 ;
        RECT 68.635 159.015 68.805 159.265 ;
        RECT 68.975 159.185 69.325 159.755 ;
        RECT 69.495 159.015 69.665 159.925 ;
        RECT 69.925 159.875 70.095 160.255 ;
        RECT 70.310 160.045 70.640 160.425 ;
        RECT 69.925 159.705 70.640 159.875 ;
        RECT 69.835 159.155 70.190 159.525 ;
        RECT 70.470 159.515 70.640 159.705 ;
        RECT 70.810 159.680 71.065 160.255 ;
        RECT 70.470 159.185 70.725 159.515 ;
        RECT 68.635 158.845 69.665 159.015 ;
        RECT 70.470 158.975 70.640 159.185 ;
        RECT 67.585 158.505 68.705 158.675 ;
        RECT 67.585 158.045 67.845 158.505 ;
        RECT 68.020 157.875 68.275 158.335 ;
        RECT 68.445 158.045 68.705 158.505 ;
        RECT 68.875 157.875 69.185 158.675 ;
        RECT 69.355 158.045 69.665 158.845 ;
        RECT 69.925 158.805 70.640 158.975 ;
        RECT 70.895 158.950 71.065 159.680 ;
        RECT 71.240 159.585 71.500 160.425 ;
        RECT 71.675 159.925 71.975 160.255 ;
        RECT 72.145 159.945 72.420 160.425 ;
        RECT 69.925 158.045 70.095 158.805 ;
        RECT 70.310 157.875 70.640 158.635 ;
        RECT 70.810 158.045 71.065 158.950 ;
        RECT 71.240 157.875 71.500 159.025 ;
        RECT 71.675 159.015 71.845 159.925 ;
        RECT 72.600 159.775 72.895 160.165 ;
        RECT 73.065 159.945 73.320 160.425 ;
        RECT 73.495 159.775 73.755 160.165 ;
        RECT 73.925 159.945 74.205 160.425 ;
        RECT 72.015 159.185 72.365 159.755 ;
        RECT 72.600 159.605 74.250 159.775 ;
        RECT 74.435 159.700 74.725 160.425 ;
        RECT 74.895 159.750 75.155 160.255 ;
        RECT 75.335 160.045 75.665 160.425 ;
        RECT 75.845 159.875 76.015 160.255 ;
        RECT 72.535 159.265 73.675 159.435 ;
        RECT 72.535 159.015 72.705 159.265 ;
        RECT 73.845 159.095 74.250 159.605 ;
        RECT 71.675 158.845 72.705 159.015 ;
        RECT 73.495 158.925 74.250 159.095 ;
        RECT 71.675 158.045 71.985 158.845 ;
        RECT 73.495 158.675 73.755 158.925 ;
        RECT 72.155 157.875 72.465 158.675 ;
        RECT 72.635 158.505 73.755 158.675 ;
        RECT 72.635 158.045 72.895 158.505 ;
        RECT 73.065 157.875 73.320 158.335 ;
        RECT 73.495 158.045 73.755 158.505 ;
        RECT 73.925 157.875 74.210 158.745 ;
        RECT 74.435 157.875 74.725 159.040 ;
        RECT 74.895 158.950 75.065 159.750 ;
        RECT 75.350 159.705 76.015 159.875 ;
        RECT 76.365 159.875 76.535 160.255 ;
        RECT 76.715 160.045 77.045 160.425 ;
        RECT 76.365 159.705 77.030 159.875 ;
        RECT 77.225 159.750 77.485 160.255 ;
        RECT 75.350 159.450 75.520 159.705 ;
        RECT 75.235 159.120 75.520 159.450 ;
        RECT 75.755 159.155 76.085 159.525 ;
        RECT 76.295 159.155 76.625 159.525 ;
        RECT 76.860 159.450 77.030 159.705 ;
        RECT 75.350 158.975 75.520 159.120 ;
        RECT 76.860 159.120 77.145 159.450 ;
        RECT 76.860 158.975 77.030 159.120 ;
        RECT 74.895 158.045 75.165 158.950 ;
        RECT 75.350 158.805 76.015 158.975 ;
        RECT 75.335 157.875 75.665 158.635 ;
        RECT 75.845 158.045 76.015 158.805 ;
        RECT 76.365 158.805 77.030 158.975 ;
        RECT 77.315 158.950 77.485 159.750 ;
        RECT 78.030 159.745 78.285 160.245 ;
        RECT 78.465 159.965 78.750 160.425 ;
        RECT 77.945 159.715 78.285 159.745 ;
        RECT 77.945 159.575 78.210 159.715 ;
        RECT 76.365 158.045 76.535 158.805 ;
        RECT 76.715 157.875 77.045 158.635 ;
        RECT 77.215 158.045 77.485 158.950 ;
        RECT 78.030 158.855 78.210 159.575 ;
        RECT 78.930 159.515 79.180 160.165 ;
        RECT 78.380 159.185 79.180 159.515 ;
        RECT 78.030 158.185 78.285 158.855 ;
        RECT 78.465 157.875 78.750 158.675 ;
        RECT 78.930 158.595 79.180 159.185 ;
        RECT 79.380 159.830 79.700 160.160 ;
        RECT 79.880 159.945 80.540 160.425 ;
        RECT 80.740 160.035 81.590 160.205 ;
        RECT 79.380 158.935 79.570 159.830 ;
        RECT 79.890 159.505 80.550 159.775 ;
        RECT 80.220 159.445 80.550 159.505 ;
        RECT 79.740 159.275 80.070 159.335 ;
        RECT 80.740 159.275 80.910 160.035 ;
        RECT 82.150 159.965 82.470 160.425 ;
        RECT 82.670 159.785 82.920 160.215 ;
        RECT 83.210 159.985 83.620 160.425 ;
        RECT 83.790 160.045 84.805 160.245 ;
        RECT 81.080 159.615 82.330 159.785 ;
        RECT 81.080 159.495 81.410 159.615 ;
        RECT 79.740 159.105 81.640 159.275 ;
        RECT 79.380 158.765 81.300 158.935 ;
        RECT 79.380 158.745 79.700 158.765 ;
        RECT 78.930 158.085 79.260 158.595 ;
        RECT 79.530 158.135 79.700 158.745 ;
        RECT 81.470 158.595 81.640 159.105 ;
        RECT 81.810 159.035 81.990 159.445 ;
        RECT 82.160 158.855 82.330 159.615 ;
        RECT 79.870 157.875 80.200 158.565 ;
        RECT 80.430 158.425 81.640 158.595 ;
        RECT 81.810 158.545 82.330 158.855 ;
        RECT 82.500 159.445 82.920 159.785 ;
        RECT 83.210 159.445 83.620 159.775 ;
        RECT 82.500 158.675 82.690 159.445 ;
        RECT 83.790 159.315 83.960 160.045 ;
        RECT 85.105 159.875 85.275 160.205 ;
        RECT 85.445 160.045 85.775 160.425 ;
        RECT 84.130 159.495 84.480 159.865 ;
        RECT 83.790 159.275 84.210 159.315 ;
        RECT 82.860 159.105 84.210 159.275 ;
        RECT 82.860 158.945 83.110 159.105 ;
        RECT 83.620 158.675 83.870 158.935 ;
        RECT 82.500 158.425 83.870 158.675 ;
        RECT 80.430 158.135 80.670 158.425 ;
        RECT 81.470 158.345 81.640 158.425 ;
        RECT 80.870 157.875 81.290 158.255 ;
        RECT 81.470 158.095 82.100 158.345 ;
        RECT 82.570 157.875 82.900 158.255 ;
        RECT 83.070 158.135 83.240 158.425 ;
        RECT 84.040 158.260 84.210 159.105 ;
        RECT 84.660 158.935 84.880 159.805 ;
        RECT 85.105 159.685 85.800 159.875 ;
        RECT 84.380 158.555 84.880 158.935 ;
        RECT 85.050 158.885 85.460 159.505 ;
        RECT 85.630 158.715 85.800 159.685 ;
        RECT 85.105 158.545 85.800 158.715 ;
        RECT 83.420 157.875 83.800 158.255 ;
        RECT 84.040 158.090 84.870 158.260 ;
        RECT 85.105 158.045 85.275 158.545 ;
        RECT 85.445 157.875 85.775 158.375 ;
        RECT 85.990 158.045 86.215 160.165 ;
        RECT 86.385 160.045 86.715 160.425 ;
        RECT 86.885 159.875 87.055 160.165 ;
        RECT 86.390 159.705 87.055 159.875 ;
        RECT 87.320 159.875 87.575 160.165 ;
        RECT 87.745 160.045 88.075 160.425 ;
        RECT 87.320 159.705 88.070 159.875 ;
        RECT 86.390 158.715 86.620 159.705 ;
        RECT 86.790 158.885 87.140 159.535 ;
        RECT 87.320 158.885 87.670 159.535 ;
        RECT 87.840 158.715 88.070 159.705 ;
        RECT 86.390 158.545 87.055 158.715 ;
        RECT 86.385 157.875 86.715 158.375 ;
        RECT 86.885 158.045 87.055 158.545 ;
        RECT 87.320 158.545 88.070 158.715 ;
        RECT 87.320 158.045 87.575 158.545 ;
        RECT 87.745 157.875 88.075 158.375 ;
        RECT 88.245 158.045 88.415 160.165 ;
        RECT 88.775 160.065 89.105 160.425 ;
        RECT 89.275 160.035 89.770 160.205 ;
        RECT 89.975 160.035 90.830 160.205 ;
        RECT 88.645 158.845 89.105 159.895 ;
        RECT 88.585 158.060 88.910 158.845 ;
        RECT 89.275 158.675 89.445 160.035 ;
        RECT 89.615 159.125 89.965 159.745 ;
        RECT 90.135 159.525 90.490 159.745 ;
        RECT 90.135 158.935 90.305 159.525 ;
        RECT 90.660 159.325 90.830 160.035 ;
        RECT 91.705 159.965 92.035 160.425 ;
        RECT 92.245 160.065 92.595 160.235 ;
        RECT 91.035 159.495 91.825 159.745 ;
        RECT 92.245 159.675 92.505 160.065 ;
        RECT 92.815 159.975 93.765 160.255 ;
        RECT 93.935 159.985 94.125 160.425 ;
        RECT 94.295 160.045 95.365 160.215 ;
        RECT 91.995 159.325 92.165 159.505 ;
        RECT 89.275 158.505 89.670 158.675 ;
        RECT 89.840 158.545 90.305 158.935 ;
        RECT 90.475 159.155 92.165 159.325 ;
        RECT 89.500 158.375 89.670 158.505 ;
        RECT 90.475 158.375 90.645 159.155 ;
        RECT 92.335 158.985 92.505 159.675 ;
        RECT 91.005 158.815 92.505 158.985 ;
        RECT 92.695 159.015 92.905 159.805 ;
        RECT 93.075 159.185 93.425 159.805 ;
        RECT 93.595 159.195 93.765 159.975 ;
        RECT 94.295 159.815 94.465 160.045 ;
        RECT 93.935 159.645 94.465 159.815 ;
        RECT 93.935 159.365 94.155 159.645 ;
        RECT 94.635 159.475 94.875 159.875 ;
        RECT 93.595 159.025 94.000 159.195 ;
        RECT 94.335 159.105 94.875 159.475 ;
        RECT 95.045 159.690 95.365 160.045 ;
        RECT 95.610 159.965 95.915 160.425 ;
        RECT 96.085 159.715 96.340 160.245 ;
        RECT 95.045 159.515 95.370 159.690 ;
        RECT 95.045 159.215 95.960 159.515 ;
        RECT 95.220 159.185 95.960 159.215 ;
        RECT 92.695 158.855 93.370 159.015 ;
        RECT 93.830 158.935 94.000 159.025 ;
        RECT 92.695 158.845 93.660 158.855 ;
        RECT 92.335 158.675 92.505 158.815 ;
        RECT 89.080 157.875 89.330 158.335 ;
        RECT 89.500 158.045 89.750 158.375 ;
        RECT 89.965 158.045 90.645 158.375 ;
        RECT 90.815 158.475 91.890 158.645 ;
        RECT 92.335 158.505 92.895 158.675 ;
        RECT 93.200 158.555 93.660 158.845 ;
        RECT 93.830 158.765 95.050 158.935 ;
        RECT 90.815 158.135 90.985 158.475 ;
        RECT 91.220 157.875 91.550 158.305 ;
        RECT 91.720 158.135 91.890 158.475 ;
        RECT 92.185 157.875 92.555 158.335 ;
        RECT 92.725 158.045 92.895 158.505 ;
        RECT 93.830 158.385 94.000 158.765 ;
        RECT 95.220 158.595 95.390 159.185 ;
        RECT 96.130 159.065 96.340 159.715 ;
        RECT 93.130 158.045 94.000 158.385 ;
        RECT 94.590 158.425 95.390 158.595 ;
        RECT 94.170 157.875 94.420 158.335 ;
        RECT 94.590 158.135 94.760 158.425 ;
        RECT 94.940 157.875 95.270 158.255 ;
        RECT 95.610 157.875 95.915 159.015 ;
        RECT 96.085 158.185 96.340 159.065 ;
        RECT 96.515 159.625 96.855 160.255 ;
        RECT 97.025 159.625 97.275 160.425 ;
        RECT 97.465 159.775 97.795 160.255 ;
        RECT 97.965 159.965 98.190 160.425 ;
        RECT 98.360 159.775 98.690 160.255 ;
        RECT 96.515 159.015 96.690 159.625 ;
        RECT 97.465 159.605 98.690 159.775 ;
        RECT 99.320 159.645 99.820 160.255 ;
        RECT 100.195 159.700 100.485 160.425 ;
        RECT 96.860 159.265 97.555 159.435 ;
        RECT 97.385 159.015 97.555 159.265 ;
        RECT 97.730 159.235 98.150 159.435 ;
        RECT 98.320 159.235 98.650 159.435 ;
        RECT 98.820 159.235 99.150 159.435 ;
        RECT 99.320 159.015 99.490 159.645 ;
        RECT 101.155 159.605 101.385 160.425 ;
        RECT 101.555 159.625 101.885 160.255 ;
        RECT 99.675 159.185 100.025 159.435 ;
        RECT 101.135 159.185 101.465 159.435 ;
        RECT 96.515 158.045 96.855 159.015 ;
        RECT 97.025 157.875 97.195 159.015 ;
        RECT 97.385 158.845 99.820 159.015 ;
        RECT 97.465 157.875 97.715 158.675 ;
        RECT 98.360 158.045 98.690 158.845 ;
        RECT 98.990 157.875 99.320 158.675 ;
        RECT 99.490 158.045 99.820 158.845 ;
        RECT 100.195 157.875 100.485 159.040 ;
        RECT 101.635 159.025 101.885 159.625 ;
        RECT 102.055 159.605 102.265 160.425 ;
        RECT 103.230 159.615 103.475 160.220 ;
        RECT 103.695 159.890 104.205 160.425 ;
        RECT 101.155 157.875 101.385 159.015 ;
        RECT 101.555 158.045 101.885 159.025 ;
        RECT 102.955 159.445 104.185 159.615 ;
        RECT 102.055 157.875 102.265 159.015 ;
        RECT 102.955 158.635 103.295 159.445 ;
        RECT 103.465 158.880 104.215 159.070 ;
        RECT 102.955 158.225 103.470 158.635 ;
        RECT 103.705 157.875 103.875 158.635 ;
        RECT 104.045 158.215 104.215 158.880 ;
        RECT 104.385 158.895 104.575 160.255 ;
        RECT 104.745 159.405 105.020 160.255 ;
        RECT 105.210 159.890 105.740 160.255 ;
        RECT 106.165 160.025 106.495 160.425 ;
        RECT 105.565 159.855 105.740 159.890 ;
        RECT 104.745 159.235 105.025 159.405 ;
        RECT 104.745 159.095 105.020 159.235 ;
        RECT 105.225 158.895 105.395 159.695 ;
        RECT 104.385 158.725 105.395 158.895 ;
        RECT 105.565 159.685 106.495 159.855 ;
        RECT 106.665 159.685 106.920 160.255 ;
        RECT 105.565 158.555 105.735 159.685 ;
        RECT 106.325 159.515 106.495 159.685 ;
        RECT 104.610 158.385 105.735 158.555 ;
        RECT 105.905 159.185 106.100 159.515 ;
        RECT 106.325 159.185 106.580 159.515 ;
        RECT 105.905 158.215 106.075 159.185 ;
        RECT 106.750 159.015 106.920 159.685 ;
        RECT 107.210 159.795 107.495 160.255 ;
        RECT 107.665 159.965 107.935 160.425 ;
        RECT 107.210 159.625 108.165 159.795 ;
        RECT 104.045 158.045 106.075 158.215 ;
        RECT 106.245 157.875 106.415 159.015 ;
        RECT 106.585 158.045 106.920 159.015 ;
        RECT 107.095 158.895 107.785 159.455 ;
        RECT 107.955 158.725 108.165 159.625 ;
        RECT 107.210 158.505 108.165 158.725 ;
        RECT 108.335 159.455 108.735 160.255 ;
        RECT 108.925 159.795 109.205 160.255 ;
        RECT 109.725 159.965 110.050 160.425 ;
        RECT 108.925 159.625 110.050 159.795 ;
        RECT 110.220 159.685 110.605 160.255 ;
        RECT 109.600 159.515 110.050 159.625 ;
        RECT 108.335 158.895 109.430 159.455 ;
        RECT 109.600 159.185 110.155 159.515 ;
        RECT 107.210 158.045 107.495 158.505 ;
        RECT 107.665 157.875 107.935 158.335 ;
        RECT 108.335 158.045 108.735 158.895 ;
        RECT 109.600 158.725 110.050 159.185 ;
        RECT 110.325 159.015 110.605 159.685 ;
        RECT 110.835 159.605 111.045 160.425 ;
        RECT 111.215 159.625 111.545 160.255 ;
        RECT 111.215 159.025 111.465 159.625 ;
        RECT 111.715 159.605 111.945 160.425 ;
        RECT 112.155 159.675 113.365 160.425 ;
        RECT 111.635 159.185 111.965 159.435 ;
        RECT 108.925 158.505 110.050 158.725 ;
        RECT 108.925 158.045 109.205 158.505 ;
        RECT 109.725 157.875 110.050 158.335 ;
        RECT 110.220 158.045 110.605 159.015 ;
        RECT 110.835 157.875 111.045 159.015 ;
        RECT 111.215 158.045 111.545 159.025 ;
        RECT 111.715 157.875 111.945 159.015 ;
        RECT 112.155 158.965 112.675 159.505 ;
        RECT 112.845 159.135 113.365 159.675 ;
        RECT 112.155 157.875 113.365 158.965 ;
        RECT 26.970 157.705 113.450 157.875 ;
        RECT 27.055 156.615 28.265 157.705 ;
        RECT 28.635 157.035 28.915 157.705 ;
        RECT 29.085 156.815 29.385 157.365 ;
        RECT 29.585 156.985 29.915 157.705 ;
        RECT 30.105 156.985 30.565 157.535 ;
        RECT 27.055 155.905 27.575 156.445 ;
        RECT 27.745 156.075 28.265 156.615 ;
        RECT 28.450 156.395 28.715 156.755 ;
        RECT 29.085 156.645 30.025 156.815 ;
        RECT 29.855 156.395 30.025 156.645 ;
        RECT 28.450 156.145 29.125 156.395 ;
        RECT 29.345 156.145 29.685 156.395 ;
        RECT 29.855 156.065 30.145 156.395 ;
        RECT 29.855 155.975 30.025 156.065 ;
        RECT 27.055 155.155 28.265 155.905 ;
        RECT 28.635 155.785 30.025 155.975 ;
        RECT 28.635 155.425 28.965 155.785 ;
        RECT 30.315 155.615 30.565 156.985 ;
        RECT 29.585 155.155 29.835 155.615 ;
        RECT 30.005 155.325 30.565 155.615 ;
        RECT 30.740 156.565 31.075 157.535 ;
        RECT 31.245 156.565 31.415 157.705 ;
        RECT 31.585 157.365 33.615 157.535 ;
        RECT 30.740 155.895 30.910 156.565 ;
        RECT 31.585 156.395 31.755 157.365 ;
        RECT 31.080 156.065 31.335 156.395 ;
        RECT 31.560 156.065 31.755 156.395 ;
        RECT 31.925 157.025 33.050 157.195 ;
        RECT 31.165 155.895 31.335 156.065 ;
        RECT 31.925 155.895 32.095 157.025 ;
        RECT 30.740 155.325 30.995 155.895 ;
        RECT 31.165 155.725 32.095 155.895 ;
        RECT 32.265 156.685 33.275 156.855 ;
        RECT 32.265 155.885 32.435 156.685 ;
        RECT 32.640 156.345 32.915 156.485 ;
        RECT 32.635 156.175 32.915 156.345 ;
        RECT 31.920 155.690 32.095 155.725 ;
        RECT 31.165 155.155 31.495 155.555 ;
        RECT 31.920 155.325 32.450 155.690 ;
        RECT 32.640 155.325 32.915 156.175 ;
        RECT 33.085 155.325 33.275 156.685 ;
        RECT 33.445 156.700 33.615 157.365 ;
        RECT 33.785 156.945 33.955 157.705 ;
        RECT 34.190 156.945 34.705 157.355 ;
        RECT 33.445 156.510 34.195 156.700 ;
        RECT 34.365 156.135 34.705 156.945 ;
        RECT 35.795 156.540 36.085 157.705 ;
        RECT 36.255 156.565 36.525 157.535 ;
        RECT 36.735 156.905 37.015 157.705 ;
        RECT 37.185 157.195 38.840 157.485 ;
        RECT 37.250 156.855 38.840 157.025 ;
        RECT 37.250 156.735 37.420 156.855 ;
        RECT 36.695 156.565 37.420 156.735 ;
        RECT 33.475 155.965 34.705 156.135 ;
        RECT 33.455 155.155 33.965 155.690 ;
        RECT 34.185 155.360 34.430 155.965 ;
        RECT 35.795 155.155 36.085 155.880 ;
        RECT 36.255 155.830 36.425 156.565 ;
        RECT 36.695 156.395 36.865 156.565 ;
        RECT 37.610 156.515 38.325 156.685 ;
        RECT 38.520 156.565 38.840 156.855 ;
        RECT 39.015 156.565 39.285 157.535 ;
        RECT 39.495 156.905 39.775 157.705 ;
        RECT 39.945 157.195 41.600 157.485 ;
        RECT 40.010 156.855 41.600 157.025 ;
        RECT 40.010 156.735 40.180 156.855 ;
        RECT 39.455 156.565 40.180 156.735 ;
        RECT 36.595 156.065 36.865 156.395 ;
        RECT 37.035 156.065 37.440 156.395 ;
        RECT 37.610 156.065 38.320 156.515 ;
        RECT 36.695 155.895 36.865 156.065 ;
        RECT 36.255 155.485 36.525 155.830 ;
        RECT 36.695 155.725 38.305 155.895 ;
        RECT 38.490 155.825 38.840 156.395 ;
        RECT 39.015 155.830 39.185 156.565 ;
        RECT 39.455 156.395 39.625 156.565 ;
        RECT 40.370 156.515 41.085 156.685 ;
        RECT 41.280 156.565 41.600 156.855 ;
        RECT 41.775 156.565 42.045 157.535 ;
        RECT 42.255 156.905 42.535 157.705 ;
        RECT 42.705 157.195 44.360 157.485 ;
        RECT 42.770 156.855 44.360 157.025 ;
        RECT 42.770 156.735 42.940 156.855 ;
        RECT 42.215 156.565 42.940 156.735 ;
        RECT 39.355 156.065 39.625 156.395 ;
        RECT 39.795 156.065 40.200 156.395 ;
        RECT 40.370 156.065 41.080 156.515 ;
        RECT 39.455 155.895 39.625 156.065 ;
        RECT 36.715 155.155 37.095 155.555 ;
        RECT 37.265 155.375 37.435 155.725 ;
        RECT 37.605 155.155 37.935 155.555 ;
        RECT 38.135 155.375 38.305 155.725 ;
        RECT 38.505 155.155 38.835 155.655 ;
        RECT 39.015 155.485 39.285 155.830 ;
        RECT 39.455 155.725 41.065 155.895 ;
        RECT 41.250 155.825 41.600 156.395 ;
        RECT 41.775 155.830 41.945 156.565 ;
        RECT 42.215 156.395 42.385 156.565 ;
        RECT 43.130 156.515 43.845 156.685 ;
        RECT 44.040 156.565 44.360 156.855 ;
        RECT 44.535 156.565 44.875 157.535 ;
        RECT 45.045 156.565 45.215 157.705 ;
        RECT 45.485 156.905 45.735 157.705 ;
        RECT 46.380 156.735 46.710 157.535 ;
        RECT 47.010 156.905 47.340 157.705 ;
        RECT 47.510 156.735 47.840 157.535 ;
        RECT 45.405 156.565 47.840 156.735 ;
        RECT 48.215 156.565 48.555 157.535 ;
        RECT 48.725 156.565 48.895 157.705 ;
        RECT 49.165 156.905 49.415 157.705 ;
        RECT 50.060 156.735 50.390 157.535 ;
        RECT 50.690 156.905 51.020 157.705 ;
        RECT 51.190 156.735 51.520 157.535 ;
        RECT 49.085 156.565 51.520 156.735 ;
        RECT 51.895 156.630 52.165 157.535 ;
        RECT 52.335 156.945 52.665 157.705 ;
        RECT 52.845 156.775 53.015 157.535 ;
        RECT 42.115 156.065 42.385 156.395 ;
        RECT 42.555 156.065 42.960 156.395 ;
        RECT 43.130 156.065 43.840 156.515 ;
        RECT 42.215 155.895 42.385 156.065 ;
        RECT 39.475 155.155 39.855 155.555 ;
        RECT 40.025 155.375 40.195 155.725 ;
        RECT 40.365 155.155 40.695 155.555 ;
        RECT 40.895 155.375 41.065 155.725 ;
        RECT 41.265 155.155 41.595 155.655 ;
        RECT 41.775 155.485 42.045 155.830 ;
        RECT 42.215 155.725 43.825 155.895 ;
        RECT 44.010 155.825 44.360 156.395 ;
        RECT 44.535 156.005 44.710 156.565 ;
        RECT 45.405 156.315 45.575 156.565 ;
        RECT 44.880 156.145 45.575 156.315 ;
        RECT 45.750 156.145 46.170 156.345 ;
        RECT 46.340 156.145 46.670 156.345 ;
        RECT 46.840 156.145 47.170 156.345 ;
        RECT 44.535 155.955 44.765 156.005 ;
        RECT 42.235 155.155 42.615 155.555 ;
        RECT 42.785 155.375 42.955 155.725 ;
        RECT 43.125 155.155 43.455 155.555 ;
        RECT 43.655 155.375 43.825 155.725 ;
        RECT 44.025 155.155 44.355 155.655 ;
        RECT 44.535 155.325 44.875 155.955 ;
        RECT 45.045 155.155 45.295 155.955 ;
        RECT 45.485 155.805 46.710 155.975 ;
        RECT 45.485 155.325 45.815 155.805 ;
        RECT 45.985 155.155 46.210 155.615 ;
        RECT 46.380 155.325 46.710 155.805 ;
        RECT 47.340 155.935 47.510 156.565 ;
        RECT 47.695 156.145 48.045 156.395 ;
        RECT 48.215 155.955 48.390 156.565 ;
        RECT 49.085 156.315 49.255 156.565 ;
        RECT 48.560 156.145 49.255 156.315 ;
        RECT 49.430 156.145 49.850 156.345 ;
        RECT 50.020 156.145 50.350 156.345 ;
        RECT 50.520 156.145 50.850 156.345 ;
        RECT 47.340 155.325 47.840 155.935 ;
        RECT 48.215 155.325 48.555 155.955 ;
        RECT 48.725 155.155 48.975 155.955 ;
        RECT 49.165 155.805 50.390 155.975 ;
        RECT 49.165 155.325 49.495 155.805 ;
        RECT 49.665 155.155 49.890 155.615 ;
        RECT 50.060 155.325 50.390 155.805 ;
        RECT 51.020 155.935 51.190 156.565 ;
        RECT 51.375 156.145 51.725 156.395 ;
        RECT 51.020 155.325 51.520 155.935 ;
        RECT 51.895 155.830 52.065 156.630 ;
        RECT 52.350 156.605 53.015 156.775 ;
        RECT 52.350 156.460 52.520 156.605 ;
        RECT 52.235 156.130 52.520 156.460 ;
        RECT 53.280 156.565 53.615 157.535 ;
        RECT 53.785 156.565 53.955 157.705 ;
        RECT 54.125 157.365 56.155 157.535 ;
        RECT 52.350 155.875 52.520 156.130 ;
        RECT 52.755 156.055 53.085 156.425 ;
        RECT 53.280 155.895 53.450 156.565 ;
        RECT 54.125 156.395 54.295 157.365 ;
        RECT 53.620 156.065 53.875 156.395 ;
        RECT 54.100 156.065 54.295 156.395 ;
        RECT 54.465 157.025 55.590 157.195 ;
        RECT 53.705 155.895 53.875 156.065 ;
        RECT 54.465 155.895 54.635 157.025 ;
        RECT 51.895 155.325 52.155 155.830 ;
        RECT 52.350 155.705 53.015 155.875 ;
        RECT 52.335 155.155 52.665 155.535 ;
        RECT 52.845 155.325 53.015 155.705 ;
        RECT 53.280 155.325 53.535 155.895 ;
        RECT 53.705 155.725 54.635 155.895 ;
        RECT 54.805 156.685 55.815 156.855 ;
        RECT 54.805 155.885 54.975 156.685 ;
        RECT 55.180 156.345 55.455 156.485 ;
        RECT 55.175 156.175 55.455 156.345 ;
        RECT 54.460 155.690 54.635 155.725 ;
        RECT 53.705 155.155 54.035 155.555 ;
        RECT 54.460 155.325 54.990 155.690 ;
        RECT 55.180 155.325 55.455 156.175 ;
        RECT 55.625 155.325 55.815 156.685 ;
        RECT 55.985 156.700 56.155 157.365 ;
        RECT 56.325 156.945 56.495 157.705 ;
        RECT 56.730 156.945 57.245 157.355 ;
        RECT 55.985 156.510 56.735 156.700 ;
        RECT 56.905 156.135 57.245 156.945 ;
        RECT 58.340 157.315 58.675 157.535 ;
        RECT 59.680 157.325 60.035 157.705 ;
        RECT 58.340 156.695 58.595 157.315 ;
        RECT 58.845 157.155 59.075 157.195 ;
        RECT 60.205 157.155 60.455 157.535 ;
        RECT 58.845 156.955 60.455 157.155 ;
        RECT 58.845 156.865 59.030 156.955 ;
        RECT 59.620 156.945 60.455 156.955 ;
        RECT 60.705 156.925 60.955 157.705 ;
        RECT 61.125 156.855 61.385 157.535 ;
        RECT 59.185 156.755 59.515 156.785 ;
        RECT 59.185 156.695 60.985 156.755 ;
        RECT 58.340 156.585 61.045 156.695 ;
        RECT 58.340 156.525 59.515 156.585 ;
        RECT 60.845 156.550 61.045 156.585 ;
        RECT 58.335 156.145 58.825 156.345 ;
        RECT 59.015 156.145 59.490 156.355 ;
        RECT 56.015 155.965 57.245 156.135 ;
        RECT 55.995 155.155 56.505 155.690 ;
        RECT 56.725 155.360 56.970 155.965 ;
        RECT 58.340 155.155 58.795 155.920 ;
        RECT 59.270 155.745 59.490 156.145 ;
        RECT 59.735 156.145 60.065 156.355 ;
        RECT 59.735 155.745 59.945 156.145 ;
        RECT 60.235 156.110 60.645 156.415 ;
        RECT 60.875 155.975 61.045 156.550 ;
        RECT 60.775 155.855 61.045 155.975 ;
        RECT 60.200 155.810 61.045 155.855 ;
        RECT 60.200 155.685 60.955 155.810 ;
        RECT 60.200 155.535 60.370 155.685 ;
        RECT 61.215 155.665 61.385 156.855 ;
        RECT 61.555 156.540 61.845 157.705 ;
        RECT 62.475 156.945 62.990 157.355 ;
        RECT 63.225 156.945 63.395 157.705 ;
        RECT 63.565 157.365 65.595 157.535 ;
        RECT 62.475 156.135 62.815 156.945 ;
        RECT 63.565 156.700 63.735 157.365 ;
        RECT 64.130 157.025 65.255 157.195 ;
        RECT 62.985 156.510 63.735 156.700 ;
        RECT 63.905 156.685 64.915 156.855 ;
        RECT 62.475 155.965 63.705 156.135 ;
        RECT 61.155 155.655 61.385 155.665 ;
        RECT 59.070 155.325 60.370 155.535 ;
        RECT 60.625 155.155 60.955 155.515 ;
        RECT 61.125 155.325 61.385 155.655 ;
        RECT 61.555 155.155 61.845 155.880 ;
        RECT 62.750 155.360 62.995 155.965 ;
        RECT 63.215 155.155 63.725 155.690 ;
        RECT 63.905 155.325 64.095 156.685 ;
        RECT 64.265 156.005 64.540 156.485 ;
        RECT 64.265 155.835 64.545 156.005 ;
        RECT 64.745 155.885 64.915 156.685 ;
        RECT 65.085 155.895 65.255 157.025 ;
        RECT 65.425 156.395 65.595 157.365 ;
        RECT 65.765 156.565 65.935 157.705 ;
        RECT 66.105 156.565 66.440 157.535 ;
        RECT 66.675 156.565 66.885 157.705 ;
        RECT 65.425 156.065 65.620 156.395 ;
        RECT 65.845 156.065 66.100 156.395 ;
        RECT 65.845 155.895 66.015 156.065 ;
        RECT 66.270 155.895 66.440 156.565 ;
        RECT 67.055 156.555 67.385 157.535 ;
        RECT 67.555 156.565 67.785 157.705 ;
        RECT 69.005 156.775 69.175 157.535 ;
        RECT 69.390 156.945 69.720 157.705 ;
        RECT 69.005 156.605 69.720 156.775 ;
        RECT 69.890 156.630 70.145 157.535 ;
        RECT 64.265 155.325 64.540 155.835 ;
        RECT 65.085 155.725 66.015 155.895 ;
        RECT 65.085 155.690 65.260 155.725 ;
        RECT 64.730 155.325 65.260 155.690 ;
        RECT 65.685 155.155 66.015 155.555 ;
        RECT 66.185 155.325 66.440 155.895 ;
        RECT 66.675 155.155 66.885 155.975 ;
        RECT 67.055 155.955 67.305 156.555 ;
        RECT 67.475 156.145 67.805 156.395 ;
        RECT 68.915 156.055 69.270 156.425 ;
        RECT 69.550 156.395 69.720 156.605 ;
        RECT 69.550 156.065 69.805 156.395 ;
        RECT 67.055 155.325 67.385 155.955 ;
        RECT 67.555 155.155 67.785 155.975 ;
        RECT 69.550 155.875 69.720 156.065 ;
        RECT 69.975 155.900 70.145 156.630 ;
        RECT 70.320 156.555 70.580 157.705 ;
        RECT 70.845 156.775 71.015 157.535 ;
        RECT 71.230 156.945 71.560 157.705 ;
        RECT 70.845 156.605 71.560 156.775 ;
        RECT 71.730 156.630 71.985 157.535 ;
        RECT 70.755 156.055 71.110 156.425 ;
        RECT 71.390 156.395 71.560 156.605 ;
        RECT 71.390 156.065 71.645 156.395 ;
        RECT 69.005 155.705 69.720 155.875 ;
        RECT 69.005 155.325 69.175 155.705 ;
        RECT 69.390 155.155 69.720 155.535 ;
        RECT 69.890 155.325 70.145 155.900 ;
        RECT 70.320 155.155 70.580 155.995 ;
        RECT 71.390 155.875 71.560 156.065 ;
        RECT 71.815 155.900 71.985 156.630 ;
        RECT 72.160 156.555 72.420 157.705 ;
        RECT 73.055 156.565 73.325 157.535 ;
        RECT 73.535 156.905 73.815 157.705 ;
        RECT 73.985 157.195 75.640 157.485 ;
        RECT 74.050 156.855 75.640 157.025 ;
        RECT 74.050 156.735 74.220 156.855 ;
        RECT 73.495 156.565 74.220 156.735 ;
        RECT 70.845 155.705 71.560 155.875 ;
        RECT 70.845 155.325 71.015 155.705 ;
        RECT 71.230 155.155 71.560 155.535 ;
        RECT 71.730 155.325 71.985 155.900 ;
        RECT 72.160 155.155 72.420 155.995 ;
        RECT 73.055 155.830 73.225 156.565 ;
        RECT 73.495 156.395 73.665 156.565 ;
        RECT 73.395 156.065 73.665 156.395 ;
        RECT 73.835 156.065 74.240 156.395 ;
        RECT 74.410 156.065 75.120 156.685 ;
        RECT 75.320 156.565 75.640 156.855 ;
        RECT 75.815 156.565 76.155 157.535 ;
        RECT 76.325 156.565 76.495 157.705 ;
        RECT 76.765 156.905 77.015 157.705 ;
        RECT 77.660 156.735 77.990 157.535 ;
        RECT 78.290 156.905 78.620 157.705 ;
        RECT 78.790 156.735 79.120 157.535 ;
        RECT 76.685 156.565 79.120 156.735 ;
        RECT 79.495 156.945 80.010 157.355 ;
        RECT 80.245 156.945 80.415 157.705 ;
        RECT 80.585 157.365 82.615 157.535 ;
        RECT 73.495 155.895 73.665 156.065 ;
        RECT 73.055 155.485 73.325 155.830 ;
        RECT 73.495 155.725 75.105 155.895 ;
        RECT 75.290 155.825 75.640 156.395 ;
        RECT 75.815 156.005 75.990 156.565 ;
        RECT 76.685 156.315 76.855 156.565 ;
        RECT 76.160 156.145 76.855 156.315 ;
        RECT 77.030 156.145 77.450 156.345 ;
        RECT 77.620 156.145 77.950 156.345 ;
        RECT 78.120 156.145 78.450 156.345 ;
        RECT 75.815 155.955 76.045 156.005 ;
        RECT 73.515 155.155 73.895 155.555 ;
        RECT 74.065 155.375 74.235 155.725 ;
        RECT 74.405 155.155 74.735 155.555 ;
        RECT 74.935 155.375 75.105 155.725 ;
        RECT 75.305 155.155 75.635 155.655 ;
        RECT 75.815 155.325 76.155 155.955 ;
        RECT 76.325 155.155 76.575 155.955 ;
        RECT 76.765 155.805 77.990 155.975 ;
        RECT 76.765 155.325 77.095 155.805 ;
        RECT 77.265 155.155 77.490 155.615 ;
        RECT 77.660 155.325 77.990 155.805 ;
        RECT 78.620 155.935 78.790 156.565 ;
        RECT 78.975 156.145 79.325 156.395 ;
        RECT 79.495 156.135 79.835 156.945 ;
        RECT 80.585 156.700 80.755 157.365 ;
        RECT 81.150 157.025 82.275 157.195 ;
        RECT 80.005 156.510 80.755 156.700 ;
        RECT 80.925 156.685 81.935 156.855 ;
        RECT 79.495 155.965 80.725 156.135 ;
        RECT 78.620 155.325 79.120 155.935 ;
        RECT 79.770 155.360 80.015 155.965 ;
        RECT 80.235 155.155 80.745 155.690 ;
        RECT 80.925 155.325 81.115 156.685 ;
        RECT 81.285 155.665 81.560 156.485 ;
        RECT 81.765 155.885 81.935 156.685 ;
        RECT 82.105 155.895 82.275 157.025 ;
        RECT 82.445 156.395 82.615 157.365 ;
        RECT 82.785 156.565 82.955 157.705 ;
        RECT 83.125 156.565 83.460 157.535 ;
        RECT 82.445 156.065 82.640 156.395 ;
        RECT 82.865 156.065 83.120 156.395 ;
        RECT 82.865 155.895 83.035 156.065 ;
        RECT 83.290 155.895 83.460 156.565 ;
        RECT 82.105 155.725 83.035 155.895 ;
        RECT 82.105 155.690 82.280 155.725 ;
        RECT 81.285 155.495 81.565 155.665 ;
        RECT 81.285 155.325 81.560 155.495 ;
        RECT 81.750 155.325 82.280 155.690 ;
        RECT 82.705 155.155 83.035 155.555 ;
        RECT 83.205 155.325 83.460 155.895 ;
        RECT 83.635 156.565 84.020 157.535 ;
        RECT 84.190 157.245 84.515 157.705 ;
        RECT 85.035 157.075 85.315 157.535 ;
        RECT 84.190 156.855 85.315 157.075 ;
        RECT 83.635 155.895 83.915 156.565 ;
        RECT 84.190 156.395 84.640 156.855 ;
        RECT 85.505 156.685 85.905 157.535 ;
        RECT 86.305 157.245 86.575 157.705 ;
        RECT 86.745 157.075 87.030 157.535 ;
        RECT 84.085 156.065 84.640 156.395 ;
        RECT 84.810 156.125 85.905 156.685 ;
        RECT 84.190 155.955 84.640 156.065 ;
        RECT 83.635 155.325 84.020 155.895 ;
        RECT 84.190 155.785 85.315 155.955 ;
        RECT 84.190 155.155 84.515 155.615 ;
        RECT 85.035 155.325 85.315 155.785 ;
        RECT 85.505 155.325 85.905 156.125 ;
        RECT 86.075 156.855 87.030 157.075 ;
        RECT 86.075 155.955 86.285 156.855 ;
        RECT 86.455 156.125 87.145 156.685 ;
        RECT 87.315 156.540 87.605 157.705 ;
        RECT 88.235 156.565 88.505 157.535 ;
        RECT 88.715 156.905 88.995 157.705 ;
        RECT 89.165 157.195 90.820 157.485 ;
        RECT 91.000 157.195 92.655 157.485 ;
        RECT 89.230 156.855 90.820 157.025 ;
        RECT 89.230 156.735 89.400 156.855 ;
        RECT 88.675 156.565 89.400 156.735 ;
        RECT 86.075 155.785 87.030 155.955 ;
        RECT 86.305 155.155 86.575 155.615 ;
        RECT 86.745 155.325 87.030 155.785 ;
        RECT 87.315 155.155 87.605 155.880 ;
        RECT 88.235 155.830 88.405 156.565 ;
        RECT 88.675 156.395 88.845 156.565 ;
        RECT 88.575 156.065 88.845 156.395 ;
        RECT 89.015 156.065 89.420 156.395 ;
        RECT 89.590 156.065 90.300 156.685 ;
        RECT 90.500 156.565 90.820 156.855 ;
        RECT 91.000 156.855 92.590 157.025 ;
        RECT 92.825 156.905 93.105 157.705 ;
        RECT 91.000 156.565 91.320 156.855 ;
        RECT 92.420 156.735 92.590 156.855 ;
        RECT 88.675 155.895 88.845 156.065 ;
        RECT 88.235 155.485 88.505 155.830 ;
        RECT 88.675 155.725 90.285 155.895 ;
        RECT 90.470 155.825 90.820 156.395 ;
        RECT 91.000 155.825 91.350 156.395 ;
        RECT 91.520 156.065 92.230 156.685 ;
        RECT 92.420 156.565 93.145 156.735 ;
        RECT 93.315 156.565 93.585 157.535 ;
        RECT 92.975 156.395 93.145 156.565 ;
        RECT 92.400 156.065 92.805 156.395 ;
        RECT 92.975 156.065 93.245 156.395 ;
        RECT 92.975 155.895 93.145 156.065 ;
        RECT 88.695 155.155 89.075 155.555 ;
        RECT 89.245 155.375 89.415 155.725 ;
        RECT 89.585 155.155 89.915 155.555 ;
        RECT 90.115 155.375 90.285 155.725 ;
        RECT 91.535 155.725 93.145 155.895 ;
        RECT 93.415 155.830 93.585 156.565 ;
        RECT 90.485 155.155 90.815 155.655 ;
        RECT 91.005 155.155 91.335 155.655 ;
        RECT 91.535 155.375 91.705 155.725 ;
        RECT 91.905 155.155 92.235 155.555 ;
        RECT 92.405 155.375 92.575 155.725 ;
        RECT 92.745 155.155 93.125 155.555 ;
        RECT 93.315 155.485 93.585 155.830 ;
        RECT 93.755 156.565 94.095 157.535 ;
        RECT 94.265 156.565 94.435 157.705 ;
        RECT 94.705 156.905 94.955 157.705 ;
        RECT 95.600 156.735 95.930 157.535 ;
        RECT 96.230 156.905 96.560 157.705 ;
        RECT 96.730 156.735 97.060 157.535 ;
        RECT 94.625 156.565 97.060 156.735 ;
        RECT 97.435 156.565 97.775 157.535 ;
        RECT 97.945 156.565 98.115 157.705 ;
        RECT 98.385 156.905 98.635 157.705 ;
        RECT 99.280 156.735 99.610 157.535 ;
        RECT 99.910 156.905 100.240 157.705 ;
        RECT 100.410 156.735 100.740 157.535 ;
        RECT 98.305 156.565 100.740 156.735 ;
        RECT 101.155 156.565 101.385 157.705 ;
        RECT 93.755 156.005 93.930 156.565 ;
        RECT 94.625 156.315 94.795 156.565 ;
        RECT 94.100 156.145 94.795 156.315 ;
        RECT 94.970 156.145 95.390 156.345 ;
        RECT 95.560 156.145 95.890 156.345 ;
        RECT 96.060 156.145 96.390 156.345 ;
        RECT 93.755 155.955 93.985 156.005 ;
        RECT 93.755 155.325 94.095 155.955 ;
        RECT 94.265 155.155 94.515 155.955 ;
        RECT 94.705 155.805 95.930 155.975 ;
        RECT 94.705 155.325 95.035 155.805 ;
        RECT 95.205 155.155 95.430 155.615 ;
        RECT 95.600 155.325 95.930 155.805 ;
        RECT 96.560 155.935 96.730 156.565 ;
        RECT 96.915 156.145 97.265 156.395 ;
        RECT 97.435 155.955 97.610 156.565 ;
        RECT 98.305 156.315 98.475 156.565 ;
        RECT 97.780 156.145 98.475 156.315 ;
        RECT 98.650 156.145 99.070 156.345 ;
        RECT 99.240 156.145 99.570 156.345 ;
        RECT 99.740 156.145 100.070 156.345 ;
        RECT 96.560 155.325 97.060 155.935 ;
        RECT 97.435 155.325 97.775 155.955 ;
        RECT 97.945 155.155 98.195 155.955 ;
        RECT 98.385 155.805 99.610 155.975 ;
        RECT 98.385 155.325 98.715 155.805 ;
        RECT 98.885 155.155 99.110 155.615 ;
        RECT 99.280 155.325 99.610 155.805 ;
        RECT 100.240 155.935 100.410 156.565 ;
        RECT 101.555 156.555 101.885 157.535 ;
        RECT 102.055 156.565 102.265 157.705 ;
        RECT 102.870 157.365 103.125 157.395 ;
        RECT 102.785 157.195 103.125 157.365 ;
        RECT 102.870 156.725 103.125 157.195 ;
        RECT 103.305 156.905 103.590 157.705 ;
        RECT 103.770 156.985 104.100 157.495 ;
        RECT 100.595 156.145 100.945 156.395 ;
        RECT 101.135 156.145 101.465 156.395 ;
        RECT 100.240 155.325 100.740 155.935 ;
        RECT 101.155 155.155 101.385 155.975 ;
        RECT 101.635 155.955 101.885 156.555 ;
        RECT 101.555 155.325 101.885 155.955 ;
        RECT 102.055 155.155 102.265 155.975 ;
        RECT 102.870 155.865 103.050 156.725 ;
        RECT 103.770 156.395 104.020 156.985 ;
        RECT 104.370 156.835 104.540 157.445 ;
        RECT 104.710 157.015 105.040 157.705 ;
        RECT 105.270 157.155 105.510 157.445 ;
        RECT 105.710 157.325 106.130 157.705 ;
        RECT 106.310 157.235 106.940 157.485 ;
        RECT 107.410 157.325 107.740 157.705 ;
        RECT 106.310 157.155 106.480 157.235 ;
        RECT 107.910 157.155 108.080 157.445 ;
        RECT 108.260 157.325 108.640 157.705 ;
        RECT 108.880 157.320 109.710 157.490 ;
        RECT 105.270 156.985 106.480 157.155 ;
        RECT 103.220 156.065 104.020 156.395 ;
        RECT 102.870 155.335 103.125 155.865 ;
        RECT 103.305 155.155 103.590 155.615 ;
        RECT 103.770 155.415 104.020 156.065 ;
        RECT 104.220 156.815 104.540 156.835 ;
        RECT 104.220 156.645 106.140 156.815 ;
        RECT 104.220 155.750 104.410 156.645 ;
        RECT 106.310 156.475 106.480 156.985 ;
        RECT 106.650 156.725 107.170 157.035 ;
        RECT 104.580 156.305 106.480 156.475 ;
        RECT 104.580 156.245 104.910 156.305 ;
        RECT 105.060 156.075 105.390 156.135 ;
        RECT 104.730 155.805 105.390 156.075 ;
        RECT 104.220 155.420 104.540 155.750 ;
        RECT 104.720 155.155 105.380 155.635 ;
        RECT 105.580 155.545 105.750 156.305 ;
        RECT 106.650 156.135 106.830 156.545 ;
        RECT 105.920 155.965 106.250 156.085 ;
        RECT 107.000 155.965 107.170 156.725 ;
        RECT 105.920 155.795 107.170 155.965 ;
        RECT 107.340 156.905 108.710 157.155 ;
        RECT 107.340 156.135 107.530 156.905 ;
        RECT 108.460 156.645 108.710 156.905 ;
        RECT 107.700 156.475 107.950 156.635 ;
        RECT 108.880 156.475 109.050 157.320 ;
        RECT 109.945 157.035 110.115 157.535 ;
        RECT 110.285 157.205 110.615 157.705 ;
        RECT 109.220 156.645 109.720 157.025 ;
        RECT 109.945 156.865 110.640 157.035 ;
        RECT 107.700 156.305 109.050 156.475 ;
        RECT 108.630 156.265 109.050 156.305 ;
        RECT 107.340 155.795 107.760 156.135 ;
        RECT 108.050 155.805 108.460 156.135 ;
        RECT 105.580 155.375 106.430 155.545 ;
        RECT 106.990 155.155 107.310 155.615 ;
        RECT 107.510 155.365 107.760 155.795 ;
        RECT 108.050 155.155 108.460 155.595 ;
        RECT 108.630 155.535 108.800 156.265 ;
        RECT 108.970 155.715 109.320 156.085 ;
        RECT 109.500 155.775 109.720 156.645 ;
        RECT 109.890 156.075 110.300 156.695 ;
        RECT 110.470 155.895 110.640 156.865 ;
        RECT 109.945 155.705 110.640 155.895 ;
        RECT 108.630 155.335 109.645 155.535 ;
        RECT 109.945 155.375 110.115 155.705 ;
        RECT 110.285 155.155 110.615 155.535 ;
        RECT 110.830 155.415 111.055 157.535 ;
        RECT 111.225 157.205 111.555 157.705 ;
        RECT 111.725 157.035 111.895 157.535 ;
        RECT 111.230 156.865 111.895 157.035 ;
        RECT 111.230 155.875 111.460 156.865 ;
        RECT 111.630 156.045 111.980 156.695 ;
        RECT 112.155 156.615 113.365 157.705 ;
        RECT 112.155 156.075 112.675 156.615 ;
        RECT 112.845 155.905 113.365 156.445 ;
        RECT 111.230 155.705 111.895 155.875 ;
        RECT 111.225 155.155 111.555 155.535 ;
        RECT 111.725 155.415 111.895 155.705 ;
        RECT 112.155 155.155 113.365 155.905 ;
        RECT 26.970 154.985 113.450 155.155 ;
        RECT 27.055 154.235 28.265 154.985 ;
        RECT 28.810 154.275 29.065 154.805 ;
        RECT 29.245 154.525 29.530 154.985 ;
        RECT 27.055 153.695 27.575 154.235 ;
        RECT 27.745 153.525 28.265 154.065 ;
        RECT 27.055 152.435 28.265 153.525 ;
        RECT 28.810 153.415 28.990 154.275 ;
        RECT 29.710 154.075 29.960 154.725 ;
        RECT 29.160 153.745 29.960 154.075 ;
        RECT 28.810 152.945 29.065 153.415 ;
        RECT 28.725 152.775 29.065 152.945 ;
        RECT 28.810 152.745 29.065 152.775 ;
        RECT 29.245 152.435 29.530 153.235 ;
        RECT 29.710 153.155 29.960 153.745 ;
        RECT 30.160 154.390 30.480 154.720 ;
        RECT 30.660 154.505 31.320 154.985 ;
        RECT 31.520 154.595 32.370 154.765 ;
        RECT 30.160 153.495 30.350 154.390 ;
        RECT 30.670 154.065 31.330 154.335 ;
        RECT 31.000 154.005 31.330 154.065 ;
        RECT 30.520 153.835 30.850 153.895 ;
        RECT 31.520 153.835 31.690 154.595 ;
        RECT 32.930 154.525 33.250 154.985 ;
        RECT 33.450 154.345 33.700 154.775 ;
        RECT 33.990 154.545 34.400 154.985 ;
        RECT 34.570 154.605 35.585 154.805 ;
        RECT 31.860 154.175 33.110 154.345 ;
        RECT 31.860 154.055 32.190 154.175 ;
        RECT 30.520 153.665 32.420 153.835 ;
        RECT 30.160 153.325 32.080 153.495 ;
        RECT 30.160 153.305 30.480 153.325 ;
        RECT 29.710 152.645 30.040 153.155 ;
        RECT 30.310 152.695 30.480 153.305 ;
        RECT 32.250 153.155 32.420 153.665 ;
        RECT 32.590 153.595 32.770 154.005 ;
        RECT 32.940 153.415 33.110 154.175 ;
        RECT 30.650 152.435 30.980 153.125 ;
        RECT 31.210 152.985 32.420 153.155 ;
        RECT 32.590 153.105 33.110 153.415 ;
        RECT 33.280 154.005 33.700 154.345 ;
        RECT 33.990 154.005 34.400 154.335 ;
        RECT 33.280 153.235 33.470 154.005 ;
        RECT 34.570 153.875 34.740 154.605 ;
        RECT 35.885 154.435 36.055 154.765 ;
        RECT 36.225 154.605 36.555 154.985 ;
        RECT 34.910 154.055 35.260 154.425 ;
        RECT 34.570 153.835 34.990 153.875 ;
        RECT 33.640 153.665 34.990 153.835 ;
        RECT 33.640 153.505 33.890 153.665 ;
        RECT 34.400 153.235 34.650 153.495 ;
        RECT 33.280 152.985 34.650 153.235 ;
        RECT 31.210 152.695 31.450 152.985 ;
        RECT 32.250 152.905 32.420 152.985 ;
        RECT 31.650 152.435 32.070 152.815 ;
        RECT 32.250 152.655 32.880 152.905 ;
        RECT 33.350 152.435 33.680 152.815 ;
        RECT 33.850 152.695 34.020 152.985 ;
        RECT 34.820 152.820 34.990 153.665 ;
        RECT 35.440 153.495 35.660 154.365 ;
        RECT 35.885 154.245 36.580 154.435 ;
        RECT 35.160 153.115 35.660 153.495 ;
        RECT 35.830 153.445 36.240 154.065 ;
        RECT 36.410 153.275 36.580 154.245 ;
        RECT 35.885 153.105 36.580 153.275 ;
        RECT 34.200 152.435 34.580 152.815 ;
        RECT 34.820 152.650 35.650 152.820 ;
        RECT 35.885 152.605 36.055 153.105 ;
        RECT 36.225 152.435 36.555 152.935 ;
        RECT 36.770 152.605 36.995 154.725 ;
        RECT 37.165 154.605 37.495 154.985 ;
        RECT 37.665 154.435 37.835 154.725 ;
        RECT 38.155 154.505 38.435 154.985 ;
        RECT 37.170 154.265 37.835 154.435 ;
        RECT 38.605 154.335 38.865 154.725 ;
        RECT 39.040 154.505 39.295 154.985 ;
        RECT 39.465 154.335 39.760 154.725 ;
        RECT 39.940 154.505 40.215 154.985 ;
        RECT 40.385 154.485 40.685 154.815 ;
        RECT 37.170 153.275 37.400 154.265 ;
        RECT 38.110 154.165 39.760 154.335 ;
        RECT 37.570 153.445 37.920 154.095 ;
        RECT 38.110 153.655 38.515 154.165 ;
        RECT 38.685 153.825 39.825 153.995 ;
        RECT 38.110 153.485 38.865 153.655 ;
        RECT 37.170 153.105 37.835 153.275 ;
        RECT 37.165 152.435 37.495 152.935 ;
        RECT 37.665 152.605 37.835 153.105 ;
        RECT 38.150 152.435 38.435 153.305 ;
        RECT 38.605 153.235 38.865 153.485 ;
        RECT 39.655 153.575 39.825 153.825 ;
        RECT 39.995 153.745 40.345 154.315 ;
        RECT 40.515 153.575 40.685 154.485 ;
        RECT 39.655 153.405 40.685 153.575 ;
        RECT 38.605 153.065 39.725 153.235 ;
        RECT 38.605 152.605 38.865 153.065 ;
        RECT 39.040 152.435 39.295 152.895 ;
        RECT 39.465 152.605 39.725 153.065 ;
        RECT 39.895 152.435 40.205 153.235 ;
        RECT 40.375 152.605 40.685 153.405 ;
        RECT 40.860 154.245 41.115 154.815 ;
        RECT 41.285 154.585 41.615 154.985 ;
        RECT 42.040 154.450 42.570 154.815 ;
        RECT 42.760 154.645 43.035 154.815 ;
        RECT 42.755 154.475 43.035 154.645 ;
        RECT 42.040 154.415 42.215 154.450 ;
        RECT 41.285 154.245 42.215 154.415 ;
        RECT 40.860 153.575 41.030 154.245 ;
        RECT 41.285 154.075 41.455 154.245 ;
        RECT 41.200 153.745 41.455 154.075 ;
        RECT 41.680 153.745 41.875 154.075 ;
        RECT 40.860 152.605 41.195 153.575 ;
        RECT 41.365 152.435 41.535 153.575 ;
        RECT 41.705 152.775 41.875 153.745 ;
        RECT 42.045 153.115 42.215 154.245 ;
        RECT 42.385 153.455 42.555 154.255 ;
        RECT 42.760 153.655 43.035 154.475 ;
        RECT 43.205 153.455 43.395 154.815 ;
        RECT 43.575 154.450 44.085 154.985 ;
        RECT 44.305 154.175 44.550 154.780 ;
        RECT 45.925 154.485 46.255 154.985 ;
        RECT 46.455 154.415 46.625 154.765 ;
        RECT 46.825 154.585 47.155 154.985 ;
        RECT 47.325 154.415 47.495 154.765 ;
        RECT 47.665 154.585 48.045 154.985 ;
        RECT 43.595 154.005 44.825 154.175 ;
        RECT 42.385 153.285 43.395 153.455 ;
        RECT 43.565 153.440 44.315 153.630 ;
        RECT 42.045 152.945 43.170 153.115 ;
        RECT 43.565 152.775 43.735 153.440 ;
        RECT 44.485 153.195 44.825 154.005 ;
        RECT 45.920 153.745 46.270 154.315 ;
        RECT 46.455 154.245 48.065 154.415 ;
        RECT 48.235 154.310 48.505 154.655 ;
        RECT 47.895 154.075 48.065 154.245 ;
        RECT 41.705 152.605 43.735 152.775 ;
        RECT 43.905 152.435 44.075 153.195 ;
        RECT 44.310 152.785 44.825 153.195 ;
        RECT 45.920 153.285 46.240 153.575 ;
        RECT 46.440 153.455 47.150 154.075 ;
        RECT 47.320 153.745 47.725 154.075 ;
        RECT 47.895 153.745 48.165 154.075 ;
        RECT 47.895 153.575 48.065 153.745 ;
        RECT 48.335 153.575 48.505 154.310 ;
        RECT 48.675 154.260 48.965 154.985 ;
        RECT 49.135 154.525 49.695 154.815 ;
        RECT 49.865 154.525 50.115 154.985 ;
        RECT 47.340 153.405 48.065 153.575 ;
        RECT 47.340 153.285 47.510 153.405 ;
        RECT 45.920 153.115 47.510 153.285 ;
        RECT 45.920 152.655 47.575 152.945 ;
        RECT 47.745 152.435 48.025 153.235 ;
        RECT 48.235 152.605 48.505 153.575 ;
        RECT 48.675 152.435 48.965 153.600 ;
        RECT 49.135 153.155 49.385 154.525 ;
        RECT 50.735 154.355 51.065 154.715 ;
        RECT 51.810 154.645 52.065 154.805 ;
        RECT 51.725 154.475 52.065 154.645 ;
        RECT 52.245 154.525 52.530 154.985 ;
        RECT 49.675 154.165 51.065 154.355 ;
        RECT 51.810 154.275 52.065 154.475 ;
        RECT 49.675 154.075 49.845 154.165 ;
        RECT 49.555 153.745 49.845 154.075 ;
        RECT 50.015 153.745 50.355 153.995 ;
        RECT 50.575 153.745 51.250 153.995 ;
        RECT 49.675 153.495 49.845 153.745 ;
        RECT 49.675 153.325 50.615 153.495 ;
        RECT 50.985 153.385 51.250 153.745 ;
        RECT 51.810 153.415 51.990 154.275 ;
        RECT 52.710 154.075 52.960 154.725 ;
        RECT 52.160 153.745 52.960 154.075 ;
        RECT 49.135 152.605 49.595 153.155 ;
        RECT 49.785 152.435 50.115 153.155 ;
        RECT 50.315 152.775 50.615 153.325 ;
        RECT 50.785 152.435 51.065 153.105 ;
        RECT 51.810 152.745 52.065 153.415 ;
        RECT 52.245 152.435 52.530 153.235 ;
        RECT 52.710 153.155 52.960 153.745 ;
        RECT 53.160 154.390 53.480 154.720 ;
        RECT 53.660 154.505 54.320 154.985 ;
        RECT 54.520 154.595 55.370 154.765 ;
        RECT 53.160 153.495 53.350 154.390 ;
        RECT 53.670 154.065 54.330 154.335 ;
        RECT 54.000 154.005 54.330 154.065 ;
        RECT 53.520 153.835 53.850 153.895 ;
        RECT 54.520 153.835 54.690 154.595 ;
        RECT 55.930 154.525 56.250 154.985 ;
        RECT 56.450 154.345 56.700 154.775 ;
        RECT 56.990 154.545 57.400 154.985 ;
        RECT 57.570 154.605 58.585 154.805 ;
        RECT 54.860 154.175 56.110 154.345 ;
        RECT 54.860 154.055 55.190 154.175 ;
        RECT 53.520 153.665 55.420 153.835 ;
        RECT 53.160 153.325 55.080 153.495 ;
        RECT 53.160 153.305 53.480 153.325 ;
        RECT 52.710 152.645 53.040 153.155 ;
        RECT 53.310 152.695 53.480 153.305 ;
        RECT 55.250 153.155 55.420 153.665 ;
        RECT 55.590 153.595 55.770 154.005 ;
        RECT 55.940 153.415 56.110 154.175 ;
        RECT 53.650 152.435 53.980 153.125 ;
        RECT 54.210 152.985 55.420 153.155 ;
        RECT 55.590 153.105 56.110 153.415 ;
        RECT 56.280 154.005 56.700 154.345 ;
        RECT 56.990 154.005 57.400 154.335 ;
        RECT 56.280 153.235 56.470 154.005 ;
        RECT 57.570 153.875 57.740 154.605 ;
        RECT 58.885 154.435 59.055 154.765 ;
        RECT 59.225 154.605 59.555 154.985 ;
        RECT 57.910 154.055 58.260 154.425 ;
        RECT 57.570 153.835 57.990 153.875 ;
        RECT 56.640 153.665 57.990 153.835 ;
        RECT 56.640 153.505 56.890 153.665 ;
        RECT 57.400 153.235 57.650 153.495 ;
        RECT 56.280 152.985 57.650 153.235 ;
        RECT 54.210 152.695 54.450 152.985 ;
        RECT 55.250 152.905 55.420 152.985 ;
        RECT 54.650 152.435 55.070 152.815 ;
        RECT 55.250 152.655 55.880 152.905 ;
        RECT 56.350 152.435 56.680 152.815 ;
        RECT 56.850 152.695 57.020 152.985 ;
        RECT 57.820 152.820 57.990 153.665 ;
        RECT 58.440 153.495 58.660 154.365 ;
        RECT 58.885 154.245 59.580 154.435 ;
        RECT 58.160 153.115 58.660 153.495 ;
        RECT 58.830 153.445 59.240 154.065 ;
        RECT 59.410 153.275 59.580 154.245 ;
        RECT 58.885 153.105 59.580 153.275 ;
        RECT 57.200 152.435 57.580 152.815 ;
        RECT 57.820 152.650 58.650 152.820 ;
        RECT 58.885 152.605 59.055 153.105 ;
        RECT 59.225 152.435 59.555 152.935 ;
        RECT 59.770 152.605 59.995 154.725 ;
        RECT 60.165 154.605 60.495 154.985 ;
        RECT 60.665 154.435 60.835 154.725 ;
        RECT 60.170 154.265 60.835 154.435 ;
        RECT 62.020 154.275 62.275 154.805 ;
        RECT 62.445 154.525 62.750 154.985 ;
        RECT 62.995 154.605 64.065 154.775 ;
        RECT 60.170 153.275 60.400 154.265 ;
        RECT 60.570 153.445 60.920 154.095 ;
        RECT 62.020 153.625 62.230 154.275 ;
        RECT 62.995 154.250 63.315 154.605 ;
        RECT 62.990 154.075 63.315 154.250 ;
        RECT 62.400 153.775 63.315 154.075 ;
        RECT 63.485 154.035 63.725 154.435 ;
        RECT 63.895 154.375 64.065 154.605 ;
        RECT 64.235 154.545 64.425 154.985 ;
        RECT 64.595 154.535 65.545 154.815 ;
        RECT 65.765 154.625 66.115 154.795 ;
        RECT 63.895 154.205 64.425 154.375 ;
        RECT 62.400 153.745 63.140 153.775 ;
        RECT 60.170 153.105 60.835 153.275 ;
        RECT 60.165 152.435 60.495 152.935 ;
        RECT 60.665 152.605 60.835 153.105 ;
        RECT 62.020 152.745 62.275 153.625 ;
        RECT 62.445 152.435 62.750 153.575 ;
        RECT 62.970 153.155 63.140 153.745 ;
        RECT 63.485 153.665 64.025 154.035 ;
        RECT 64.205 153.925 64.425 154.205 ;
        RECT 64.595 153.755 64.765 154.535 ;
        RECT 64.360 153.585 64.765 153.755 ;
        RECT 64.935 153.745 65.285 154.365 ;
        RECT 64.360 153.495 64.530 153.585 ;
        RECT 65.455 153.575 65.665 154.365 ;
        RECT 63.310 153.325 64.530 153.495 ;
        RECT 64.990 153.415 65.665 153.575 ;
        RECT 62.970 152.985 63.770 153.155 ;
        RECT 63.090 152.435 63.420 152.815 ;
        RECT 63.600 152.695 63.770 152.985 ;
        RECT 64.360 152.945 64.530 153.325 ;
        RECT 64.700 153.405 65.665 153.415 ;
        RECT 65.855 154.235 66.115 154.625 ;
        RECT 66.325 154.525 66.655 154.985 ;
        RECT 67.530 154.595 68.385 154.765 ;
        RECT 68.590 154.595 69.085 154.765 ;
        RECT 69.255 154.625 69.585 154.985 ;
        RECT 65.855 153.545 66.025 154.235 ;
        RECT 66.195 153.885 66.365 154.065 ;
        RECT 66.535 154.055 67.325 154.305 ;
        RECT 67.530 153.885 67.700 154.595 ;
        RECT 67.870 154.085 68.225 154.305 ;
        RECT 66.195 153.715 67.885 153.885 ;
        RECT 64.700 153.115 65.160 153.405 ;
        RECT 65.855 153.375 67.355 153.545 ;
        RECT 65.855 153.235 66.025 153.375 ;
        RECT 65.465 153.065 66.025 153.235 ;
        RECT 63.940 152.435 64.190 152.895 ;
        RECT 64.360 152.605 65.230 152.945 ;
        RECT 65.465 152.605 65.635 153.065 ;
        RECT 66.470 153.035 67.545 153.205 ;
        RECT 65.805 152.435 66.175 152.895 ;
        RECT 66.470 152.695 66.640 153.035 ;
        RECT 66.810 152.435 67.140 152.865 ;
        RECT 67.375 152.695 67.545 153.035 ;
        RECT 67.715 152.935 67.885 153.715 ;
        RECT 68.055 153.495 68.225 154.085 ;
        RECT 68.395 153.685 68.745 154.305 ;
        RECT 68.055 153.105 68.520 153.495 ;
        RECT 68.915 153.235 69.085 154.595 ;
        RECT 69.255 153.405 69.715 154.455 ;
        RECT 68.690 153.065 69.085 153.235 ;
        RECT 68.690 152.935 68.860 153.065 ;
        RECT 67.715 152.605 68.395 152.935 ;
        RECT 68.610 152.605 68.860 152.935 ;
        RECT 69.030 152.435 69.280 152.895 ;
        RECT 69.450 152.620 69.775 153.405 ;
        RECT 69.945 152.605 70.115 154.725 ;
        RECT 70.285 154.605 70.615 154.985 ;
        RECT 70.785 154.435 71.040 154.725 ;
        RECT 70.290 154.265 71.040 154.435 ;
        RECT 71.675 154.310 71.945 154.655 ;
        RECT 72.135 154.585 72.515 154.985 ;
        RECT 72.685 154.415 72.855 154.765 ;
        RECT 73.025 154.585 73.355 154.985 ;
        RECT 73.555 154.415 73.725 154.765 ;
        RECT 73.925 154.485 74.255 154.985 ;
        RECT 70.290 153.275 70.520 154.265 ;
        RECT 70.690 153.445 71.040 154.095 ;
        RECT 71.675 153.575 71.845 154.310 ;
        RECT 72.115 154.245 73.725 154.415 ;
        RECT 72.115 154.075 72.285 154.245 ;
        RECT 72.015 153.745 72.285 154.075 ;
        RECT 72.455 153.745 72.860 154.075 ;
        RECT 72.115 153.575 72.285 153.745 ;
        RECT 73.030 153.625 73.740 154.075 ;
        RECT 73.910 153.745 74.260 154.315 ;
        RECT 74.435 154.260 74.725 154.985 ;
        RECT 74.895 154.185 75.235 154.815 ;
        RECT 75.405 154.185 75.655 154.985 ;
        RECT 75.845 154.335 76.175 154.815 ;
        RECT 76.345 154.525 76.570 154.985 ;
        RECT 76.740 154.335 77.070 154.815 ;
        RECT 74.895 154.135 75.125 154.185 ;
        RECT 75.845 154.165 77.070 154.335 ;
        RECT 77.700 154.205 78.200 154.815 ;
        RECT 78.950 154.275 79.205 154.805 ;
        RECT 79.385 154.525 79.670 154.985 ;
        RECT 70.290 153.105 71.040 153.275 ;
        RECT 70.285 152.435 70.615 152.935 ;
        RECT 70.785 152.605 71.040 153.105 ;
        RECT 71.675 152.605 71.945 153.575 ;
        RECT 72.115 153.405 72.840 153.575 ;
        RECT 73.030 153.455 73.745 153.625 ;
        RECT 72.670 153.285 72.840 153.405 ;
        RECT 73.940 153.285 74.260 153.575 ;
        RECT 72.155 152.435 72.435 153.235 ;
        RECT 72.670 153.115 74.260 153.285 ;
        RECT 72.605 152.655 74.260 152.945 ;
        RECT 74.435 152.435 74.725 153.600 ;
        RECT 74.895 153.575 75.070 154.135 ;
        RECT 75.240 153.825 75.935 153.995 ;
        RECT 75.765 153.575 75.935 153.825 ;
        RECT 76.110 153.795 76.530 153.995 ;
        RECT 76.700 153.795 77.030 153.995 ;
        RECT 77.200 153.795 77.530 153.995 ;
        RECT 77.700 153.575 77.870 154.205 ;
        RECT 78.055 153.745 78.405 153.995 ;
        RECT 74.895 152.605 75.235 153.575 ;
        RECT 75.405 152.435 75.575 153.575 ;
        RECT 75.765 153.405 78.200 153.575 ;
        RECT 75.845 152.435 76.095 153.235 ;
        RECT 76.740 152.605 77.070 153.405 ;
        RECT 77.370 152.435 77.700 153.235 ;
        RECT 77.870 152.605 78.200 153.405 ;
        RECT 78.950 153.415 79.130 154.275 ;
        RECT 79.850 154.075 80.100 154.725 ;
        RECT 79.300 153.745 80.100 154.075 ;
        RECT 78.950 152.945 79.205 153.415 ;
        RECT 78.865 152.775 79.205 152.945 ;
        RECT 78.950 152.745 79.205 152.775 ;
        RECT 79.385 152.435 79.670 153.235 ;
        RECT 79.850 153.155 80.100 153.745 ;
        RECT 80.300 154.390 80.620 154.720 ;
        RECT 80.800 154.505 81.460 154.985 ;
        RECT 81.660 154.595 82.510 154.765 ;
        RECT 80.300 153.495 80.490 154.390 ;
        RECT 80.810 154.065 81.470 154.335 ;
        RECT 81.140 154.005 81.470 154.065 ;
        RECT 80.660 153.835 80.990 153.895 ;
        RECT 81.660 153.835 81.830 154.595 ;
        RECT 83.070 154.525 83.390 154.985 ;
        RECT 83.590 154.345 83.840 154.775 ;
        RECT 84.130 154.545 84.540 154.985 ;
        RECT 84.710 154.605 85.725 154.805 ;
        RECT 82.000 154.175 83.250 154.345 ;
        RECT 82.000 154.055 82.330 154.175 ;
        RECT 80.660 153.665 82.560 153.835 ;
        RECT 80.300 153.325 82.220 153.495 ;
        RECT 80.300 153.305 80.620 153.325 ;
        RECT 79.850 152.645 80.180 153.155 ;
        RECT 80.450 152.695 80.620 153.305 ;
        RECT 82.390 153.155 82.560 153.665 ;
        RECT 82.730 153.595 82.910 154.005 ;
        RECT 83.080 153.415 83.250 154.175 ;
        RECT 80.790 152.435 81.120 153.125 ;
        RECT 81.350 152.985 82.560 153.155 ;
        RECT 82.730 153.105 83.250 153.415 ;
        RECT 83.420 154.005 83.840 154.345 ;
        RECT 84.130 154.005 84.540 154.335 ;
        RECT 83.420 153.235 83.610 154.005 ;
        RECT 84.710 153.875 84.880 154.605 ;
        RECT 86.025 154.435 86.195 154.765 ;
        RECT 86.365 154.605 86.695 154.985 ;
        RECT 85.050 154.055 85.400 154.425 ;
        RECT 84.710 153.835 85.130 153.875 ;
        RECT 83.780 153.665 85.130 153.835 ;
        RECT 83.780 153.505 84.030 153.665 ;
        RECT 84.540 153.235 84.790 153.495 ;
        RECT 83.420 152.985 84.790 153.235 ;
        RECT 81.350 152.695 81.590 152.985 ;
        RECT 82.390 152.905 82.560 152.985 ;
        RECT 81.790 152.435 82.210 152.815 ;
        RECT 82.390 152.655 83.020 152.905 ;
        RECT 83.490 152.435 83.820 152.815 ;
        RECT 83.990 152.695 84.160 152.985 ;
        RECT 84.960 152.820 85.130 153.665 ;
        RECT 85.580 153.495 85.800 154.365 ;
        RECT 86.025 154.245 86.720 154.435 ;
        RECT 85.300 153.115 85.800 153.495 ;
        RECT 85.970 153.445 86.380 154.065 ;
        RECT 86.550 153.275 86.720 154.245 ;
        RECT 86.025 153.105 86.720 153.275 ;
        RECT 84.340 152.435 84.720 152.815 ;
        RECT 84.960 152.650 85.790 152.820 ;
        RECT 86.025 152.605 86.195 153.105 ;
        RECT 86.365 152.435 86.695 152.935 ;
        RECT 86.910 152.605 87.135 154.725 ;
        RECT 87.305 154.605 87.635 154.985 ;
        RECT 87.805 154.435 87.975 154.725 ;
        RECT 87.310 154.265 87.975 154.435 ;
        RECT 88.235 154.310 88.495 154.815 ;
        RECT 88.675 154.605 89.005 154.985 ;
        RECT 89.185 154.435 89.355 154.815 ;
        RECT 89.625 154.485 89.955 154.985 ;
        RECT 87.310 153.275 87.540 154.265 ;
        RECT 87.710 153.445 88.060 154.095 ;
        RECT 88.235 153.510 88.405 154.310 ;
        RECT 88.690 154.265 89.355 154.435 ;
        RECT 90.155 154.415 90.325 154.765 ;
        RECT 90.525 154.585 90.855 154.985 ;
        RECT 91.025 154.415 91.195 154.765 ;
        RECT 91.365 154.585 91.745 154.985 ;
        RECT 88.690 154.010 88.860 154.265 ;
        RECT 88.575 153.680 88.860 154.010 ;
        RECT 89.095 153.715 89.425 154.085 ;
        RECT 89.620 153.745 89.970 154.315 ;
        RECT 90.155 154.245 91.765 154.415 ;
        RECT 91.935 154.310 92.205 154.655 ;
        RECT 91.595 154.075 91.765 154.245 ;
        RECT 88.690 153.535 88.860 153.680 ;
        RECT 87.310 153.105 87.975 153.275 ;
        RECT 87.305 152.435 87.635 152.935 ;
        RECT 87.805 152.605 87.975 153.105 ;
        RECT 88.235 152.605 88.505 153.510 ;
        RECT 88.690 153.365 89.355 153.535 ;
        RECT 88.675 152.435 89.005 153.195 ;
        RECT 89.185 152.605 89.355 153.365 ;
        RECT 89.620 153.285 89.940 153.575 ;
        RECT 90.140 153.455 90.850 154.075 ;
        RECT 91.020 153.745 91.425 154.075 ;
        RECT 91.595 153.745 91.865 154.075 ;
        RECT 91.595 153.575 91.765 153.745 ;
        RECT 92.035 153.575 92.205 154.310 ;
        RECT 91.040 153.405 91.765 153.575 ;
        RECT 91.040 153.285 91.210 153.405 ;
        RECT 89.620 153.115 91.210 153.285 ;
        RECT 89.620 152.655 91.275 152.945 ;
        RECT 91.445 152.435 91.725 153.235 ;
        RECT 91.935 152.605 92.205 153.575 ;
        RECT 92.375 154.185 92.715 154.815 ;
        RECT 92.885 154.185 93.135 154.985 ;
        RECT 93.325 154.335 93.655 154.815 ;
        RECT 93.825 154.525 94.050 154.985 ;
        RECT 94.220 154.335 94.550 154.815 ;
        RECT 92.375 154.135 92.605 154.185 ;
        RECT 93.325 154.165 94.550 154.335 ;
        RECT 95.180 154.205 95.680 154.815 ;
        RECT 92.375 153.575 92.550 154.135 ;
        RECT 92.720 153.825 93.415 153.995 ;
        RECT 93.245 153.575 93.415 153.825 ;
        RECT 93.590 153.795 94.010 153.995 ;
        RECT 94.180 153.795 94.510 153.995 ;
        RECT 94.680 153.795 95.010 153.995 ;
        RECT 95.180 153.575 95.350 154.205 ;
        RECT 96.330 154.175 96.575 154.780 ;
        RECT 96.795 154.450 97.305 154.985 ;
        RECT 96.055 154.005 97.285 154.175 ;
        RECT 95.535 153.745 95.885 153.995 ;
        RECT 92.375 152.605 92.715 153.575 ;
        RECT 92.885 152.435 93.055 153.575 ;
        RECT 93.245 153.405 95.680 153.575 ;
        RECT 93.325 152.435 93.575 153.235 ;
        RECT 94.220 152.605 94.550 153.405 ;
        RECT 94.850 152.435 95.180 153.235 ;
        RECT 95.350 152.605 95.680 153.405 ;
        RECT 96.055 153.195 96.395 154.005 ;
        RECT 96.565 153.440 97.315 153.630 ;
        RECT 96.055 152.785 96.570 153.195 ;
        RECT 96.805 152.435 96.975 153.195 ;
        RECT 97.145 152.775 97.315 153.440 ;
        RECT 97.485 153.455 97.675 154.815 ;
        RECT 97.845 154.645 98.120 154.815 ;
        RECT 97.845 154.475 98.125 154.645 ;
        RECT 97.845 153.655 98.120 154.475 ;
        RECT 98.310 154.450 98.840 154.815 ;
        RECT 99.265 154.585 99.595 154.985 ;
        RECT 98.665 154.415 98.840 154.450 ;
        RECT 98.325 153.455 98.495 154.255 ;
        RECT 97.485 153.285 98.495 153.455 ;
        RECT 98.665 154.245 99.595 154.415 ;
        RECT 99.765 154.245 100.020 154.815 ;
        RECT 100.195 154.260 100.485 154.985 ;
        RECT 101.205 154.435 101.375 154.815 ;
        RECT 101.555 154.605 101.885 154.985 ;
        RECT 101.205 154.265 101.870 154.435 ;
        RECT 102.065 154.310 102.325 154.815 ;
        RECT 98.665 153.115 98.835 154.245 ;
        RECT 99.425 154.075 99.595 154.245 ;
        RECT 97.710 152.945 98.835 153.115 ;
        RECT 99.005 153.745 99.200 154.075 ;
        RECT 99.425 153.745 99.680 154.075 ;
        RECT 99.005 152.775 99.175 153.745 ;
        RECT 99.850 153.575 100.020 154.245 ;
        RECT 101.135 153.715 101.465 154.085 ;
        RECT 101.700 154.010 101.870 154.265 ;
        RECT 101.700 153.680 101.985 154.010 ;
        RECT 97.145 152.605 99.175 152.775 ;
        RECT 99.345 152.435 99.515 153.575 ;
        RECT 99.685 152.605 100.020 153.575 ;
        RECT 100.195 152.435 100.485 153.600 ;
        RECT 101.700 153.535 101.870 153.680 ;
        RECT 101.205 153.365 101.870 153.535 ;
        RECT 102.155 153.510 102.325 154.310 ;
        RECT 101.205 152.605 101.375 153.365 ;
        RECT 101.555 152.435 101.885 153.195 ;
        RECT 102.055 152.605 102.325 153.510 ;
        RECT 102.870 154.275 103.125 154.805 ;
        RECT 103.305 154.525 103.590 154.985 ;
        RECT 102.870 153.415 103.050 154.275 ;
        RECT 103.770 154.075 104.020 154.725 ;
        RECT 103.220 153.745 104.020 154.075 ;
        RECT 102.870 152.945 103.125 153.415 ;
        RECT 102.785 152.775 103.125 152.945 ;
        RECT 102.870 152.745 103.125 152.775 ;
        RECT 103.305 152.435 103.590 153.235 ;
        RECT 103.770 153.155 104.020 153.745 ;
        RECT 104.220 154.390 104.540 154.720 ;
        RECT 104.720 154.505 105.380 154.985 ;
        RECT 105.580 154.595 106.430 154.765 ;
        RECT 104.220 153.495 104.410 154.390 ;
        RECT 104.730 154.065 105.390 154.335 ;
        RECT 105.060 154.005 105.390 154.065 ;
        RECT 104.580 153.835 104.910 153.895 ;
        RECT 105.580 153.835 105.750 154.595 ;
        RECT 106.990 154.525 107.310 154.985 ;
        RECT 107.510 154.345 107.760 154.775 ;
        RECT 108.050 154.545 108.460 154.985 ;
        RECT 108.630 154.605 109.645 154.805 ;
        RECT 105.920 154.175 107.170 154.345 ;
        RECT 105.920 154.055 106.250 154.175 ;
        RECT 104.580 153.665 106.480 153.835 ;
        RECT 104.220 153.325 106.140 153.495 ;
        RECT 104.220 153.305 104.540 153.325 ;
        RECT 103.770 152.645 104.100 153.155 ;
        RECT 104.370 152.695 104.540 153.305 ;
        RECT 106.310 153.155 106.480 153.665 ;
        RECT 106.650 153.595 106.830 154.005 ;
        RECT 107.000 153.415 107.170 154.175 ;
        RECT 104.710 152.435 105.040 153.125 ;
        RECT 105.270 152.985 106.480 153.155 ;
        RECT 106.650 153.105 107.170 153.415 ;
        RECT 107.340 154.005 107.760 154.345 ;
        RECT 108.050 154.005 108.460 154.335 ;
        RECT 107.340 153.235 107.530 154.005 ;
        RECT 108.630 153.875 108.800 154.605 ;
        RECT 109.945 154.435 110.115 154.765 ;
        RECT 110.285 154.605 110.615 154.985 ;
        RECT 108.970 154.055 109.320 154.425 ;
        RECT 108.630 153.835 109.050 153.875 ;
        RECT 107.700 153.665 109.050 153.835 ;
        RECT 107.700 153.505 107.950 153.665 ;
        RECT 108.460 153.235 108.710 153.495 ;
        RECT 107.340 152.985 108.710 153.235 ;
        RECT 105.270 152.695 105.510 152.985 ;
        RECT 106.310 152.905 106.480 152.985 ;
        RECT 105.710 152.435 106.130 152.815 ;
        RECT 106.310 152.655 106.940 152.905 ;
        RECT 107.410 152.435 107.740 152.815 ;
        RECT 107.910 152.695 108.080 152.985 ;
        RECT 108.880 152.820 109.050 153.665 ;
        RECT 109.500 153.495 109.720 154.365 ;
        RECT 109.945 154.245 110.640 154.435 ;
        RECT 109.220 153.115 109.720 153.495 ;
        RECT 109.890 153.445 110.300 154.065 ;
        RECT 110.470 153.275 110.640 154.245 ;
        RECT 109.945 153.105 110.640 153.275 ;
        RECT 108.260 152.435 108.640 152.815 ;
        RECT 108.880 152.650 109.710 152.820 ;
        RECT 109.945 152.605 110.115 153.105 ;
        RECT 110.285 152.435 110.615 152.935 ;
        RECT 110.830 152.605 111.055 154.725 ;
        RECT 111.225 154.605 111.555 154.985 ;
        RECT 111.725 154.435 111.895 154.725 ;
        RECT 111.230 154.265 111.895 154.435 ;
        RECT 111.230 153.275 111.460 154.265 ;
        RECT 112.155 154.235 113.365 154.985 ;
        RECT 111.630 153.445 111.980 154.095 ;
        RECT 112.155 153.525 112.675 154.065 ;
        RECT 112.845 153.695 113.365 154.235 ;
        RECT 111.230 153.105 111.895 153.275 ;
        RECT 111.225 152.435 111.555 152.935 ;
        RECT 111.725 152.605 111.895 153.105 ;
        RECT 112.155 152.435 113.365 153.525 ;
        RECT 26.970 152.265 113.450 152.435 ;
        RECT 27.055 151.175 28.265 152.265 ;
        RECT 29.555 151.595 29.835 152.265 ;
        RECT 30.005 151.375 30.305 151.925 ;
        RECT 30.505 151.545 30.835 152.265 ;
        RECT 31.025 151.545 31.485 152.095 ;
        RECT 27.055 150.465 27.575 151.005 ;
        RECT 27.745 150.635 28.265 151.175 ;
        RECT 29.370 150.955 29.635 151.315 ;
        RECT 30.005 151.205 30.945 151.375 ;
        RECT 30.775 150.955 30.945 151.205 ;
        RECT 29.370 150.705 30.045 150.955 ;
        RECT 30.265 150.705 30.605 150.955 ;
        RECT 30.775 150.625 31.065 150.955 ;
        RECT 30.775 150.535 30.945 150.625 ;
        RECT 27.055 149.715 28.265 150.465 ;
        RECT 29.555 150.345 30.945 150.535 ;
        RECT 29.555 149.985 29.885 150.345 ;
        RECT 31.235 150.175 31.485 151.545 ;
        RECT 30.505 149.715 30.755 150.175 ;
        RECT 30.925 149.885 31.485 150.175 ;
        RECT 31.660 151.125 31.995 152.095 ;
        RECT 32.165 151.125 32.335 152.265 ;
        RECT 32.505 151.925 34.535 152.095 ;
        RECT 31.660 150.455 31.830 151.125 ;
        RECT 32.505 150.955 32.675 151.925 ;
        RECT 32.000 150.625 32.255 150.955 ;
        RECT 32.480 150.625 32.675 150.955 ;
        RECT 32.845 151.585 33.970 151.755 ;
        RECT 32.085 150.455 32.255 150.625 ;
        RECT 32.845 150.455 33.015 151.585 ;
        RECT 31.660 149.885 31.915 150.455 ;
        RECT 32.085 150.285 33.015 150.455 ;
        RECT 33.185 151.245 34.195 151.415 ;
        RECT 33.185 150.445 33.355 151.245 ;
        RECT 33.560 150.905 33.835 151.045 ;
        RECT 33.555 150.735 33.835 150.905 ;
        RECT 32.840 150.250 33.015 150.285 ;
        RECT 32.085 149.715 32.415 150.115 ;
        RECT 32.840 149.885 33.370 150.250 ;
        RECT 33.560 149.885 33.835 150.735 ;
        RECT 34.005 149.885 34.195 151.245 ;
        RECT 34.365 151.260 34.535 151.925 ;
        RECT 34.705 151.505 34.875 152.265 ;
        RECT 35.110 151.505 35.625 151.915 ;
        RECT 34.365 151.070 35.115 151.260 ;
        RECT 35.285 150.695 35.625 151.505 ;
        RECT 35.795 151.100 36.085 152.265 ;
        RECT 36.345 151.595 36.515 152.095 ;
        RECT 36.685 151.765 37.015 152.265 ;
        RECT 36.345 151.425 37.010 151.595 ;
        RECT 34.395 150.525 35.625 150.695 ;
        RECT 36.260 150.605 36.610 151.255 ;
        RECT 34.375 149.715 34.885 150.250 ;
        RECT 35.105 149.920 35.350 150.525 ;
        RECT 35.795 149.715 36.085 150.440 ;
        RECT 36.780 150.435 37.010 151.425 ;
        RECT 36.345 150.265 37.010 150.435 ;
        RECT 36.345 149.975 36.515 150.265 ;
        RECT 36.685 149.715 37.015 150.095 ;
        RECT 37.185 149.975 37.410 152.095 ;
        RECT 37.625 151.765 37.955 152.265 ;
        RECT 38.125 151.595 38.295 152.095 ;
        RECT 38.530 151.880 39.360 152.050 ;
        RECT 39.600 151.885 39.980 152.265 ;
        RECT 37.600 151.425 38.295 151.595 ;
        RECT 37.600 150.455 37.770 151.425 ;
        RECT 37.940 150.635 38.350 151.255 ;
        RECT 38.520 151.205 39.020 151.585 ;
        RECT 37.600 150.265 38.295 150.455 ;
        RECT 38.520 150.335 38.740 151.205 ;
        RECT 39.190 151.035 39.360 151.880 ;
        RECT 40.160 151.715 40.330 152.005 ;
        RECT 40.500 151.885 40.830 152.265 ;
        RECT 41.300 151.795 41.930 152.045 ;
        RECT 42.110 151.885 42.530 152.265 ;
        RECT 41.760 151.715 41.930 151.795 ;
        RECT 42.730 151.715 42.970 152.005 ;
        RECT 39.530 151.465 40.900 151.715 ;
        RECT 39.530 151.205 39.780 151.465 ;
        RECT 40.290 151.035 40.540 151.195 ;
        RECT 39.190 150.865 40.540 151.035 ;
        RECT 39.190 150.825 39.610 150.865 ;
        RECT 38.920 150.275 39.270 150.645 ;
        RECT 37.625 149.715 37.955 150.095 ;
        RECT 38.125 149.935 38.295 150.265 ;
        RECT 39.440 150.095 39.610 150.825 ;
        RECT 40.710 150.695 40.900 151.465 ;
        RECT 39.780 150.365 40.190 150.695 ;
        RECT 40.480 150.355 40.900 150.695 ;
        RECT 41.070 151.285 41.590 151.595 ;
        RECT 41.760 151.545 42.970 151.715 ;
        RECT 43.200 151.575 43.530 152.265 ;
        RECT 41.070 150.525 41.240 151.285 ;
        RECT 41.410 150.695 41.590 151.105 ;
        RECT 41.760 151.035 41.930 151.545 ;
        RECT 43.700 151.395 43.870 152.005 ;
        RECT 44.140 151.545 44.470 152.055 ;
        RECT 43.700 151.375 44.020 151.395 ;
        RECT 42.100 151.205 44.020 151.375 ;
        RECT 41.760 150.865 43.660 151.035 ;
        RECT 41.990 150.525 42.320 150.645 ;
        RECT 41.070 150.355 42.320 150.525 ;
        RECT 38.595 149.895 39.610 150.095 ;
        RECT 39.780 149.715 40.190 150.155 ;
        RECT 40.480 149.925 40.730 150.355 ;
        RECT 40.930 149.715 41.250 150.175 ;
        RECT 42.490 150.105 42.660 150.865 ;
        RECT 43.330 150.805 43.660 150.865 ;
        RECT 42.850 150.635 43.180 150.695 ;
        RECT 42.850 150.365 43.510 150.635 ;
        RECT 43.830 150.310 44.020 151.205 ;
        RECT 41.810 149.935 42.660 150.105 ;
        RECT 42.860 149.715 43.520 150.195 ;
        RECT 43.700 149.980 44.020 150.310 ;
        RECT 44.220 150.955 44.470 151.545 ;
        RECT 44.650 151.465 44.935 152.265 ;
        RECT 45.115 151.285 45.370 151.955 ;
        RECT 45.190 151.245 45.370 151.285 ;
        RECT 45.190 151.075 45.455 151.245 ;
        RECT 45.955 151.125 46.185 152.265 ;
        RECT 46.355 151.115 46.685 152.095 ;
        RECT 46.855 151.125 47.065 152.265 ;
        RECT 47.760 151.755 49.415 152.045 ;
        RECT 47.760 151.415 49.350 151.585 ;
        RECT 49.585 151.465 49.865 152.265 ;
        RECT 47.760 151.125 48.080 151.415 ;
        RECT 49.180 151.295 49.350 151.415 ;
        RECT 44.220 150.625 45.020 150.955 ;
        RECT 44.220 149.975 44.470 150.625 ;
        RECT 45.190 150.425 45.370 151.075 ;
        RECT 45.935 150.705 46.265 150.955 ;
        RECT 44.650 149.715 44.935 150.175 ;
        RECT 45.115 149.895 45.370 150.425 ;
        RECT 45.955 149.715 46.185 150.535 ;
        RECT 46.435 150.515 46.685 151.115 ;
        RECT 46.355 149.885 46.685 150.515 ;
        RECT 46.855 149.715 47.065 150.535 ;
        RECT 47.760 150.385 48.110 150.955 ;
        RECT 48.280 150.625 48.990 151.245 ;
        RECT 49.180 151.125 49.905 151.295 ;
        RECT 50.075 151.125 50.345 152.095 ;
        RECT 50.630 151.635 50.915 152.095 ;
        RECT 51.085 151.805 51.355 152.265 ;
        RECT 50.630 151.415 51.585 151.635 ;
        RECT 49.735 150.955 49.905 151.125 ;
        RECT 49.160 150.625 49.565 150.955 ;
        RECT 49.735 150.625 50.005 150.955 ;
        RECT 49.735 150.455 49.905 150.625 ;
        RECT 48.295 150.285 49.905 150.455 ;
        RECT 50.175 150.390 50.345 151.125 ;
        RECT 50.515 150.685 51.205 151.245 ;
        RECT 51.375 150.515 51.585 151.415 ;
        RECT 47.765 149.715 48.095 150.215 ;
        RECT 48.295 149.935 48.465 150.285 ;
        RECT 48.665 149.715 48.995 150.115 ;
        RECT 49.165 149.935 49.335 150.285 ;
        RECT 49.505 149.715 49.885 150.115 ;
        RECT 50.075 150.045 50.345 150.390 ;
        RECT 50.630 150.345 51.585 150.515 ;
        RECT 51.755 151.245 52.155 152.095 ;
        RECT 52.345 151.635 52.625 152.095 ;
        RECT 53.145 151.805 53.470 152.265 ;
        RECT 52.345 151.415 53.470 151.635 ;
        RECT 51.755 150.685 52.850 151.245 ;
        RECT 53.020 150.955 53.470 151.415 ;
        RECT 53.640 151.125 54.025 152.095 ;
        RECT 50.630 149.885 50.915 150.345 ;
        RECT 51.085 149.715 51.355 150.175 ;
        RECT 51.755 149.885 52.155 150.685 ;
        RECT 53.020 150.625 53.575 150.955 ;
        RECT 53.020 150.515 53.470 150.625 ;
        RECT 52.345 150.345 53.470 150.515 ;
        RECT 53.745 150.455 54.025 151.125 ;
        RECT 52.345 149.885 52.625 150.345 ;
        RECT 53.145 149.715 53.470 150.175 ;
        RECT 53.640 149.885 54.025 150.455 ;
        RECT 54.195 151.125 54.535 152.095 ;
        RECT 54.705 151.125 54.875 152.265 ;
        RECT 55.145 151.465 55.395 152.265 ;
        RECT 56.040 151.295 56.370 152.095 ;
        RECT 56.670 151.465 57.000 152.265 ;
        RECT 57.170 151.295 57.500 152.095 ;
        RECT 57.990 151.635 58.275 152.095 ;
        RECT 58.445 151.805 58.715 152.265 ;
        RECT 57.990 151.415 58.945 151.635 ;
        RECT 55.065 151.125 57.500 151.295 ;
        RECT 54.195 150.565 54.370 151.125 ;
        RECT 55.065 150.875 55.235 151.125 ;
        RECT 54.540 150.705 55.235 150.875 ;
        RECT 55.410 150.705 55.830 150.905 ;
        RECT 56.000 150.705 56.330 150.905 ;
        RECT 56.500 150.705 56.830 150.905 ;
        RECT 54.195 150.515 54.425 150.565 ;
        RECT 54.195 149.885 54.535 150.515 ;
        RECT 54.705 149.715 54.955 150.515 ;
        RECT 55.145 150.365 56.370 150.535 ;
        RECT 55.145 149.885 55.475 150.365 ;
        RECT 55.645 149.715 55.870 150.175 ;
        RECT 56.040 149.885 56.370 150.365 ;
        RECT 57.000 150.495 57.170 151.125 ;
        RECT 57.355 150.705 57.705 150.955 ;
        RECT 57.875 150.685 58.565 151.245 ;
        RECT 58.735 150.515 58.945 151.415 ;
        RECT 57.000 149.885 57.500 150.495 ;
        RECT 57.990 150.345 58.945 150.515 ;
        RECT 59.115 151.245 59.515 152.095 ;
        RECT 59.705 151.635 59.985 152.095 ;
        RECT 60.505 151.805 60.830 152.265 ;
        RECT 59.705 151.415 60.830 151.635 ;
        RECT 59.115 150.685 60.210 151.245 ;
        RECT 60.380 150.955 60.830 151.415 ;
        RECT 61.000 151.125 61.385 152.095 ;
        RECT 57.990 149.885 58.275 150.345 ;
        RECT 58.445 149.715 58.715 150.175 ;
        RECT 59.115 149.885 59.515 150.685 ;
        RECT 60.380 150.625 60.935 150.955 ;
        RECT 60.380 150.515 60.830 150.625 ;
        RECT 59.705 150.345 60.830 150.515 ;
        RECT 61.105 150.455 61.385 151.125 ;
        RECT 61.555 151.100 61.845 152.265 ;
        RECT 63.310 151.285 63.565 151.955 ;
        RECT 63.745 151.465 64.030 152.265 ;
        RECT 64.210 151.545 64.540 152.055 ;
        RECT 63.310 150.905 63.490 151.285 ;
        RECT 64.210 150.955 64.460 151.545 ;
        RECT 64.810 151.395 64.980 152.005 ;
        RECT 65.150 151.575 65.480 152.265 ;
        RECT 65.710 151.715 65.950 152.005 ;
        RECT 66.150 151.885 66.570 152.265 ;
        RECT 66.750 151.795 67.380 152.045 ;
        RECT 67.850 151.885 68.180 152.265 ;
        RECT 66.750 151.715 66.920 151.795 ;
        RECT 68.350 151.715 68.520 152.005 ;
        RECT 68.700 151.885 69.080 152.265 ;
        RECT 69.320 151.880 70.150 152.050 ;
        RECT 65.710 151.545 66.920 151.715 ;
        RECT 63.225 150.735 63.490 150.905 ;
        RECT 59.705 149.885 59.985 150.345 ;
        RECT 60.505 149.715 60.830 150.175 ;
        RECT 61.000 149.885 61.385 150.455 ;
        RECT 61.555 149.715 61.845 150.440 ;
        RECT 63.310 150.425 63.490 150.735 ;
        RECT 63.660 150.625 64.460 150.955 ;
        RECT 63.310 149.895 63.565 150.425 ;
        RECT 63.745 149.715 64.030 150.175 ;
        RECT 64.210 149.975 64.460 150.625 ;
        RECT 64.660 151.375 64.980 151.395 ;
        RECT 64.660 151.205 66.580 151.375 ;
        RECT 64.660 150.310 64.850 151.205 ;
        RECT 66.750 151.035 66.920 151.545 ;
        RECT 67.090 151.285 67.610 151.595 ;
        RECT 65.020 150.865 66.920 151.035 ;
        RECT 65.020 150.805 65.350 150.865 ;
        RECT 65.500 150.635 65.830 150.695 ;
        RECT 65.170 150.365 65.830 150.635 ;
        RECT 64.660 149.980 64.980 150.310 ;
        RECT 65.160 149.715 65.820 150.195 ;
        RECT 66.020 150.105 66.190 150.865 ;
        RECT 67.090 150.695 67.270 151.105 ;
        RECT 66.360 150.525 66.690 150.645 ;
        RECT 67.440 150.525 67.610 151.285 ;
        RECT 66.360 150.355 67.610 150.525 ;
        RECT 67.780 151.465 69.150 151.715 ;
        RECT 67.780 150.695 67.970 151.465 ;
        RECT 68.900 151.205 69.150 151.465 ;
        RECT 68.140 151.035 68.390 151.195 ;
        RECT 69.320 151.035 69.490 151.880 ;
        RECT 70.385 151.595 70.555 152.095 ;
        RECT 70.725 151.765 71.055 152.265 ;
        RECT 69.660 151.205 70.160 151.585 ;
        RECT 70.385 151.425 71.080 151.595 ;
        RECT 68.140 150.865 69.490 151.035 ;
        RECT 69.070 150.825 69.490 150.865 ;
        RECT 67.780 150.355 68.200 150.695 ;
        RECT 68.490 150.365 68.900 150.695 ;
        RECT 66.020 149.935 66.870 150.105 ;
        RECT 67.430 149.715 67.750 150.175 ;
        RECT 67.950 149.925 68.200 150.355 ;
        RECT 68.490 149.715 68.900 150.155 ;
        RECT 69.070 150.095 69.240 150.825 ;
        RECT 69.410 150.275 69.760 150.645 ;
        RECT 69.940 150.335 70.160 151.205 ;
        RECT 70.330 150.635 70.740 151.255 ;
        RECT 70.910 150.455 71.080 151.425 ;
        RECT 70.385 150.265 71.080 150.455 ;
        RECT 69.070 149.895 70.085 150.095 ;
        RECT 70.385 149.935 70.555 150.265 ;
        RECT 70.725 149.715 71.055 150.095 ;
        RECT 71.270 149.975 71.495 152.095 ;
        RECT 71.665 151.765 71.995 152.265 ;
        RECT 72.165 151.595 72.335 152.095 ;
        RECT 71.670 151.425 72.335 151.595 ;
        RECT 71.670 150.435 71.900 151.425 ;
        RECT 72.070 150.605 72.420 151.255 ;
        RECT 72.635 151.125 72.865 152.265 ;
        RECT 73.035 151.115 73.365 152.095 ;
        RECT 73.535 151.125 73.745 152.265 ;
        RECT 73.975 151.190 74.245 152.095 ;
        RECT 74.415 151.505 74.745 152.265 ;
        RECT 74.925 151.335 75.095 152.095 ;
        RECT 72.615 150.705 72.945 150.955 ;
        RECT 71.670 150.265 72.335 150.435 ;
        RECT 71.665 149.715 71.995 150.095 ;
        RECT 72.165 149.975 72.335 150.265 ;
        RECT 72.635 149.715 72.865 150.535 ;
        RECT 73.115 150.515 73.365 151.115 ;
        RECT 73.035 149.885 73.365 150.515 ;
        RECT 73.535 149.715 73.745 150.535 ;
        RECT 73.975 150.390 74.145 151.190 ;
        RECT 74.430 151.165 75.095 151.335 ;
        RECT 75.355 151.175 77.945 152.265 ;
        RECT 78.205 151.335 78.375 152.095 ;
        RECT 78.555 151.505 78.885 152.265 ;
        RECT 74.430 151.020 74.600 151.165 ;
        RECT 74.315 150.690 74.600 151.020 ;
        RECT 74.430 150.435 74.600 150.690 ;
        RECT 74.835 150.615 75.165 150.985 ;
        RECT 75.355 150.655 76.565 151.175 ;
        RECT 78.205 151.165 78.870 151.335 ;
        RECT 79.055 151.190 79.325 152.095 ;
        RECT 78.700 151.020 78.870 151.165 ;
        RECT 76.735 150.485 77.945 151.005 ;
        RECT 78.135 150.615 78.465 150.985 ;
        RECT 78.700 150.690 78.985 151.020 ;
        RECT 73.975 149.885 74.235 150.390 ;
        RECT 74.430 150.265 75.095 150.435 ;
        RECT 74.415 149.715 74.745 150.095 ;
        RECT 74.925 149.885 75.095 150.265 ;
        RECT 75.355 149.715 77.945 150.485 ;
        RECT 78.700 150.435 78.870 150.690 ;
        RECT 78.205 150.265 78.870 150.435 ;
        RECT 79.155 150.390 79.325 151.190 ;
        RECT 78.205 149.885 78.375 150.265 ;
        RECT 78.555 149.715 78.885 150.095 ;
        RECT 79.065 149.885 79.325 150.390 ;
        RECT 79.500 151.125 79.835 152.095 ;
        RECT 80.005 151.125 80.175 152.265 ;
        RECT 80.345 151.925 82.375 152.095 ;
        RECT 79.500 150.455 79.670 151.125 ;
        RECT 80.345 150.955 80.515 151.925 ;
        RECT 79.840 150.625 80.095 150.955 ;
        RECT 80.320 150.625 80.515 150.955 ;
        RECT 80.685 151.585 81.810 151.755 ;
        RECT 79.925 150.455 80.095 150.625 ;
        RECT 80.685 150.455 80.855 151.585 ;
        RECT 79.500 149.885 79.755 150.455 ;
        RECT 79.925 150.285 80.855 150.455 ;
        RECT 81.025 151.245 82.035 151.415 ;
        RECT 81.025 150.445 81.195 151.245 ;
        RECT 80.680 150.250 80.855 150.285 ;
        RECT 79.925 149.715 80.255 150.115 ;
        RECT 80.680 149.885 81.210 150.250 ;
        RECT 81.400 150.225 81.675 151.045 ;
        RECT 81.395 150.055 81.675 150.225 ;
        RECT 81.400 149.885 81.675 150.055 ;
        RECT 81.845 149.885 82.035 151.245 ;
        RECT 82.205 151.260 82.375 151.925 ;
        RECT 82.545 151.505 82.715 152.265 ;
        RECT 82.950 151.505 83.465 151.915 ;
        RECT 82.205 151.070 82.955 151.260 ;
        RECT 83.125 150.695 83.465 151.505 ;
        RECT 83.695 151.125 83.905 152.265 ;
        RECT 82.235 150.525 83.465 150.695 ;
        RECT 84.075 151.115 84.405 152.095 ;
        RECT 84.575 151.125 84.805 152.265 ;
        RECT 85.105 151.335 85.275 152.095 ;
        RECT 85.455 151.505 85.785 152.265 ;
        RECT 85.105 151.165 85.770 151.335 ;
        RECT 85.955 151.190 86.225 152.095 ;
        RECT 82.215 149.715 82.725 150.250 ;
        RECT 82.945 149.920 83.190 150.525 ;
        RECT 83.695 149.715 83.905 150.535 ;
        RECT 84.075 150.515 84.325 151.115 ;
        RECT 85.600 151.020 85.770 151.165 ;
        RECT 84.495 150.705 84.825 150.955 ;
        RECT 85.035 150.615 85.365 150.985 ;
        RECT 85.600 150.690 85.885 151.020 ;
        RECT 84.075 149.885 84.405 150.515 ;
        RECT 84.575 149.715 84.805 150.535 ;
        RECT 85.600 150.435 85.770 150.690 ;
        RECT 85.105 150.265 85.770 150.435 ;
        RECT 86.055 150.390 86.225 151.190 ;
        RECT 87.315 151.100 87.605 152.265 ;
        RECT 88.895 151.595 89.175 152.265 ;
        RECT 89.345 151.375 89.645 151.925 ;
        RECT 89.845 151.545 90.175 152.265 ;
        RECT 90.365 151.545 90.825 152.095 ;
        RECT 88.710 150.955 88.975 151.315 ;
        RECT 89.345 151.205 90.285 151.375 ;
        RECT 90.115 150.955 90.285 151.205 ;
        RECT 88.710 150.705 89.385 150.955 ;
        RECT 89.605 150.705 89.945 150.955 ;
        RECT 90.115 150.625 90.405 150.955 ;
        RECT 90.115 150.535 90.285 150.625 ;
        RECT 85.105 149.885 85.275 150.265 ;
        RECT 85.455 149.715 85.785 150.095 ;
        RECT 85.965 149.885 86.225 150.390 ;
        RECT 87.315 149.715 87.605 150.440 ;
        RECT 88.895 150.345 90.285 150.535 ;
        RECT 88.895 149.985 89.225 150.345 ;
        RECT 90.575 150.175 90.825 151.545 ;
        RECT 90.995 151.505 91.510 151.915 ;
        RECT 91.745 151.505 91.915 152.265 ;
        RECT 92.085 151.925 94.115 152.095 ;
        RECT 90.995 150.695 91.335 151.505 ;
        RECT 92.085 151.260 92.255 151.925 ;
        RECT 92.650 151.585 93.775 151.755 ;
        RECT 91.505 151.070 92.255 151.260 ;
        RECT 92.425 151.245 93.435 151.415 ;
        RECT 90.995 150.525 92.225 150.695 ;
        RECT 89.845 149.715 90.095 150.175 ;
        RECT 90.265 149.885 90.825 150.175 ;
        RECT 91.270 149.920 91.515 150.525 ;
        RECT 91.735 149.715 92.245 150.250 ;
        RECT 92.425 149.885 92.615 151.245 ;
        RECT 92.785 150.565 93.060 151.045 ;
        RECT 92.785 150.395 93.065 150.565 ;
        RECT 93.265 150.445 93.435 151.245 ;
        RECT 93.605 150.455 93.775 151.585 ;
        RECT 93.945 150.955 94.115 151.925 ;
        RECT 94.285 151.125 94.455 152.265 ;
        RECT 94.625 151.125 94.960 152.095 ;
        RECT 93.945 150.625 94.140 150.955 ;
        RECT 94.365 150.625 94.620 150.955 ;
        RECT 94.365 150.455 94.535 150.625 ;
        RECT 94.790 150.455 94.960 151.125 ;
        RECT 92.785 149.885 93.060 150.395 ;
        RECT 93.605 150.285 94.535 150.455 ;
        RECT 93.605 150.250 93.780 150.285 ;
        RECT 93.250 149.885 93.780 150.250 ;
        RECT 94.205 149.715 94.535 150.115 ;
        RECT 94.705 149.885 94.960 150.455 ;
        RECT 95.135 151.125 95.405 152.095 ;
        RECT 95.615 151.465 95.895 152.265 ;
        RECT 96.065 151.755 97.720 152.045 ;
        RECT 96.130 151.415 97.720 151.585 ;
        RECT 96.130 151.295 96.300 151.415 ;
        RECT 95.575 151.125 96.300 151.295 ;
        RECT 95.135 150.390 95.305 151.125 ;
        RECT 95.575 150.955 95.745 151.125 ;
        RECT 96.490 151.075 97.205 151.245 ;
        RECT 97.400 151.125 97.720 151.415 ;
        RECT 97.895 151.545 98.355 152.095 ;
        RECT 98.545 151.545 98.875 152.265 ;
        RECT 95.475 150.625 95.745 150.955 ;
        RECT 95.915 150.625 96.320 150.955 ;
        RECT 96.490 150.625 97.200 151.075 ;
        RECT 95.575 150.455 95.745 150.625 ;
        RECT 95.135 150.045 95.405 150.390 ;
        RECT 95.575 150.285 97.185 150.455 ;
        RECT 97.370 150.385 97.720 150.955 ;
        RECT 95.595 149.715 95.975 150.115 ;
        RECT 96.145 149.935 96.315 150.285 ;
        RECT 96.485 149.715 96.815 150.115 ;
        RECT 97.015 149.935 97.185 150.285 ;
        RECT 97.385 149.715 97.715 150.215 ;
        RECT 97.895 150.175 98.145 151.545 ;
        RECT 99.075 151.375 99.375 151.925 ;
        RECT 99.545 151.595 99.825 152.265 ;
        RECT 98.435 151.205 99.375 151.375 ;
        RECT 98.435 150.955 98.605 151.205 ;
        RECT 99.745 150.955 100.010 151.315 ;
        RECT 100.235 151.125 100.465 152.265 ;
        RECT 100.635 151.115 100.965 152.095 ;
        RECT 101.135 151.125 101.345 152.265 ;
        RECT 101.575 151.505 102.090 151.915 ;
        RECT 102.325 151.505 102.495 152.265 ;
        RECT 102.665 151.925 104.695 152.095 ;
        RECT 98.315 150.625 98.605 150.955 ;
        RECT 98.775 150.705 99.115 150.955 ;
        RECT 99.335 150.705 100.010 150.955 ;
        RECT 100.215 150.705 100.545 150.955 ;
        RECT 98.435 150.535 98.605 150.625 ;
        RECT 98.435 150.345 99.825 150.535 ;
        RECT 97.895 149.885 98.455 150.175 ;
        RECT 98.625 149.715 98.875 150.175 ;
        RECT 99.495 149.985 99.825 150.345 ;
        RECT 100.235 149.715 100.465 150.535 ;
        RECT 100.715 150.515 100.965 151.115 ;
        RECT 101.575 150.695 101.915 151.505 ;
        RECT 102.665 151.260 102.835 151.925 ;
        RECT 103.230 151.585 104.355 151.755 ;
        RECT 102.085 151.070 102.835 151.260 ;
        RECT 103.005 151.245 104.015 151.415 ;
        RECT 100.635 149.885 100.965 150.515 ;
        RECT 101.135 149.715 101.345 150.535 ;
        RECT 101.575 150.525 102.805 150.695 ;
        RECT 101.850 149.920 102.095 150.525 ;
        RECT 102.315 149.715 102.825 150.250 ;
        RECT 103.005 149.885 103.195 151.245 ;
        RECT 103.365 150.905 103.640 151.045 ;
        RECT 103.365 150.735 103.645 150.905 ;
        RECT 103.365 149.885 103.640 150.735 ;
        RECT 103.845 150.445 104.015 151.245 ;
        RECT 104.185 150.455 104.355 151.585 ;
        RECT 104.525 150.955 104.695 151.925 ;
        RECT 104.865 151.125 105.035 152.265 ;
        RECT 105.205 151.125 105.540 152.095 ;
        RECT 106.725 151.335 106.895 152.095 ;
        RECT 107.075 151.505 107.405 152.265 ;
        RECT 106.725 151.165 107.390 151.335 ;
        RECT 107.575 151.190 107.845 152.095 ;
        RECT 104.525 150.625 104.720 150.955 ;
        RECT 104.945 150.625 105.200 150.955 ;
        RECT 104.945 150.455 105.115 150.625 ;
        RECT 105.370 150.455 105.540 151.125 ;
        RECT 107.220 151.020 107.390 151.165 ;
        RECT 106.655 150.615 106.985 150.985 ;
        RECT 107.220 150.690 107.505 151.020 ;
        RECT 104.185 150.285 105.115 150.455 ;
        RECT 104.185 150.250 104.360 150.285 ;
        RECT 103.830 149.885 104.360 150.250 ;
        RECT 104.785 149.715 105.115 150.115 ;
        RECT 105.285 149.885 105.540 150.455 ;
        RECT 107.220 150.435 107.390 150.690 ;
        RECT 106.725 150.265 107.390 150.435 ;
        RECT 107.675 150.390 107.845 151.190 ;
        RECT 108.565 151.335 108.735 152.095 ;
        RECT 108.915 151.505 109.245 152.265 ;
        RECT 108.565 151.165 109.230 151.335 ;
        RECT 109.415 151.190 109.685 152.095 ;
        RECT 109.060 151.020 109.230 151.165 ;
        RECT 108.495 150.615 108.825 150.985 ;
        RECT 109.060 150.690 109.345 151.020 ;
        RECT 109.060 150.435 109.230 150.690 ;
        RECT 106.725 149.885 106.895 150.265 ;
        RECT 107.075 149.715 107.405 150.095 ;
        RECT 107.585 149.885 107.845 150.390 ;
        RECT 108.565 150.265 109.230 150.435 ;
        RECT 109.515 150.390 109.685 151.190 ;
        RECT 109.945 151.335 110.115 152.095 ;
        RECT 110.295 151.505 110.625 152.265 ;
        RECT 109.945 151.165 110.610 151.335 ;
        RECT 110.795 151.190 111.065 152.095 ;
        RECT 110.440 151.020 110.610 151.165 ;
        RECT 109.875 150.615 110.205 150.985 ;
        RECT 110.440 150.690 110.725 151.020 ;
        RECT 110.440 150.435 110.610 150.690 ;
        RECT 108.565 149.885 108.735 150.265 ;
        RECT 108.915 149.715 109.245 150.095 ;
        RECT 109.425 149.885 109.685 150.390 ;
        RECT 109.945 150.265 110.610 150.435 ;
        RECT 110.895 150.390 111.065 151.190 ;
        RECT 112.155 151.175 113.365 152.265 ;
        RECT 112.155 150.635 112.675 151.175 ;
        RECT 112.845 150.465 113.365 151.005 ;
        RECT 109.945 149.885 110.115 150.265 ;
        RECT 110.295 149.715 110.625 150.095 ;
        RECT 110.805 149.885 111.065 150.390 ;
        RECT 112.155 149.715 113.365 150.465 ;
        RECT 26.970 149.545 113.450 149.715 ;
        RECT 27.055 148.795 28.265 149.545 ;
        RECT 28.810 148.835 29.065 149.365 ;
        RECT 29.245 149.085 29.530 149.545 ;
        RECT 27.055 148.255 27.575 148.795 ;
        RECT 27.745 148.085 28.265 148.625 ;
        RECT 27.055 146.995 28.265 148.085 ;
        RECT 28.810 147.975 28.990 148.835 ;
        RECT 29.710 148.635 29.960 149.285 ;
        RECT 29.160 148.305 29.960 148.635 ;
        RECT 28.810 147.505 29.065 147.975 ;
        RECT 28.725 147.335 29.065 147.505 ;
        RECT 28.810 147.305 29.065 147.335 ;
        RECT 29.245 146.995 29.530 147.795 ;
        RECT 29.710 147.715 29.960 148.305 ;
        RECT 30.160 148.950 30.480 149.280 ;
        RECT 30.660 149.065 31.320 149.545 ;
        RECT 31.520 149.155 32.370 149.325 ;
        RECT 30.160 148.055 30.350 148.950 ;
        RECT 30.670 148.625 31.330 148.895 ;
        RECT 31.000 148.565 31.330 148.625 ;
        RECT 30.520 148.395 30.850 148.455 ;
        RECT 31.520 148.395 31.690 149.155 ;
        RECT 32.930 149.085 33.250 149.545 ;
        RECT 33.450 148.905 33.700 149.335 ;
        RECT 33.990 149.105 34.400 149.545 ;
        RECT 34.570 149.165 35.585 149.365 ;
        RECT 31.860 148.735 33.110 148.905 ;
        RECT 31.860 148.615 32.190 148.735 ;
        RECT 30.520 148.225 32.420 148.395 ;
        RECT 30.160 147.885 32.080 148.055 ;
        RECT 30.160 147.865 30.480 147.885 ;
        RECT 29.710 147.205 30.040 147.715 ;
        RECT 30.310 147.255 30.480 147.865 ;
        RECT 32.250 147.715 32.420 148.225 ;
        RECT 32.590 148.155 32.770 148.565 ;
        RECT 32.940 147.975 33.110 148.735 ;
        RECT 30.650 146.995 30.980 147.685 ;
        RECT 31.210 147.545 32.420 147.715 ;
        RECT 32.590 147.665 33.110 147.975 ;
        RECT 33.280 148.565 33.700 148.905 ;
        RECT 33.990 148.565 34.400 148.895 ;
        RECT 33.280 147.795 33.470 148.565 ;
        RECT 34.570 148.435 34.740 149.165 ;
        RECT 35.885 148.995 36.055 149.325 ;
        RECT 36.225 149.165 36.555 149.545 ;
        RECT 34.910 148.615 35.260 148.985 ;
        RECT 34.570 148.395 34.990 148.435 ;
        RECT 33.640 148.225 34.990 148.395 ;
        RECT 33.640 148.065 33.890 148.225 ;
        RECT 34.400 147.795 34.650 148.055 ;
        RECT 33.280 147.545 34.650 147.795 ;
        RECT 31.210 147.255 31.450 147.545 ;
        RECT 32.250 147.465 32.420 147.545 ;
        RECT 31.650 146.995 32.070 147.375 ;
        RECT 32.250 147.215 32.880 147.465 ;
        RECT 33.350 146.995 33.680 147.375 ;
        RECT 33.850 147.255 34.020 147.545 ;
        RECT 34.820 147.380 34.990 148.225 ;
        RECT 35.440 148.055 35.660 148.925 ;
        RECT 35.885 148.805 36.580 148.995 ;
        RECT 35.160 147.675 35.660 148.055 ;
        RECT 35.830 148.005 36.240 148.625 ;
        RECT 36.410 147.835 36.580 148.805 ;
        RECT 35.885 147.665 36.580 147.835 ;
        RECT 34.200 146.995 34.580 147.375 ;
        RECT 34.820 147.210 35.650 147.380 ;
        RECT 35.885 147.165 36.055 147.665 ;
        RECT 36.225 146.995 36.555 147.495 ;
        RECT 36.770 147.165 36.995 149.285 ;
        RECT 37.165 149.165 37.495 149.545 ;
        RECT 37.665 148.995 37.835 149.285 ;
        RECT 38.185 149.065 38.485 149.545 ;
        RECT 37.170 148.825 37.835 148.995 ;
        RECT 38.655 148.895 38.915 149.350 ;
        RECT 39.085 149.065 39.345 149.545 ;
        RECT 39.525 148.895 39.785 149.350 ;
        RECT 39.955 149.065 40.205 149.545 ;
        RECT 40.385 148.895 40.645 149.350 ;
        RECT 40.815 149.065 41.065 149.545 ;
        RECT 41.245 148.895 41.505 149.350 ;
        RECT 41.675 149.065 41.920 149.545 ;
        RECT 42.090 148.895 42.365 149.350 ;
        RECT 42.535 149.065 42.780 149.545 ;
        RECT 42.950 148.895 43.210 149.350 ;
        RECT 43.380 149.065 43.640 149.545 ;
        RECT 43.810 148.895 44.070 149.350 ;
        RECT 44.240 149.065 44.500 149.545 ;
        RECT 44.670 148.895 44.930 149.350 ;
        RECT 45.100 148.985 45.360 149.545 ;
        RECT 37.170 147.835 37.400 148.825 ;
        RECT 38.185 148.725 44.930 148.895 ;
        RECT 37.570 148.005 37.920 148.655 ;
        RECT 38.185 148.135 39.350 148.725 ;
        RECT 45.530 148.555 45.780 149.365 ;
        RECT 45.960 149.020 46.220 149.545 ;
        RECT 46.390 148.555 46.640 149.365 ;
        RECT 46.820 149.035 47.125 149.545 ;
        RECT 47.385 148.995 47.555 149.375 ;
        RECT 47.735 149.165 48.065 149.545 ;
        RECT 39.520 148.305 46.640 148.555 ;
        RECT 46.810 148.305 47.125 148.865 ;
        RECT 47.385 148.825 48.050 148.995 ;
        RECT 48.245 148.870 48.505 149.375 ;
        RECT 38.185 147.910 44.930 148.135 ;
        RECT 37.170 147.665 37.835 147.835 ;
        RECT 37.165 146.995 37.495 147.495 ;
        RECT 37.665 147.165 37.835 147.665 ;
        RECT 38.185 146.995 38.455 147.740 ;
        RECT 38.625 147.170 38.915 147.910 ;
        RECT 39.525 147.895 44.930 147.910 ;
        RECT 39.085 147.000 39.340 147.725 ;
        RECT 39.525 147.170 39.785 147.895 ;
        RECT 39.955 147.000 40.200 147.725 ;
        RECT 40.385 147.170 40.645 147.895 ;
        RECT 40.815 147.000 41.060 147.725 ;
        RECT 41.245 147.170 41.505 147.895 ;
        RECT 41.675 147.000 41.920 147.725 ;
        RECT 42.090 147.170 42.350 147.895 ;
        RECT 42.520 147.000 42.780 147.725 ;
        RECT 42.950 147.170 43.210 147.895 ;
        RECT 43.380 147.000 43.640 147.725 ;
        RECT 43.810 147.170 44.070 147.895 ;
        RECT 44.240 147.000 44.500 147.725 ;
        RECT 44.670 147.170 44.930 147.895 ;
        RECT 45.100 147.000 45.360 147.795 ;
        RECT 45.530 147.170 45.780 148.305 ;
        RECT 39.085 146.995 45.360 147.000 ;
        RECT 45.960 146.995 46.220 147.805 ;
        RECT 46.395 147.165 46.640 148.305 ;
        RECT 47.315 148.275 47.645 148.645 ;
        RECT 47.880 148.570 48.050 148.825 ;
        RECT 47.880 148.240 48.165 148.570 ;
        RECT 47.880 148.095 48.050 148.240 ;
        RECT 47.385 147.925 48.050 148.095 ;
        RECT 48.335 148.070 48.505 148.870 ;
        RECT 48.675 148.820 48.965 149.545 ;
        RECT 49.605 149.045 49.935 149.545 ;
        RECT 50.135 148.975 50.305 149.325 ;
        RECT 50.505 149.145 50.835 149.545 ;
        RECT 51.005 148.975 51.175 149.325 ;
        RECT 51.345 149.145 51.725 149.545 ;
        RECT 49.600 148.305 49.950 148.875 ;
        RECT 50.135 148.805 51.745 148.975 ;
        RECT 51.915 148.870 52.185 149.215 ;
        RECT 51.575 148.635 51.745 148.805 ;
        RECT 46.820 146.995 47.115 147.805 ;
        RECT 47.385 147.165 47.555 147.925 ;
        RECT 47.735 146.995 48.065 147.755 ;
        RECT 48.235 147.165 48.505 148.070 ;
        RECT 48.675 146.995 48.965 148.160 ;
        RECT 49.600 147.845 49.920 148.135 ;
        RECT 50.120 148.015 50.830 148.635 ;
        RECT 51.000 148.305 51.405 148.635 ;
        RECT 51.575 148.305 51.845 148.635 ;
        RECT 51.575 148.135 51.745 148.305 ;
        RECT 52.015 148.135 52.185 148.870 ;
        RECT 51.020 147.965 51.745 148.135 ;
        RECT 51.020 147.845 51.190 147.965 ;
        RECT 49.600 147.675 51.190 147.845 ;
        RECT 49.600 147.215 51.255 147.505 ;
        RECT 51.425 146.995 51.705 147.795 ;
        RECT 51.915 147.165 52.185 148.135 ;
        RECT 52.355 148.745 52.695 149.375 ;
        RECT 52.865 148.745 53.115 149.545 ;
        RECT 53.305 148.895 53.635 149.375 ;
        RECT 53.805 149.085 54.030 149.545 ;
        RECT 54.200 148.895 54.530 149.375 ;
        RECT 52.355 148.695 52.585 148.745 ;
        RECT 53.305 148.725 54.530 148.895 ;
        RECT 55.160 148.765 55.660 149.375 ;
        RECT 52.355 148.135 52.530 148.695 ;
        RECT 52.700 148.385 53.395 148.555 ;
        RECT 53.225 148.135 53.395 148.385 ;
        RECT 53.570 148.355 53.990 148.555 ;
        RECT 54.160 148.355 54.490 148.555 ;
        RECT 54.660 148.355 54.990 148.555 ;
        RECT 55.160 148.135 55.330 148.765 ;
        RECT 56.035 148.745 56.375 149.375 ;
        RECT 56.545 148.745 56.795 149.545 ;
        RECT 56.985 148.895 57.315 149.375 ;
        RECT 57.485 149.085 57.710 149.545 ;
        RECT 57.880 148.895 58.210 149.375 ;
        RECT 55.515 148.305 55.865 148.555 ;
        RECT 56.035 148.135 56.210 148.745 ;
        RECT 56.985 148.725 58.210 148.895 ;
        RECT 58.840 148.765 59.340 149.375 ;
        RECT 56.380 148.385 57.075 148.555 ;
        RECT 56.905 148.135 57.075 148.385 ;
        RECT 57.250 148.355 57.670 148.555 ;
        RECT 57.840 148.355 58.170 148.555 ;
        RECT 58.340 148.355 58.670 148.555 ;
        RECT 58.840 148.135 59.010 148.765 ;
        RECT 60.175 148.745 60.515 149.375 ;
        RECT 60.685 148.745 60.935 149.545 ;
        RECT 61.125 148.895 61.455 149.375 ;
        RECT 61.625 149.085 61.850 149.545 ;
        RECT 62.020 148.895 62.350 149.375 ;
        RECT 59.195 148.305 59.545 148.555 ;
        RECT 60.175 148.135 60.350 148.745 ;
        RECT 61.125 148.725 62.350 148.895 ;
        RECT 62.980 148.765 63.480 149.375 ;
        RECT 60.520 148.385 61.215 148.555 ;
        RECT 61.045 148.135 61.215 148.385 ;
        RECT 61.390 148.355 61.810 148.555 ;
        RECT 61.980 148.355 62.310 148.555 ;
        RECT 62.480 148.355 62.810 148.555 ;
        RECT 62.980 148.135 63.150 148.765 ;
        RECT 64.130 148.735 64.375 149.340 ;
        RECT 64.595 149.010 65.105 149.545 ;
        RECT 63.855 148.565 65.085 148.735 ;
        RECT 63.335 148.305 63.685 148.555 ;
        RECT 52.355 147.165 52.695 148.135 ;
        RECT 52.865 146.995 53.035 148.135 ;
        RECT 53.225 147.965 55.660 148.135 ;
        RECT 53.305 146.995 53.555 147.795 ;
        RECT 54.200 147.165 54.530 147.965 ;
        RECT 54.830 146.995 55.160 147.795 ;
        RECT 55.330 147.165 55.660 147.965 ;
        RECT 56.035 147.165 56.375 148.135 ;
        RECT 56.545 146.995 56.715 148.135 ;
        RECT 56.905 147.965 59.340 148.135 ;
        RECT 56.985 146.995 57.235 147.795 ;
        RECT 57.880 147.165 58.210 147.965 ;
        RECT 58.510 146.995 58.840 147.795 ;
        RECT 59.010 147.165 59.340 147.965 ;
        RECT 60.175 147.165 60.515 148.135 ;
        RECT 60.685 146.995 60.855 148.135 ;
        RECT 61.045 147.965 63.480 148.135 ;
        RECT 61.125 146.995 61.375 147.795 ;
        RECT 62.020 147.165 62.350 147.965 ;
        RECT 62.650 146.995 62.980 147.795 ;
        RECT 63.150 147.165 63.480 147.965 ;
        RECT 63.855 147.755 64.195 148.565 ;
        RECT 64.365 148.000 65.115 148.190 ;
        RECT 63.855 147.345 64.370 147.755 ;
        RECT 64.605 146.995 64.775 147.755 ;
        RECT 64.945 147.335 65.115 148.000 ;
        RECT 65.285 148.015 65.475 149.375 ;
        RECT 65.645 149.205 65.920 149.375 ;
        RECT 65.645 149.035 65.925 149.205 ;
        RECT 65.645 148.215 65.920 149.035 ;
        RECT 66.110 149.010 66.640 149.375 ;
        RECT 67.065 149.145 67.395 149.545 ;
        RECT 66.465 148.975 66.640 149.010 ;
        RECT 66.125 148.015 66.295 148.815 ;
        RECT 65.285 147.845 66.295 148.015 ;
        RECT 66.465 148.805 67.395 148.975 ;
        RECT 67.565 148.805 67.820 149.375 ;
        RECT 68.000 149.145 68.335 149.545 ;
        RECT 68.505 148.975 68.710 149.375 ;
        RECT 68.920 149.065 69.195 149.545 ;
        RECT 69.405 149.045 69.665 149.375 ;
        RECT 66.465 147.675 66.635 148.805 ;
        RECT 67.225 148.635 67.395 148.805 ;
        RECT 65.510 147.505 66.635 147.675 ;
        RECT 66.805 148.305 67.000 148.635 ;
        RECT 67.225 148.305 67.480 148.635 ;
        RECT 66.805 147.335 66.975 148.305 ;
        RECT 67.650 148.135 67.820 148.805 ;
        RECT 64.945 147.165 66.975 147.335 ;
        RECT 67.145 146.995 67.315 148.135 ;
        RECT 67.485 147.165 67.820 148.135 ;
        RECT 68.025 148.805 68.710 148.975 ;
        RECT 68.025 147.775 68.365 148.805 ;
        RECT 68.535 148.135 68.785 148.635 ;
        RECT 68.965 148.305 69.325 148.885 ;
        RECT 69.495 148.135 69.665 149.045 ;
        RECT 68.535 147.965 69.665 148.135 ;
        RECT 68.025 147.600 68.690 147.775 ;
        RECT 68.000 146.995 68.335 147.420 ;
        RECT 68.505 147.195 68.690 147.600 ;
        RECT 68.895 146.995 69.225 147.775 ;
        RECT 69.395 147.195 69.665 147.965 ;
        RECT 69.835 149.045 70.095 149.375 ;
        RECT 70.305 149.065 70.580 149.545 ;
        RECT 69.835 148.135 70.005 149.045 ;
        RECT 70.790 148.975 70.995 149.375 ;
        RECT 71.165 149.145 71.500 149.545 ;
        RECT 70.175 148.305 70.535 148.885 ;
        RECT 70.790 148.805 71.475 148.975 ;
        RECT 70.715 148.135 70.965 148.635 ;
        RECT 69.835 147.965 70.965 148.135 ;
        RECT 69.835 147.195 70.105 147.965 ;
        RECT 71.135 147.775 71.475 148.805 ;
        RECT 70.275 146.995 70.605 147.775 ;
        RECT 70.810 147.600 71.475 147.775 ;
        RECT 71.675 148.870 71.945 149.215 ;
        RECT 72.135 149.145 72.515 149.545 ;
        RECT 72.685 148.975 72.855 149.325 ;
        RECT 73.025 149.145 73.355 149.545 ;
        RECT 73.555 148.975 73.725 149.325 ;
        RECT 73.925 149.045 74.255 149.545 ;
        RECT 71.675 148.135 71.845 148.870 ;
        RECT 72.115 148.805 73.725 148.975 ;
        RECT 72.115 148.635 72.285 148.805 ;
        RECT 72.015 148.305 72.285 148.635 ;
        RECT 72.455 148.305 72.860 148.635 ;
        RECT 72.115 148.135 72.285 148.305 ;
        RECT 70.810 147.195 70.995 147.600 ;
        RECT 71.165 146.995 71.500 147.420 ;
        RECT 71.675 147.165 71.945 148.135 ;
        RECT 72.115 147.965 72.840 148.135 ;
        RECT 73.030 148.015 73.740 148.635 ;
        RECT 73.910 148.305 74.260 148.875 ;
        RECT 74.435 148.820 74.725 149.545 ;
        RECT 75.355 148.745 75.695 149.375 ;
        RECT 75.865 148.745 76.115 149.545 ;
        RECT 76.305 148.895 76.635 149.375 ;
        RECT 76.805 149.085 77.030 149.545 ;
        RECT 77.200 148.895 77.530 149.375 ;
        RECT 75.355 148.695 75.585 148.745 ;
        RECT 76.305 148.725 77.530 148.895 ;
        RECT 78.160 148.765 78.660 149.375 ;
        RECT 79.410 148.835 79.665 149.365 ;
        RECT 79.845 149.085 80.130 149.545 ;
        RECT 72.670 147.845 72.840 147.965 ;
        RECT 73.940 147.845 74.260 148.135 ;
        RECT 72.155 146.995 72.435 147.795 ;
        RECT 72.670 147.675 74.260 147.845 ;
        RECT 72.605 147.215 74.260 147.505 ;
        RECT 74.435 146.995 74.725 148.160 ;
        RECT 75.355 148.135 75.530 148.695 ;
        RECT 75.700 148.385 76.395 148.555 ;
        RECT 76.225 148.135 76.395 148.385 ;
        RECT 76.570 148.355 76.990 148.555 ;
        RECT 77.160 148.355 77.490 148.555 ;
        RECT 77.660 148.355 77.990 148.555 ;
        RECT 78.160 148.135 78.330 148.765 ;
        RECT 78.515 148.305 78.865 148.555 ;
        RECT 75.355 147.165 75.695 148.135 ;
        RECT 75.865 146.995 76.035 148.135 ;
        RECT 76.225 147.965 78.660 148.135 ;
        RECT 76.305 146.995 76.555 147.795 ;
        RECT 77.200 147.165 77.530 147.965 ;
        RECT 77.830 146.995 78.160 147.795 ;
        RECT 78.330 147.165 78.660 147.965 ;
        RECT 79.410 147.975 79.590 148.835 ;
        RECT 80.310 148.635 80.560 149.285 ;
        RECT 79.760 148.305 80.560 148.635 ;
        RECT 79.410 147.505 79.665 147.975 ;
        RECT 79.325 147.335 79.665 147.505 ;
        RECT 79.410 147.305 79.665 147.335 ;
        RECT 79.845 146.995 80.130 147.795 ;
        RECT 80.310 147.715 80.560 148.305 ;
        RECT 80.760 148.950 81.080 149.280 ;
        RECT 81.260 149.065 81.920 149.545 ;
        RECT 82.120 149.155 82.970 149.325 ;
        RECT 80.760 148.055 80.950 148.950 ;
        RECT 81.270 148.625 81.930 148.895 ;
        RECT 81.600 148.565 81.930 148.625 ;
        RECT 81.120 148.395 81.450 148.455 ;
        RECT 82.120 148.395 82.290 149.155 ;
        RECT 83.530 149.085 83.850 149.545 ;
        RECT 84.050 148.905 84.300 149.335 ;
        RECT 84.590 149.105 85.000 149.545 ;
        RECT 85.170 149.165 86.185 149.365 ;
        RECT 82.460 148.735 83.710 148.905 ;
        RECT 82.460 148.615 82.790 148.735 ;
        RECT 81.120 148.225 83.020 148.395 ;
        RECT 80.760 147.885 82.680 148.055 ;
        RECT 80.760 147.865 81.080 147.885 ;
        RECT 80.310 147.205 80.640 147.715 ;
        RECT 80.910 147.255 81.080 147.865 ;
        RECT 82.850 147.715 83.020 148.225 ;
        RECT 83.190 148.155 83.370 148.565 ;
        RECT 83.540 147.975 83.710 148.735 ;
        RECT 81.250 146.995 81.580 147.685 ;
        RECT 81.810 147.545 83.020 147.715 ;
        RECT 83.190 147.665 83.710 147.975 ;
        RECT 83.880 148.565 84.300 148.905 ;
        RECT 84.590 148.565 85.000 148.895 ;
        RECT 83.880 147.795 84.070 148.565 ;
        RECT 85.170 148.435 85.340 149.165 ;
        RECT 86.485 148.995 86.655 149.325 ;
        RECT 86.825 149.165 87.155 149.545 ;
        RECT 85.510 148.615 85.860 148.985 ;
        RECT 85.170 148.395 85.590 148.435 ;
        RECT 84.240 148.225 85.590 148.395 ;
        RECT 84.240 148.065 84.490 148.225 ;
        RECT 85.000 147.795 85.250 148.055 ;
        RECT 83.880 147.545 85.250 147.795 ;
        RECT 81.810 147.255 82.050 147.545 ;
        RECT 82.850 147.465 83.020 147.545 ;
        RECT 82.250 146.995 82.670 147.375 ;
        RECT 82.850 147.215 83.480 147.465 ;
        RECT 83.950 146.995 84.280 147.375 ;
        RECT 84.450 147.255 84.620 147.545 ;
        RECT 85.420 147.380 85.590 148.225 ;
        RECT 86.040 148.055 86.260 148.925 ;
        RECT 86.485 148.805 87.180 148.995 ;
        RECT 85.760 147.675 86.260 148.055 ;
        RECT 86.430 148.005 86.840 148.625 ;
        RECT 87.010 147.835 87.180 148.805 ;
        RECT 86.485 147.665 87.180 147.835 ;
        RECT 84.800 146.995 85.180 147.375 ;
        RECT 85.420 147.210 86.250 147.380 ;
        RECT 86.485 147.165 86.655 147.665 ;
        RECT 86.825 146.995 87.155 147.495 ;
        RECT 87.370 147.165 87.595 149.285 ;
        RECT 87.765 149.165 88.095 149.545 ;
        RECT 88.265 148.995 88.435 149.285 ;
        RECT 87.770 148.825 88.435 148.995 ;
        RECT 89.070 148.835 89.325 149.365 ;
        RECT 89.505 149.085 89.790 149.545 ;
        RECT 87.770 147.835 88.000 148.825 ;
        RECT 88.170 148.005 88.520 148.655 ;
        RECT 89.070 147.975 89.250 148.835 ;
        RECT 89.970 148.635 90.220 149.285 ;
        RECT 89.420 148.305 90.220 148.635 ;
        RECT 87.770 147.665 88.435 147.835 ;
        RECT 87.765 146.995 88.095 147.495 ;
        RECT 88.265 147.165 88.435 147.665 ;
        RECT 89.070 147.505 89.325 147.975 ;
        RECT 88.985 147.335 89.325 147.505 ;
        RECT 89.070 147.305 89.325 147.335 ;
        RECT 89.505 146.995 89.790 147.795 ;
        RECT 89.970 147.715 90.220 148.305 ;
        RECT 90.420 148.950 90.740 149.280 ;
        RECT 90.920 149.065 91.580 149.545 ;
        RECT 91.780 149.155 92.630 149.325 ;
        RECT 90.420 148.055 90.610 148.950 ;
        RECT 90.930 148.625 91.590 148.895 ;
        RECT 91.260 148.565 91.590 148.625 ;
        RECT 90.780 148.395 91.110 148.455 ;
        RECT 91.780 148.395 91.950 149.155 ;
        RECT 93.190 149.085 93.510 149.545 ;
        RECT 93.710 148.905 93.960 149.335 ;
        RECT 94.250 149.105 94.660 149.545 ;
        RECT 94.830 149.165 95.845 149.365 ;
        RECT 92.120 148.735 93.370 148.905 ;
        RECT 92.120 148.615 92.450 148.735 ;
        RECT 90.780 148.225 92.680 148.395 ;
        RECT 90.420 147.885 92.340 148.055 ;
        RECT 90.420 147.865 90.740 147.885 ;
        RECT 89.970 147.205 90.300 147.715 ;
        RECT 90.570 147.255 90.740 147.865 ;
        RECT 92.510 147.715 92.680 148.225 ;
        RECT 92.850 148.155 93.030 148.565 ;
        RECT 93.200 147.975 93.370 148.735 ;
        RECT 90.910 146.995 91.240 147.685 ;
        RECT 91.470 147.545 92.680 147.715 ;
        RECT 92.850 147.665 93.370 147.975 ;
        RECT 93.540 148.565 93.960 148.905 ;
        RECT 94.250 148.565 94.660 148.895 ;
        RECT 93.540 147.795 93.730 148.565 ;
        RECT 94.830 148.435 95.000 149.165 ;
        RECT 96.145 148.995 96.315 149.325 ;
        RECT 96.485 149.165 96.815 149.545 ;
        RECT 95.170 148.615 95.520 148.985 ;
        RECT 94.830 148.395 95.250 148.435 ;
        RECT 93.900 148.225 95.250 148.395 ;
        RECT 93.900 148.065 94.150 148.225 ;
        RECT 94.660 147.795 94.910 148.055 ;
        RECT 93.540 147.545 94.910 147.795 ;
        RECT 91.470 147.255 91.710 147.545 ;
        RECT 92.510 147.465 92.680 147.545 ;
        RECT 91.910 146.995 92.330 147.375 ;
        RECT 92.510 147.215 93.140 147.465 ;
        RECT 93.610 146.995 93.940 147.375 ;
        RECT 94.110 147.255 94.280 147.545 ;
        RECT 95.080 147.380 95.250 148.225 ;
        RECT 95.700 148.055 95.920 148.925 ;
        RECT 96.145 148.805 96.840 148.995 ;
        RECT 95.420 147.675 95.920 148.055 ;
        RECT 96.090 148.005 96.500 148.625 ;
        RECT 96.670 147.835 96.840 148.805 ;
        RECT 96.145 147.665 96.840 147.835 ;
        RECT 94.460 146.995 94.840 147.375 ;
        RECT 95.080 147.210 95.910 147.380 ;
        RECT 96.145 147.165 96.315 147.665 ;
        RECT 96.485 146.995 96.815 147.495 ;
        RECT 97.030 147.165 97.255 149.285 ;
        RECT 97.425 149.165 97.755 149.545 ;
        RECT 97.925 148.995 98.095 149.285 ;
        RECT 97.430 148.825 98.095 148.995 ;
        RECT 97.430 147.835 97.660 148.825 ;
        RECT 98.395 148.725 98.625 149.545 ;
        RECT 98.795 148.745 99.125 149.375 ;
        RECT 97.830 148.005 98.180 148.655 ;
        RECT 98.375 148.305 98.705 148.555 ;
        RECT 98.875 148.145 99.125 148.745 ;
        RECT 99.295 148.725 99.505 149.545 ;
        RECT 100.195 148.820 100.485 149.545 ;
        RECT 101.490 149.205 101.745 149.365 ;
        RECT 101.405 149.035 101.745 149.205 ;
        RECT 101.925 149.085 102.210 149.545 ;
        RECT 101.490 148.835 101.745 149.035 ;
        RECT 97.430 147.665 98.095 147.835 ;
        RECT 97.425 146.995 97.755 147.495 ;
        RECT 97.925 147.165 98.095 147.665 ;
        RECT 98.395 146.995 98.625 148.135 ;
        RECT 98.795 147.165 99.125 148.145 ;
        RECT 99.295 146.995 99.505 148.135 ;
        RECT 100.195 146.995 100.485 148.160 ;
        RECT 101.490 147.975 101.670 148.835 ;
        RECT 102.390 148.635 102.640 149.285 ;
        RECT 101.840 148.305 102.640 148.635 ;
        RECT 101.490 147.305 101.745 147.975 ;
        RECT 101.925 146.995 102.210 147.795 ;
        RECT 102.390 147.715 102.640 148.305 ;
        RECT 102.840 148.950 103.160 149.280 ;
        RECT 103.340 149.065 104.000 149.545 ;
        RECT 104.200 149.155 105.050 149.325 ;
        RECT 102.840 148.055 103.030 148.950 ;
        RECT 103.350 148.625 104.010 148.895 ;
        RECT 103.680 148.565 104.010 148.625 ;
        RECT 103.200 148.395 103.530 148.455 ;
        RECT 104.200 148.395 104.370 149.155 ;
        RECT 105.610 149.085 105.930 149.545 ;
        RECT 106.130 148.905 106.380 149.335 ;
        RECT 106.670 149.105 107.080 149.545 ;
        RECT 107.250 149.165 108.265 149.365 ;
        RECT 104.540 148.735 105.790 148.905 ;
        RECT 104.540 148.615 104.870 148.735 ;
        RECT 103.200 148.225 105.100 148.395 ;
        RECT 102.840 147.885 104.760 148.055 ;
        RECT 102.840 147.865 103.160 147.885 ;
        RECT 102.390 147.205 102.720 147.715 ;
        RECT 102.990 147.255 103.160 147.865 ;
        RECT 104.930 147.715 105.100 148.225 ;
        RECT 105.270 148.155 105.450 148.565 ;
        RECT 105.620 147.975 105.790 148.735 ;
        RECT 103.330 146.995 103.660 147.685 ;
        RECT 103.890 147.545 105.100 147.715 ;
        RECT 105.270 147.665 105.790 147.975 ;
        RECT 105.960 148.565 106.380 148.905 ;
        RECT 106.670 148.565 107.080 148.895 ;
        RECT 105.960 147.795 106.150 148.565 ;
        RECT 107.250 148.435 107.420 149.165 ;
        RECT 108.565 148.995 108.735 149.325 ;
        RECT 108.905 149.165 109.235 149.545 ;
        RECT 107.590 148.615 107.940 148.985 ;
        RECT 107.250 148.395 107.670 148.435 ;
        RECT 106.320 148.225 107.670 148.395 ;
        RECT 106.320 148.065 106.570 148.225 ;
        RECT 107.080 147.795 107.330 148.055 ;
        RECT 105.960 147.545 107.330 147.795 ;
        RECT 103.890 147.255 104.130 147.545 ;
        RECT 104.930 147.465 105.100 147.545 ;
        RECT 104.330 146.995 104.750 147.375 ;
        RECT 104.930 147.215 105.560 147.465 ;
        RECT 106.030 146.995 106.360 147.375 ;
        RECT 106.530 147.255 106.700 147.545 ;
        RECT 107.500 147.380 107.670 148.225 ;
        RECT 108.120 148.055 108.340 148.925 ;
        RECT 108.565 148.805 109.260 148.995 ;
        RECT 107.840 147.675 108.340 148.055 ;
        RECT 108.510 148.005 108.920 148.625 ;
        RECT 109.090 147.835 109.260 148.805 ;
        RECT 108.565 147.665 109.260 147.835 ;
        RECT 106.880 146.995 107.260 147.375 ;
        RECT 107.500 147.210 108.330 147.380 ;
        RECT 108.565 147.165 108.735 147.665 ;
        RECT 108.905 146.995 109.235 147.495 ;
        RECT 109.450 147.165 109.675 149.285 ;
        RECT 109.845 149.165 110.175 149.545 ;
        RECT 110.345 148.995 110.515 149.285 ;
        RECT 109.850 148.825 110.515 148.995 ;
        RECT 109.850 147.835 110.080 148.825 ;
        RECT 110.815 148.725 111.045 149.545 ;
        RECT 111.215 148.745 111.545 149.375 ;
        RECT 110.250 148.005 110.600 148.655 ;
        RECT 110.795 148.305 111.125 148.555 ;
        RECT 111.295 148.145 111.545 148.745 ;
        RECT 111.715 148.725 111.925 149.545 ;
        RECT 112.155 148.795 113.365 149.545 ;
        RECT 109.850 147.665 110.515 147.835 ;
        RECT 109.845 146.995 110.175 147.495 ;
        RECT 110.345 147.165 110.515 147.665 ;
        RECT 110.815 146.995 111.045 148.135 ;
        RECT 111.215 147.165 111.545 148.145 ;
        RECT 111.715 146.995 111.925 148.135 ;
        RECT 112.155 148.085 112.675 148.625 ;
        RECT 112.845 148.255 113.365 148.795 ;
        RECT 112.155 146.995 113.365 148.085 ;
        RECT 26.970 146.825 113.450 146.995 ;
        RECT 27.055 145.735 28.265 146.825 ;
        RECT 29.555 146.155 29.835 146.825 ;
        RECT 30.005 145.935 30.305 146.485 ;
        RECT 30.505 146.105 30.835 146.825 ;
        RECT 31.025 146.105 31.485 146.655 ;
        RECT 27.055 145.025 27.575 145.565 ;
        RECT 27.745 145.195 28.265 145.735 ;
        RECT 29.370 145.515 29.635 145.875 ;
        RECT 30.005 145.765 30.945 145.935 ;
        RECT 30.775 145.515 30.945 145.765 ;
        RECT 29.370 145.265 30.045 145.515 ;
        RECT 30.265 145.265 30.605 145.515 ;
        RECT 30.775 145.185 31.065 145.515 ;
        RECT 30.775 145.095 30.945 145.185 ;
        RECT 27.055 144.275 28.265 145.025 ;
        RECT 29.555 144.905 30.945 145.095 ;
        RECT 29.555 144.545 29.885 144.905 ;
        RECT 31.235 144.735 31.485 146.105 ;
        RECT 30.505 144.275 30.755 144.735 ;
        RECT 30.925 144.445 31.485 144.735 ;
        RECT 31.660 145.685 31.995 146.655 ;
        RECT 32.165 145.685 32.335 146.825 ;
        RECT 32.505 146.485 34.535 146.655 ;
        RECT 31.660 145.015 31.830 145.685 ;
        RECT 32.505 145.515 32.675 146.485 ;
        RECT 32.000 145.185 32.255 145.515 ;
        RECT 32.480 145.185 32.675 145.515 ;
        RECT 32.845 146.145 33.970 146.315 ;
        RECT 32.085 145.015 32.255 145.185 ;
        RECT 32.845 145.015 33.015 146.145 ;
        RECT 31.660 144.445 31.915 145.015 ;
        RECT 32.085 144.845 33.015 145.015 ;
        RECT 33.185 145.805 34.195 145.975 ;
        RECT 33.185 145.005 33.355 145.805 ;
        RECT 33.560 145.465 33.835 145.605 ;
        RECT 33.555 145.295 33.835 145.465 ;
        RECT 32.840 144.810 33.015 144.845 ;
        RECT 32.085 144.275 32.415 144.675 ;
        RECT 32.840 144.445 33.370 144.810 ;
        RECT 33.560 144.445 33.835 145.295 ;
        RECT 34.005 144.445 34.195 145.805 ;
        RECT 34.365 145.820 34.535 146.485 ;
        RECT 34.705 146.065 34.875 146.825 ;
        RECT 35.110 146.065 35.625 146.475 ;
        RECT 34.365 145.630 35.115 145.820 ;
        RECT 35.285 145.255 35.625 146.065 ;
        RECT 35.795 145.660 36.085 146.825 ;
        RECT 36.255 146.065 36.770 146.475 ;
        RECT 37.005 146.065 37.175 146.825 ;
        RECT 37.345 146.485 39.375 146.655 ;
        RECT 34.395 145.085 35.625 145.255 ;
        RECT 36.255 145.255 36.595 146.065 ;
        RECT 37.345 145.820 37.515 146.485 ;
        RECT 37.910 146.145 39.035 146.315 ;
        RECT 36.765 145.630 37.515 145.820 ;
        RECT 37.685 145.805 38.695 145.975 ;
        RECT 36.255 145.085 37.485 145.255 ;
        RECT 34.375 144.275 34.885 144.810 ;
        RECT 35.105 144.480 35.350 145.085 ;
        RECT 35.795 144.275 36.085 145.000 ;
        RECT 36.530 144.480 36.775 145.085 ;
        RECT 36.995 144.275 37.505 144.810 ;
        RECT 37.685 144.445 37.875 145.805 ;
        RECT 38.045 145.125 38.320 145.605 ;
        RECT 38.045 144.955 38.325 145.125 ;
        RECT 38.525 145.005 38.695 145.805 ;
        RECT 38.865 145.015 39.035 146.145 ;
        RECT 39.205 145.515 39.375 146.485 ;
        RECT 39.545 145.685 39.715 146.825 ;
        RECT 39.885 145.685 40.220 146.655 ;
        RECT 39.205 145.185 39.400 145.515 ;
        RECT 39.625 145.185 39.880 145.515 ;
        RECT 39.625 145.015 39.795 145.185 ;
        RECT 40.050 145.015 40.220 145.685 ;
        RECT 40.770 145.845 41.025 146.515 ;
        RECT 41.205 146.025 41.490 146.825 ;
        RECT 41.670 146.105 42.000 146.615 ;
        RECT 40.770 145.125 40.950 145.845 ;
        RECT 41.670 145.515 41.920 146.105 ;
        RECT 42.270 145.955 42.440 146.565 ;
        RECT 42.610 146.135 42.940 146.825 ;
        RECT 43.170 146.275 43.410 146.565 ;
        RECT 43.610 146.445 44.030 146.825 ;
        RECT 44.210 146.355 44.840 146.605 ;
        RECT 45.310 146.445 45.640 146.825 ;
        RECT 44.210 146.275 44.380 146.355 ;
        RECT 45.810 146.275 45.980 146.565 ;
        RECT 46.160 146.445 46.540 146.825 ;
        RECT 46.780 146.440 47.610 146.610 ;
        RECT 43.170 146.105 44.380 146.275 ;
        RECT 41.120 145.185 41.920 145.515 ;
        RECT 38.045 144.445 38.320 144.955 ;
        RECT 38.865 144.845 39.795 145.015 ;
        RECT 38.865 144.810 39.040 144.845 ;
        RECT 38.510 144.445 39.040 144.810 ;
        RECT 39.465 144.275 39.795 144.675 ;
        RECT 39.965 144.445 40.220 145.015 ;
        RECT 40.685 144.985 40.950 145.125 ;
        RECT 40.685 144.955 41.025 144.985 ;
        RECT 40.770 144.455 41.025 144.955 ;
        RECT 41.205 144.275 41.490 144.735 ;
        RECT 41.670 144.535 41.920 145.185 ;
        RECT 42.120 145.935 42.440 145.955 ;
        RECT 42.120 145.765 44.040 145.935 ;
        RECT 42.120 144.870 42.310 145.765 ;
        RECT 44.210 145.595 44.380 146.105 ;
        RECT 44.550 145.845 45.070 146.155 ;
        RECT 42.480 145.425 44.380 145.595 ;
        RECT 42.480 145.365 42.810 145.425 ;
        RECT 42.960 145.195 43.290 145.255 ;
        RECT 42.630 144.925 43.290 145.195 ;
        RECT 42.120 144.540 42.440 144.870 ;
        RECT 42.620 144.275 43.280 144.755 ;
        RECT 43.480 144.665 43.650 145.425 ;
        RECT 44.550 145.255 44.730 145.665 ;
        RECT 43.820 145.085 44.150 145.205 ;
        RECT 44.900 145.085 45.070 145.845 ;
        RECT 43.820 144.915 45.070 145.085 ;
        RECT 45.240 146.025 46.610 146.275 ;
        RECT 45.240 145.255 45.430 146.025 ;
        RECT 46.360 145.765 46.610 146.025 ;
        RECT 45.600 145.595 45.850 145.755 ;
        RECT 46.780 145.595 46.950 146.440 ;
        RECT 47.845 146.155 48.015 146.655 ;
        RECT 48.185 146.325 48.515 146.825 ;
        RECT 47.120 145.765 47.620 146.145 ;
        RECT 47.845 145.985 48.540 146.155 ;
        RECT 45.600 145.425 46.950 145.595 ;
        RECT 46.530 145.385 46.950 145.425 ;
        RECT 45.240 144.915 45.660 145.255 ;
        RECT 45.950 144.925 46.360 145.255 ;
        RECT 43.480 144.495 44.330 144.665 ;
        RECT 44.890 144.275 45.210 144.735 ;
        RECT 45.410 144.485 45.660 144.915 ;
        RECT 45.950 144.275 46.360 144.715 ;
        RECT 46.530 144.655 46.700 145.385 ;
        RECT 46.870 144.835 47.220 145.205 ;
        RECT 47.400 144.895 47.620 145.765 ;
        RECT 47.790 145.195 48.200 145.815 ;
        RECT 48.370 145.015 48.540 145.985 ;
        RECT 47.845 144.825 48.540 145.015 ;
        RECT 46.530 144.455 47.545 144.655 ;
        RECT 47.845 144.495 48.015 144.825 ;
        RECT 48.185 144.275 48.515 144.655 ;
        RECT 48.730 144.535 48.955 146.655 ;
        RECT 49.125 146.325 49.455 146.825 ;
        RECT 49.625 146.155 49.795 146.655 ;
        RECT 49.130 145.985 49.795 146.155 ;
        RECT 50.055 146.065 50.570 146.475 ;
        RECT 50.805 146.065 50.975 146.825 ;
        RECT 51.145 146.485 53.175 146.655 ;
        RECT 49.130 144.995 49.360 145.985 ;
        RECT 49.530 145.165 49.880 145.815 ;
        RECT 50.055 145.255 50.395 146.065 ;
        RECT 51.145 145.820 51.315 146.485 ;
        RECT 51.710 146.145 52.835 146.315 ;
        RECT 50.565 145.630 51.315 145.820 ;
        RECT 51.485 145.805 52.495 145.975 ;
        RECT 50.055 145.085 51.285 145.255 ;
        RECT 49.130 144.825 49.795 144.995 ;
        RECT 49.125 144.275 49.455 144.655 ;
        RECT 49.625 144.535 49.795 144.825 ;
        RECT 50.330 144.480 50.575 145.085 ;
        RECT 50.795 144.275 51.305 144.810 ;
        RECT 51.485 144.445 51.675 145.805 ;
        RECT 51.845 144.785 52.120 145.605 ;
        RECT 52.325 145.005 52.495 145.805 ;
        RECT 52.665 145.015 52.835 146.145 ;
        RECT 53.005 145.515 53.175 146.485 ;
        RECT 53.345 145.685 53.515 146.825 ;
        RECT 53.685 145.685 54.020 146.655 ;
        RECT 54.400 145.855 54.730 146.655 ;
        RECT 54.900 146.025 55.230 146.825 ;
        RECT 55.530 145.855 55.860 146.655 ;
        RECT 56.505 146.025 56.755 146.825 ;
        RECT 54.400 145.685 56.835 145.855 ;
        RECT 57.025 145.685 57.195 146.825 ;
        RECT 57.365 145.685 57.705 146.655 ;
        RECT 53.005 145.185 53.200 145.515 ;
        RECT 53.425 145.185 53.680 145.515 ;
        RECT 53.425 145.015 53.595 145.185 ;
        RECT 53.850 145.015 54.020 145.685 ;
        RECT 54.195 145.265 54.545 145.515 ;
        RECT 54.730 145.055 54.900 145.685 ;
        RECT 55.070 145.265 55.400 145.465 ;
        RECT 55.570 145.265 55.900 145.465 ;
        RECT 56.070 145.265 56.490 145.465 ;
        RECT 56.665 145.435 56.835 145.685 ;
        RECT 56.665 145.265 57.360 145.435 ;
        RECT 52.665 144.845 53.595 145.015 ;
        RECT 52.665 144.810 52.840 144.845 ;
        RECT 51.845 144.615 52.125 144.785 ;
        RECT 51.845 144.445 52.120 144.615 ;
        RECT 52.310 144.445 52.840 144.810 ;
        RECT 53.265 144.275 53.595 144.675 ;
        RECT 53.765 144.445 54.020 145.015 ;
        RECT 54.400 144.445 54.900 145.055 ;
        RECT 55.530 144.925 56.755 145.095 ;
        RECT 57.530 145.075 57.705 145.685 ;
        RECT 55.530 144.445 55.860 144.925 ;
        RECT 56.030 144.275 56.255 144.735 ;
        RECT 56.425 144.445 56.755 144.925 ;
        RECT 56.945 144.275 57.195 145.075 ;
        RECT 57.365 144.445 57.705 145.075 ;
        RECT 57.875 145.685 58.215 146.655 ;
        RECT 58.385 145.685 58.555 146.825 ;
        RECT 58.825 146.025 59.075 146.825 ;
        RECT 59.720 145.855 60.050 146.655 ;
        RECT 60.350 146.025 60.680 146.825 ;
        RECT 60.850 145.855 61.180 146.655 ;
        RECT 58.745 145.685 61.180 145.855 ;
        RECT 57.875 145.075 58.050 145.685 ;
        RECT 58.745 145.435 58.915 145.685 ;
        RECT 58.220 145.265 58.915 145.435 ;
        RECT 59.090 145.265 59.510 145.465 ;
        RECT 59.680 145.265 60.010 145.465 ;
        RECT 60.180 145.265 60.510 145.465 ;
        RECT 57.875 144.445 58.215 145.075 ;
        RECT 58.385 144.275 58.635 145.075 ;
        RECT 58.825 144.925 60.050 145.095 ;
        RECT 58.825 144.445 59.155 144.925 ;
        RECT 59.325 144.275 59.550 144.735 ;
        RECT 59.720 144.445 60.050 144.925 ;
        RECT 60.680 145.055 60.850 145.685 ;
        RECT 61.555 145.660 61.845 146.825 ;
        RECT 62.975 145.685 63.205 146.825 ;
        RECT 63.375 145.675 63.705 146.655 ;
        RECT 63.875 145.685 64.085 146.825 ;
        RECT 64.315 146.065 64.830 146.475 ;
        RECT 65.065 146.065 65.235 146.825 ;
        RECT 65.405 146.485 67.435 146.655 ;
        RECT 61.035 145.265 61.385 145.515 ;
        RECT 62.955 145.265 63.285 145.515 ;
        RECT 60.680 144.445 61.180 145.055 ;
        RECT 61.555 144.275 61.845 145.000 ;
        RECT 62.975 144.275 63.205 145.095 ;
        RECT 63.455 145.075 63.705 145.675 ;
        RECT 64.315 145.255 64.655 146.065 ;
        RECT 65.405 145.820 65.575 146.485 ;
        RECT 65.970 146.145 67.095 146.315 ;
        RECT 64.825 145.630 65.575 145.820 ;
        RECT 65.745 145.805 66.755 145.975 ;
        RECT 63.375 144.445 63.705 145.075 ;
        RECT 63.875 144.275 64.085 145.095 ;
        RECT 64.315 145.085 65.545 145.255 ;
        RECT 64.590 144.480 64.835 145.085 ;
        RECT 65.055 144.275 65.565 144.810 ;
        RECT 65.745 144.445 65.935 145.805 ;
        RECT 66.105 145.125 66.380 145.605 ;
        RECT 66.105 144.955 66.385 145.125 ;
        RECT 66.585 145.005 66.755 145.805 ;
        RECT 66.925 145.015 67.095 146.145 ;
        RECT 67.265 145.515 67.435 146.485 ;
        RECT 67.605 145.685 67.775 146.825 ;
        RECT 67.945 145.685 68.280 146.655 ;
        RECT 69.115 146.155 69.395 146.825 ;
        RECT 69.565 145.935 69.865 146.485 ;
        RECT 70.065 146.105 70.395 146.825 ;
        RECT 70.585 146.105 71.045 146.655 ;
        RECT 67.265 145.185 67.460 145.515 ;
        RECT 67.685 145.185 67.940 145.515 ;
        RECT 67.685 145.015 67.855 145.185 ;
        RECT 68.110 145.015 68.280 145.685 ;
        RECT 68.930 145.515 69.195 145.875 ;
        RECT 69.565 145.765 70.505 145.935 ;
        RECT 70.335 145.515 70.505 145.765 ;
        RECT 68.930 145.265 69.605 145.515 ;
        RECT 69.825 145.265 70.165 145.515 ;
        RECT 70.335 145.185 70.625 145.515 ;
        RECT 70.335 145.095 70.505 145.185 ;
        RECT 66.105 144.445 66.380 144.955 ;
        RECT 66.925 144.845 67.855 145.015 ;
        RECT 66.925 144.810 67.100 144.845 ;
        RECT 66.570 144.445 67.100 144.810 ;
        RECT 67.525 144.275 67.855 144.675 ;
        RECT 68.025 144.445 68.280 145.015 ;
        RECT 69.115 144.905 70.505 145.095 ;
        RECT 69.115 144.545 69.445 144.905 ;
        RECT 70.795 144.735 71.045 146.105 ;
        RECT 70.065 144.275 70.315 144.735 ;
        RECT 70.485 144.445 71.045 144.735 ;
        RECT 71.215 145.855 71.525 146.655 ;
        RECT 71.695 146.025 72.005 146.825 ;
        RECT 72.175 146.195 72.435 146.655 ;
        RECT 72.605 146.365 72.860 146.825 ;
        RECT 73.035 146.195 73.295 146.655 ;
        RECT 72.175 146.025 73.295 146.195 ;
        RECT 71.215 145.685 72.245 145.855 ;
        RECT 71.215 144.775 71.385 145.685 ;
        RECT 71.555 144.945 71.905 145.515 ;
        RECT 72.075 145.435 72.245 145.685 ;
        RECT 73.035 145.775 73.295 146.025 ;
        RECT 73.465 145.955 73.750 146.825 ;
        RECT 73.035 145.605 73.790 145.775 ;
        RECT 72.075 145.265 73.215 145.435 ;
        RECT 73.385 145.095 73.790 145.605 ;
        RECT 72.140 144.925 73.790 145.095 ;
        RECT 73.975 145.685 74.245 146.655 ;
        RECT 74.455 146.025 74.735 146.825 ;
        RECT 74.905 146.315 76.560 146.605 ;
        RECT 74.970 145.975 76.560 146.145 ;
        RECT 74.970 145.855 75.140 145.975 ;
        RECT 74.415 145.685 75.140 145.855 ;
        RECT 73.975 144.950 74.145 145.685 ;
        RECT 74.415 145.515 74.585 145.685 ;
        RECT 74.315 145.185 74.585 145.515 ;
        RECT 74.755 145.185 75.160 145.515 ;
        RECT 75.330 145.185 76.040 145.805 ;
        RECT 76.240 145.685 76.560 145.975 ;
        RECT 76.735 145.685 77.075 146.655 ;
        RECT 77.245 145.685 77.415 146.825 ;
        RECT 77.685 146.025 77.935 146.825 ;
        RECT 78.580 145.855 78.910 146.655 ;
        RECT 79.210 146.025 79.540 146.825 ;
        RECT 79.710 145.855 80.040 146.655 ;
        RECT 77.605 145.685 80.040 145.855 ;
        RECT 80.875 146.065 81.390 146.475 ;
        RECT 81.625 146.065 81.795 146.825 ;
        RECT 81.965 146.485 83.995 146.655 ;
        RECT 74.415 145.015 74.585 145.185 ;
        RECT 71.215 144.445 71.515 144.775 ;
        RECT 71.685 144.275 71.960 144.755 ;
        RECT 72.140 144.535 72.435 144.925 ;
        RECT 72.605 144.275 72.860 144.755 ;
        RECT 73.035 144.535 73.295 144.925 ;
        RECT 73.465 144.275 73.745 144.755 ;
        RECT 73.975 144.605 74.245 144.950 ;
        RECT 74.415 144.845 76.025 145.015 ;
        RECT 76.210 144.945 76.560 145.515 ;
        RECT 76.735 145.125 76.910 145.685 ;
        RECT 77.605 145.435 77.775 145.685 ;
        RECT 77.080 145.265 77.775 145.435 ;
        RECT 77.950 145.265 78.370 145.465 ;
        RECT 78.540 145.265 78.870 145.465 ;
        RECT 79.040 145.265 79.370 145.465 ;
        RECT 76.735 145.075 76.965 145.125 ;
        RECT 74.435 144.275 74.815 144.675 ;
        RECT 74.985 144.495 75.155 144.845 ;
        RECT 75.325 144.275 75.655 144.675 ;
        RECT 75.855 144.495 76.025 144.845 ;
        RECT 76.225 144.275 76.555 144.775 ;
        RECT 76.735 144.445 77.075 145.075 ;
        RECT 77.245 144.275 77.495 145.075 ;
        RECT 77.685 144.925 78.910 145.095 ;
        RECT 77.685 144.445 78.015 144.925 ;
        RECT 78.185 144.275 78.410 144.735 ;
        RECT 78.580 144.445 78.910 144.925 ;
        RECT 79.540 145.055 79.710 145.685 ;
        RECT 79.895 145.265 80.245 145.515 ;
        RECT 80.875 145.255 81.215 146.065 ;
        RECT 81.965 145.820 82.135 146.485 ;
        RECT 82.530 146.145 83.655 146.315 ;
        RECT 81.385 145.630 82.135 145.820 ;
        RECT 82.305 145.805 83.315 145.975 ;
        RECT 80.875 145.085 82.105 145.255 ;
        RECT 79.540 144.445 80.040 145.055 ;
        RECT 81.150 144.480 81.395 145.085 ;
        RECT 81.615 144.275 82.125 144.810 ;
        RECT 82.305 144.445 82.495 145.805 ;
        RECT 82.665 145.465 82.940 145.605 ;
        RECT 82.665 145.295 82.945 145.465 ;
        RECT 82.665 144.445 82.940 145.295 ;
        RECT 83.145 145.005 83.315 145.805 ;
        RECT 83.485 145.015 83.655 146.145 ;
        RECT 83.825 145.515 83.995 146.485 ;
        RECT 84.165 145.685 84.335 146.825 ;
        RECT 84.505 145.685 84.840 146.655 ;
        RECT 85.105 145.895 85.275 146.655 ;
        RECT 85.455 146.065 85.785 146.825 ;
        RECT 85.105 145.725 85.770 145.895 ;
        RECT 85.955 145.750 86.225 146.655 ;
        RECT 83.825 145.185 84.020 145.515 ;
        RECT 84.245 145.185 84.500 145.515 ;
        RECT 84.245 145.015 84.415 145.185 ;
        RECT 84.670 145.015 84.840 145.685 ;
        RECT 85.600 145.580 85.770 145.725 ;
        RECT 85.035 145.175 85.365 145.545 ;
        RECT 85.600 145.250 85.885 145.580 ;
        RECT 83.485 144.845 84.415 145.015 ;
        RECT 83.485 144.810 83.660 144.845 ;
        RECT 83.130 144.445 83.660 144.810 ;
        RECT 84.085 144.275 84.415 144.675 ;
        RECT 84.585 144.445 84.840 145.015 ;
        RECT 85.600 144.995 85.770 145.250 ;
        RECT 85.105 144.825 85.770 144.995 ;
        RECT 86.055 144.950 86.225 145.750 ;
        RECT 87.315 145.660 87.605 146.825 ;
        RECT 87.775 146.065 88.290 146.475 ;
        RECT 88.525 146.065 88.695 146.825 ;
        RECT 88.865 146.485 90.895 146.655 ;
        RECT 87.775 145.255 88.115 146.065 ;
        RECT 88.865 145.820 89.035 146.485 ;
        RECT 89.430 146.145 90.555 146.315 ;
        RECT 88.285 145.630 89.035 145.820 ;
        RECT 89.205 145.805 90.215 145.975 ;
        RECT 87.775 145.085 89.005 145.255 ;
        RECT 85.105 144.445 85.275 144.825 ;
        RECT 85.455 144.275 85.785 144.655 ;
        RECT 85.965 144.445 86.225 144.950 ;
        RECT 87.315 144.275 87.605 145.000 ;
        RECT 88.050 144.480 88.295 145.085 ;
        RECT 88.515 144.275 89.025 144.810 ;
        RECT 89.205 144.445 89.395 145.805 ;
        RECT 89.565 144.785 89.840 145.605 ;
        RECT 90.045 145.005 90.215 145.805 ;
        RECT 90.385 145.015 90.555 146.145 ;
        RECT 90.725 145.515 90.895 146.485 ;
        RECT 91.065 145.685 91.235 146.825 ;
        RECT 91.405 145.685 91.740 146.655 ;
        RECT 91.955 145.685 92.185 146.825 ;
        RECT 90.725 145.185 90.920 145.515 ;
        RECT 91.145 145.185 91.400 145.515 ;
        RECT 91.145 145.015 91.315 145.185 ;
        RECT 91.570 145.015 91.740 145.685 ;
        RECT 92.355 145.675 92.685 146.655 ;
        RECT 92.855 145.685 93.065 146.825 ;
        RECT 93.295 146.105 93.755 146.655 ;
        RECT 93.945 146.105 94.275 146.825 ;
        RECT 91.935 145.265 92.265 145.515 ;
        RECT 90.385 144.845 91.315 145.015 ;
        RECT 90.385 144.810 90.560 144.845 ;
        RECT 89.565 144.615 89.845 144.785 ;
        RECT 89.565 144.445 89.840 144.615 ;
        RECT 90.030 144.445 90.560 144.810 ;
        RECT 90.985 144.275 91.315 144.675 ;
        RECT 91.485 144.445 91.740 145.015 ;
        RECT 91.955 144.275 92.185 145.095 ;
        RECT 92.435 145.075 92.685 145.675 ;
        RECT 92.355 144.445 92.685 145.075 ;
        RECT 92.855 144.275 93.065 145.095 ;
        RECT 93.295 144.735 93.545 146.105 ;
        RECT 94.475 145.935 94.775 146.485 ;
        RECT 94.945 146.155 95.225 146.825 ;
        RECT 95.795 146.155 96.075 146.825 ;
        RECT 93.835 145.765 94.775 145.935 ;
        RECT 96.245 145.935 96.545 146.485 ;
        RECT 96.745 146.105 97.075 146.825 ;
        RECT 97.265 146.105 97.725 146.655 ;
        RECT 93.835 145.515 94.005 145.765 ;
        RECT 95.145 145.515 95.410 145.875 ;
        RECT 93.715 145.185 94.005 145.515 ;
        RECT 94.175 145.265 94.515 145.515 ;
        RECT 94.735 145.265 95.410 145.515 ;
        RECT 95.610 145.515 95.875 145.875 ;
        RECT 96.245 145.765 97.185 145.935 ;
        RECT 97.015 145.515 97.185 145.765 ;
        RECT 95.610 145.265 96.285 145.515 ;
        RECT 96.505 145.265 96.845 145.515 ;
        RECT 93.835 145.095 94.005 145.185 ;
        RECT 97.015 145.185 97.305 145.515 ;
        RECT 97.015 145.095 97.185 145.185 ;
        RECT 93.835 144.905 95.225 145.095 ;
        RECT 93.295 144.445 93.855 144.735 ;
        RECT 94.025 144.275 94.275 144.735 ;
        RECT 94.895 144.545 95.225 144.905 ;
        RECT 95.795 144.905 97.185 145.095 ;
        RECT 95.795 144.545 96.125 144.905 ;
        RECT 97.475 144.735 97.725 146.105 ;
        RECT 96.745 144.275 96.995 144.735 ;
        RECT 97.165 144.445 97.725 144.735 ;
        RECT 98.355 146.105 98.815 146.655 ;
        RECT 99.005 146.105 99.335 146.825 ;
        RECT 98.355 144.735 98.605 146.105 ;
        RECT 99.535 145.935 99.835 146.485 ;
        RECT 100.005 146.155 100.285 146.825 ;
        RECT 98.895 145.765 99.835 145.935 ;
        RECT 100.655 146.105 101.115 146.655 ;
        RECT 101.305 146.105 101.635 146.825 ;
        RECT 98.895 145.515 99.065 145.765 ;
        RECT 100.205 145.515 100.470 145.875 ;
        RECT 98.775 145.185 99.065 145.515 ;
        RECT 99.235 145.265 99.575 145.515 ;
        RECT 99.795 145.265 100.470 145.515 ;
        RECT 98.895 145.095 99.065 145.185 ;
        RECT 98.895 144.905 100.285 145.095 ;
        RECT 98.355 144.445 98.915 144.735 ;
        RECT 99.085 144.275 99.335 144.735 ;
        RECT 99.955 144.545 100.285 144.905 ;
        RECT 100.655 144.735 100.905 146.105 ;
        RECT 101.835 145.935 102.135 146.485 ;
        RECT 102.305 146.155 102.585 146.825 ;
        RECT 101.195 145.765 102.135 145.935 ;
        RECT 101.195 145.515 101.365 145.765 ;
        RECT 102.505 145.515 102.770 145.875 ;
        RECT 102.995 145.685 103.225 146.825 ;
        RECT 103.395 145.675 103.725 146.655 ;
        RECT 103.895 145.685 104.105 146.825 ;
        RECT 104.375 145.685 104.605 146.825 ;
        RECT 104.775 145.675 105.105 146.655 ;
        RECT 105.275 145.685 105.485 146.825 ;
        RECT 106.725 145.895 106.895 146.655 ;
        RECT 107.075 146.065 107.405 146.825 ;
        RECT 106.725 145.725 107.390 145.895 ;
        RECT 107.575 145.750 107.845 146.655 ;
        RECT 101.075 145.185 101.365 145.515 ;
        RECT 101.535 145.265 101.875 145.515 ;
        RECT 102.095 145.265 102.770 145.515 ;
        RECT 102.975 145.265 103.305 145.515 ;
        RECT 101.195 145.095 101.365 145.185 ;
        RECT 101.195 144.905 102.585 145.095 ;
        RECT 100.655 144.445 101.215 144.735 ;
        RECT 101.385 144.275 101.635 144.735 ;
        RECT 102.255 144.545 102.585 144.905 ;
        RECT 102.995 144.275 103.225 145.095 ;
        RECT 103.475 145.075 103.725 145.675 ;
        RECT 104.355 145.265 104.685 145.515 ;
        RECT 103.395 144.445 103.725 145.075 ;
        RECT 103.895 144.275 104.105 145.095 ;
        RECT 104.375 144.275 104.605 145.095 ;
        RECT 104.855 145.075 105.105 145.675 ;
        RECT 107.220 145.580 107.390 145.725 ;
        RECT 106.655 145.175 106.985 145.545 ;
        RECT 107.220 145.250 107.505 145.580 ;
        RECT 104.775 144.445 105.105 145.075 ;
        RECT 105.275 144.275 105.485 145.095 ;
        RECT 107.220 144.995 107.390 145.250 ;
        RECT 106.725 144.825 107.390 144.995 ;
        RECT 107.675 144.950 107.845 145.750 ;
        RECT 108.075 145.685 108.285 146.825 ;
        RECT 108.455 145.675 108.785 146.655 ;
        RECT 108.955 145.685 109.185 146.825 ;
        RECT 109.485 145.895 109.655 146.655 ;
        RECT 109.835 146.065 110.165 146.825 ;
        RECT 109.485 145.725 110.150 145.895 ;
        RECT 110.335 145.750 110.605 146.655 ;
        RECT 106.725 144.445 106.895 144.825 ;
        RECT 107.075 144.275 107.405 144.655 ;
        RECT 107.585 144.445 107.845 144.950 ;
        RECT 108.075 144.275 108.285 145.095 ;
        RECT 108.455 145.075 108.705 145.675 ;
        RECT 109.980 145.580 110.150 145.725 ;
        RECT 108.875 145.265 109.205 145.515 ;
        RECT 109.415 145.175 109.745 145.545 ;
        RECT 109.980 145.250 110.265 145.580 ;
        RECT 108.455 144.445 108.785 145.075 ;
        RECT 108.955 144.275 109.185 145.095 ;
        RECT 109.980 144.995 110.150 145.250 ;
        RECT 109.485 144.825 110.150 144.995 ;
        RECT 110.435 144.950 110.605 145.750 ;
        RECT 109.485 144.445 109.655 144.825 ;
        RECT 109.835 144.275 110.165 144.655 ;
        RECT 110.345 144.445 110.605 144.950 ;
        RECT 110.775 145.750 111.045 146.655 ;
        RECT 111.215 146.065 111.545 146.825 ;
        RECT 111.725 145.895 111.895 146.655 ;
        RECT 110.775 144.950 110.945 145.750 ;
        RECT 111.230 145.725 111.895 145.895 ;
        RECT 112.155 145.735 113.365 146.825 ;
        RECT 111.230 145.580 111.400 145.725 ;
        RECT 111.115 145.250 111.400 145.580 ;
        RECT 111.230 144.995 111.400 145.250 ;
        RECT 111.635 145.175 111.965 145.545 ;
        RECT 112.155 145.195 112.675 145.735 ;
        RECT 112.845 145.025 113.365 145.565 ;
        RECT 110.775 144.445 111.035 144.950 ;
        RECT 111.230 144.825 111.895 144.995 ;
        RECT 111.215 144.275 111.545 144.655 ;
        RECT 111.725 144.445 111.895 144.825 ;
        RECT 112.155 144.275 113.365 145.025 ;
        RECT 26.970 144.105 113.450 144.275 ;
        RECT 27.055 143.355 28.265 144.105 ;
        RECT 29.730 143.765 29.985 143.925 ;
        RECT 29.645 143.595 29.985 143.765 ;
        RECT 30.165 143.645 30.450 144.105 ;
        RECT 29.730 143.395 29.985 143.595 ;
        RECT 27.055 142.815 27.575 143.355 ;
        RECT 27.745 142.645 28.265 143.185 ;
        RECT 27.055 141.555 28.265 142.645 ;
        RECT 29.730 142.535 29.910 143.395 ;
        RECT 30.630 143.195 30.880 143.845 ;
        RECT 30.080 142.865 30.880 143.195 ;
        RECT 29.730 141.865 29.985 142.535 ;
        RECT 30.165 141.555 30.450 142.355 ;
        RECT 30.630 142.275 30.880 142.865 ;
        RECT 31.080 143.510 31.400 143.840 ;
        RECT 31.580 143.625 32.240 144.105 ;
        RECT 32.440 143.715 33.290 143.885 ;
        RECT 31.080 142.615 31.270 143.510 ;
        RECT 31.590 143.185 32.250 143.455 ;
        RECT 31.920 143.125 32.250 143.185 ;
        RECT 31.440 142.955 31.770 143.015 ;
        RECT 32.440 142.955 32.610 143.715 ;
        RECT 33.850 143.645 34.170 144.105 ;
        RECT 34.370 143.465 34.620 143.895 ;
        RECT 34.910 143.665 35.320 144.105 ;
        RECT 35.490 143.725 36.505 143.925 ;
        RECT 32.780 143.295 34.030 143.465 ;
        RECT 32.780 143.175 33.110 143.295 ;
        RECT 31.440 142.785 33.340 142.955 ;
        RECT 31.080 142.445 33.000 142.615 ;
        RECT 31.080 142.425 31.400 142.445 ;
        RECT 30.630 141.765 30.960 142.275 ;
        RECT 31.230 141.815 31.400 142.425 ;
        RECT 33.170 142.275 33.340 142.785 ;
        RECT 33.510 142.715 33.690 143.125 ;
        RECT 33.860 142.535 34.030 143.295 ;
        RECT 31.570 141.555 31.900 142.245 ;
        RECT 32.130 142.105 33.340 142.275 ;
        RECT 33.510 142.225 34.030 142.535 ;
        RECT 34.200 143.125 34.620 143.465 ;
        RECT 34.910 143.125 35.320 143.455 ;
        RECT 34.200 142.355 34.390 143.125 ;
        RECT 35.490 142.995 35.660 143.725 ;
        RECT 36.805 143.555 36.975 143.885 ;
        RECT 37.145 143.725 37.475 144.105 ;
        RECT 35.830 143.175 36.180 143.545 ;
        RECT 35.490 142.955 35.910 142.995 ;
        RECT 34.560 142.785 35.910 142.955 ;
        RECT 34.560 142.625 34.810 142.785 ;
        RECT 35.320 142.355 35.570 142.615 ;
        RECT 34.200 142.105 35.570 142.355 ;
        RECT 32.130 141.815 32.370 142.105 ;
        RECT 33.170 142.025 33.340 142.105 ;
        RECT 32.570 141.555 32.990 141.935 ;
        RECT 33.170 141.775 33.800 142.025 ;
        RECT 34.270 141.555 34.600 141.935 ;
        RECT 34.770 141.815 34.940 142.105 ;
        RECT 35.740 141.940 35.910 142.785 ;
        RECT 36.360 142.615 36.580 143.485 ;
        RECT 36.805 143.365 37.500 143.555 ;
        RECT 36.080 142.235 36.580 142.615 ;
        RECT 36.750 142.565 37.160 143.185 ;
        RECT 37.330 142.395 37.500 143.365 ;
        RECT 36.805 142.225 37.500 142.395 ;
        RECT 35.120 141.555 35.500 141.935 ;
        RECT 35.740 141.770 36.570 141.940 ;
        RECT 36.805 141.725 36.975 142.225 ;
        RECT 37.145 141.555 37.475 142.055 ;
        RECT 37.690 141.725 37.915 143.845 ;
        RECT 38.085 143.725 38.415 144.105 ;
        RECT 38.585 143.555 38.755 143.845 ;
        RECT 38.090 143.385 38.755 143.555 ;
        RECT 39.390 143.395 39.645 143.925 ;
        RECT 39.825 143.645 40.110 144.105 ;
        RECT 38.090 142.395 38.320 143.385 ;
        RECT 38.490 142.565 38.840 143.215 ;
        RECT 39.390 142.535 39.570 143.395 ;
        RECT 40.290 143.195 40.540 143.845 ;
        RECT 39.740 142.865 40.540 143.195 ;
        RECT 38.090 142.225 38.755 142.395 ;
        RECT 38.085 141.555 38.415 142.055 ;
        RECT 38.585 141.725 38.755 142.225 ;
        RECT 39.390 142.065 39.645 142.535 ;
        RECT 39.305 141.895 39.645 142.065 ;
        RECT 39.390 141.865 39.645 141.895 ;
        RECT 39.825 141.555 40.110 142.355 ;
        RECT 40.290 142.275 40.540 142.865 ;
        RECT 40.740 143.510 41.060 143.840 ;
        RECT 41.240 143.625 41.900 144.105 ;
        RECT 42.100 143.715 42.950 143.885 ;
        RECT 40.740 142.615 40.930 143.510 ;
        RECT 41.250 143.185 41.910 143.455 ;
        RECT 41.580 143.125 41.910 143.185 ;
        RECT 41.100 142.955 41.430 143.015 ;
        RECT 42.100 142.955 42.270 143.715 ;
        RECT 43.510 143.645 43.830 144.105 ;
        RECT 44.030 143.465 44.280 143.895 ;
        RECT 44.570 143.665 44.980 144.105 ;
        RECT 45.150 143.725 46.165 143.925 ;
        RECT 42.440 143.295 43.690 143.465 ;
        RECT 42.440 143.175 42.770 143.295 ;
        RECT 41.100 142.785 43.000 142.955 ;
        RECT 40.740 142.445 42.660 142.615 ;
        RECT 40.740 142.425 41.060 142.445 ;
        RECT 40.290 141.765 40.620 142.275 ;
        RECT 40.890 141.815 41.060 142.425 ;
        RECT 42.830 142.275 43.000 142.785 ;
        RECT 43.170 142.715 43.350 143.125 ;
        RECT 43.520 142.535 43.690 143.295 ;
        RECT 41.230 141.555 41.560 142.245 ;
        RECT 41.790 142.105 43.000 142.275 ;
        RECT 43.170 142.225 43.690 142.535 ;
        RECT 43.860 143.125 44.280 143.465 ;
        RECT 44.570 143.125 44.980 143.455 ;
        RECT 43.860 142.355 44.050 143.125 ;
        RECT 45.150 142.995 45.320 143.725 ;
        RECT 46.465 143.555 46.635 143.885 ;
        RECT 46.805 143.725 47.135 144.105 ;
        RECT 45.490 143.175 45.840 143.545 ;
        RECT 45.150 142.955 45.570 142.995 ;
        RECT 44.220 142.785 45.570 142.955 ;
        RECT 44.220 142.625 44.470 142.785 ;
        RECT 44.980 142.355 45.230 142.615 ;
        RECT 43.860 142.105 45.230 142.355 ;
        RECT 41.790 141.815 42.030 142.105 ;
        RECT 42.830 142.025 43.000 142.105 ;
        RECT 42.230 141.555 42.650 141.935 ;
        RECT 42.830 141.775 43.460 142.025 ;
        RECT 43.930 141.555 44.260 141.935 ;
        RECT 44.430 141.815 44.600 142.105 ;
        RECT 45.400 141.940 45.570 142.785 ;
        RECT 46.020 142.615 46.240 143.485 ;
        RECT 46.465 143.365 47.160 143.555 ;
        RECT 45.740 142.235 46.240 142.615 ;
        RECT 46.410 142.565 46.820 143.185 ;
        RECT 46.990 142.395 47.160 143.365 ;
        RECT 46.465 142.225 47.160 142.395 ;
        RECT 44.780 141.555 45.160 141.935 ;
        RECT 45.400 141.770 46.230 141.940 ;
        RECT 46.465 141.725 46.635 142.225 ;
        RECT 46.805 141.555 47.135 142.055 ;
        RECT 47.350 141.725 47.575 143.845 ;
        RECT 47.745 143.725 48.075 144.105 ;
        RECT 48.245 143.555 48.415 143.845 ;
        RECT 47.750 143.385 48.415 143.555 ;
        RECT 47.750 142.395 47.980 143.385 ;
        RECT 48.675 143.380 48.965 144.105 ;
        RECT 50.685 143.665 51.015 144.105 ;
        RECT 51.185 143.495 51.375 143.910 ;
        RECT 51.545 143.665 51.875 144.105 ;
        RECT 52.045 143.495 52.235 143.910 ;
        RECT 52.405 143.665 52.735 144.105 ;
        RECT 52.905 143.495 53.095 143.910 ;
        RECT 53.265 143.665 53.595 144.105 ;
        RECT 53.765 143.495 53.955 143.910 ;
        RECT 54.125 143.665 54.455 144.105 ;
        RECT 50.050 143.325 55.375 143.495 ;
        RECT 48.150 142.565 48.500 143.215 ;
        RECT 50.050 142.730 50.320 143.325 ;
        RECT 50.625 142.900 55.035 143.155 ;
        RECT 55.205 142.730 55.375 143.325 ;
        RECT 47.750 142.225 48.415 142.395 ;
        RECT 47.745 141.555 48.075 142.055 ;
        RECT 48.245 141.725 48.415 142.225 ;
        RECT 48.675 141.555 48.965 142.720 ;
        RECT 50.050 142.560 55.375 142.730 ;
        RECT 55.575 143.430 55.835 143.935 ;
        RECT 56.015 143.725 56.345 144.105 ;
        RECT 56.525 143.555 56.695 143.935 ;
        RECT 55.575 142.630 55.745 143.430 ;
        RECT 56.030 143.385 56.695 143.555 ;
        RECT 56.030 143.130 56.200 143.385 ;
        RECT 57.690 143.295 57.935 143.900 ;
        RECT 58.155 143.570 58.665 144.105 ;
        RECT 55.915 142.800 56.200 143.130 ;
        RECT 56.435 142.835 56.765 143.205 ;
        RECT 57.415 143.125 58.645 143.295 ;
        RECT 56.030 142.655 56.200 142.800 ;
        RECT 50.060 141.555 50.315 142.390 ;
        RECT 50.485 141.755 50.725 142.560 ;
        RECT 50.895 141.555 51.145 142.390 ;
        RECT 51.315 141.755 51.570 142.560 ;
        RECT 51.740 141.555 51.995 142.390 ;
        RECT 52.165 141.755 52.410 142.560 ;
        RECT 52.580 141.555 52.825 142.390 ;
        RECT 52.995 141.755 53.245 142.560 ;
        RECT 53.415 141.555 53.675 142.390 ;
        RECT 53.845 141.755 54.085 142.560 ;
        RECT 54.255 141.555 54.515 142.390 ;
        RECT 54.685 141.755 54.925 142.560 ;
        RECT 55.095 141.555 55.355 142.390 ;
        RECT 55.575 141.725 55.845 142.630 ;
        RECT 56.030 142.485 56.695 142.655 ;
        RECT 56.015 141.555 56.345 142.315 ;
        RECT 56.525 141.725 56.695 142.485 ;
        RECT 57.415 142.315 57.755 143.125 ;
        RECT 57.925 142.560 58.675 142.750 ;
        RECT 57.415 141.905 57.930 142.315 ;
        RECT 58.165 141.555 58.335 142.315 ;
        RECT 58.505 141.895 58.675 142.560 ;
        RECT 58.845 142.575 59.035 143.935 ;
        RECT 59.205 143.085 59.480 143.935 ;
        RECT 59.670 143.570 60.200 143.935 ;
        RECT 60.625 143.705 60.955 144.105 ;
        RECT 60.025 143.535 60.200 143.570 ;
        RECT 59.205 142.915 59.485 143.085 ;
        RECT 59.205 142.775 59.480 142.915 ;
        RECT 59.685 142.575 59.855 143.375 ;
        RECT 58.845 142.405 59.855 142.575 ;
        RECT 60.025 143.365 60.955 143.535 ;
        RECT 61.125 143.365 61.380 143.935 ;
        RECT 60.025 142.235 60.195 143.365 ;
        RECT 60.785 143.195 60.955 143.365 ;
        RECT 59.070 142.065 60.195 142.235 ;
        RECT 60.365 142.865 60.560 143.195 ;
        RECT 60.785 142.865 61.040 143.195 ;
        RECT 60.365 141.895 60.535 142.865 ;
        RECT 61.210 142.695 61.380 143.365 ;
        RECT 61.555 143.355 62.765 144.105 ;
        RECT 63.310 143.765 63.565 143.925 ;
        RECT 63.225 143.595 63.565 143.765 ;
        RECT 63.745 143.645 64.030 144.105 ;
        RECT 58.505 141.725 60.535 141.895 ;
        RECT 60.705 141.555 60.875 142.695 ;
        RECT 61.045 141.725 61.380 142.695 ;
        RECT 61.555 142.645 62.075 143.185 ;
        RECT 62.245 142.815 62.765 143.355 ;
        RECT 63.310 143.395 63.565 143.595 ;
        RECT 61.555 141.555 62.765 142.645 ;
        RECT 63.310 142.535 63.490 143.395 ;
        RECT 64.210 143.195 64.460 143.845 ;
        RECT 63.660 142.865 64.460 143.195 ;
        RECT 63.310 141.865 63.565 142.535 ;
        RECT 63.745 141.555 64.030 142.355 ;
        RECT 64.210 142.275 64.460 142.865 ;
        RECT 64.660 143.510 64.980 143.840 ;
        RECT 65.160 143.625 65.820 144.105 ;
        RECT 66.020 143.715 66.870 143.885 ;
        RECT 64.660 142.615 64.850 143.510 ;
        RECT 65.170 143.185 65.830 143.455 ;
        RECT 65.500 143.125 65.830 143.185 ;
        RECT 65.020 142.955 65.350 143.015 ;
        RECT 66.020 142.955 66.190 143.715 ;
        RECT 67.430 143.645 67.750 144.105 ;
        RECT 67.950 143.465 68.200 143.895 ;
        RECT 68.490 143.665 68.900 144.105 ;
        RECT 69.070 143.725 70.085 143.925 ;
        RECT 66.360 143.295 67.610 143.465 ;
        RECT 66.360 143.175 66.690 143.295 ;
        RECT 65.020 142.785 66.920 142.955 ;
        RECT 64.660 142.445 66.580 142.615 ;
        RECT 64.660 142.425 64.980 142.445 ;
        RECT 64.210 141.765 64.540 142.275 ;
        RECT 64.810 141.815 64.980 142.425 ;
        RECT 66.750 142.275 66.920 142.785 ;
        RECT 67.090 142.715 67.270 143.125 ;
        RECT 67.440 142.535 67.610 143.295 ;
        RECT 65.150 141.555 65.480 142.245 ;
        RECT 65.710 142.105 66.920 142.275 ;
        RECT 67.090 142.225 67.610 142.535 ;
        RECT 67.780 143.125 68.200 143.465 ;
        RECT 68.490 143.125 68.900 143.455 ;
        RECT 67.780 142.355 67.970 143.125 ;
        RECT 69.070 142.995 69.240 143.725 ;
        RECT 70.385 143.555 70.555 143.885 ;
        RECT 70.725 143.725 71.055 144.105 ;
        RECT 69.410 143.175 69.760 143.545 ;
        RECT 69.070 142.955 69.490 142.995 ;
        RECT 68.140 142.785 69.490 142.955 ;
        RECT 68.140 142.625 68.390 142.785 ;
        RECT 68.900 142.355 69.150 142.615 ;
        RECT 67.780 142.105 69.150 142.355 ;
        RECT 65.710 141.815 65.950 142.105 ;
        RECT 66.750 142.025 66.920 142.105 ;
        RECT 66.150 141.555 66.570 141.935 ;
        RECT 66.750 141.775 67.380 142.025 ;
        RECT 67.850 141.555 68.180 141.935 ;
        RECT 68.350 141.815 68.520 142.105 ;
        RECT 69.320 141.940 69.490 142.785 ;
        RECT 69.940 142.615 70.160 143.485 ;
        RECT 70.385 143.365 71.080 143.555 ;
        RECT 69.660 142.235 70.160 142.615 ;
        RECT 70.330 142.565 70.740 143.185 ;
        RECT 70.910 142.395 71.080 143.365 ;
        RECT 70.385 142.225 71.080 142.395 ;
        RECT 68.700 141.555 69.080 141.935 ;
        RECT 69.320 141.770 70.150 141.940 ;
        RECT 70.385 141.725 70.555 142.225 ;
        RECT 70.725 141.555 71.055 142.055 ;
        RECT 71.270 141.725 71.495 143.845 ;
        RECT 71.665 143.725 71.995 144.105 ;
        RECT 72.165 143.555 72.335 143.845 ;
        RECT 71.670 143.385 72.335 143.555 ;
        RECT 72.595 143.430 72.855 143.935 ;
        RECT 73.035 143.725 73.365 144.105 ;
        RECT 73.545 143.555 73.715 143.935 ;
        RECT 71.670 142.395 71.900 143.385 ;
        RECT 72.070 142.565 72.420 143.215 ;
        RECT 72.595 142.630 72.765 143.430 ;
        RECT 73.050 143.385 73.715 143.555 ;
        RECT 73.050 143.130 73.220 143.385 ;
        RECT 74.435 143.380 74.725 144.105 ;
        RECT 74.995 143.640 75.245 144.105 ;
        RECT 75.415 143.465 75.585 143.935 ;
        RECT 75.835 143.645 76.005 144.105 ;
        RECT 76.255 143.465 76.425 143.935 ;
        RECT 76.675 143.645 76.845 144.105 ;
        RECT 77.095 143.465 77.265 143.935 ;
        RECT 77.635 143.645 77.900 144.105 ;
        RECT 74.895 143.285 77.265 143.465 ;
        RECT 78.390 143.295 78.635 143.900 ;
        RECT 78.855 143.570 79.365 144.105 ;
        RECT 72.935 142.800 73.220 143.130 ;
        RECT 73.455 142.835 73.785 143.205 ;
        RECT 73.050 142.655 73.220 142.800 ;
        RECT 71.670 142.225 72.335 142.395 ;
        RECT 71.665 141.555 71.995 142.055 ;
        RECT 72.165 141.725 72.335 142.225 ;
        RECT 72.595 141.725 72.865 142.630 ;
        RECT 73.050 142.485 73.715 142.655 ;
        RECT 73.035 141.555 73.365 142.315 ;
        RECT 73.545 141.725 73.715 142.485 ;
        RECT 74.435 141.555 74.725 142.720 ;
        RECT 74.895 142.695 75.245 143.285 ;
        RECT 78.115 143.125 79.345 143.295 ;
        RECT 75.415 142.865 77.925 143.115 ;
        RECT 74.895 142.525 77.345 142.695 ;
        RECT 74.895 142.505 75.665 142.525 ;
        RECT 74.995 141.555 75.165 142.015 ;
        RECT 75.335 141.725 75.665 142.505 ;
        RECT 75.835 141.555 76.005 142.355 ;
        RECT 76.175 141.725 76.505 142.525 ;
        RECT 76.675 141.555 76.845 142.355 ;
        RECT 77.015 141.725 77.345 142.525 ;
        RECT 77.605 141.555 77.900 142.695 ;
        RECT 78.115 142.315 78.455 143.125 ;
        RECT 78.625 142.560 79.375 142.750 ;
        RECT 78.115 141.905 78.630 142.315 ;
        RECT 78.865 141.555 79.035 142.315 ;
        RECT 79.205 141.895 79.375 142.560 ;
        RECT 79.545 142.575 79.735 143.935 ;
        RECT 79.905 143.765 80.180 143.935 ;
        RECT 79.905 143.595 80.185 143.765 ;
        RECT 79.905 142.775 80.180 143.595 ;
        RECT 80.370 143.570 80.900 143.935 ;
        RECT 81.325 143.705 81.655 144.105 ;
        RECT 80.725 143.535 80.900 143.570 ;
        RECT 80.385 142.575 80.555 143.375 ;
        RECT 79.545 142.405 80.555 142.575 ;
        RECT 80.725 143.365 81.655 143.535 ;
        RECT 81.825 143.365 82.080 143.935 ;
        RECT 80.725 142.235 80.895 143.365 ;
        RECT 81.485 143.195 81.655 143.365 ;
        RECT 79.770 142.065 80.895 142.235 ;
        RECT 81.065 142.865 81.260 143.195 ;
        RECT 81.485 142.865 81.740 143.195 ;
        RECT 81.065 141.895 81.235 142.865 ;
        RECT 81.910 142.695 82.080 143.365 ;
        RECT 79.205 141.725 81.235 141.895 ;
        RECT 81.405 141.555 81.575 142.695 ;
        RECT 81.745 141.725 82.080 142.695 ;
        RECT 82.255 143.645 82.815 143.935 ;
        RECT 82.985 143.645 83.235 144.105 ;
        RECT 82.255 142.275 82.505 143.645 ;
        RECT 83.855 143.475 84.185 143.835 ;
        RECT 84.645 143.625 84.945 144.105 ;
        RECT 82.795 143.285 84.185 143.475 ;
        RECT 85.115 143.455 85.375 143.910 ;
        RECT 85.545 143.625 85.805 144.105 ;
        RECT 85.985 143.455 86.245 143.910 ;
        RECT 86.415 143.625 86.665 144.105 ;
        RECT 86.845 143.455 87.105 143.910 ;
        RECT 87.275 143.625 87.525 144.105 ;
        RECT 87.705 143.455 87.965 143.910 ;
        RECT 88.135 143.625 88.380 144.105 ;
        RECT 88.550 143.455 88.825 143.910 ;
        RECT 88.995 143.625 89.240 144.105 ;
        RECT 89.410 143.455 89.670 143.910 ;
        RECT 89.840 143.625 90.100 144.105 ;
        RECT 90.270 143.455 90.530 143.910 ;
        RECT 90.700 143.625 90.960 144.105 ;
        RECT 91.130 143.455 91.390 143.910 ;
        RECT 91.560 143.545 91.820 144.105 ;
        RECT 84.645 143.285 91.390 143.455 ;
        RECT 82.795 143.195 82.965 143.285 ;
        RECT 82.675 142.865 82.965 143.195 ;
        RECT 83.135 142.865 83.475 143.115 ;
        RECT 83.695 142.865 84.370 143.115 ;
        RECT 82.795 142.615 82.965 142.865 ;
        RECT 82.795 142.445 83.735 142.615 ;
        RECT 84.105 142.505 84.370 142.865 ;
        RECT 84.645 142.695 85.810 143.285 ;
        RECT 91.990 143.115 92.240 143.925 ;
        RECT 92.420 143.580 92.680 144.105 ;
        RECT 92.850 143.115 93.100 143.925 ;
        RECT 93.280 143.595 93.585 144.105 ;
        RECT 93.845 143.555 94.015 143.935 ;
        RECT 94.195 143.725 94.525 144.105 ;
        RECT 85.980 142.865 93.100 143.115 ;
        RECT 93.270 142.865 93.585 143.425 ;
        RECT 93.845 143.385 94.510 143.555 ;
        RECT 94.705 143.430 94.965 143.935 ;
        RECT 84.645 142.470 91.390 142.695 ;
        RECT 82.255 141.725 82.715 142.275 ;
        RECT 82.905 141.555 83.235 142.275 ;
        RECT 83.435 141.895 83.735 142.445 ;
        RECT 83.905 141.555 84.185 142.225 ;
        RECT 84.645 141.555 84.915 142.300 ;
        RECT 85.085 141.730 85.375 142.470 ;
        RECT 85.985 142.455 91.390 142.470 ;
        RECT 85.545 141.560 85.800 142.285 ;
        RECT 85.985 141.730 86.245 142.455 ;
        RECT 86.415 141.560 86.660 142.285 ;
        RECT 86.845 141.730 87.105 142.455 ;
        RECT 87.275 141.560 87.520 142.285 ;
        RECT 87.705 141.730 87.965 142.455 ;
        RECT 88.135 141.560 88.380 142.285 ;
        RECT 88.550 141.730 88.810 142.455 ;
        RECT 88.980 141.560 89.240 142.285 ;
        RECT 89.410 141.730 89.670 142.455 ;
        RECT 89.840 141.560 90.100 142.285 ;
        RECT 90.270 141.730 90.530 142.455 ;
        RECT 90.700 141.560 90.960 142.285 ;
        RECT 91.130 141.730 91.390 142.455 ;
        RECT 91.560 141.560 91.820 142.355 ;
        RECT 91.990 141.730 92.240 142.865 ;
        RECT 85.545 141.555 91.820 141.560 ;
        RECT 92.420 141.555 92.680 142.365 ;
        RECT 92.855 141.725 93.100 142.865 ;
        RECT 93.775 142.835 94.105 143.205 ;
        RECT 94.340 143.130 94.510 143.385 ;
        RECT 94.340 142.800 94.625 143.130 ;
        RECT 94.340 142.655 94.510 142.800 ;
        RECT 93.845 142.485 94.510 142.655 ;
        RECT 94.795 142.630 94.965 143.430 ;
        RECT 96.330 143.295 96.575 143.900 ;
        RECT 96.795 143.570 97.305 144.105 ;
        RECT 93.280 141.555 93.575 142.365 ;
        RECT 93.845 141.725 94.015 142.485 ;
        RECT 94.195 141.555 94.525 142.315 ;
        RECT 94.695 141.725 94.965 142.630 ;
        RECT 96.055 143.125 97.285 143.295 ;
        RECT 96.055 142.315 96.395 143.125 ;
        RECT 96.565 142.560 97.315 142.750 ;
        RECT 96.055 141.905 96.570 142.315 ;
        RECT 96.805 141.555 96.975 142.315 ;
        RECT 97.145 141.895 97.315 142.560 ;
        RECT 97.485 142.575 97.675 143.935 ;
        RECT 97.845 143.085 98.120 143.935 ;
        RECT 98.310 143.570 98.840 143.935 ;
        RECT 99.265 143.705 99.595 144.105 ;
        RECT 98.665 143.535 98.840 143.570 ;
        RECT 97.845 142.915 98.125 143.085 ;
        RECT 97.845 142.775 98.120 142.915 ;
        RECT 98.325 142.575 98.495 143.375 ;
        RECT 97.485 142.405 98.495 142.575 ;
        RECT 98.665 143.365 99.595 143.535 ;
        RECT 99.765 143.365 100.020 143.935 ;
        RECT 100.195 143.380 100.485 144.105 ;
        RECT 100.655 143.430 100.915 143.935 ;
        RECT 101.095 143.725 101.425 144.105 ;
        RECT 101.605 143.555 101.775 143.935 ;
        RECT 98.665 142.235 98.835 143.365 ;
        RECT 99.425 143.195 99.595 143.365 ;
        RECT 97.710 142.065 98.835 142.235 ;
        RECT 99.005 142.865 99.200 143.195 ;
        RECT 99.425 142.865 99.680 143.195 ;
        RECT 99.005 141.895 99.175 142.865 ;
        RECT 99.850 142.695 100.020 143.365 ;
        RECT 97.145 141.725 99.175 141.895 ;
        RECT 99.345 141.555 99.515 142.695 ;
        RECT 99.685 141.725 100.020 142.695 ;
        RECT 100.195 141.555 100.485 142.720 ;
        RECT 100.655 142.630 100.825 143.430 ;
        RECT 101.110 143.385 101.775 143.555 ;
        RECT 102.410 143.425 102.665 143.925 ;
        RECT 102.845 143.645 103.130 144.105 ;
        RECT 102.325 143.395 102.665 143.425 ;
        RECT 101.110 143.130 101.280 143.385 ;
        RECT 102.325 143.255 102.590 143.395 ;
        RECT 100.995 142.800 101.280 143.130 ;
        RECT 101.515 142.835 101.845 143.205 ;
        RECT 101.110 142.655 101.280 142.800 ;
        RECT 100.655 141.725 100.925 142.630 ;
        RECT 101.110 142.485 101.775 142.655 ;
        RECT 101.095 141.555 101.425 142.315 ;
        RECT 101.605 141.725 101.775 142.485 ;
        RECT 102.410 142.535 102.590 143.255 ;
        RECT 103.310 143.195 103.560 143.845 ;
        RECT 102.760 142.865 103.560 143.195 ;
        RECT 102.410 141.865 102.665 142.535 ;
        RECT 102.845 141.555 103.130 142.355 ;
        RECT 103.310 142.275 103.560 142.865 ;
        RECT 103.760 143.510 104.080 143.840 ;
        RECT 104.260 143.625 104.920 144.105 ;
        RECT 105.120 143.715 105.970 143.885 ;
        RECT 103.760 142.615 103.950 143.510 ;
        RECT 104.270 143.185 104.930 143.455 ;
        RECT 104.600 143.125 104.930 143.185 ;
        RECT 104.120 142.955 104.450 143.015 ;
        RECT 105.120 142.955 105.290 143.715 ;
        RECT 106.530 143.645 106.850 144.105 ;
        RECT 107.050 143.465 107.300 143.895 ;
        RECT 107.590 143.665 108.000 144.105 ;
        RECT 108.170 143.725 109.185 143.925 ;
        RECT 105.460 143.295 106.710 143.465 ;
        RECT 105.460 143.175 105.790 143.295 ;
        RECT 104.120 142.785 106.020 142.955 ;
        RECT 103.760 142.445 105.680 142.615 ;
        RECT 103.760 142.425 104.080 142.445 ;
        RECT 103.310 141.765 103.640 142.275 ;
        RECT 103.910 141.815 104.080 142.425 ;
        RECT 105.850 142.275 106.020 142.785 ;
        RECT 106.190 142.715 106.370 143.125 ;
        RECT 106.540 142.535 106.710 143.295 ;
        RECT 104.250 141.555 104.580 142.245 ;
        RECT 104.810 142.105 106.020 142.275 ;
        RECT 106.190 142.225 106.710 142.535 ;
        RECT 106.880 143.125 107.300 143.465 ;
        RECT 107.590 143.125 108.000 143.455 ;
        RECT 106.880 142.355 107.070 143.125 ;
        RECT 108.170 142.995 108.340 143.725 ;
        RECT 109.485 143.555 109.655 143.885 ;
        RECT 109.825 143.725 110.155 144.105 ;
        RECT 108.510 143.175 108.860 143.545 ;
        RECT 108.170 142.955 108.590 142.995 ;
        RECT 107.240 142.785 108.590 142.955 ;
        RECT 107.240 142.625 107.490 142.785 ;
        RECT 108.000 142.355 108.250 142.615 ;
        RECT 106.880 142.105 108.250 142.355 ;
        RECT 104.810 141.815 105.050 142.105 ;
        RECT 105.850 142.025 106.020 142.105 ;
        RECT 105.250 141.555 105.670 141.935 ;
        RECT 105.850 141.775 106.480 142.025 ;
        RECT 106.950 141.555 107.280 141.935 ;
        RECT 107.450 141.815 107.620 142.105 ;
        RECT 108.420 141.940 108.590 142.785 ;
        RECT 109.040 142.615 109.260 143.485 ;
        RECT 109.485 143.365 110.180 143.555 ;
        RECT 108.760 142.235 109.260 142.615 ;
        RECT 109.430 142.565 109.840 143.185 ;
        RECT 110.010 142.395 110.180 143.365 ;
        RECT 109.485 142.225 110.180 142.395 ;
        RECT 107.800 141.555 108.180 141.935 ;
        RECT 108.420 141.770 109.250 141.940 ;
        RECT 109.485 141.725 109.655 142.225 ;
        RECT 109.825 141.555 110.155 142.055 ;
        RECT 110.370 141.725 110.595 143.845 ;
        RECT 110.765 143.725 111.095 144.105 ;
        RECT 111.265 143.555 111.435 143.845 ;
        RECT 110.770 143.385 111.435 143.555 ;
        RECT 110.770 142.395 111.000 143.385 ;
        RECT 112.155 143.355 113.365 144.105 ;
        RECT 111.170 142.565 111.520 143.215 ;
        RECT 112.155 142.645 112.675 143.185 ;
        RECT 112.845 142.815 113.365 143.355 ;
        RECT 110.770 142.225 111.435 142.395 ;
        RECT 110.765 141.555 111.095 142.055 ;
        RECT 111.265 141.725 111.435 142.225 ;
        RECT 112.155 141.555 113.365 142.645 ;
        RECT 26.970 141.385 113.450 141.555 ;
        RECT 27.055 140.295 28.265 141.385 ;
        RECT 29.555 140.715 29.835 141.385 ;
        RECT 30.005 140.495 30.305 141.045 ;
        RECT 30.505 140.665 30.835 141.385 ;
        RECT 31.025 140.665 31.485 141.215 ;
        RECT 27.055 139.585 27.575 140.125 ;
        RECT 27.745 139.755 28.265 140.295 ;
        RECT 29.370 140.075 29.635 140.435 ;
        RECT 30.005 140.325 30.945 140.495 ;
        RECT 30.775 140.075 30.945 140.325 ;
        RECT 29.370 139.825 30.045 140.075 ;
        RECT 30.265 139.825 30.605 140.075 ;
        RECT 30.775 139.745 31.065 140.075 ;
        RECT 30.775 139.655 30.945 139.745 ;
        RECT 27.055 138.835 28.265 139.585 ;
        RECT 29.555 139.465 30.945 139.655 ;
        RECT 29.555 139.105 29.885 139.465 ;
        RECT 31.235 139.295 31.485 140.665 ;
        RECT 30.505 138.835 30.755 139.295 ;
        RECT 30.925 139.005 31.485 139.295 ;
        RECT 31.660 140.245 31.995 141.215 ;
        RECT 32.165 140.245 32.335 141.385 ;
        RECT 32.505 141.045 34.535 141.215 ;
        RECT 31.660 139.575 31.830 140.245 ;
        RECT 32.505 140.075 32.675 141.045 ;
        RECT 32.000 139.745 32.255 140.075 ;
        RECT 32.480 139.745 32.675 140.075 ;
        RECT 32.845 140.705 33.970 140.875 ;
        RECT 32.085 139.575 32.255 139.745 ;
        RECT 32.845 139.575 33.015 140.705 ;
        RECT 31.660 139.005 31.915 139.575 ;
        RECT 32.085 139.405 33.015 139.575 ;
        RECT 33.185 140.365 34.195 140.535 ;
        RECT 33.185 139.565 33.355 140.365 ;
        RECT 33.560 140.025 33.835 140.165 ;
        RECT 33.555 139.855 33.835 140.025 ;
        RECT 32.840 139.370 33.015 139.405 ;
        RECT 32.085 138.835 32.415 139.235 ;
        RECT 32.840 139.005 33.370 139.370 ;
        RECT 33.560 139.005 33.835 139.855 ;
        RECT 34.005 139.005 34.195 140.365 ;
        RECT 34.365 140.380 34.535 141.045 ;
        RECT 34.705 140.625 34.875 141.385 ;
        RECT 35.110 140.625 35.625 141.035 ;
        RECT 34.365 140.190 35.115 140.380 ;
        RECT 35.285 139.815 35.625 140.625 ;
        RECT 35.795 140.220 36.085 141.385 ;
        RECT 36.355 140.925 36.525 141.385 ;
        RECT 36.695 140.435 37.025 141.215 ;
        RECT 37.195 140.585 37.365 141.385 ;
        RECT 36.255 140.415 37.025 140.435 ;
        RECT 37.535 140.415 37.865 141.215 ;
        RECT 38.035 140.585 38.205 141.385 ;
        RECT 38.375 140.415 38.705 141.215 ;
        RECT 36.255 140.245 38.705 140.415 ;
        RECT 38.965 140.245 39.260 141.385 ;
        RECT 39.850 141.045 40.105 141.075 ;
        RECT 39.765 140.875 40.105 141.045 ;
        RECT 39.850 140.405 40.105 140.875 ;
        RECT 40.285 140.585 40.570 141.385 ;
        RECT 40.750 140.665 41.080 141.175 ;
        RECT 34.395 139.645 35.625 139.815 ;
        RECT 36.255 139.655 36.605 140.245 ;
        RECT 36.775 139.825 39.285 140.075 ;
        RECT 34.375 138.835 34.885 139.370 ;
        RECT 35.105 139.040 35.350 139.645 ;
        RECT 35.795 138.835 36.085 139.560 ;
        RECT 36.255 139.475 38.625 139.655 ;
        RECT 36.355 138.835 36.605 139.300 ;
        RECT 36.775 139.005 36.945 139.475 ;
        RECT 37.195 138.835 37.365 139.295 ;
        RECT 37.615 139.005 37.785 139.475 ;
        RECT 38.035 138.835 38.205 139.295 ;
        RECT 38.455 139.005 38.625 139.475 ;
        RECT 39.850 139.545 40.030 140.405 ;
        RECT 40.750 140.075 41.000 140.665 ;
        RECT 41.350 140.515 41.520 141.125 ;
        RECT 41.690 140.695 42.020 141.385 ;
        RECT 42.250 140.835 42.490 141.125 ;
        RECT 42.690 141.005 43.110 141.385 ;
        RECT 43.290 140.915 43.920 141.165 ;
        RECT 44.390 141.005 44.720 141.385 ;
        RECT 43.290 140.835 43.460 140.915 ;
        RECT 44.890 140.835 45.060 141.125 ;
        RECT 45.240 141.005 45.620 141.385 ;
        RECT 45.860 141.000 46.690 141.170 ;
        RECT 42.250 140.665 43.460 140.835 ;
        RECT 40.200 139.745 41.000 140.075 ;
        RECT 38.995 138.835 39.260 139.295 ;
        RECT 39.850 139.015 40.105 139.545 ;
        RECT 40.285 138.835 40.570 139.295 ;
        RECT 40.750 139.095 41.000 139.745 ;
        RECT 41.200 140.495 41.520 140.515 ;
        RECT 41.200 140.325 43.120 140.495 ;
        RECT 41.200 139.430 41.390 140.325 ;
        RECT 43.290 140.155 43.460 140.665 ;
        RECT 43.630 140.405 44.150 140.715 ;
        RECT 41.560 139.985 43.460 140.155 ;
        RECT 41.560 139.925 41.890 139.985 ;
        RECT 42.040 139.755 42.370 139.815 ;
        RECT 41.710 139.485 42.370 139.755 ;
        RECT 41.200 139.100 41.520 139.430 ;
        RECT 41.700 138.835 42.360 139.315 ;
        RECT 42.560 139.225 42.730 139.985 ;
        RECT 43.630 139.815 43.810 140.225 ;
        RECT 42.900 139.645 43.230 139.765 ;
        RECT 43.980 139.645 44.150 140.405 ;
        RECT 42.900 139.475 44.150 139.645 ;
        RECT 44.320 140.585 45.690 140.835 ;
        RECT 44.320 139.815 44.510 140.585 ;
        RECT 45.440 140.325 45.690 140.585 ;
        RECT 44.680 140.155 44.930 140.315 ;
        RECT 45.860 140.155 46.030 141.000 ;
        RECT 46.925 140.715 47.095 141.215 ;
        RECT 47.265 140.885 47.595 141.385 ;
        RECT 46.200 140.325 46.700 140.705 ;
        RECT 46.925 140.545 47.620 140.715 ;
        RECT 44.680 139.985 46.030 140.155 ;
        RECT 45.610 139.945 46.030 139.985 ;
        RECT 44.320 139.475 44.740 139.815 ;
        RECT 45.030 139.485 45.440 139.815 ;
        RECT 42.560 139.055 43.410 139.225 ;
        RECT 43.970 138.835 44.290 139.295 ;
        RECT 44.490 139.045 44.740 139.475 ;
        RECT 45.030 138.835 45.440 139.275 ;
        RECT 45.610 139.215 45.780 139.945 ;
        RECT 45.950 139.395 46.300 139.765 ;
        RECT 46.480 139.455 46.700 140.325 ;
        RECT 46.870 139.755 47.280 140.375 ;
        RECT 47.450 139.575 47.620 140.545 ;
        RECT 46.925 139.385 47.620 139.575 ;
        RECT 45.610 139.015 46.625 139.215 ;
        RECT 46.925 139.055 47.095 139.385 ;
        RECT 47.265 138.835 47.595 139.215 ;
        RECT 47.810 139.095 48.035 141.215 ;
        RECT 48.205 140.885 48.535 141.385 ;
        RECT 48.705 140.715 48.875 141.215 ;
        RECT 48.210 140.545 48.875 140.715 ;
        RECT 49.145 140.575 49.440 141.385 ;
        RECT 48.210 139.555 48.440 140.545 ;
        RECT 48.610 139.725 48.960 140.375 ;
        RECT 49.620 140.075 49.865 141.215 ;
        RECT 50.040 140.575 50.300 141.385 ;
        RECT 50.900 141.380 57.175 141.385 ;
        RECT 50.480 140.075 50.730 141.210 ;
        RECT 50.900 140.585 51.160 141.380 ;
        RECT 51.330 140.485 51.590 141.210 ;
        RECT 51.760 140.655 52.020 141.380 ;
        RECT 52.190 140.485 52.450 141.210 ;
        RECT 52.620 140.655 52.880 141.380 ;
        RECT 53.050 140.485 53.310 141.210 ;
        RECT 53.480 140.655 53.740 141.380 ;
        RECT 53.910 140.485 54.170 141.210 ;
        RECT 54.340 140.655 54.585 141.380 ;
        RECT 54.755 140.485 55.015 141.210 ;
        RECT 55.200 140.655 55.445 141.380 ;
        RECT 55.615 140.485 55.875 141.210 ;
        RECT 56.060 140.655 56.305 141.380 ;
        RECT 56.475 140.485 56.735 141.210 ;
        RECT 56.920 140.655 57.175 141.380 ;
        RECT 51.330 140.470 56.735 140.485 ;
        RECT 57.345 140.470 57.635 141.210 ;
        RECT 57.805 140.640 58.075 141.385 ;
        RECT 58.340 140.875 59.995 141.165 ;
        RECT 58.340 140.535 59.930 140.705 ;
        RECT 60.165 140.585 60.445 141.385 ;
        RECT 51.330 140.245 58.075 140.470 ;
        RECT 58.340 140.245 58.660 140.535 ;
        RECT 59.760 140.415 59.930 140.535 ;
        RECT 48.210 139.385 48.875 139.555 ;
        RECT 49.135 139.515 49.450 140.075 ;
        RECT 49.620 139.825 56.740 140.075 ;
        RECT 48.205 138.835 48.535 139.215 ;
        RECT 48.705 139.095 48.875 139.385 ;
        RECT 49.135 138.835 49.440 139.345 ;
        RECT 49.620 139.015 49.870 139.825 ;
        RECT 50.040 138.835 50.300 139.360 ;
        RECT 50.480 139.015 50.730 139.825 ;
        RECT 56.910 139.655 58.075 140.245 ;
        RECT 58.855 140.195 59.570 140.365 ;
        RECT 59.760 140.245 60.485 140.415 ;
        RECT 60.655 140.245 60.925 141.215 ;
        RECT 51.330 139.485 58.075 139.655 ;
        RECT 58.340 139.505 58.690 140.075 ;
        RECT 58.860 139.745 59.570 140.195 ;
        RECT 60.315 140.075 60.485 140.245 ;
        RECT 59.740 139.745 60.145 140.075 ;
        RECT 60.315 139.745 60.585 140.075 ;
        RECT 60.315 139.575 60.485 139.745 ;
        RECT 50.900 138.835 51.160 139.395 ;
        RECT 51.330 139.030 51.590 139.485 ;
        RECT 51.760 138.835 52.020 139.315 ;
        RECT 52.190 139.030 52.450 139.485 ;
        RECT 52.620 138.835 52.880 139.315 ;
        RECT 53.050 139.030 53.310 139.485 ;
        RECT 53.480 138.835 53.725 139.315 ;
        RECT 53.895 139.030 54.170 139.485 ;
        RECT 54.340 138.835 54.585 139.315 ;
        RECT 54.755 139.030 55.015 139.485 ;
        RECT 55.195 138.835 55.445 139.315 ;
        RECT 55.615 139.030 55.875 139.485 ;
        RECT 56.055 138.835 56.305 139.315 ;
        RECT 56.475 139.030 56.735 139.485 ;
        RECT 56.915 138.835 57.175 139.315 ;
        RECT 57.345 139.030 57.605 139.485 ;
        RECT 58.875 139.405 60.485 139.575 ;
        RECT 60.755 139.510 60.925 140.245 ;
        RECT 61.555 140.220 61.845 141.385 ;
        RECT 62.055 140.245 62.285 141.385 ;
        RECT 62.455 140.235 62.785 141.215 ;
        RECT 62.955 140.245 63.165 141.385 ;
        RECT 63.395 140.625 63.910 141.035 ;
        RECT 64.145 140.625 64.315 141.385 ;
        RECT 64.485 141.045 66.515 141.215 ;
        RECT 62.035 139.825 62.365 140.075 ;
        RECT 57.775 138.835 58.075 139.315 ;
        RECT 58.345 138.835 58.675 139.335 ;
        RECT 58.875 139.055 59.045 139.405 ;
        RECT 59.245 138.835 59.575 139.235 ;
        RECT 59.745 139.055 59.915 139.405 ;
        RECT 60.085 138.835 60.465 139.235 ;
        RECT 60.655 139.165 60.925 139.510 ;
        RECT 61.555 138.835 61.845 139.560 ;
        RECT 62.055 138.835 62.285 139.655 ;
        RECT 62.535 139.635 62.785 140.235 ;
        RECT 63.395 139.815 63.735 140.625 ;
        RECT 64.485 140.380 64.655 141.045 ;
        RECT 65.050 140.705 66.175 140.875 ;
        RECT 63.905 140.190 64.655 140.380 ;
        RECT 64.825 140.365 65.835 140.535 ;
        RECT 62.455 139.005 62.785 139.635 ;
        RECT 62.955 138.835 63.165 139.655 ;
        RECT 63.395 139.645 64.625 139.815 ;
        RECT 63.670 139.040 63.915 139.645 ;
        RECT 64.135 138.835 64.645 139.370 ;
        RECT 64.825 139.005 65.015 140.365 ;
        RECT 65.185 140.025 65.460 140.165 ;
        RECT 65.185 139.855 65.465 140.025 ;
        RECT 65.185 139.005 65.460 139.855 ;
        RECT 65.665 139.565 65.835 140.365 ;
        RECT 66.005 139.575 66.175 140.705 ;
        RECT 66.345 140.075 66.515 141.045 ;
        RECT 66.685 140.245 66.855 141.385 ;
        RECT 67.025 140.245 67.360 141.215 ;
        RECT 68.465 140.575 68.760 141.385 ;
        RECT 66.345 139.745 66.540 140.075 ;
        RECT 66.765 139.745 67.020 140.075 ;
        RECT 66.765 139.575 66.935 139.745 ;
        RECT 67.190 139.575 67.360 140.245 ;
        RECT 68.940 140.075 69.185 141.215 ;
        RECT 69.360 140.575 69.620 141.385 ;
        RECT 70.220 141.380 76.495 141.385 ;
        RECT 69.800 140.075 70.050 141.210 ;
        RECT 70.220 140.585 70.480 141.380 ;
        RECT 70.650 140.485 70.910 141.210 ;
        RECT 71.080 140.655 71.340 141.380 ;
        RECT 71.510 140.485 71.770 141.210 ;
        RECT 71.940 140.655 72.200 141.380 ;
        RECT 72.370 140.485 72.630 141.210 ;
        RECT 72.800 140.655 73.060 141.380 ;
        RECT 73.230 140.485 73.490 141.210 ;
        RECT 73.660 140.655 73.905 141.380 ;
        RECT 74.075 140.485 74.335 141.210 ;
        RECT 74.520 140.655 74.765 141.380 ;
        RECT 74.935 140.485 75.195 141.210 ;
        RECT 75.380 140.655 75.625 141.380 ;
        RECT 75.795 140.485 76.055 141.210 ;
        RECT 76.240 140.655 76.495 141.380 ;
        RECT 70.650 140.470 76.055 140.485 ;
        RECT 76.665 140.470 76.955 141.210 ;
        RECT 77.125 140.640 77.395 141.385 ;
        RECT 70.650 140.245 77.395 140.470 ;
        RECT 78.030 140.405 78.285 141.075 ;
        RECT 78.465 140.585 78.750 141.385 ;
        RECT 78.930 140.665 79.260 141.175 ;
        RECT 78.030 140.365 78.210 140.405 ;
        RECT 66.005 139.405 66.935 139.575 ;
        RECT 66.005 139.370 66.180 139.405 ;
        RECT 65.650 139.005 66.180 139.370 ;
        RECT 66.605 138.835 66.935 139.235 ;
        RECT 67.105 139.005 67.360 139.575 ;
        RECT 68.455 139.515 68.770 140.075 ;
        RECT 68.940 139.825 76.060 140.075 ;
        RECT 68.455 138.835 68.760 139.345 ;
        RECT 68.940 139.015 69.190 139.825 ;
        RECT 69.360 138.835 69.620 139.360 ;
        RECT 69.800 139.015 70.050 139.825 ;
        RECT 76.230 139.655 77.395 140.245 ;
        RECT 77.945 140.195 78.210 140.365 ;
        RECT 70.650 139.485 77.395 139.655 ;
        RECT 78.030 139.545 78.210 140.195 ;
        RECT 78.930 140.075 79.180 140.665 ;
        RECT 79.530 140.515 79.700 141.125 ;
        RECT 79.870 140.695 80.200 141.385 ;
        RECT 80.430 140.835 80.670 141.125 ;
        RECT 80.870 141.005 81.290 141.385 ;
        RECT 81.470 140.915 82.100 141.165 ;
        RECT 82.570 141.005 82.900 141.385 ;
        RECT 81.470 140.835 81.640 140.915 ;
        RECT 83.070 140.835 83.240 141.125 ;
        RECT 83.420 141.005 83.800 141.385 ;
        RECT 84.040 141.000 84.870 141.170 ;
        RECT 80.430 140.665 81.640 140.835 ;
        RECT 78.380 139.745 79.180 140.075 ;
        RECT 70.220 138.835 70.480 139.395 ;
        RECT 70.650 139.030 70.910 139.485 ;
        RECT 71.080 138.835 71.340 139.315 ;
        RECT 71.510 139.030 71.770 139.485 ;
        RECT 71.940 138.835 72.200 139.315 ;
        RECT 72.370 139.030 72.630 139.485 ;
        RECT 72.800 138.835 73.045 139.315 ;
        RECT 73.215 139.030 73.490 139.485 ;
        RECT 73.660 138.835 73.905 139.315 ;
        RECT 74.075 139.030 74.335 139.485 ;
        RECT 74.515 138.835 74.765 139.315 ;
        RECT 74.935 139.030 75.195 139.485 ;
        RECT 75.375 138.835 75.625 139.315 ;
        RECT 75.795 139.030 76.055 139.485 ;
        RECT 76.235 138.835 76.495 139.315 ;
        RECT 76.665 139.030 76.925 139.485 ;
        RECT 77.095 138.835 77.395 139.315 ;
        RECT 78.030 139.015 78.285 139.545 ;
        RECT 78.465 138.835 78.750 139.295 ;
        RECT 78.930 139.095 79.180 139.745 ;
        RECT 79.380 140.495 79.700 140.515 ;
        RECT 79.380 140.325 81.300 140.495 ;
        RECT 79.380 139.430 79.570 140.325 ;
        RECT 81.470 140.155 81.640 140.665 ;
        RECT 81.810 140.405 82.330 140.715 ;
        RECT 79.740 139.985 81.640 140.155 ;
        RECT 79.740 139.925 80.070 139.985 ;
        RECT 80.220 139.755 80.550 139.815 ;
        RECT 79.890 139.485 80.550 139.755 ;
        RECT 79.380 139.100 79.700 139.430 ;
        RECT 79.880 138.835 80.540 139.315 ;
        RECT 80.740 139.225 80.910 139.985 ;
        RECT 81.810 139.815 81.990 140.225 ;
        RECT 81.080 139.645 81.410 139.765 ;
        RECT 82.160 139.645 82.330 140.405 ;
        RECT 81.080 139.475 82.330 139.645 ;
        RECT 82.500 140.585 83.870 140.835 ;
        RECT 82.500 139.815 82.690 140.585 ;
        RECT 83.620 140.325 83.870 140.585 ;
        RECT 82.860 140.155 83.110 140.315 ;
        RECT 84.040 140.155 84.210 141.000 ;
        RECT 85.105 140.715 85.275 141.215 ;
        RECT 85.445 140.885 85.775 141.385 ;
        RECT 84.380 140.325 84.880 140.705 ;
        RECT 85.105 140.545 85.800 140.715 ;
        RECT 82.860 139.985 84.210 140.155 ;
        RECT 83.790 139.945 84.210 139.985 ;
        RECT 82.500 139.475 82.920 139.815 ;
        RECT 83.210 139.485 83.620 139.815 ;
        RECT 80.740 139.055 81.590 139.225 ;
        RECT 82.150 138.835 82.470 139.295 ;
        RECT 82.670 139.045 82.920 139.475 ;
        RECT 83.210 138.835 83.620 139.275 ;
        RECT 83.790 139.215 83.960 139.945 ;
        RECT 84.130 139.395 84.480 139.765 ;
        RECT 84.660 139.455 84.880 140.325 ;
        RECT 85.050 139.755 85.460 140.375 ;
        RECT 85.630 139.575 85.800 140.545 ;
        RECT 85.105 139.385 85.800 139.575 ;
        RECT 83.790 139.015 84.805 139.215 ;
        RECT 85.105 139.055 85.275 139.385 ;
        RECT 85.445 138.835 85.775 139.215 ;
        RECT 85.990 139.095 86.215 141.215 ;
        RECT 86.385 140.885 86.715 141.385 ;
        RECT 86.885 140.715 87.055 141.215 ;
        RECT 86.390 140.545 87.055 140.715 ;
        RECT 86.390 139.555 86.620 140.545 ;
        RECT 86.790 139.725 87.140 140.375 ;
        RECT 87.315 140.220 87.605 141.385 ;
        RECT 88.150 141.045 88.405 141.075 ;
        RECT 88.065 140.875 88.405 141.045 ;
        RECT 88.150 140.405 88.405 140.875 ;
        RECT 88.585 140.585 88.870 141.385 ;
        RECT 89.050 140.665 89.380 141.175 ;
        RECT 86.390 139.385 87.055 139.555 ;
        RECT 86.385 138.835 86.715 139.215 ;
        RECT 86.885 139.095 87.055 139.385 ;
        RECT 87.315 138.835 87.605 139.560 ;
        RECT 88.150 139.545 88.330 140.405 ;
        RECT 89.050 140.075 89.300 140.665 ;
        RECT 89.650 140.515 89.820 141.125 ;
        RECT 89.990 140.695 90.320 141.385 ;
        RECT 90.550 140.835 90.790 141.125 ;
        RECT 90.990 141.005 91.410 141.385 ;
        RECT 91.590 140.915 92.220 141.165 ;
        RECT 92.690 141.005 93.020 141.385 ;
        RECT 91.590 140.835 91.760 140.915 ;
        RECT 93.190 140.835 93.360 141.125 ;
        RECT 93.540 141.005 93.920 141.385 ;
        RECT 94.160 141.000 94.990 141.170 ;
        RECT 90.550 140.665 91.760 140.835 ;
        RECT 88.500 139.745 89.300 140.075 ;
        RECT 88.150 139.015 88.405 139.545 ;
        RECT 88.585 138.835 88.870 139.295 ;
        RECT 89.050 139.095 89.300 139.745 ;
        RECT 89.500 140.495 89.820 140.515 ;
        RECT 89.500 140.325 91.420 140.495 ;
        RECT 89.500 139.430 89.690 140.325 ;
        RECT 91.590 140.155 91.760 140.665 ;
        RECT 91.930 140.405 92.450 140.715 ;
        RECT 89.860 139.985 91.760 140.155 ;
        RECT 89.860 139.925 90.190 139.985 ;
        RECT 90.340 139.755 90.670 139.815 ;
        RECT 90.010 139.485 90.670 139.755 ;
        RECT 89.500 139.100 89.820 139.430 ;
        RECT 90.000 138.835 90.660 139.315 ;
        RECT 90.860 139.225 91.030 139.985 ;
        RECT 91.930 139.815 92.110 140.225 ;
        RECT 91.200 139.645 91.530 139.765 ;
        RECT 92.280 139.645 92.450 140.405 ;
        RECT 91.200 139.475 92.450 139.645 ;
        RECT 92.620 140.585 93.990 140.835 ;
        RECT 92.620 139.815 92.810 140.585 ;
        RECT 93.740 140.325 93.990 140.585 ;
        RECT 92.980 140.155 93.230 140.315 ;
        RECT 94.160 140.155 94.330 141.000 ;
        RECT 95.225 140.715 95.395 141.215 ;
        RECT 95.565 140.885 95.895 141.385 ;
        RECT 94.500 140.325 95.000 140.705 ;
        RECT 95.225 140.545 95.920 140.715 ;
        RECT 92.980 139.985 94.330 140.155 ;
        RECT 93.910 139.945 94.330 139.985 ;
        RECT 92.620 139.475 93.040 139.815 ;
        RECT 93.330 139.485 93.740 139.815 ;
        RECT 90.860 139.055 91.710 139.225 ;
        RECT 92.270 138.835 92.590 139.295 ;
        RECT 92.790 139.045 93.040 139.475 ;
        RECT 93.330 138.835 93.740 139.275 ;
        RECT 93.910 139.215 94.080 139.945 ;
        RECT 94.250 139.395 94.600 139.765 ;
        RECT 94.780 139.455 95.000 140.325 ;
        RECT 95.170 139.755 95.580 140.375 ;
        RECT 95.750 139.575 95.920 140.545 ;
        RECT 95.225 139.385 95.920 139.575 ;
        RECT 93.910 139.015 94.925 139.215 ;
        RECT 95.225 139.055 95.395 139.385 ;
        RECT 95.565 138.835 95.895 139.215 ;
        RECT 96.110 139.095 96.335 141.215 ;
        RECT 96.505 140.885 96.835 141.385 ;
        RECT 97.005 140.715 97.175 141.215 ;
        RECT 96.510 140.545 97.175 140.715 ;
        RECT 97.895 140.625 98.410 141.035 ;
        RECT 98.645 140.625 98.815 141.385 ;
        RECT 98.985 141.045 101.015 141.215 ;
        RECT 96.510 139.555 96.740 140.545 ;
        RECT 96.910 139.725 97.260 140.375 ;
        RECT 97.895 139.815 98.235 140.625 ;
        RECT 98.985 140.380 99.155 141.045 ;
        RECT 99.550 140.705 100.675 140.875 ;
        RECT 98.405 140.190 99.155 140.380 ;
        RECT 99.325 140.365 100.335 140.535 ;
        RECT 97.895 139.645 99.125 139.815 ;
        RECT 96.510 139.385 97.175 139.555 ;
        RECT 96.505 138.835 96.835 139.215 ;
        RECT 97.005 139.095 97.175 139.385 ;
        RECT 98.170 139.040 98.415 139.645 ;
        RECT 98.635 138.835 99.145 139.370 ;
        RECT 99.325 139.005 99.515 140.365 ;
        RECT 99.685 139.345 99.960 140.165 ;
        RECT 100.165 139.565 100.335 140.365 ;
        RECT 100.505 139.575 100.675 140.705 ;
        RECT 100.845 140.075 101.015 141.045 ;
        RECT 101.185 140.245 101.355 141.385 ;
        RECT 101.525 140.245 101.860 141.215 ;
        RECT 100.845 139.745 101.040 140.075 ;
        RECT 101.265 139.745 101.520 140.075 ;
        RECT 101.265 139.575 101.435 139.745 ;
        RECT 101.690 139.575 101.860 140.245 ;
        RECT 102.410 140.405 102.665 141.075 ;
        RECT 102.845 140.585 103.130 141.385 ;
        RECT 103.310 140.665 103.640 141.175 ;
        RECT 102.410 139.685 102.590 140.405 ;
        RECT 103.310 140.075 103.560 140.665 ;
        RECT 103.910 140.515 104.080 141.125 ;
        RECT 104.250 140.695 104.580 141.385 ;
        RECT 104.810 140.835 105.050 141.125 ;
        RECT 105.250 141.005 105.670 141.385 ;
        RECT 105.850 140.915 106.480 141.165 ;
        RECT 106.950 141.005 107.280 141.385 ;
        RECT 105.850 140.835 106.020 140.915 ;
        RECT 107.450 140.835 107.620 141.125 ;
        RECT 107.800 141.005 108.180 141.385 ;
        RECT 108.420 141.000 109.250 141.170 ;
        RECT 104.810 140.665 106.020 140.835 ;
        RECT 102.760 139.745 103.560 140.075 ;
        RECT 100.505 139.405 101.435 139.575 ;
        RECT 100.505 139.370 100.680 139.405 ;
        RECT 99.685 139.175 99.965 139.345 ;
        RECT 99.685 139.005 99.960 139.175 ;
        RECT 100.150 139.005 100.680 139.370 ;
        RECT 101.105 138.835 101.435 139.235 ;
        RECT 101.605 139.005 101.860 139.575 ;
        RECT 102.325 139.545 102.590 139.685 ;
        RECT 102.325 139.515 102.665 139.545 ;
        RECT 102.410 139.015 102.665 139.515 ;
        RECT 102.845 138.835 103.130 139.295 ;
        RECT 103.310 139.095 103.560 139.745 ;
        RECT 103.760 140.495 104.080 140.515 ;
        RECT 103.760 140.325 105.680 140.495 ;
        RECT 103.760 139.430 103.950 140.325 ;
        RECT 105.850 140.155 106.020 140.665 ;
        RECT 106.190 140.405 106.710 140.715 ;
        RECT 104.120 139.985 106.020 140.155 ;
        RECT 104.120 139.925 104.450 139.985 ;
        RECT 104.600 139.755 104.930 139.815 ;
        RECT 104.270 139.485 104.930 139.755 ;
        RECT 103.760 139.100 104.080 139.430 ;
        RECT 104.260 138.835 104.920 139.315 ;
        RECT 105.120 139.225 105.290 139.985 ;
        RECT 106.190 139.815 106.370 140.225 ;
        RECT 105.460 139.645 105.790 139.765 ;
        RECT 106.540 139.645 106.710 140.405 ;
        RECT 105.460 139.475 106.710 139.645 ;
        RECT 106.880 140.585 108.250 140.835 ;
        RECT 106.880 139.815 107.070 140.585 ;
        RECT 108.000 140.325 108.250 140.585 ;
        RECT 107.240 140.155 107.490 140.315 ;
        RECT 108.420 140.155 108.590 141.000 ;
        RECT 109.485 140.715 109.655 141.215 ;
        RECT 109.825 140.885 110.155 141.385 ;
        RECT 108.760 140.325 109.260 140.705 ;
        RECT 109.485 140.545 110.180 140.715 ;
        RECT 107.240 139.985 108.590 140.155 ;
        RECT 108.170 139.945 108.590 139.985 ;
        RECT 106.880 139.475 107.300 139.815 ;
        RECT 107.590 139.485 108.000 139.815 ;
        RECT 105.120 139.055 105.970 139.225 ;
        RECT 106.530 138.835 106.850 139.295 ;
        RECT 107.050 139.045 107.300 139.475 ;
        RECT 107.590 138.835 108.000 139.275 ;
        RECT 108.170 139.215 108.340 139.945 ;
        RECT 108.510 139.395 108.860 139.765 ;
        RECT 109.040 139.455 109.260 140.325 ;
        RECT 109.430 139.755 109.840 140.375 ;
        RECT 110.010 139.575 110.180 140.545 ;
        RECT 109.485 139.385 110.180 139.575 ;
        RECT 108.170 139.015 109.185 139.215 ;
        RECT 109.485 139.055 109.655 139.385 ;
        RECT 109.825 138.835 110.155 139.215 ;
        RECT 110.370 139.095 110.595 141.215 ;
        RECT 110.765 140.885 111.095 141.385 ;
        RECT 111.265 140.715 111.435 141.215 ;
        RECT 110.770 140.545 111.435 140.715 ;
        RECT 110.770 139.555 111.000 140.545 ;
        RECT 111.170 139.725 111.520 140.375 ;
        RECT 112.155 140.295 113.365 141.385 ;
        RECT 112.155 139.755 112.675 140.295 ;
        RECT 112.845 139.585 113.365 140.125 ;
        RECT 110.770 139.385 111.435 139.555 ;
        RECT 110.765 138.835 111.095 139.215 ;
        RECT 111.265 139.095 111.435 139.385 ;
        RECT 112.155 138.835 113.365 139.585 ;
        RECT 26.970 138.665 113.450 138.835 ;
        RECT 27.055 137.915 28.265 138.665 ;
        RECT 28.745 138.195 28.915 138.665 ;
        RECT 29.085 138.015 29.415 138.495 ;
        RECT 29.585 138.195 29.755 138.665 ;
        RECT 29.925 138.015 30.255 138.495 ;
        RECT 27.055 137.375 27.575 137.915 ;
        RECT 28.490 137.845 30.255 138.015 ;
        RECT 30.425 137.855 30.595 138.665 ;
        RECT 30.795 138.285 31.865 138.455 ;
        RECT 30.795 137.930 31.115 138.285 ;
        RECT 27.745 137.205 28.265 137.745 ;
        RECT 27.055 136.115 28.265 137.205 ;
        RECT 28.490 137.295 28.900 137.845 ;
        RECT 30.790 137.675 31.115 137.930 ;
        RECT 29.085 137.465 31.115 137.675 ;
        RECT 30.770 137.455 31.115 137.465 ;
        RECT 31.285 137.715 31.525 138.115 ;
        RECT 31.695 138.055 31.865 138.285 ;
        RECT 32.035 138.225 32.225 138.665 ;
        RECT 32.395 138.215 33.345 138.495 ;
        RECT 33.565 138.305 33.915 138.475 ;
        RECT 31.695 137.885 32.225 138.055 ;
        RECT 28.490 137.125 30.215 137.295 ;
        RECT 28.745 136.115 28.915 136.955 ;
        RECT 29.125 136.285 29.375 137.125 ;
        RECT 29.585 136.115 29.755 136.955 ;
        RECT 29.925 136.285 30.215 137.125 ;
        RECT 30.425 136.115 30.595 137.175 ;
        RECT 30.770 136.835 30.940 137.455 ;
        RECT 31.285 137.345 31.825 137.715 ;
        RECT 32.005 137.605 32.225 137.885 ;
        RECT 32.395 137.435 32.565 138.215 ;
        RECT 32.160 137.265 32.565 137.435 ;
        RECT 32.735 137.425 33.085 138.045 ;
        RECT 32.160 137.175 32.330 137.265 ;
        RECT 33.255 137.255 33.465 138.045 ;
        RECT 31.110 137.005 32.330 137.175 ;
        RECT 32.790 137.095 33.465 137.255 ;
        RECT 30.770 136.665 31.570 136.835 ;
        RECT 30.890 136.115 31.220 136.495 ;
        RECT 31.400 136.375 31.570 136.665 ;
        RECT 32.160 136.625 32.330 137.005 ;
        RECT 32.500 137.085 33.465 137.095 ;
        RECT 33.655 137.915 33.915 138.305 ;
        RECT 34.125 138.205 34.455 138.665 ;
        RECT 35.330 138.275 36.185 138.445 ;
        RECT 36.390 138.275 36.885 138.445 ;
        RECT 37.055 138.305 37.385 138.665 ;
        RECT 33.655 137.225 33.825 137.915 ;
        RECT 33.995 137.565 34.165 137.745 ;
        RECT 34.335 137.735 35.125 137.985 ;
        RECT 35.330 137.565 35.500 138.275 ;
        RECT 35.670 137.765 36.025 137.985 ;
        RECT 33.995 137.395 35.685 137.565 ;
        RECT 32.500 136.795 32.960 137.085 ;
        RECT 33.655 137.055 35.155 137.225 ;
        RECT 33.655 136.915 33.825 137.055 ;
        RECT 33.265 136.745 33.825 136.915 ;
        RECT 31.740 136.115 31.990 136.575 ;
        RECT 32.160 136.285 33.030 136.625 ;
        RECT 33.265 136.285 33.435 136.745 ;
        RECT 34.270 136.715 35.345 136.885 ;
        RECT 33.605 136.115 33.975 136.575 ;
        RECT 34.270 136.375 34.440 136.715 ;
        RECT 34.610 136.115 34.940 136.545 ;
        RECT 35.175 136.375 35.345 136.715 ;
        RECT 35.515 136.615 35.685 137.395 ;
        RECT 35.855 137.175 36.025 137.765 ;
        RECT 36.195 137.365 36.545 137.985 ;
        RECT 35.855 136.785 36.320 137.175 ;
        RECT 36.715 136.915 36.885 138.275 ;
        RECT 37.055 137.085 37.515 138.135 ;
        RECT 36.490 136.745 36.885 136.915 ;
        RECT 36.490 136.615 36.660 136.745 ;
        RECT 35.515 136.285 36.195 136.615 ;
        RECT 36.410 136.285 36.660 136.615 ;
        RECT 36.830 136.115 37.080 136.575 ;
        RECT 37.250 136.300 37.575 137.085 ;
        RECT 37.745 136.285 37.915 138.405 ;
        RECT 38.085 138.285 38.415 138.665 ;
        RECT 38.585 138.115 38.840 138.405 ;
        RECT 38.090 137.945 38.840 138.115 ;
        RECT 39.105 138.115 39.275 138.405 ;
        RECT 39.445 138.285 39.775 138.665 ;
        RECT 39.105 137.945 39.770 138.115 ;
        RECT 38.090 136.955 38.320 137.945 ;
        RECT 38.490 137.125 38.840 137.775 ;
        RECT 39.020 137.125 39.370 137.775 ;
        RECT 39.540 136.955 39.770 137.945 ;
        RECT 38.090 136.785 38.840 136.955 ;
        RECT 38.085 136.115 38.415 136.615 ;
        RECT 38.585 136.285 38.840 136.785 ;
        RECT 39.105 136.785 39.770 136.955 ;
        RECT 39.105 136.285 39.275 136.785 ;
        RECT 39.445 136.115 39.775 136.615 ;
        RECT 39.945 136.285 40.170 138.405 ;
        RECT 40.385 138.285 40.715 138.665 ;
        RECT 40.885 138.115 41.055 138.445 ;
        RECT 41.355 138.285 42.370 138.485 ;
        RECT 40.360 137.925 41.055 138.115 ;
        RECT 40.360 136.955 40.530 137.925 ;
        RECT 40.700 137.125 41.110 137.745 ;
        RECT 41.280 137.175 41.500 138.045 ;
        RECT 41.680 137.735 42.030 138.105 ;
        RECT 42.200 137.555 42.370 138.285 ;
        RECT 42.540 138.225 42.950 138.665 ;
        RECT 43.240 138.025 43.490 138.455 ;
        RECT 43.690 138.205 44.010 138.665 ;
        RECT 44.570 138.275 45.420 138.445 ;
        RECT 42.540 137.685 42.950 138.015 ;
        RECT 43.240 137.685 43.660 138.025 ;
        RECT 41.950 137.515 42.370 137.555 ;
        RECT 41.950 137.345 43.300 137.515 ;
        RECT 40.360 136.785 41.055 136.955 ;
        RECT 41.280 136.795 41.780 137.175 ;
        RECT 40.385 136.115 40.715 136.615 ;
        RECT 40.885 136.285 41.055 136.785 ;
        RECT 41.950 136.500 42.120 137.345 ;
        RECT 43.050 137.185 43.300 137.345 ;
        RECT 42.290 136.915 42.540 137.175 ;
        RECT 43.470 136.915 43.660 137.685 ;
        RECT 42.290 136.665 43.660 136.915 ;
        RECT 43.830 137.855 45.080 138.025 ;
        RECT 43.830 137.095 44.000 137.855 ;
        RECT 44.750 137.735 45.080 137.855 ;
        RECT 44.170 137.275 44.350 137.685 ;
        RECT 45.250 137.515 45.420 138.275 ;
        RECT 45.620 138.185 46.280 138.665 ;
        RECT 46.460 138.070 46.780 138.400 ;
        RECT 45.610 137.745 46.270 138.015 ;
        RECT 45.610 137.685 45.940 137.745 ;
        RECT 46.090 137.515 46.420 137.575 ;
        RECT 44.520 137.345 46.420 137.515 ;
        RECT 43.830 136.785 44.350 137.095 ;
        RECT 44.520 136.835 44.690 137.345 ;
        RECT 46.590 137.175 46.780 138.070 ;
        RECT 44.860 137.005 46.780 137.175 ;
        RECT 46.460 136.985 46.780 137.005 ;
        RECT 46.980 137.755 47.230 138.405 ;
        RECT 47.410 138.205 47.695 138.665 ;
        RECT 47.875 137.955 48.130 138.485 ;
        RECT 46.980 137.425 47.780 137.755 ;
        RECT 44.520 136.665 45.730 136.835 ;
        RECT 41.290 136.330 42.120 136.500 ;
        RECT 42.360 136.115 42.740 136.495 ;
        RECT 42.920 136.375 43.090 136.665 ;
        RECT 44.520 136.585 44.690 136.665 ;
        RECT 43.260 136.115 43.590 136.495 ;
        RECT 44.060 136.335 44.690 136.585 ;
        RECT 44.870 136.115 45.290 136.495 ;
        RECT 45.490 136.375 45.730 136.665 ;
        RECT 45.960 136.115 46.290 136.805 ;
        RECT 46.460 136.375 46.630 136.985 ;
        RECT 46.980 136.835 47.230 137.425 ;
        RECT 47.950 137.095 48.130 137.955 ;
        RECT 48.675 137.940 48.965 138.665 ;
        RECT 49.225 138.115 49.395 138.405 ;
        RECT 49.565 138.285 49.895 138.665 ;
        RECT 49.225 137.945 49.890 138.115 ;
        RECT 46.900 136.325 47.230 136.835 ;
        RECT 47.410 136.115 47.695 136.915 ;
        RECT 47.875 136.625 48.130 137.095 ;
        RECT 47.875 136.455 48.215 136.625 ;
        RECT 47.875 136.425 48.130 136.455 ;
        RECT 48.675 136.115 48.965 137.280 ;
        RECT 49.140 137.125 49.490 137.775 ;
        RECT 49.660 136.955 49.890 137.945 ;
        RECT 49.225 136.785 49.890 136.955 ;
        RECT 49.225 136.285 49.395 136.785 ;
        RECT 49.565 136.115 49.895 136.615 ;
        RECT 50.065 136.285 50.290 138.405 ;
        RECT 50.505 138.285 50.835 138.665 ;
        RECT 51.005 138.115 51.175 138.445 ;
        RECT 51.475 138.285 52.490 138.485 ;
        RECT 50.480 137.925 51.175 138.115 ;
        RECT 50.480 136.955 50.650 137.925 ;
        RECT 50.820 137.125 51.230 137.745 ;
        RECT 51.400 137.175 51.620 138.045 ;
        RECT 51.800 137.735 52.150 138.105 ;
        RECT 52.320 137.555 52.490 138.285 ;
        RECT 52.660 138.225 53.070 138.665 ;
        RECT 53.360 138.025 53.610 138.455 ;
        RECT 53.810 138.205 54.130 138.665 ;
        RECT 54.690 138.275 55.540 138.445 ;
        RECT 52.660 137.685 53.070 138.015 ;
        RECT 53.360 137.685 53.780 138.025 ;
        RECT 52.070 137.515 52.490 137.555 ;
        RECT 52.070 137.345 53.420 137.515 ;
        RECT 50.480 136.785 51.175 136.955 ;
        RECT 51.400 136.795 51.900 137.175 ;
        RECT 50.505 136.115 50.835 136.615 ;
        RECT 51.005 136.285 51.175 136.785 ;
        RECT 52.070 136.500 52.240 137.345 ;
        RECT 53.170 137.185 53.420 137.345 ;
        RECT 52.410 136.915 52.660 137.175 ;
        RECT 53.590 136.915 53.780 137.685 ;
        RECT 52.410 136.665 53.780 136.915 ;
        RECT 53.950 137.855 55.200 138.025 ;
        RECT 53.950 137.095 54.120 137.855 ;
        RECT 54.870 137.735 55.200 137.855 ;
        RECT 54.290 137.275 54.470 137.685 ;
        RECT 55.370 137.515 55.540 138.275 ;
        RECT 55.740 138.185 56.400 138.665 ;
        RECT 56.580 138.070 56.900 138.400 ;
        RECT 55.730 137.745 56.390 138.015 ;
        RECT 55.730 137.685 56.060 137.745 ;
        RECT 56.210 137.515 56.540 137.575 ;
        RECT 54.640 137.345 56.540 137.515 ;
        RECT 53.950 136.785 54.470 137.095 ;
        RECT 54.640 136.835 54.810 137.345 ;
        RECT 56.710 137.175 56.900 138.070 ;
        RECT 54.980 137.005 56.900 137.175 ;
        RECT 56.580 136.985 56.900 137.005 ;
        RECT 57.100 137.755 57.350 138.405 ;
        RECT 57.530 138.205 57.815 138.665 ;
        RECT 57.995 137.955 58.250 138.485 ;
        RECT 57.100 137.425 57.900 137.755 ;
        RECT 54.640 136.665 55.850 136.835 ;
        RECT 51.410 136.330 52.240 136.500 ;
        RECT 52.480 136.115 52.860 136.495 ;
        RECT 53.040 136.375 53.210 136.665 ;
        RECT 54.640 136.585 54.810 136.665 ;
        RECT 53.380 136.115 53.710 136.495 ;
        RECT 54.180 136.335 54.810 136.585 ;
        RECT 54.990 136.115 55.410 136.495 ;
        RECT 55.610 136.375 55.850 136.665 ;
        RECT 56.080 136.115 56.410 136.805 ;
        RECT 56.580 136.375 56.750 136.985 ;
        RECT 57.100 136.835 57.350 137.425 ;
        RECT 58.070 137.095 58.250 137.955 ;
        RECT 59.345 138.115 59.515 138.495 ;
        RECT 59.695 138.285 60.025 138.665 ;
        RECT 59.345 137.945 60.010 138.115 ;
        RECT 60.205 137.990 60.465 138.495 ;
        RECT 61.010 138.325 61.265 138.485 ;
        RECT 60.925 138.155 61.265 138.325 ;
        RECT 61.445 138.205 61.730 138.665 ;
        RECT 59.275 137.395 59.605 137.765 ;
        RECT 59.840 137.690 60.010 137.945 ;
        RECT 59.840 137.360 60.125 137.690 ;
        RECT 59.840 137.215 60.010 137.360 ;
        RECT 57.020 136.325 57.350 136.835 ;
        RECT 57.530 136.115 57.815 136.915 ;
        RECT 57.995 136.625 58.250 137.095 ;
        RECT 59.345 137.045 60.010 137.215 ;
        RECT 60.295 137.190 60.465 137.990 ;
        RECT 57.995 136.455 58.335 136.625 ;
        RECT 57.995 136.425 58.250 136.455 ;
        RECT 59.345 136.285 59.515 137.045 ;
        RECT 59.695 136.115 60.025 136.875 ;
        RECT 60.195 136.285 60.465 137.190 ;
        RECT 61.010 137.955 61.265 138.155 ;
        RECT 61.010 137.095 61.190 137.955 ;
        RECT 61.910 137.755 62.160 138.405 ;
        RECT 61.360 137.425 62.160 137.755 ;
        RECT 61.010 136.425 61.265 137.095 ;
        RECT 61.445 136.115 61.730 136.915 ;
        RECT 61.910 136.835 62.160 137.425 ;
        RECT 62.360 138.070 62.680 138.400 ;
        RECT 62.860 138.185 63.520 138.665 ;
        RECT 63.720 138.275 64.570 138.445 ;
        RECT 62.360 137.175 62.550 138.070 ;
        RECT 62.870 137.745 63.530 138.015 ;
        RECT 63.200 137.685 63.530 137.745 ;
        RECT 62.720 137.515 63.050 137.575 ;
        RECT 63.720 137.515 63.890 138.275 ;
        RECT 65.130 138.205 65.450 138.665 ;
        RECT 65.650 138.025 65.900 138.455 ;
        RECT 66.190 138.225 66.600 138.665 ;
        RECT 66.770 138.285 67.785 138.485 ;
        RECT 64.060 137.855 65.310 138.025 ;
        RECT 64.060 137.735 64.390 137.855 ;
        RECT 62.720 137.345 64.620 137.515 ;
        RECT 62.360 137.005 64.280 137.175 ;
        RECT 62.360 136.985 62.680 137.005 ;
        RECT 61.910 136.325 62.240 136.835 ;
        RECT 62.510 136.375 62.680 136.985 ;
        RECT 64.450 136.835 64.620 137.345 ;
        RECT 64.790 137.275 64.970 137.685 ;
        RECT 65.140 137.095 65.310 137.855 ;
        RECT 62.850 136.115 63.180 136.805 ;
        RECT 63.410 136.665 64.620 136.835 ;
        RECT 64.790 136.785 65.310 137.095 ;
        RECT 65.480 137.685 65.900 138.025 ;
        RECT 66.190 137.685 66.600 138.015 ;
        RECT 65.480 136.915 65.670 137.685 ;
        RECT 66.770 137.555 66.940 138.285 ;
        RECT 68.085 138.115 68.255 138.445 ;
        RECT 68.425 138.285 68.755 138.665 ;
        RECT 67.110 137.735 67.460 138.105 ;
        RECT 66.770 137.515 67.190 137.555 ;
        RECT 65.840 137.345 67.190 137.515 ;
        RECT 65.840 137.185 66.090 137.345 ;
        RECT 66.600 136.915 66.850 137.175 ;
        RECT 65.480 136.665 66.850 136.915 ;
        RECT 63.410 136.375 63.650 136.665 ;
        RECT 64.450 136.585 64.620 136.665 ;
        RECT 63.850 136.115 64.270 136.495 ;
        RECT 64.450 136.335 65.080 136.585 ;
        RECT 65.550 136.115 65.880 136.495 ;
        RECT 66.050 136.375 66.220 136.665 ;
        RECT 67.020 136.500 67.190 137.345 ;
        RECT 67.640 137.175 67.860 138.045 ;
        RECT 68.085 137.925 68.780 138.115 ;
        RECT 67.360 136.795 67.860 137.175 ;
        RECT 68.030 137.125 68.440 137.745 ;
        RECT 68.610 136.955 68.780 137.925 ;
        RECT 68.085 136.785 68.780 136.955 ;
        RECT 66.400 136.115 66.780 136.495 ;
        RECT 67.020 136.330 67.850 136.500 ;
        RECT 68.085 136.285 68.255 136.785 ;
        RECT 68.425 136.115 68.755 136.615 ;
        RECT 68.970 136.285 69.195 138.405 ;
        RECT 69.365 138.285 69.695 138.665 ;
        RECT 69.865 138.115 70.035 138.405 ;
        RECT 69.370 137.945 70.035 138.115 ;
        RECT 70.955 138.035 71.285 138.395 ;
        RECT 71.905 138.205 72.155 138.665 ;
        RECT 72.325 138.205 72.885 138.495 ;
        RECT 69.370 136.955 69.600 137.945 ;
        RECT 70.955 137.845 72.345 138.035 ;
        RECT 69.770 137.125 70.120 137.775 ;
        RECT 72.175 137.755 72.345 137.845 ;
        RECT 70.770 137.425 71.445 137.675 ;
        RECT 71.665 137.425 72.005 137.675 ;
        RECT 72.175 137.425 72.465 137.755 ;
        RECT 70.770 137.065 71.035 137.425 ;
        RECT 72.175 137.175 72.345 137.425 ;
        RECT 71.405 137.005 72.345 137.175 ;
        RECT 69.370 136.785 70.035 136.955 ;
        RECT 69.365 136.115 69.695 136.615 ;
        RECT 69.865 136.285 70.035 136.785 ;
        RECT 70.955 136.115 71.235 136.785 ;
        RECT 71.405 136.455 71.705 137.005 ;
        RECT 72.635 136.835 72.885 138.205 ;
        RECT 71.905 136.115 72.235 136.835 ;
        RECT 72.425 136.285 72.885 136.835 ;
        RECT 73.055 137.990 73.315 138.495 ;
        RECT 73.495 138.285 73.825 138.665 ;
        RECT 74.005 138.115 74.175 138.495 ;
        RECT 73.055 137.190 73.225 137.990 ;
        RECT 73.510 137.945 74.175 138.115 ;
        RECT 73.510 137.690 73.680 137.945 ;
        RECT 74.435 137.940 74.725 138.665 ;
        RECT 75.170 137.855 75.415 138.460 ;
        RECT 75.635 138.130 76.145 138.665 ;
        RECT 73.395 137.360 73.680 137.690 ;
        RECT 73.915 137.395 74.245 137.765 ;
        RECT 74.895 137.685 76.125 137.855 ;
        RECT 73.510 137.215 73.680 137.360 ;
        RECT 73.055 136.285 73.325 137.190 ;
        RECT 73.510 137.045 74.175 137.215 ;
        RECT 73.495 136.115 73.825 136.875 ;
        RECT 74.005 136.285 74.175 137.045 ;
        RECT 74.435 136.115 74.725 137.280 ;
        RECT 74.895 136.875 75.235 137.685 ;
        RECT 75.405 137.120 76.155 137.310 ;
        RECT 74.895 136.465 75.410 136.875 ;
        RECT 75.645 136.115 75.815 136.875 ;
        RECT 75.985 136.455 76.155 137.120 ;
        RECT 76.325 137.135 76.515 138.495 ;
        RECT 76.685 137.645 76.960 138.495 ;
        RECT 77.150 138.130 77.680 138.495 ;
        RECT 78.105 138.265 78.435 138.665 ;
        RECT 77.505 138.095 77.680 138.130 ;
        RECT 76.685 137.475 76.965 137.645 ;
        RECT 76.685 137.335 76.960 137.475 ;
        RECT 77.165 137.135 77.335 137.935 ;
        RECT 76.325 136.965 77.335 137.135 ;
        RECT 77.505 137.925 78.435 138.095 ;
        RECT 78.605 137.925 78.860 138.495 ;
        RECT 77.505 136.795 77.675 137.925 ;
        RECT 78.265 137.755 78.435 137.925 ;
        RECT 76.550 136.625 77.675 136.795 ;
        RECT 77.845 137.425 78.040 137.755 ;
        RECT 78.265 137.425 78.520 137.755 ;
        RECT 77.845 136.455 78.015 137.425 ;
        RECT 78.690 137.255 78.860 137.925 ;
        RECT 75.985 136.285 78.015 136.455 ;
        RECT 78.185 136.115 78.355 137.255 ;
        RECT 78.525 136.285 78.860 137.255 ;
        RECT 79.035 138.205 79.595 138.495 ;
        RECT 79.765 138.205 80.015 138.665 ;
        RECT 79.035 136.835 79.285 138.205 ;
        RECT 80.635 138.035 80.965 138.395 ;
        RECT 79.575 137.845 80.965 138.035 ;
        RECT 81.335 138.205 81.895 138.495 ;
        RECT 82.065 138.205 82.315 138.665 ;
        RECT 79.575 137.755 79.745 137.845 ;
        RECT 79.455 137.425 79.745 137.755 ;
        RECT 79.915 137.425 80.255 137.675 ;
        RECT 80.475 137.425 81.150 137.675 ;
        RECT 79.575 137.175 79.745 137.425 ;
        RECT 79.575 137.005 80.515 137.175 ;
        RECT 80.885 137.065 81.150 137.425 ;
        RECT 79.035 136.285 79.495 136.835 ;
        RECT 79.685 136.115 80.015 136.835 ;
        RECT 80.215 136.455 80.515 137.005 ;
        RECT 81.335 136.835 81.585 138.205 ;
        RECT 82.935 138.035 83.265 138.395 ;
        RECT 81.875 137.845 83.265 138.035 ;
        RECT 84.830 137.855 85.075 138.460 ;
        RECT 85.295 138.130 85.805 138.665 ;
        RECT 81.875 137.755 82.045 137.845 ;
        RECT 81.755 137.425 82.045 137.755 ;
        RECT 84.555 137.685 85.785 137.855 ;
        RECT 82.215 137.425 82.555 137.675 ;
        RECT 82.775 137.425 83.450 137.675 ;
        RECT 81.875 137.175 82.045 137.425 ;
        RECT 81.875 137.005 82.815 137.175 ;
        RECT 83.185 137.065 83.450 137.425 ;
        RECT 80.685 136.115 80.965 136.785 ;
        RECT 81.335 136.285 81.795 136.835 ;
        RECT 81.985 136.115 82.315 136.835 ;
        RECT 82.515 136.455 82.815 137.005 ;
        RECT 84.555 136.875 84.895 137.685 ;
        RECT 85.065 137.120 85.815 137.310 ;
        RECT 82.985 136.115 83.265 136.785 ;
        RECT 84.555 136.465 85.070 136.875 ;
        RECT 85.305 136.115 85.475 136.875 ;
        RECT 85.645 136.455 85.815 137.120 ;
        RECT 85.985 137.135 86.175 138.495 ;
        RECT 86.345 137.645 86.620 138.495 ;
        RECT 86.810 138.130 87.340 138.495 ;
        RECT 87.765 138.265 88.095 138.665 ;
        RECT 87.165 138.095 87.340 138.130 ;
        RECT 86.345 137.475 86.625 137.645 ;
        RECT 86.345 137.335 86.620 137.475 ;
        RECT 86.825 137.135 86.995 137.935 ;
        RECT 85.985 136.965 86.995 137.135 ;
        RECT 87.165 137.925 88.095 138.095 ;
        RECT 88.265 137.925 88.520 138.495 ;
        RECT 87.165 136.795 87.335 137.925 ;
        RECT 87.925 137.755 88.095 137.925 ;
        RECT 86.210 136.625 87.335 136.795 ;
        RECT 87.505 137.425 87.700 137.755 ;
        RECT 87.925 137.425 88.180 137.755 ;
        RECT 87.505 136.455 87.675 137.425 ;
        RECT 88.350 137.255 88.520 137.925 ;
        RECT 88.755 137.845 88.965 138.665 ;
        RECT 89.135 137.865 89.465 138.495 ;
        RECT 89.135 137.265 89.385 137.865 ;
        RECT 89.635 137.845 89.865 138.665 ;
        RECT 90.115 137.845 90.345 138.665 ;
        RECT 90.515 137.865 90.845 138.495 ;
        RECT 89.555 137.425 89.885 137.675 ;
        RECT 90.095 137.425 90.425 137.675 ;
        RECT 90.595 137.265 90.845 137.865 ;
        RECT 91.015 137.845 91.225 138.665 ;
        RECT 92.190 137.855 92.435 138.460 ;
        RECT 92.655 138.130 93.165 138.665 ;
        RECT 85.645 136.285 87.675 136.455 ;
        RECT 87.845 136.115 88.015 137.255 ;
        RECT 88.185 136.285 88.520 137.255 ;
        RECT 88.755 136.115 88.965 137.255 ;
        RECT 89.135 136.285 89.465 137.265 ;
        RECT 89.635 136.115 89.865 137.255 ;
        RECT 90.115 136.115 90.345 137.255 ;
        RECT 90.515 136.285 90.845 137.265 ;
        RECT 91.915 137.685 93.145 137.855 ;
        RECT 91.015 136.115 91.225 137.255 ;
        RECT 91.915 136.875 92.255 137.685 ;
        RECT 92.425 137.120 93.175 137.310 ;
        RECT 91.915 136.465 92.430 136.875 ;
        RECT 92.665 136.115 92.835 136.875 ;
        RECT 93.005 136.455 93.175 137.120 ;
        RECT 93.345 137.135 93.535 138.495 ;
        RECT 93.705 138.325 93.980 138.495 ;
        RECT 93.705 138.155 93.985 138.325 ;
        RECT 93.705 137.335 93.980 138.155 ;
        RECT 94.170 138.130 94.700 138.495 ;
        RECT 95.125 138.265 95.455 138.665 ;
        RECT 94.525 138.095 94.700 138.130 ;
        RECT 94.185 137.135 94.355 137.935 ;
        RECT 93.345 136.965 94.355 137.135 ;
        RECT 94.525 137.925 95.455 138.095 ;
        RECT 95.625 137.925 95.880 138.495 ;
        RECT 94.525 136.795 94.695 137.925 ;
        RECT 95.285 137.755 95.455 137.925 ;
        RECT 93.570 136.625 94.695 136.795 ;
        RECT 94.865 137.425 95.060 137.755 ;
        RECT 95.285 137.425 95.540 137.755 ;
        RECT 94.865 136.455 95.035 137.425 ;
        RECT 95.710 137.255 95.880 137.925 ;
        RECT 96.330 137.855 96.575 138.460 ;
        RECT 96.795 138.130 97.305 138.665 ;
        RECT 93.005 136.285 95.035 136.455 ;
        RECT 95.205 136.115 95.375 137.255 ;
        RECT 95.545 136.285 95.880 137.255 ;
        RECT 96.055 137.685 97.285 137.855 ;
        RECT 96.055 136.875 96.395 137.685 ;
        RECT 96.565 137.120 97.315 137.310 ;
        RECT 96.055 136.465 96.570 136.875 ;
        RECT 96.805 136.115 96.975 136.875 ;
        RECT 97.145 136.455 97.315 137.120 ;
        RECT 97.485 137.135 97.675 138.495 ;
        RECT 97.845 137.645 98.120 138.495 ;
        RECT 98.310 138.130 98.840 138.495 ;
        RECT 99.265 138.265 99.595 138.665 ;
        RECT 98.665 138.095 98.840 138.130 ;
        RECT 97.845 137.475 98.125 137.645 ;
        RECT 97.845 137.335 98.120 137.475 ;
        RECT 98.325 137.135 98.495 137.935 ;
        RECT 97.485 136.965 98.495 137.135 ;
        RECT 98.665 137.925 99.595 138.095 ;
        RECT 99.765 137.925 100.020 138.495 ;
        RECT 100.195 137.940 100.485 138.665 ;
        RECT 101.030 138.325 101.285 138.485 ;
        RECT 100.945 138.155 101.285 138.325 ;
        RECT 101.465 138.205 101.750 138.665 ;
        RECT 101.030 137.955 101.285 138.155 ;
        RECT 98.665 136.795 98.835 137.925 ;
        RECT 99.425 137.755 99.595 137.925 ;
        RECT 97.710 136.625 98.835 136.795 ;
        RECT 99.005 137.425 99.200 137.755 ;
        RECT 99.425 137.425 99.680 137.755 ;
        RECT 99.005 136.455 99.175 137.425 ;
        RECT 99.850 137.255 100.020 137.925 ;
        RECT 97.145 136.285 99.175 136.455 ;
        RECT 99.345 136.115 99.515 137.255 ;
        RECT 99.685 136.285 100.020 137.255 ;
        RECT 100.195 136.115 100.485 137.280 ;
        RECT 101.030 137.095 101.210 137.955 ;
        RECT 101.930 137.755 102.180 138.405 ;
        RECT 101.380 137.425 102.180 137.755 ;
        RECT 101.030 136.425 101.285 137.095 ;
        RECT 101.465 136.115 101.750 136.915 ;
        RECT 101.930 136.835 102.180 137.425 ;
        RECT 102.380 138.070 102.700 138.400 ;
        RECT 102.880 138.185 103.540 138.665 ;
        RECT 103.740 138.275 104.590 138.445 ;
        RECT 102.380 137.175 102.570 138.070 ;
        RECT 102.890 137.745 103.550 138.015 ;
        RECT 103.220 137.685 103.550 137.745 ;
        RECT 102.740 137.515 103.070 137.575 ;
        RECT 103.740 137.515 103.910 138.275 ;
        RECT 105.150 138.205 105.470 138.665 ;
        RECT 105.670 138.025 105.920 138.455 ;
        RECT 106.210 138.225 106.620 138.665 ;
        RECT 106.790 138.285 107.805 138.485 ;
        RECT 104.080 137.855 105.330 138.025 ;
        RECT 104.080 137.735 104.410 137.855 ;
        RECT 102.740 137.345 104.640 137.515 ;
        RECT 102.380 137.005 104.300 137.175 ;
        RECT 102.380 136.985 102.700 137.005 ;
        RECT 101.930 136.325 102.260 136.835 ;
        RECT 102.530 136.375 102.700 136.985 ;
        RECT 104.470 136.835 104.640 137.345 ;
        RECT 104.810 137.275 104.990 137.685 ;
        RECT 105.160 137.095 105.330 137.855 ;
        RECT 102.870 136.115 103.200 136.805 ;
        RECT 103.430 136.665 104.640 136.835 ;
        RECT 104.810 136.785 105.330 137.095 ;
        RECT 105.500 137.685 105.920 138.025 ;
        RECT 106.210 137.685 106.620 138.015 ;
        RECT 105.500 136.915 105.690 137.685 ;
        RECT 106.790 137.555 106.960 138.285 ;
        RECT 108.105 138.115 108.275 138.445 ;
        RECT 108.445 138.285 108.775 138.665 ;
        RECT 107.130 137.735 107.480 138.105 ;
        RECT 106.790 137.515 107.210 137.555 ;
        RECT 105.860 137.345 107.210 137.515 ;
        RECT 105.860 137.185 106.110 137.345 ;
        RECT 106.620 136.915 106.870 137.175 ;
        RECT 105.500 136.665 106.870 136.915 ;
        RECT 103.430 136.375 103.670 136.665 ;
        RECT 104.470 136.585 104.640 136.665 ;
        RECT 103.870 136.115 104.290 136.495 ;
        RECT 104.470 136.335 105.100 136.585 ;
        RECT 105.570 136.115 105.900 136.495 ;
        RECT 106.070 136.375 106.240 136.665 ;
        RECT 107.040 136.500 107.210 137.345 ;
        RECT 107.660 137.175 107.880 138.045 ;
        RECT 108.105 137.925 108.800 138.115 ;
        RECT 107.380 136.795 107.880 137.175 ;
        RECT 108.050 137.125 108.460 137.745 ;
        RECT 108.630 136.955 108.800 137.925 ;
        RECT 108.105 136.785 108.800 136.955 ;
        RECT 106.420 136.115 106.800 136.495 ;
        RECT 107.040 136.330 107.870 136.500 ;
        RECT 108.105 136.285 108.275 136.785 ;
        RECT 108.445 136.115 108.775 136.615 ;
        RECT 108.990 136.285 109.215 138.405 ;
        RECT 109.385 138.285 109.715 138.665 ;
        RECT 109.885 138.115 110.055 138.405 ;
        RECT 109.390 137.945 110.055 138.115 ;
        RECT 110.315 137.990 110.575 138.495 ;
        RECT 110.755 138.285 111.085 138.665 ;
        RECT 111.265 138.115 111.435 138.495 ;
        RECT 109.390 136.955 109.620 137.945 ;
        RECT 109.790 137.125 110.140 137.775 ;
        RECT 110.315 137.190 110.485 137.990 ;
        RECT 110.770 137.945 111.435 138.115 ;
        RECT 110.770 137.690 110.940 137.945 ;
        RECT 112.155 137.915 113.365 138.665 ;
        RECT 110.655 137.360 110.940 137.690 ;
        RECT 111.175 137.395 111.505 137.765 ;
        RECT 110.770 137.215 110.940 137.360 ;
        RECT 109.390 136.785 110.055 136.955 ;
        RECT 109.385 136.115 109.715 136.615 ;
        RECT 109.885 136.285 110.055 136.785 ;
        RECT 110.315 136.285 110.585 137.190 ;
        RECT 110.770 137.045 111.435 137.215 ;
        RECT 110.755 136.115 111.085 136.875 ;
        RECT 111.265 136.285 111.435 137.045 ;
        RECT 112.155 137.205 112.675 137.745 ;
        RECT 112.845 137.375 113.365 137.915 ;
        RECT 112.155 136.115 113.365 137.205 ;
        RECT 26.970 135.945 113.450 136.115 ;
        RECT 27.055 134.855 28.265 135.945 ;
        RECT 27.055 134.145 27.575 134.685 ;
        RECT 27.745 134.315 28.265 134.855 ;
        RECT 28.525 135.015 28.695 135.775 ;
        RECT 28.875 135.185 29.205 135.945 ;
        RECT 28.525 134.845 29.190 135.015 ;
        RECT 29.375 134.870 29.645 135.775 ;
        RECT 29.020 134.700 29.190 134.845 ;
        RECT 28.455 134.295 28.785 134.665 ;
        RECT 29.020 134.370 29.305 134.700 ;
        RECT 27.055 133.395 28.265 134.145 ;
        RECT 29.020 134.115 29.190 134.370 ;
        RECT 28.525 133.945 29.190 134.115 ;
        RECT 29.475 134.070 29.645 134.870 ;
        RECT 29.855 134.805 30.085 135.945 ;
        RECT 30.255 134.795 30.585 135.775 ;
        RECT 30.755 134.805 30.965 135.945 ;
        RECT 31.195 135.185 31.710 135.595 ;
        RECT 31.945 135.185 32.115 135.945 ;
        RECT 32.285 135.605 34.315 135.775 ;
        RECT 29.835 134.385 30.165 134.635 ;
        RECT 28.525 133.565 28.695 133.945 ;
        RECT 28.875 133.395 29.205 133.775 ;
        RECT 29.385 133.565 29.645 134.070 ;
        RECT 29.855 133.395 30.085 134.215 ;
        RECT 30.335 134.195 30.585 134.795 ;
        RECT 31.195 134.375 31.535 135.185 ;
        RECT 32.285 134.940 32.455 135.605 ;
        RECT 32.850 135.265 33.975 135.435 ;
        RECT 31.705 134.750 32.455 134.940 ;
        RECT 32.625 134.925 33.635 135.095 ;
        RECT 30.255 133.565 30.585 134.195 ;
        RECT 30.755 133.395 30.965 134.215 ;
        RECT 31.195 134.205 32.425 134.375 ;
        RECT 31.470 133.600 31.715 134.205 ;
        RECT 31.935 133.395 32.445 133.930 ;
        RECT 32.625 133.565 32.815 134.925 ;
        RECT 32.985 134.245 33.260 134.725 ;
        RECT 32.985 134.075 33.265 134.245 ;
        RECT 33.465 134.125 33.635 134.925 ;
        RECT 33.805 134.135 33.975 135.265 ;
        RECT 34.145 134.635 34.315 135.605 ;
        RECT 34.485 134.805 34.655 135.945 ;
        RECT 34.825 134.805 35.160 135.775 ;
        RECT 34.145 134.305 34.340 134.635 ;
        RECT 34.565 134.305 34.820 134.635 ;
        RECT 34.565 134.135 34.735 134.305 ;
        RECT 34.990 134.135 35.160 134.805 ;
        RECT 35.795 134.780 36.085 135.945 ;
        RECT 36.405 134.795 36.735 135.945 ;
        RECT 36.905 134.925 37.075 135.775 ;
        RECT 37.245 135.145 37.575 135.945 ;
        RECT 37.745 134.925 37.915 135.775 ;
        RECT 38.095 135.145 38.335 135.945 ;
        RECT 38.505 134.965 38.835 135.775 ;
        RECT 39.105 135.275 39.275 135.775 ;
        RECT 39.445 135.445 39.775 135.945 ;
        RECT 39.105 135.105 39.770 135.275 ;
        RECT 36.905 134.755 37.915 134.925 ;
        RECT 38.120 134.795 38.835 134.965 ;
        RECT 36.905 134.215 37.400 134.755 ;
        RECT 38.120 134.555 38.290 134.795 ;
        RECT 37.790 134.385 38.290 134.555 ;
        RECT 38.460 134.385 38.840 134.625 ;
        RECT 38.120 134.215 38.290 134.385 ;
        RECT 39.020 134.285 39.370 134.935 ;
        RECT 32.985 133.565 33.260 134.075 ;
        RECT 33.805 133.965 34.735 134.135 ;
        RECT 33.805 133.930 33.980 133.965 ;
        RECT 33.450 133.565 33.980 133.930 ;
        RECT 34.405 133.395 34.735 133.795 ;
        RECT 34.905 133.565 35.160 134.135 ;
        RECT 35.795 133.395 36.085 134.120 ;
        RECT 36.405 133.395 36.735 134.195 ;
        RECT 36.905 134.045 37.915 134.215 ;
        RECT 38.120 134.045 38.755 134.215 ;
        RECT 39.540 134.115 39.770 135.105 ;
        RECT 36.905 133.565 37.075 134.045 ;
        RECT 37.245 133.395 37.575 133.875 ;
        RECT 37.745 133.565 37.915 134.045 ;
        RECT 38.165 133.395 38.405 133.875 ;
        RECT 38.585 133.565 38.755 134.045 ;
        RECT 39.105 133.945 39.770 134.115 ;
        RECT 39.105 133.655 39.275 133.945 ;
        RECT 39.445 133.395 39.775 133.775 ;
        RECT 39.945 133.655 40.170 135.775 ;
        RECT 40.385 135.445 40.715 135.945 ;
        RECT 40.885 135.275 41.055 135.775 ;
        RECT 41.290 135.560 42.120 135.730 ;
        RECT 42.360 135.565 42.740 135.945 ;
        RECT 40.360 135.105 41.055 135.275 ;
        RECT 40.360 134.135 40.530 135.105 ;
        RECT 40.700 134.315 41.110 134.935 ;
        RECT 41.280 134.885 41.780 135.265 ;
        RECT 40.360 133.945 41.055 134.135 ;
        RECT 41.280 134.015 41.500 134.885 ;
        RECT 41.950 134.715 42.120 135.560 ;
        RECT 42.920 135.395 43.090 135.685 ;
        RECT 43.260 135.565 43.590 135.945 ;
        RECT 44.060 135.475 44.690 135.725 ;
        RECT 44.870 135.565 45.290 135.945 ;
        RECT 44.520 135.395 44.690 135.475 ;
        RECT 45.490 135.395 45.730 135.685 ;
        RECT 42.290 135.145 43.660 135.395 ;
        RECT 42.290 134.885 42.540 135.145 ;
        RECT 43.050 134.715 43.300 134.875 ;
        RECT 41.950 134.545 43.300 134.715 ;
        RECT 41.950 134.505 42.370 134.545 ;
        RECT 41.680 133.955 42.030 134.325 ;
        RECT 40.385 133.395 40.715 133.775 ;
        RECT 40.885 133.615 41.055 133.945 ;
        RECT 42.200 133.775 42.370 134.505 ;
        RECT 43.470 134.375 43.660 135.145 ;
        RECT 42.540 134.045 42.950 134.375 ;
        RECT 43.240 134.035 43.660 134.375 ;
        RECT 43.830 134.965 44.350 135.275 ;
        RECT 44.520 135.225 45.730 135.395 ;
        RECT 45.960 135.255 46.290 135.945 ;
        RECT 43.830 134.205 44.000 134.965 ;
        RECT 44.170 134.375 44.350 134.785 ;
        RECT 44.520 134.715 44.690 135.225 ;
        RECT 46.460 135.075 46.630 135.685 ;
        RECT 46.900 135.225 47.230 135.735 ;
        RECT 46.460 135.055 46.780 135.075 ;
        RECT 44.860 134.885 46.780 135.055 ;
        RECT 44.520 134.545 46.420 134.715 ;
        RECT 44.750 134.205 45.080 134.325 ;
        RECT 43.830 134.035 45.080 134.205 ;
        RECT 41.355 133.575 42.370 133.775 ;
        RECT 42.540 133.395 42.950 133.835 ;
        RECT 43.240 133.605 43.490 134.035 ;
        RECT 43.690 133.395 44.010 133.855 ;
        RECT 45.250 133.785 45.420 134.545 ;
        RECT 46.090 134.485 46.420 134.545 ;
        RECT 45.610 134.315 45.940 134.375 ;
        RECT 45.610 134.045 46.270 134.315 ;
        RECT 46.590 133.990 46.780 134.885 ;
        RECT 44.570 133.615 45.420 133.785 ;
        RECT 45.620 133.395 46.280 133.875 ;
        RECT 46.460 133.660 46.780 133.990 ;
        RECT 46.980 134.635 47.230 135.225 ;
        RECT 47.410 135.145 47.695 135.945 ;
        RECT 47.875 135.605 48.130 135.635 ;
        RECT 47.875 135.435 48.215 135.605 ;
        RECT 47.875 134.965 48.130 135.435 ;
        RECT 46.980 134.305 47.780 134.635 ;
        RECT 46.980 133.655 47.230 134.305 ;
        RECT 47.950 134.105 48.130 134.965 ;
        RECT 49.050 134.965 49.305 135.635 ;
        RECT 49.485 135.145 49.770 135.945 ;
        RECT 49.950 135.225 50.280 135.735 ;
        RECT 49.050 134.925 49.230 134.965 ;
        RECT 48.965 134.755 49.230 134.925 ;
        RECT 47.410 133.395 47.695 133.855 ;
        RECT 47.875 133.575 48.130 134.105 ;
        RECT 49.050 134.105 49.230 134.755 ;
        RECT 49.950 134.635 50.200 135.225 ;
        RECT 50.550 135.075 50.720 135.685 ;
        RECT 50.890 135.255 51.220 135.945 ;
        RECT 51.450 135.395 51.690 135.685 ;
        RECT 51.890 135.565 52.310 135.945 ;
        RECT 52.490 135.475 53.120 135.725 ;
        RECT 53.590 135.565 53.920 135.945 ;
        RECT 52.490 135.395 52.660 135.475 ;
        RECT 54.090 135.395 54.260 135.685 ;
        RECT 54.440 135.565 54.820 135.945 ;
        RECT 55.060 135.560 55.890 135.730 ;
        RECT 51.450 135.225 52.660 135.395 ;
        RECT 49.400 134.305 50.200 134.635 ;
        RECT 49.050 133.575 49.305 134.105 ;
        RECT 49.485 133.395 49.770 133.855 ;
        RECT 49.950 133.655 50.200 134.305 ;
        RECT 50.400 135.055 50.720 135.075 ;
        RECT 50.400 134.885 52.320 135.055 ;
        RECT 50.400 133.990 50.590 134.885 ;
        RECT 52.490 134.715 52.660 135.225 ;
        RECT 52.830 134.965 53.350 135.275 ;
        RECT 50.760 134.545 52.660 134.715 ;
        RECT 50.760 134.485 51.090 134.545 ;
        RECT 51.240 134.315 51.570 134.375 ;
        RECT 50.910 134.045 51.570 134.315 ;
        RECT 50.400 133.660 50.720 133.990 ;
        RECT 50.900 133.395 51.560 133.875 ;
        RECT 51.760 133.785 51.930 134.545 ;
        RECT 52.830 134.375 53.010 134.785 ;
        RECT 52.100 134.205 52.430 134.325 ;
        RECT 53.180 134.205 53.350 134.965 ;
        RECT 52.100 134.035 53.350 134.205 ;
        RECT 53.520 135.145 54.890 135.395 ;
        RECT 53.520 134.375 53.710 135.145 ;
        RECT 54.640 134.885 54.890 135.145 ;
        RECT 53.880 134.715 54.130 134.875 ;
        RECT 55.060 134.715 55.230 135.560 ;
        RECT 56.125 135.275 56.295 135.775 ;
        RECT 56.465 135.445 56.795 135.945 ;
        RECT 55.400 134.885 55.900 135.265 ;
        RECT 56.125 135.105 56.820 135.275 ;
        RECT 53.880 134.545 55.230 134.715 ;
        RECT 54.810 134.505 55.230 134.545 ;
        RECT 53.520 134.035 53.940 134.375 ;
        RECT 54.230 134.045 54.640 134.375 ;
        RECT 51.760 133.615 52.610 133.785 ;
        RECT 53.170 133.395 53.490 133.855 ;
        RECT 53.690 133.605 53.940 134.035 ;
        RECT 54.230 133.395 54.640 133.835 ;
        RECT 54.810 133.775 54.980 134.505 ;
        RECT 55.150 133.955 55.500 134.325 ;
        RECT 55.680 134.015 55.900 134.885 ;
        RECT 56.070 134.315 56.480 134.935 ;
        RECT 56.650 134.135 56.820 135.105 ;
        RECT 56.125 133.945 56.820 134.135 ;
        RECT 54.810 133.575 55.825 133.775 ;
        RECT 56.125 133.615 56.295 133.945 ;
        RECT 56.465 133.395 56.795 133.775 ;
        RECT 57.010 133.655 57.235 135.775 ;
        RECT 57.405 135.445 57.735 135.945 ;
        RECT 57.905 135.275 58.075 135.775 ;
        RECT 57.410 135.105 58.075 135.275 ;
        RECT 57.410 134.115 57.640 135.105 ;
        RECT 57.810 134.285 58.160 134.935 ;
        RECT 58.335 134.805 58.605 135.775 ;
        RECT 58.815 135.145 59.095 135.945 ;
        RECT 59.265 135.435 60.920 135.725 ;
        RECT 59.330 135.095 60.920 135.265 ;
        RECT 59.330 134.975 59.500 135.095 ;
        RECT 58.775 134.805 59.500 134.975 ;
        RECT 57.410 133.945 58.075 134.115 ;
        RECT 57.405 133.395 57.735 133.775 ;
        RECT 57.905 133.655 58.075 133.945 ;
        RECT 58.335 134.070 58.505 134.805 ;
        RECT 58.775 134.635 58.945 134.805 ;
        RECT 59.690 134.755 60.405 134.925 ;
        RECT 60.600 134.805 60.920 135.095 ;
        RECT 61.555 134.780 61.845 135.945 ;
        RECT 62.390 135.605 62.645 135.635 ;
        RECT 62.305 135.435 62.645 135.605 ;
        RECT 62.390 134.965 62.645 135.435 ;
        RECT 62.825 135.145 63.110 135.945 ;
        RECT 63.290 135.225 63.620 135.735 ;
        RECT 58.675 134.305 58.945 134.635 ;
        RECT 59.115 134.305 59.520 134.635 ;
        RECT 59.690 134.305 60.400 134.755 ;
        RECT 58.775 134.135 58.945 134.305 ;
        RECT 58.335 133.725 58.605 134.070 ;
        RECT 58.775 133.965 60.385 134.135 ;
        RECT 60.570 134.065 60.920 134.635 ;
        RECT 58.795 133.395 59.175 133.795 ;
        RECT 59.345 133.615 59.515 133.965 ;
        RECT 59.685 133.395 60.015 133.795 ;
        RECT 60.215 133.615 60.385 133.965 ;
        RECT 60.585 133.395 60.915 133.895 ;
        RECT 61.555 133.395 61.845 134.120 ;
        RECT 62.390 134.105 62.570 134.965 ;
        RECT 63.290 134.635 63.540 135.225 ;
        RECT 63.890 135.075 64.060 135.685 ;
        RECT 64.230 135.255 64.560 135.945 ;
        RECT 64.790 135.395 65.030 135.685 ;
        RECT 65.230 135.565 65.650 135.945 ;
        RECT 65.830 135.475 66.460 135.725 ;
        RECT 66.930 135.565 67.260 135.945 ;
        RECT 65.830 135.395 66.000 135.475 ;
        RECT 67.430 135.395 67.600 135.685 ;
        RECT 67.780 135.565 68.160 135.945 ;
        RECT 68.400 135.560 69.230 135.730 ;
        RECT 64.790 135.225 66.000 135.395 ;
        RECT 62.740 134.305 63.540 134.635 ;
        RECT 62.390 133.575 62.645 134.105 ;
        RECT 62.825 133.395 63.110 133.855 ;
        RECT 63.290 133.655 63.540 134.305 ;
        RECT 63.740 135.055 64.060 135.075 ;
        RECT 63.740 134.885 65.660 135.055 ;
        RECT 63.740 133.990 63.930 134.885 ;
        RECT 65.830 134.715 66.000 135.225 ;
        RECT 66.170 134.965 66.690 135.275 ;
        RECT 64.100 134.545 66.000 134.715 ;
        RECT 64.100 134.485 64.430 134.545 ;
        RECT 64.580 134.315 64.910 134.375 ;
        RECT 64.250 134.045 64.910 134.315 ;
        RECT 63.740 133.660 64.060 133.990 ;
        RECT 64.240 133.395 64.900 133.875 ;
        RECT 65.100 133.785 65.270 134.545 ;
        RECT 66.170 134.375 66.350 134.785 ;
        RECT 65.440 134.205 65.770 134.325 ;
        RECT 66.520 134.205 66.690 134.965 ;
        RECT 65.440 134.035 66.690 134.205 ;
        RECT 66.860 135.145 68.230 135.395 ;
        RECT 66.860 134.375 67.050 135.145 ;
        RECT 67.980 134.885 68.230 135.145 ;
        RECT 67.220 134.715 67.470 134.875 ;
        RECT 68.400 134.715 68.570 135.560 ;
        RECT 69.465 135.275 69.635 135.775 ;
        RECT 69.805 135.445 70.135 135.945 ;
        RECT 68.740 134.885 69.240 135.265 ;
        RECT 69.465 135.105 70.160 135.275 ;
        RECT 67.220 134.545 68.570 134.715 ;
        RECT 68.150 134.505 68.570 134.545 ;
        RECT 66.860 134.035 67.280 134.375 ;
        RECT 67.570 134.045 67.980 134.375 ;
        RECT 65.100 133.615 65.950 133.785 ;
        RECT 66.510 133.395 66.830 133.855 ;
        RECT 67.030 133.605 67.280 134.035 ;
        RECT 67.570 133.395 67.980 133.835 ;
        RECT 68.150 133.775 68.320 134.505 ;
        RECT 68.490 133.955 68.840 134.325 ;
        RECT 69.020 134.015 69.240 134.885 ;
        RECT 69.410 134.315 69.820 134.935 ;
        RECT 69.990 134.135 70.160 135.105 ;
        RECT 69.465 133.945 70.160 134.135 ;
        RECT 68.150 133.575 69.165 133.775 ;
        RECT 69.465 133.615 69.635 133.945 ;
        RECT 69.805 133.395 70.135 133.775 ;
        RECT 70.350 133.655 70.575 135.775 ;
        RECT 70.745 135.445 71.075 135.945 ;
        RECT 71.245 135.275 71.415 135.775 ;
        RECT 72.050 135.605 72.305 135.635 ;
        RECT 71.965 135.435 72.305 135.605 ;
        RECT 70.750 135.105 71.415 135.275 ;
        RECT 70.750 134.115 70.980 135.105 ;
        RECT 72.050 134.965 72.305 135.435 ;
        RECT 72.485 135.145 72.770 135.945 ;
        RECT 72.950 135.225 73.280 135.735 ;
        RECT 71.150 134.285 71.500 134.935 ;
        RECT 70.750 133.945 71.415 134.115 ;
        RECT 70.745 133.395 71.075 133.775 ;
        RECT 71.245 133.655 71.415 133.945 ;
        RECT 72.050 134.105 72.230 134.965 ;
        RECT 72.950 134.635 73.200 135.225 ;
        RECT 73.550 135.075 73.720 135.685 ;
        RECT 73.890 135.255 74.220 135.945 ;
        RECT 74.450 135.395 74.690 135.685 ;
        RECT 74.890 135.565 75.310 135.945 ;
        RECT 75.490 135.475 76.120 135.725 ;
        RECT 76.590 135.565 76.920 135.945 ;
        RECT 75.490 135.395 75.660 135.475 ;
        RECT 77.090 135.395 77.260 135.685 ;
        RECT 77.440 135.565 77.820 135.945 ;
        RECT 78.060 135.560 78.890 135.730 ;
        RECT 74.450 135.225 75.660 135.395 ;
        RECT 72.400 134.305 73.200 134.635 ;
        RECT 72.050 133.575 72.305 134.105 ;
        RECT 72.485 133.395 72.770 133.855 ;
        RECT 72.950 133.655 73.200 134.305 ;
        RECT 73.400 135.055 73.720 135.075 ;
        RECT 73.400 134.885 75.320 135.055 ;
        RECT 73.400 133.990 73.590 134.885 ;
        RECT 75.490 134.715 75.660 135.225 ;
        RECT 75.830 134.965 76.350 135.275 ;
        RECT 73.760 134.545 75.660 134.715 ;
        RECT 73.760 134.485 74.090 134.545 ;
        RECT 74.240 134.315 74.570 134.375 ;
        RECT 73.910 134.045 74.570 134.315 ;
        RECT 73.400 133.660 73.720 133.990 ;
        RECT 73.900 133.395 74.560 133.875 ;
        RECT 74.760 133.785 74.930 134.545 ;
        RECT 75.830 134.375 76.010 134.785 ;
        RECT 75.100 134.205 75.430 134.325 ;
        RECT 76.180 134.205 76.350 134.965 ;
        RECT 75.100 134.035 76.350 134.205 ;
        RECT 76.520 135.145 77.890 135.395 ;
        RECT 76.520 134.375 76.710 135.145 ;
        RECT 77.640 134.885 77.890 135.145 ;
        RECT 76.880 134.715 77.130 134.875 ;
        RECT 78.060 134.715 78.230 135.560 ;
        RECT 79.125 135.275 79.295 135.775 ;
        RECT 79.465 135.445 79.795 135.945 ;
        RECT 78.400 134.885 78.900 135.265 ;
        RECT 79.125 135.105 79.820 135.275 ;
        RECT 76.880 134.545 78.230 134.715 ;
        RECT 77.810 134.505 78.230 134.545 ;
        RECT 76.520 134.035 76.940 134.375 ;
        RECT 77.230 134.045 77.640 134.375 ;
        RECT 74.760 133.615 75.610 133.785 ;
        RECT 76.170 133.395 76.490 133.855 ;
        RECT 76.690 133.605 76.940 134.035 ;
        RECT 77.230 133.395 77.640 133.835 ;
        RECT 77.810 133.775 77.980 134.505 ;
        RECT 78.150 133.955 78.500 134.325 ;
        RECT 78.680 134.015 78.900 134.885 ;
        RECT 79.070 134.315 79.480 134.935 ;
        RECT 79.650 134.135 79.820 135.105 ;
        RECT 79.125 133.945 79.820 134.135 ;
        RECT 77.810 133.575 78.825 133.775 ;
        RECT 79.125 133.615 79.295 133.945 ;
        RECT 79.465 133.395 79.795 133.775 ;
        RECT 80.010 133.655 80.235 135.775 ;
        RECT 80.405 135.445 80.735 135.945 ;
        RECT 80.905 135.275 81.075 135.775 ;
        RECT 80.410 135.105 81.075 135.275 ;
        RECT 80.410 134.115 80.640 135.105 ;
        RECT 80.810 134.285 81.160 134.935 ;
        RECT 81.340 134.805 81.675 135.775 ;
        RECT 81.845 134.805 82.015 135.945 ;
        RECT 82.185 135.605 84.215 135.775 ;
        RECT 81.340 134.135 81.510 134.805 ;
        RECT 82.185 134.635 82.355 135.605 ;
        RECT 81.680 134.305 81.935 134.635 ;
        RECT 82.160 134.305 82.355 134.635 ;
        RECT 82.525 135.265 83.650 135.435 ;
        RECT 81.765 134.135 81.935 134.305 ;
        RECT 82.525 134.135 82.695 135.265 ;
        RECT 80.410 133.945 81.075 134.115 ;
        RECT 80.405 133.395 80.735 133.775 ;
        RECT 80.905 133.655 81.075 133.945 ;
        RECT 81.340 133.565 81.595 134.135 ;
        RECT 81.765 133.965 82.695 134.135 ;
        RECT 82.865 134.925 83.875 135.095 ;
        RECT 82.865 134.125 83.035 134.925 ;
        RECT 82.520 133.930 82.695 133.965 ;
        RECT 81.765 133.395 82.095 133.795 ;
        RECT 82.520 133.565 83.050 133.930 ;
        RECT 83.240 133.905 83.515 134.725 ;
        RECT 83.235 133.735 83.515 133.905 ;
        RECT 83.240 133.565 83.515 133.735 ;
        RECT 83.685 133.565 83.875 134.925 ;
        RECT 84.045 134.940 84.215 135.605 ;
        RECT 84.385 135.185 84.555 135.945 ;
        RECT 84.790 135.185 85.305 135.595 ;
        RECT 84.045 134.750 84.795 134.940 ;
        RECT 84.965 134.375 85.305 135.185 ;
        RECT 84.075 134.205 85.305 134.375 ;
        RECT 85.475 134.870 85.745 135.775 ;
        RECT 85.915 135.185 86.245 135.945 ;
        RECT 86.425 135.015 86.595 135.775 ;
        RECT 84.055 133.395 84.565 133.930 ;
        RECT 84.785 133.600 85.030 134.205 ;
        RECT 85.475 134.070 85.645 134.870 ;
        RECT 85.930 134.845 86.595 135.015 ;
        RECT 85.930 134.700 86.100 134.845 ;
        RECT 87.315 134.780 87.605 135.945 ;
        RECT 88.150 135.605 88.405 135.635 ;
        RECT 88.065 135.435 88.405 135.605 ;
        RECT 88.150 134.965 88.405 135.435 ;
        RECT 88.585 135.145 88.870 135.945 ;
        RECT 89.050 135.225 89.380 135.735 ;
        RECT 85.815 134.370 86.100 134.700 ;
        RECT 85.930 134.115 86.100 134.370 ;
        RECT 86.335 134.295 86.665 134.665 ;
        RECT 85.475 133.565 85.735 134.070 ;
        RECT 85.930 133.945 86.595 134.115 ;
        RECT 85.915 133.395 86.245 133.775 ;
        RECT 86.425 133.565 86.595 133.945 ;
        RECT 87.315 133.395 87.605 134.120 ;
        RECT 88.150 134.105 88.330 134.965 ;
        RECT 89.050 134.635 89.300 135.225 ;
        RECT 89.650 135.075 89.820 135.685 ;
        RECT 89.990 135.255 90.320 135.945 ;
        RECT 90.550 135.395 90.790 135.685 ;
        RECT 90.990 135.565 91.410 135.945 ;
        RECT 91.590 135.475 92.220 135.725 ;
        RECT 92.690 135.565 93.020 135.945 ;
        RECT 91.590 135.395 91.760 135.475 ;
        RECT 93.190 135.395 93.360 135.685 ;
        RECT 93.540 135.565 93.920 135.945 ;
        RECT 94.160 135.560 94.990 135.730 ;
        RECT 90.550 135.225 91.760 135.395 ;
        RECT 88.500 134.305 89.300 134.635 ;
        RECT 88.150 133.575 88.405 134.105 ;
        RECT 88.585 133.395 88.870 133.855 ;
        RECT 89.050 133.655 89.300 134.305 ;
        RECT 89.500 135.055 89.820 135.075 ;
        RECT 89.500 134.885 91.420 135.055 ;
        RECT 89.500 133.990 89.690 134.885 ;
        RECT 91.590 134.715 91.760 135.225 ;
        RECT 91.930 134.965 92.450 135.275 ;
        RECT 89.860 134.545 91.760 134.715 ;
        RECT 89.860 134.485 90.190 134.545 ;
        RECT 90.340 134.315 90.670 134.375 ;
        RECT 90.010 134.045 90.670 134.315 ;
        RECT 89.500 133.660 89.820 133.990 ;
        RECT 90.000 133.395 90.660 133.875 ;
        RECT 90.860 133.785 91.030 134.545 ;
        RECT 91.930 134.375 92.110 134.785 ;
        RECT 91.200 134.205 91.530 134.325 ;
        RECT 92.280 134.205 92.450 134.965 ;
        RECT 91.200 134.035 92.450 134.205 ;
        RECT 92.620 135.145 93.990 135.395 ;
        RECT 92.620 134.375 92.810 135.145 ;
        RECT 93.740 134.885 93.990 135.145 ;
        RECT 92.980 134.715 93.230 134.875 ;
        RECT 94.160 134.715 94.330 135.560 ;
        RECT 95.225 135.275 95.395 135.775 ;
        RECT 95.565 135.445 95.895 135.945 ;
        RECT 94.500 134.885 95.000 135.265 ;
        RECT 95.225 135.105 95.920 135.275 ;
        RECT 92.980 134.545 94.330 134.715 ;
        RECT 93.910 134.505 94.330 134.545 ;
        RECT 92.620 134.035 93.040 134.375 ;
        RECT 93.330 134.045 93.740 134.375 ;
        RECT 90.860 133.615 91.710 133.785 ;
        RECT 92.270 133.395 92.590 133.855 ;
        RECT 92.790 133.605 93.040 134.035 ;
        RECT 93.330 133.395 93.740 133.835 ;
        RECT 93.910 133.775 94.080 134.505 ;
        RECT 94.250 133.955 94.600 134.325 ;
        RECT 94.780 134.015 95.000 134.885 ;
        RECT 95.170 134.315 95.580 134.935 ;
        RECT 95.750 134.135 95.920 135.105 ;
        RECT 95.225 133.945 95.920 134.135 ;
        RECT 93.910 133.575 94.925 133.775 ;
        RECT 95.225 133.615 95.395 133.945 ;
        RECT 95.565 133.395 95.895 133.775 ;
        RECT 96.110 133.655 96.335 135.775 ;
        RECT 96.505 135.445 96.835 135.945 ;
        RECT 97.005 135.275 97.175 135.775 ;
        RECT 97.810 135.605 98.065 135.635 ;
        RECT 97.725 135.435 98.065 135.605 ;
        RECT 96.510 135.105 97.175 135.275 ;
        RECT 96.510 134.115 96.740 135.105 ;
        RECT 97.810 134.965 98.065 135.435 ;
        RECT 98.245 135.145 98.530 135.945 ;
        RECT 98.710 135.225 99.040 135.735 ;
        RECT 96.910 134.285 97.260 134.935 ;
        RECT 96.510 133.945 97.175 134.115 ;
        RECT 96.505 133.395 96.835 133.775 ;
        RECT 97.005 133.655 97.175 133.945 ;
        RECT 97.810 134.105 97.990 134.965 ;
        RECT 98.710 134.635 98.960 135.225 ;
        RECT 99.310 135.075 99.480 135.685 ;
        RECT 99.650 135.255 99.980 135.945 ;
        RECT 100.210 135.395 100.450 135.685 ;
        RECT 100.650 135.565 101.070 135.945 ;
        RECT 101.250 135.475 101.880 135.725 ;
        RECT 102.350 135.565 102.680 135.945 ;
        RECT 101.250 135.395 101.420 135.475 ;
        RECT 102.850 135.395 103.020 135.685 ;
        RECT 103.200 135.565 103.580 135.945 ;
        RECT 103.820 135.560 104.650 135.730 ;
        RECT 100.210 135.225 101.420 135.395 ;
        RECT 98.160 134.305 98.960 134.635 ;
        RECT 97.810 133.575 98.065 134.105 ;
        RECT 98.245 133.395 98.530 133.855 ;
        RECT 98.710 133.655 98.960 134.305 ;
        RECT 99.160 135.055 99.480 135.075 ;
        RECT 99.160 134.885 101.080 135.055 ;
        RECT 99.160 133.990 99.350 134.885 ;
        RECT 101.250 134.715 101.420 135.225 ;
        RECT 101.590 134.965 102.110 135.275 ;
        RECT 99.520 134.545 101.420 134.715 ;
        RECT 99.520 134.485 99.850 134.545 ;
        RECT 100.000 134.315 100.330 134.375 ;
        RECT 99.670 134.045 100.330 134.315 ;
        RECT 99.160 133.660 99.480 133.990 ;
        RECT 99.660 133.395 100.320 133.875 ;
        RECT 100.520 133.785 100.690 134.545 ;
        RECT 101.590 134.375 101.770 134.785 ;
        RECT 100.860 134.205 101.190 134.325 ;
        RECT 101.940 134.205 102.110 134.965 ;
        RECT 100.860 134.035 102.110 134.205 ;
        RECT 102.280 135.145 103.650 135.395 ;
        RECT 102.280 134.375 102.470 135.145 ;
        RECT 103.400 134.885 103.650 135.145 ;
        RECT 102.640 134.715 102.890 134.875 ;
        RECT 103.820 134.715 103.990 135.560 ;
        RECT 104.885 135.275 105.055 135.775 ;
        RECT 105.225 135.445 105.555 135.945 ;
        RECT 104.160 134.885 104.660 135.265 ;
        RECT 104.885 135.105 105.580 135.275 ;
        RECT 102.640 134.545 103.990 134.715 ;
        RECT 103.570 134.505 103.990 134.545 ;
        RECT 102.280 134.035 102.700 134.375 ;
        RECT 102.990 134.045 103.400 134.375 ;
        RECT 100.520 133.615 101.370 133.785 ;
        RECT 101.930 133.395 102.250 133.855 ;
        RECT 102.450 133.605 102.700 134.035 ;
        RECT 102.990 133.395 103.400 133.835 ;
        RECT 103.570 133.775 103.740 134.505 ;
        RECT 103.910 133.955 104.260 134.325 ;
        RECT 104.440 134.015 104.660 134.885 ;
        RECT 104.830 134.315 105.240 134.935 ;
        RECT 105.410 134.135 105.580 135.105 ;
        RECT 104.885 133.945 105.580 134.135 ;
        RECT 103.570 133.575 104.585 133.775 ;
        RECT 104.885 133.615 105.055 133.945 ;
        RECT 105.225 133.395 105.555 133.775 ;
        RECT 105.770 133.655 105.995 135.775 ;
        RECT 106.165 135.445 106.495 135.945 ;
        RECT 106.665 135.275 106.835 135.775 ;
        RECT 106.170 135.105 106.835 135.275 ;
        RECT 106.170 134.115 106.400 135.105 ;
        RECT 106.570 134.285 106.920 134.935 ;
        RECT 107.135 134.805 107.365 135.945 ;
        RECT 107.535 134.795 107.865 135.775 ;
        RECT 108.035 134.805 108.245 135.945 ;
        RECT 108.935 134.855 110.605 135.945 ;
        RECT 110.775 134.870 111.045 135.775 ;
        RECT 111.215 135.185 111.545 135.945 ;
        RECT 111.725 135.015 111.905 135.775 ;
        RECT 107.115 134.385 107.445 134.635 ;
        RECT 106.170 133.945 106.835 134.115 ;
        RECT 106.165 133.395 106.495 133.775 ;
        RECT 106.665 133.655 106.835 133.945 ;
        RECT 107.135 133.395 107.365 134.215 ;
        RECT 107.615 134.195 107.865 134.795 ;
        RECT 108.935 134.335 109.685 134.855 ;
        RECT 107.535 133.565 107.865 134.195 ;
        RECT 108.035 133.395 108.245 134.215 ;
        RECT 109.855 134.165 110.605 134.685 ;
        RECT 108.935 133.395 110.605 134.165 ;
        RECT 110.775 134.070 110.955 134.870 ;
        RECT 111.230 134.845 111.905 135.015 ;
        RECT 112.155 134.855 113.365 135.945 ;
        RECT 111.230 134.700 111.400 134.845 ;
        RECT 111.125 134.370 111.400 134.700 ;
        RECT 111.230 134.115 111.400 134.370 ;
        RECT 111.625 134.295 111.965 134.665 ;
        RECT 112.155 134.315 112.675 134.855 ;
        RECT 112.845 134.145 113.365 134.685 ;
        RECT 110.775 133.565 111.035 134.070 ;
        RECT 111.230 133.945 111.895 134.115 ;
        RECT 111.215 133.395 111.545 133.775 ;
        RECT 111.725 133.565 111.895 133.945 ;
        RECT 112.155 133.395 113.365 134.145 ;
        RECT 26.970 133.225 113.450 133.395 ;
        RECT 27.055 132.475 28.265 133.225 ;
        RECT 28.525 132.675 28.695 133.055 ;
        RECT 28.875 132.845 29.205 133.225 ;
        RECT 28.525 132.505 29.190 132.675 ;
        RECT 29.385 132.550 29.645 133.055 ;
        RECT 30.125 132.755 30.295 133.225 ;
        RECT 30.465 132.575 30.795 133.055 ;
        RECT 30.965 132.755 31.135 133.225 ;
        RECT 31.305 132.575 31.635 133.055 ;
        RECT 27.055 131.935 27.575 132.475 ;
        RECT 27.745 131.765 28.265 132.305 ;
        RECT 28.455 131.955 28.785 132.325 ;
        RECT 29.020 132.250 29.190 132.505 ;
        RECT 29.020 131.920 29.305 132.250 ;
        RECT 29.020 131.775 29.190 131.920 ;
        RECT 27.055 130.675 28.265 131.765 ;
        RECT 28.525 131.605 29.190 131.775 ;
        RECT 29.475 131.750 29.645 132.550 ;
        RECT 28.525 130.845 28.695 131.605 ;
        RECT 28.875 130.675 29.205 131.435 ;
        RECT 29.375 130.845 29.645 131.750 ;
        RECT 29.870 132.405 31.635 132.575 ;
        RECT 31.805 132.415 31.975 133.225 ;
        RECT 32.175 132.845 33.245 133.015 ;
        RECT 32.175 132.490 32.495 132.845 ;
        RECT 29.870 131.855 30.280 132.405 ;
        RECT 32.170 132.235 32.495 132.490 ;
        RECT 30.465 132.025 32.495 132.235 ;
        RECT 32.150 132.015 32.495 132.025 ;
        RECT 32.665 132.275 32.905 132.675 ;
        RECT 33.075 132.615 33.245 132.845 ;
        RECT 33.415 132.785 33.605 133.225 ;
        RECT 33.775 132.775 34.725 133.055 ;
        RECT 34.945 132.865 35.295 133.035 ;
        RECT 33.075 132.445 33.605 132.615 ;
        RECT 29.870 131.685 31.595 131.855 ;
        RECT 30.125 130.675 30.295 131.515 ;
        RECT 30.505 130.845 30.755 131.685 ;
        RECT 30.965 130.675 31.135 131.515 ;
        RECT 31.305 130.845 31.595 131.685 ;
        RECT 31.805 130.675 31.975 131.735 ;
        RECT 32.150 131.395 32.320 132.015 ;
        RECT 32.665 131.905 33.205 132.275 ;
        RECT 33.385 132.165 33.605 132.445 ;
        RECT 33.775 131.995 33.945 132.775 ;
        RECT 33.540 131.825 33.945 131.995 ;
        RECT 34.115 131.985 34.465 132.605 ;
        RECT 33.540 131.735 33.710 131.825 ;
        RECT 34.635 131.815 34.845 132.605 ;
        RECT 32.490 131.565 33.710 131.735 ;
        RECT 34.170 131.655 34.845 131.815 ;
        RECT 32.150 131.225 32.950 131.395 ;
        RECT 32.270 130.675 32.600 131.055 ;
        RECT 32.780 130.935 32.950 131.225 ;
        RECT 33.540 131.185 33.710 131.565 ;
        RECT 33.880 131.645 34.845 131.655 ;
        RECT 35.035 132.475 35.295 132.865 ;
        RECT 35.505 132.765 35.835 133.225 ;
        RECT 36.710 132.835 37.565 133.005 ;
        RECT 37.770 132.835 38.265 133.005 ;
        RECT 38.435 132.865 38.765 133.225 ;
        RECT 35.035 131.785 35.205 132.475 ;
        RECT 35.375 132.125 35.545 132.305 ;
        RECT 35.715 132.295 36.505 132.545 ;
        RECT 36.710 132.125 36.880 132.835 ;
        RECT 37.050 132.325 37.405 132.545 ;
        RECT 35.375 131.955 37.065 132.125 ;
        RECT 33.880 131.355 34.340 131.645 ;
        RECT 35.035 131.615 36.535 131.785 ;
        RECT 35.035 131.475 35.205 131.615 ;
        RECT 34.645 131.305 35.205 131.475 ;
        RECT 33.120 130.675 33.370 131.135 ;
        RECT 33.540 130.845 34.410 131.185 ;
        RECT 34.645 130.845 34.815 131.305 ;
        RECT 35.650 131.275 36.725 131.445 ;
        RECT 34.985 130.675 35.355 131.135 ;
        RECT 35.650 130.935 35.820 131.275 ;
        RECT 35.990 130.675 36.320 131.105 ;
        RECT 36.555 130.935 36.725 131.275 ;
        RECT 36.895 131.175 37.065 131.955 ;
        RECT 37.235 131.735 37.405 132.325 ;
        RECT 37.575 131.925 37.925 132.545 ;
        RECT 37.235 131.345 37.700 131.735 ;
        RECT 38.095 131.475 38.265 132.835 ;
        RECT 38.435 131.645 38.895 132.695 ;
        RECT 37.870 131.305 38.265 131.475 ;
        RECT 37.870 131.175 38.040 131.305 ;
        RECT 36.895 130.845 37.575 131.175 ;
        RECT 37.790 130.845 38.040 131.175 ;
        RECT 38.210 130.675 38.460 131.135 ;
        RECT 38.630 130.860 38.955 131.645 ;
        RECT 39.125 130.845 39.295 132.965 ;
        RECT 39.465 132.845 39.795 133.225 ;
        RECT 39.965 132.675 40.220 132.965 ;
        RECT 39.470 132.505 40.220 132.675 ;
        RECT 39.470 131.515 39.700 132.505 ;
        RECT 40.400 132.485 40.655 133.055 ;
        RECT 40.825 132.825 41.155 133.225 ;
        RECT 41.580 132.690 42.110 133.055 ;
        RECT 42.300 132.885 42.575 133.055 ;
        RECT 42.295 132.715 42.575 132.885 ;
        RECT 41.580 132.655 41.755 132.690 ;
        RECT 40.825 132.485 41.755 132.655 ;
        RECT 39.870 131.685 40.220 132.335 ;
        RECT 40.400 131.815 40.570 132.485 ;
        RECT 40.825 132.315 40.995 132.485 ;
        RECT 40.740 131.985 40.995 132.315 ;
        RECT 41.220 131.985 41.415 132.315 ;
        RECT 39.470 131.345 40.220 131.515 ;
        RECT 39.465 130.675 39.795 131.175 ;
        RECT 39.965 130.845 40.220 131.345 ;
        RECT 40.400 130.845 40.735 131.815 ;
        RECT 40.905 130.675 41.075 131.815 ;
        RECT 41.245 131.015 41.415 131.985 ;
        RECT 41.585 131.355 41.755 132.485 ;
        RECT 41.925 131.695 42.095 132.495 ;
        RECT 42.300 131.895 42.575 132.715 ;
        RECT 42.745 131.695 42.935 133.055 ;
        RECT 43.115 132.690 43.625 133.225 ;
        RECT 43.845 132.415 44.090 133.020 ;
        RECT 44.540 132.485 44.795 133.055 ;
        RECT 44.965 132.825 45.295 133.225 ;
        RECT 45.720 132.690 46.250 133.055 ;
        RECT 46.440 132.885 46.715 133.055 ;
        RECT 46.435 132.715 46.715 132.885 ;
        RECT 45.720 132.655 45.895 132.690 ;
        RECT 44.965 132.485 45.895 132.655 ;
        RECT 43.135 132.245 44.365 132.415 ;
        RECT 41.925 131.525 42.935 131.695 ;
        RECT 43.105 131.680 43.855 131.870 ;
        RECT 41.585 131.185 42.710 131.355 ;
        RECT 43.105 131.015 43.275 131.680 ;
        RECT 44.025 131.435 44.365 132.245 ;
        RECT 41.245 130.845 43.275 131.015 ;
        RECT 43.445 130.675 43.615 131.435 ;
        RECT 43.850 131.025 44.365 131.435 ;
        RECT 44.540 131.815 44.710 132.485 ;
        RECT 44.965 132.315 45.135 132.485 ;
        RECT 44.880 131.985 45.135 132.315 ;
        RECT 45.360 131.985 45.555 132.315 ;
        RECT 44.540 130.845 44.875 131.815 ;
        RECT 45.045 130.675 45.215 131.815 ;
        RECT 45.385 131.015 45.555 131.985 ;
        RECT 45.725 131.355 45.895 132.485 ;
        RECT 46.065 131.695 46.235 132.495 ;
        RECT 46.440 131.895 46.715 132.715 ;
        RECT 46.885 131.695 47.075 133.055 ;
        RECT 47.255 132.690 47.765 133.225 ;
        RECT 47.985 132.415 48.230 133.020 ;
        RECT 48.675 132.500 48.965 133.225 ;
        RECT 49.410 132.415 49.655 133.020 ;
        RECT 49.875 132.690 50.385 133.225 ;
        RECT 47.275 132.245 48.505 132.415 ;
        RECT 46.065 131.525 47.075 131.695 ;
        RECT 47.245 131.680 47.995 131.870 ;
        RECT 45.725 131.185 46.850 131.355 ;
        RECT 47.245 131.015 47.415 131.680 ;
        RECT 48.165 131.435 48.505 132.245 ;
        RECT 49.135 132.245 50.365 132.415 ;
        RECT 45.385 130.845 47.415 131.015 ;
        RECT 47.585 130.675 47.755 131.435 ;
        RECT 47.990 131.025 48.505 131.435 ;
        RECT 48.675 130.675 48.965 131.840 ;
        RECT 49.135 131.435 49.475 132.245 ;
        RECT 49.645 131.680 50.395 131.870 ;
        RECT 49.135 131.025 49.650 131.435 ;
        RECT 49.885 130.675 50.055 131.435 ;
        RECT 50.225 131.015 50.395 131.680 ;
        RECT 50.565 131.695 50.755 133.055 ;
        RECT 50.925 132.885 51.200 133.055 ;
        RECT 50.925 132.715 51.205 132.885 ;
        RECT 50.925 131.895 51.200 132.715 ;
        RECT 51.390 132.690 51.920 133.055 ;
        RECT 52.345 132.825 52.675 133.225 ;
        RECT 51.745 132.655 51.920 132.690 ;
        RECT 51.405 131.695 51.575 132.495 ;
        RECT 50.565 131.525 51.575 131.695 ;
        RECT 51.745 132.485 52.675 132.655 ;
        RECT 52.845 132.485 53.100 133.055 ;
        RECT 53.650 132.885 53.905 133.045 ;
        RECT 53.565 132.715 53.905 132.885 ;
        RECT 54.085 132.765 54.370 133.225 ;
        RECT 51.745 131.355 51.915 132.485 ;
        RECT 52.505 132.315 52.675 132.485 ;
        RECT 50.790 131.185 51.915 131.355 ;
        RECT 52.085 131.985 52.280 132.315 ;
        RECT 52.505 131.985 52.760 132.315 ;
        RECT 52.085 131.015 52.255 131.985 ;
        RECT 52.930 131.815 53.100 132.485 ;
        RECT 50.225 130.845 52.255 131.015 ;
        RECT 52.425 130.675 52.595 131.815 ;
        RECT 52.765 130.845 53.100 131.815 ;
        RECT 53.650 132.515 53.905 132.715 ;
        RECT 53.650 131.655 53.830 132.515 ;
        RECT 54.550 132.315 54.800 132.965 ;
        RECT 54.000 131.985 54.800 132.315 ;
        RECT 53.650 130.985 53.905 131.655 ;
        RECT 54.085 130.675 54.370 131.475 ;
        RECT 54.550 131.395 54.800 131.985 ;
        RECT 55.000 132.630 55.320 132.960 ;
        RECT 55.500 132.745 56.160 133.225 ;
        RECT 56.360 132.835 57.210 133.005 ;
        RECT 55.000 131.735 55.190 132.630 ;
        RECT 55.510 132.305 56.170 132.575 ;
        RECT 55.840 132.245 56.170 132.305 ;
        RECT 55.360 132.075 55.690 132.135 ;
        RECT 56.360 132.075 56.530 132.835 ;
        RECT 57.770 132.765 58.090 133.225 ;
        RECT 58.290 132.585 58.540 133.015 ;
        RECT 58.830 132.785 59.240 133.225 ;
        RECT 59.410 132.845 60.425 133.045 ;
        RECT 56.700 132.415 57.950 132.585 ;
        RECT 56.700 132.295 57.030 132.415 ;
        RECT 55.360 131.905 57.260 132.075 ;
        RECT 55.000 131.565 56.920 131.735 ;
        RECT 55.000 131.545 55.320 131.565 ;
        RECT 54.550 130.885 54.880 131.395 ;
        RECT 55.150 130.935 55.320 131.545 ;
        RECT 57.090 131.395 57.260 131.905 ;
        RECT 57.430 131.835 57.610 132.245 ;
        RECT 57.780 131.655 57.950 132.415 ;
        RECT 55.490 130.675 55.820 131.365 ;
        RECT 56.050 131.225 57.260 131.395 ;
        RECT 57.430 131.345 57.950 131.655 ;
        RECT 58.120 132.245 58.540 132.585 ;
        RECT 58.830 132.245 59.240 132.575 ;
        RECT 58.120 131.475 58.310 132.245 ;
        RECT 59.410 132.115 59.580 132.845 ;
        RECT 60.725 132.675 60.895 133.005 ;
        RECT 61.065 132.845 61.395 133.225 ;
        RECT 59.750 132.295 60.100 132.665 ;
        RECT 59.410 132.075 59.830 132.115 ;
        RECT 58.480 131.905 59.830 132.075 ;
        RECT 58.480 131.745 58.730 131.905 ;
        RECT 59.240 131.475 59.490 131.735 ;
        RECT 58.120 131.225 59.490 131.475 ;
        RECT 56.050 130.935 56.290 131.225 ;
        RECT 57.090 131.145 57.260 131.225 ;
        RECT 56.490 130.675 56.910 131.055 ;
        RECT 57.090 130.895 57.720 131.145 ;
        RECT 58.190 130.675 58.520 131.055 ;
        RECT 58.690 130.935 58.860 131.225 ;
        RECT 59.660 131.060 59.830 131.905 ;
        RECT 60.280 131.735 60.500 132.605 ;
        RECT 60.725 132.485 61.420 132.675 ;
        RECT 60.000 131.355 60.500 131.735 ;
        RECT 60.670 131.685 61.080 132.305 ;
        RECT 61.250 131.515 61.420 132.485 ;
        RECT 60.725 131.345 61.420 131.515 ;
        RECT 59.040 130.675 59.420 131.055 ;
        RECT 59.660 130.890 60.490 131.060 ;
        RECT 60.725 130.845 60.895 131.345 ;
        RECT 61.065 130.675 61.395 131.175 ;
        RECT 61.610 130.845 61.835 132.965 ;
        RECT 62.005 132.845 62.335 133.225 ;
        RECT 62.505 132.675 62.675 132.965 ;
        RECT 62.010 132.505 62.675 132.675 ;
        RECT 62.010 131.515 62.240 132.505 ;
        RECT 63.210 132.415 63.455 133.020 ;
        RECT 63.675 132.690 64.185 133.225 ;
        RECT 62.410 131.685 62.760 132.335 ;
        RECT 62.935 132.245 64.165 132.415 ;
        RECT 62.010 131.345 62.675 131.515 ;
        RECT 62.005 130.675 62.335 131.175 ;
        RECT 62.505 130.845 62.675 131.345 ;
        RECT 62.935 131.435 63.275 132.245 ;
        RECT 63.445 131.680 64.195 131.870 ;
        RECT 62.935 131.025 63.450 131.435 ;
        RECT 63.685 130.675 63.855 131.435 ;
        RECT 64.025 131.015 64.195 131.680 ;
        RECT 64.365 131.695 64.555 133.055 ;
        RECT 64.725 132.885 65.000 133.055 ;
        RECT 64.725 132.715 65.005 132.885 ;
        RECT 64.725 131.895 65.000 132.715 ;
        RECT 65.190 132.690 65.720 133.055 ;
        RECT 66.145 132.825 66.475 133.225 ;
        RECT 65.545 132.655 65.720 132.690 ;
        RECT 65.205 131.695 65.375 132.495 ;
        RECT 64.365 131.525 65.375 131.695 ;
        RECT 65.545 132.485 66.475 132.655 ;
        RECT 66.645 132.485 66.900 133.055 ;
        RECT 67.165 132.675 67.335 133.055 ;
        RECT 67.515 132.845 67.845 133.225 ;
        RECT 67.165 132.505 67.830 132.675 ;
        RECT 68.025 132.550 68.285 133.055 ;
        RECT 65.545 131.355 65.715 132.485 ;
        RECT 66.305 132.315 66.475 132.485 ;
        RECT 64.590 131.185 65.715 131.355 ;
        RECT 65.885 131.985 66.080 132.315 ;
        RECT 66.305 131.985 66.560 132.315 ;
        RECT 65.885 131.015 66.055 131.985 ;
        RECT 66.730 131.815 66.900 132.485 ;
        RECT 67.095 131.955 67.425 132.325 ;
        RECT 67.660 132.250 67.830 132.505 ;
        RECT 64.025 130.845 66.055 131.015 ;
        RECT 66.225 130.675 66.395 131.815 ;
        RECT 66.565 130.845 66.900 131.815 ;
        RECT 67.660 131.920 67.945 132.250 ;
        RECT 67.660 131.775 67.830 131.920 ;
        RECT 67.165 131.605 67.830 131.775 ;
        RECT 68.115 131.750 68.285 132.550 ;
        RECT 68.915 132.455 71.505 133.225 ;
        RECT 67.165 130.845 67.335 131.605 ;
        RECT 67.515 130.675 67.845 131.435 ;
        RECT 68.015 130.845 68.285 131.750 ;
        RECT 68.915 131.765 70.125 132.285 ;
        RECT 70.295 131.935 71.505 132.455 ;
        RECT 71.715 132.405 71.945 133.225 ;
        RECT 72.115 132.425 72.445 133.055 ;
        RECT 71.695 131.985 72.025 132.235 ;
        RECT 72.195 131.825 72.445 132.425 ;
        RECT 72.615 132.405 72.825 133.225 ;
        RECT 73.095 132.405 73.325 133.225 ;
        RECT 73.495 132.425 73.825 133.055 ;
        RECT 73.075 131.985 73.405 132.235 ;
        RECT 73.575 131.825 73.825 132.425 ;
        RECT 73.995 132.405 74.205 133.225 ;
        RECT 74.435 132.500 74.725 133.225 ;
        RECT 74.985 132.675 75.155 132.965 ;
        RECT 75.325 132.845 75.655 133.225 ;
        RECT 74.985 132.505 75.650 132.675 ;
        RECT 68.915 130.675 71.505 131.765 ;
        RECT 71.715 130.675 71.945 131.815 ;
        RECT 72.115 130.845 72.445 131.825 ;
        RECT 72.615 130.675 72.825 131.815 ;
        RECT 73.095 130.675 73.325 131.815 ;
        RECT 73.495 130.845 73.825 131.825 ;
        RECT 73.995 130.675 74.205 131.815 ;
        RECT 74.435 130.675 74.725 131.840 ;
        RECT 74.900 131.685 75.250 132.335 ;
        RECT 75.420 131.515 75.650 132.505 ;
        RECT 74.985 131.345 75.650 131.515 ;
        RECT 74.985 130.845 75.155 131.345 ;
        RECT 75.325 130.675 75.655 131.175 ;
        RECT 75.825 130.845 76.050 132.965 ;
        RECT 76.265 132.845 76.595 133.225 ;
        RECT 76.765 132.675 76.935 133.005 ;
        RECT 77.235 132.845 78.250 133.045 ;
        RECT 76.240 132.485 76.935 132.675 ;
        RECT 76.240 131.515 76.410 132.485 ;
        RECT 76.580 131.685 76.990 132.305 ;
        RECT 77.160 131.735 77.380 132.605 ;
        RECT 77.560 132.295 77.910 132.665 ;
        RECT 78.080 132.115 78.250 132.845 ;
        RECT 78.420 132.785 78.830 133.225 ;
        RECT 79.120 132.585 79.370 133.015 ;
        RECT 79.570 132.765 79.890 133.225 ;
        RECT 80.450 132.835 81.300 133.005 ;
        RECT 78.420 132.245 78.830 132.575 ;
        RECT 79.120 132.245 79.540 132.585 ;
        RECT 77.830 132.075 78.250 132.115 ;
        RECT 77.830 131.905 79.180 132.075 ;
        RECT 76.240 131.345 76.935 131.515 ;
        RECT 77.160 131.355 77.660 131.735 ;
        RECT 76.265 130.675 76.595 131.175 ;
        RECT 76.765 130.845 76.935 131.345 ;
        RECT 77.830 131.060 78.000 131.905 ;
        RECT 78.930 131.745 79.180 131.905 ;
        RECT 78.170 131.475 78.420 131.735 ;
        RECT 79.350 131.475 79.540 132.245 ;
        RECT 78.170 131.225 79.540 131.475 ;
        RECT 79.710 132.415 80.960 132.585 ;
        RECT 79.710 131.655 79.880 132.415 ;
        RECT 80.630 132.295 80.960 132.415 ;
        RECT 80.050 131.835 80.230 132.245 ;
        RECT 81.130 132.075 81.300 132.835 ;
        RECT 81.500 132.745 82.160 133.225 ;
        RECT 82.340 132.630 82.660 132.960 ;
        RECT 81.490 132.305 82.150 132.575 ;
        RECT 81.490 132.245 81.820 132.305 ;
        RECT 81.970 132.075 82.300 132.135 ;
        RECT 80.400 131.905 82.300 132.075 ;
        RECT 79.710 131.345 80.230 131.655 ;
        RECT 80.400 131.395 80.570 131.905 ;
        RECT 82.470 131.735 82.660 132.630 ;
        RECT 80.740 131.565 82.660 131.735 ;
        RECT 82.340 131.545 82.660 131.565 ;
        RECT 82.860 132.315 83.110 132.965 ;
        RECT 83.290 132.765 83.575 133.225 ;
        RECT 83.755 132.885 84.010 133.045 ;
        RECT 84.930 132.885 85.185 133.045 ;
        RECT 83.755 132.715 84.095 132.885 ;
        RECT 84.845 132.715 85.185 132.885 ;
        RECT 85.365 132.765 85.650 133.225 ;
        RECT 83.755 132.515 84.010 132.715 ;
        RECT 82.860 131.985 83.660 132.315 ;
        RECT 80.400 131.225 81.610 131.395 ;
        RECT 77.170 130.890 78.000 131.060 ;
        RECT 78.240 130.675 78.620 131.055 ;
        RECT 78.800 130.935 78.970 131.225 ;
        RECT 80.400 131.145 80.570 131.225 ;
        RECT 79.140 130.675 79.470 131.055 ;
        RECT 79.940 130.895 80.570 131.145 ;
        RECT 80.750 130.675 81.170 131.055 ;
        RECT 81.370 130.935 81.610 131.225 ;
        RECT 81.840 130.675 82.170 131.365 ;
        RECT 82.340 130.935 82.510 131.545 ;
        RECT 82.860 131.395 83.110 131.985 ;
        RECT 83.830 131.655 84.010 132.515 ;
        RECT 82.780 130.885 83.110 131.395 ;
        RECT 83.290 130.675 83.575 131.475 ;
        RECT 83.755 130.985 84.010 131.655 ;
        RECT 84.930 132.515 85.185 132.715 ;
        RECT 84.930 131.655 85.110 132.515 ;
        RECT 85.830 132.315 86.080 132.965 ;
        RECT 85.280 131.985 86.080 132.315 ;
        RECT 84.930 130.985 85.185 131.655 ;
        RECT 85.365 130.675 85.650 131.475 ;
        RECT 85.830 131.395 86.080 131.985 ;
        RECT 86.280 132.630 86.600 132.960 ;
        RECT 86.780 132.745 87.440 133.225 ;
        RECT 87.640 132.835 88.490 133.005 ;
        RECT 86.280 131.735 86.470 132.630 ;
        RECT 86.790 132.305 87.450 132.575 ;
        RECT 87.120 132.245 87.450 132.305 ;
        RECT 86.640 132.075 86.970 132.135 ;
        RECT 87.640 132.075 87.810 132.835 ;
        RECT 89.050 132.765 89.370 133.225 ;
        RECT 89.570 132.585 89.820 133.015 ;
        RECT 90.110 132.785 90.520 133.225 ;
        RECT 90.690 132.845 91.705 133.045 ;
        RECT 87.980 132.415 89.230 132.585 ;
        RECT 87.980 132.295 88.310 132.415 ;
        RECT 86.640 131.905 88.540 132.075 ;
        RECT 86.280 131.565 88.200 131.735 ;
        RECT 86.280 131.545 86.600 131.565 ;
        RECT 85.830 130.885 86.160 131.395 ;
        RECT 86.430 130.935 86.600 131.545 ;
        RECT 88.370 131.395 88.540 131.905 ;
        RECT 88.710 131.835 88.890 132.245 ;
        RECT 89.060 131.655 89.230 132.415 ;
        RECT 86.770 130.675 87.100 131.365 ;
        RECT 87.330 131.225 88.540 131.395 ;
        RECT 88.710 131.345 89.230 131.655 ;
        RECT 89.400 132.245 89.820 132.585 ;
        RECT 90.110 132.245 90.520 132.575 ;
        RECT 89.400 131.475 89.590 132.245 ;
        RECT 90.690 132.115 90.860 132.845 ;
        RECT 92.005 132.675 92.175 133.005 ;
        RECT 92.345 132.845 92.675 133.225 ;
        RECT 91.030 132.295 91.380 132.665 ;
        RECT 90.690 132.075 91.110 132.115 ;
        RECT 89.760 131.905 91.110 132.075 ;
        RECT 89.760 131.745 90.010 131.905 ;
        RECT 90.520 131.475 90.770 131.735 ;
        RECT 89.400 131.225 90.770 131.475 ;
        RECT 87.330 130.935 87.570 131.225 ;
        RECT 88.370 131.145 88.540 131.225 ;
        RECT 87.770 130.675 88.190 131.055 ;
        RECT 88.370 130.895 89.000 131.145 ;
        RECT 89.470 130.675 89.800 131.055 ;
        RECT 89.970 130.935 90.140 131.225 ;
        RECT 90.940 131.060 91.110 131.905 ;
        RECT 91.560 131.735 91.780 132.605 ;
        RECT 92.005 132.485 92.700 132.675 ;
        RECT 91.280 131.355 91.780 131.735 ;
        RECT 91.950 131.685 92.360 132.305 ;
        RECT 92.530 131.515 92.700 132.485 ;
        RECT 92.005 131.345 92.700 131.515 ;
        RECT 90.320 130.675 90.700 131.055 ;
        RECT 90.940 130.890 91.770 131.060 ;
        RECT 92.005 130.845 92.175 131.345 ;
        RECT 92.345 130.675 92.675 131.175 ;
        RECT 92.890 130.845 93.115 132.965 ;
        RECT 93.285 132.845 93.615 133.225 ;
        RECT 93.785 132.675 93.955 132.965 ;
        RECT 93.290 132.505 93.955 132.675 ;
        RECT 94.305 132.675 94.475 133.055 ;
        RECT 94.655 132.845 94.985 133.225 ;
        RECT 94.305 132.505 94.970 132.675 ;
        RECT 95.165 132.550 95.425 133.055 ;
        RECT 93.290 131.515 93.520 132.505 ;
        RECT 93.690 131.685 94.040 132.335 ;
        RECT 94.235 131.955 94.565 132.325 ;
        RECT 94.800 132.250 94.970 132.505 ;
        RECT 94.800 131.920 95.085 132.250 ;
        RECT 94.800 131.775 94.970 131.920 ;
        RECT 94.305 131.605 94.970 131.775 ;
        RECT 95.255 131.750 95.425 132.550 ;
        RECT 96.330 132.415 96.575 133.020 ;
        RECT 96.795 132.690 97.305 133.225 ;
        RECT 93.290 131.345 93.955 131.515 ;
        RECT 93.285 130.675 93.615 131.175 ;
        RECT 93.785 130.845 93.955 131.345 ;
        RECT 94.305 130.845 94.475 131.605 ;
        RECT 94.655 130.675 94.985 131.435 ;
        RECT 95.155 130.845 95.425 131.750 ;
        RECT 96.055 132.245 97.285 132.415 ;
        RECT 96.055 131.435 96.395 132.245 ;
        RECT 96.565 131.680 97.315 131.870 ;
        RECT 96.055 131.025 96.570 131.435 ;
        RECT 96.805 130.675 96.975 131.435 ;
        RECT 97.145 131.015 97.315 131.680 ;
        RECT 97.485 131.695 97.675 133.055 ;
        RECT 97.845 132.885 98.120 133.055 ;
        RECT 97.845 132.715 98.125 132.885 ;
        RECT 97.845 131.895 98.120 132.715 ;
        RECT 98.310 132.690 98.840 133.055 ;
        RECT 99.265 132.825 99.595 133.225 ;
        RECT 98.665 132.655 98.840 132.690 ;
        RECT 98.325 131.695 98.495 132.495 ;
        RECT 97.485 131.525 98.495 131.695 ;
        RECT 98.665 132.485 99.595 132.655 ;
        RECT 99.765 132.485 100.020 133.055 ;
        RECT 100.195 132.500 100.485 133.225 ;
        RECT 100.745 132.675 100.915 133.055 ;
        RECT 101.095 132.845 101.425 133.225 ;
        RECT 100.745 132.505 101.410 132.675 ;
        RECT 101.605 132.550 101.865 133.055 ;
        RECT 98.665 131.355 98.835 132.485 ;
        RECT 99.425 132.315 99.595 132.485 ;
        RECT 97.710 131.185 98.835 131.355 ;
        RECT 99.005 131.985 99.200 132.315 ;
        RECT 99.425 131.985 99.680 132.315 ;
        RECT 99.005 131.015 99.175 131.985 ;
        RECT 99.850 131.815 100.020 132.485 ;
        RECT 100.675 131.955 101.005 132.325 ;
        RECT 101.240 132.250 101.410 132.505 ;
        RECT 101.240 131.920 101.525 132.250 ;
        RECT 97.145 130.845 99.175 131.015 ;
        RECT 99.345 130.675 99.515 131.815 ;
        RECT 99.685 130.845 100.020 131.815 ;
        RECT 100.195 130.675 100.485 131.840 ;
        RECT 101.240 131.775 101.410 131.920 ;
        RECT 100.745 131.605 101.410 131.775 ;
        RECT 101.695 131.750 101.865 132.550 ;
        RECT 102.995 132.405 103.225 133.225 ;
        RECT 103.395 132.425 103.725 133.055 ;
        RECT 102.975 131.985 103.305 132.235 ;
        RECT 103.475 131.825 103.725 132.425 ;
        RECT 103.895 132.405 104.105 133.225 ;
        RECT 105.345 132.675 105.515 133.055 ;
        RECT 105.695 132.845 106.025 133.225 ;
        RECT 105.345 132.505 106.010 132.675 ;
        RECT 106.205 132.550 106.465 133.055 ;
        RECT 105.275 131.955 105.605 132.325 ;
        RECT 105.840 132.250 106.010 132.505 ;
        RECT 100.745 130.845 100.915 131.605 ;
        RECT 101.095 130.675 101.425 131.435 ;
        RECT 101.595 130.845 101.865 131.750 ;
        RECT 102.995 130.675 103.225 131.815 ;
        RECT 103.395 130.845 103.725 131.825 ;
        RECT 105.840 131.920 106.125 132.250 ;
        RECT 103.895 130.675 104.105 131.815 ;
        RECT 105.840 131.775 106.010 131.920 ;
        RECT 105.345 131.605 106.010 131.775 ;
        RECT 106.295 131.750 106.465 132.550 ;
        RECT 106.675 132.405 106.905 133.225 ;
        RECT 107.075 132.425 107.405 133.055 ;
        RECT 106.655 131.985 106.985 132.235 ;
        RECT 107.155 131.825 107.405 132.425 ;
        RECT 107.575 132.405 107.785 133.225 ;
        RECT 108.935 132.550 109.195 133.055 ;
        RECT 109.375 132.845 109.705 133.225 ;
        RECT 109.885 132.675 110.055 133.055 ;
        RECT 105.345 130.845 105.515 131.605 ;
        RECT 105.695 130.675 106.025 131.435 ;
        RECT 106.195 130.845 106.465 131.750 ;
        RECT 106.675 130.675 106.905 131.815 ;
        RECT 107.075 130.845 107.405 131.825 ;
        RECT 107.575 130.675 107.785 131.815 ;
        RECT 108.935 131.750 109.105 132.550 ;
        RECT 109.390 132.505 110.055 132.675 ;
        RECT 109.390 132.250 109.560 132.505 ;
        RECT 110.355 132.405 110.585 133.225 ;
        RECT 110.755 132.425 111.085 133.055 ;
        RECT 109.275 131.920 109.560 132.250 ;
        RECT 109.795 131.955 110.125 132.325 ;
        RECT 110.335 131.985 110.665 132.235 ;
        RECT 109.390 131.775 109.560 131.920 ;
        RECT 110.835 131.825 111.085 132.425 ;
        RECT 111.255 132.405 111.465 133.225 ;
        RECT 112.155 132.475 113.365 133.225 ;
        RECT 108.935 130.845 109.205 131.750 ;
        RECT 109.390 131.605 110.055 131.775 ;
        RECT 109.375 130.675 109.705 131.435 ;
        RECT 109.885 130.845 110.055 131.605 ;
        RECT 110.355 130.675 110.585 131.815 ;
        RECT 110.755 130.845 111.085 131.825 ;
        RECT 111.255 130.675 111.465 131.815 ;
        RECT 112.155 131.765 112.675 132.305 ;
        RECT 112.845 131.935 113.365 132.475 ;
        RECT 112.155 130.675 113.365 131.765 ;
        RECT 26.970 130.505 113.450 130.675 ;
        RECT 27.055 129.415 28.265 130.505 ;
        RECT 27.055 128.705 27.575 129.245 ;
        RECT 27.745 128.875 28.265 129.415 ;
        RECT 28.525 129.575 28.695 130.335 ;
        RECT 28.875 129.745 29.205 130.505 ;
        RECT 28.525 129.405 29.190 129.575 ;
        RECT 29.375 129.430 29.645 130.335 ;
        RECT 29.020 129.260 29.190 129.405 ;
        RECT 28.455 128.855 28.785 129.225 ;
        RECT 29.020 128.930 29.305 129.260 ;
        RECT 27.055 127.955 28.265 128.705 ;
        RECT 29.020 128.675 29.190 128.930 ;
        RECT 28.525 128.505 29.190 128.675 ;
        RECT 29.475 128.630 29.645 129.430 ;
        RECT 29.855 129.365 30.085 130.505 ;
        RECT 30.255 129.355 30.585 130.335 ;
        RECT 30.755 129.365 30.965 130.505 ;
        RECT 31.695 129.365 31.925 130.505 ;
        RECT 32.095 129.355 32.425 130.335 ;
        RECT 32.595 129.365 32.805 130.505 ;
        RECT 34.045 129.575 34.215 130.335 ;
        RECT 34.395 129.745 34.725 130.505 ;
        RECT 34.045 129.405 34.710 129.575 ;
        RECT 34.895 129.430 35.165 130.335 ;
        RECT 29.835 128.945 30.165 129.195 ;
        RECT 28.525 128.125 28.695 128.505 ;
        RECT 28.875 127.955 29.205 128.335 ;
        RECT 29.385 128.125 29.645 128.630 ;
        RECT 29.855 127.955 30.085 128.775 ;
        RECT 30.335 128.755 30.585 129.355 ;
        RECT 31.675 128.945 32.005 129.195 ;
        RECT 30.255 128.125 30.585 128.755 ;
        RECT 30.755 127.955 30.965 128.775 ;
        RECT 31.695 127.955 31.925 128.775 ;
        RECT 32.175 128.755 32.425 129.355 ;
        RECT 34.540 129.260 34.710 129.405 ;
        RECT 33.975 128.855 34.305 129.225 ;
        RECT 34.540 128.930 34.825 129.260 ;
        RECT 32.095 128.125 32.425 128.755 ;
        RECT 32.595 127.955 32.805 128.775 ;
        RECT 34.540 128.675 34.710 128.930 ;
        RECT 34.045 128.505 34.710 128.675 ;
        RECT 34.995 128.630 35.165 129.430 ;
        RECT 35.795 129.340 36.085 130.505 ;
        RECT 37.215 129.365 37.445 130.505 ;
        RECT 37.615 129.355 37.945 130.335 ;
        RECT 38.115 129.365 38.325 130.505 ;
        RECT 38.645 129.575 38.815 130.335 ;
        RECT 38.995 129.745 39.325 130.505 ;
        RECT 38.645 129.405 39.310 129.575 ;
        RECT 39.495 129.430 39.765 130.335 ;
        RECT 37.195 128.945 37.525 129.195 ;
        RECT 34.045 128.125 34.215 128.505 ;
        RECT 34.395 127.955 34.725 128.335 ;
        RECT 34.905 128.125 35.165 128.630 ;
        RECT 35.795 127.955 36.085 128.680 ;
        RECT 37.215 127.955 37.445 128.775 ;
        RECT 37.695 128.755 37.945 129.355 ;
        RECT 39.140 129.260 39.310 129.405 ;
        RECT 38.575 128.855 38.905 129.225 ;
        RECT 39.140 128.930 39.425 129.260 ;
        RECT 37.615 128.125 37.945 128.755 ;
        RECT 38.115 127.955 38.325 128.775 ;
        RECT 39.140 128.675 39.310 128.930 ;
        RECT 38.645 128.505 39.310 128.675 ;
        RECT 39.595 128.630 39.765 129.430 ;
        RECT 39.975 129.365 40.205 130.505 ;
        RECT 40.375 129.355 40.705 130.335 ;
        RECT 40.875 129.365 41.085 130.505 ;
        RECT 41.315 129.430 41.585 130.335 ;
        RECT 41.755 129.745 42.085 130.505 ;
        RECT 42.265 129.575 42.435 130.335 ;
        RECT 43.005 129.665 43.175 130.505 ;
        RECT 39.955 128.945 40.285 129.195 ;
        RECT 38.645 128.125 38.815 128.505 ;
        RECT 38.995 127.955 39.325 128.335 ;
        RECT 39.505 128.125 39.765 128.630 ;
        RECT 39.975 127.955 40.205 128.775 ;
        RECT 40.455 128.755 40.705 129.355 ;
        RECT 40.375 128.125 40.705 128.755 ;
        RECT 40.875 127.955 41.085 128.775 ;
        RECT 41.315 128.630 41.485 129.430 ;
        RECT 41.770 129.405 42.435 129.575 ;
        RECT 43.385 129.495 43.635 130.335 ;
        RECT 43.845 129.665 44.015 130.505 ;
        RECT 44.185 129.495 44.475 130.335 ;
        RECT 41.770 129.260 41.940 129.405 ;
        RECT 41.655 128.930 41.940 129.260 ;
        RECT 42.750 129.325 44.475 129.495 ;
        RECT 44.685 129.445 44.855 130.505 ;
        RECT 45.150 130.125 45.480 130.505 ;
        RECT 45.660 129.955 45.830 130.245 ;
        RECT 46.000 130.045 46.250 130.505 ;
        RECT 45.030 129.785 45.830 129.955 ;
        RECT 46.420 129.995 47.290 130.335 ;
        RECT 41.770 128.675 41.940 128.930 ;
        RECT 42.175 128.855 42.505 129.225 ;
        RECT 42.750 128.775 43.160 129.325 ;
        RECT 45.030 129.165 45.200 129.785 ;
        RECT 46.420 129.615 46.590 129.995 ;
        RECT 47.525 129.875 47.695 130.335 ;
        RECT 47.865 130.045 48.235 130.505 ;
        RECT 48.530 129.905 48.700 130.245 ;
        RECT 48.870 130.075 49.200 130.505 ;
        RECT 49.435 129.905 49.605 130.245 ;
        RECT 45.370 129.445 46.590 129.615 ;
        RECT 46.760 129.535 47.220 129.825 ;
        RECT 47.525 129.705 48.085 129.875 ;
        RECT 48.530 129.735 49.605 129.905 ;
        RECT 49.775 130.005 50.455 130.335 ;
        RECT 50.670 130.005 50.920 130.335 ;
        RECT 51.090 130.045 51.340 130.505 ;
        RECT 47.915 129.565 48.085 129.705 ;
        RECT 46.760 129.525 47.725 129.535 ;
        RECT 46.420 129.355 46.590 129.445 ;
        RECT 47.050 129.365 47.725 129.525 ;
        RECT 45.030 129.155 45.375 129.165 ;
        RECT 43.345 128.945 45.375 129.155 ;
        RECT 41.315 128.125 41.575 128.630 ;
        RECT 41.770 128.505 42.435 128.675 ;
        RECT 42.750 128.605 44.515 128.775 ;
        RECT 41.755 127.955 42.085 128.335 ;
        RECT 42.265 128.125 42.435 128.505 ;
        RECT 43.005 127.955 43.175 128.425 ;
        RECT 43.345 128.125 43.675 128.605 ;
        RECT 43.845 127.955 44.015 128.425 ;
        RECT 44.185 128.125 44.515 128.605 ;
        RECT 44.685 127.955 44.855 128.765 ;
        RECT 45.050 128.690 45.375 128.945 ;
        RECT 45.055 128.335 45.375 128.690 ;
        RECT 45.545 128.905 46.085 129.275 ;
        RECT 46.420 129.185 46.825 129.355 ;
        RECT 45.545 128.505 45.785 128.905 ;
        RECT 46.265 128.735 46.485 129.015 ;
        RECT 45.955 128.565 46.485 128.735 ;
        RECT 45.955 128.335 46.125 128.565 ;
        RECT 46.655 128.405 46.825 129.185 ;
        RECT 46.995 128.575 47.345 129.195 ;
        RECT 47.515 128.575 47.725 129.365 ;
        RECT 47.915 129.395 49.415 129.565 ;
        RECT 47.915 128.705 48.085 129.395 ;
        RECT 49.775 129.225 49.945 130.005 ;
        RECT 50.750 129.875 50.920 130.005 ;
        RECT 48.255 129.055 49.945 129.225 ;
        RECT 50.115 129.445 50.580 129.835 ;
        RECT 50.750 129.705 51.145 129.875 ;
        RECT 48.255 128.875 48.425 129.055 ;
        RECT 45.055 128.165 46.125 128.335 ;
        RECT 46.295 127.955 46.485 128.395 ;
        RECT 46.655 128.125 47.605 128.405 ;
        RECT 47.915 128.315 48.175 128.705 ;
        RECT 48.595 128.635 49.385 128.885 ;
        RECT 47.825 128.145 48.175 128.315 ;
        RECT 48.385 127.955 48.715 128.415 ;
        RECT 49.590 128.345 49.760 129.055 ;
        RECT 50.115 128.855 50.285 129.445 ;
        RECT 49.930 128.635 50.285 128.855 ;
        RECT 50.455 128.635 50.805 129.255 ;
        RECT 50.975 128.345 51.145 129.705 ;
        RECT 51.510 129.535 51.835 130.320 ;
        RECT 51.315 128.485 51.775 129.535 ;
        RECT 49.590 128.175 50.445 128.345 ;
        RECT 50.650 128.175 51.145 128.345 ;
        RECT 51.315 127.955 51.645 128.315 ;
        RECT 52.005 128.215 52.175 130.335 ;
        RECT 52.345 130.005 52.675 130.505 ;
        RECT 52.845 129.835 53.100 130.335 ;
        RECT 52.350 129.665 53.100 129.835 ;
        RECT 52.350 128.675 52.580 129.665 ;
        RECT 52.750 128.845 53.100 129.495 ;
        RECT 54.235 129.365 54.465 130.505 ;
        RECT 54.635 129.355 54.965 130.335 ;
        RECT 55.135 129.365 55.345 130.505 ;
        RECT 55.665 129.575 55.835 130.335 ;
        RECT 56.015 129.745 56.345 130.505 ;
        RECT 55.665 129.405 56.330 129.575 ;
        RECT 56.515 129.430 56.785 130.335 ;
        RECT 54.215 128.945 54.545 129.195 ;
        RECT 52.350 128.505 53.100 128.675 ;
        RECT 52.345 127.955 52.675 128.335 ;
        RECT 52.845 128.215 53.100 128.505 ;
        RECT 54.235 127.955 54.465 128.775 ;
        RECT 54.715 128.755 54.965 129.355 ;
        RECT 56.160 129.260 56.330 129.405 ;
        RECT 55.595 128.855 55.925 129.225 ;
        RECT 56.160 128.930 56.445 129.260 ;
        RECT 54.635 128.125 54.965 128.755 ;
        RECT 55.135 127.955 55.345 128.775 ;
        RECT 56.160 128.675 56.330 128.930 ;
        RECT 55.665 128.505 56.330 128.675 ;
        RECT 56.615 128.630 56.785 129.430 ;
        RECT 57.045 129.575 57.215 130.335 ;
        RECT 57.395 129.745 57.725 130.505 ;
        RECT 57.045 129.405 57.710 129.575 ;
        RECT 57.895 129.430 58.165 130.335 ;
        RECT 58.535 129.835 58.815 130.505 ;
        RECT 58.985 129.615 59.285 130.165 ;
        RECT 59.485 129.785 59.815 130.505 ;
        RECT 60.005 129.785 60.465 130.335 ;
        RECT 57.540 129.260 57.710 129.405 ;
        RECT 56.975 128.855 57.305 129.225 ;
        RECT 57.540 128.930 57.825 129.260 ;
        RECT 57.540 128.675 57.710 128.930 ;
        RECT 55.665 128.125 55.835 128.505 ;
        RECT 56.015 127.955 56.345 128.335 ;
        RECT 56.525 128.125 56.785 128.630 ;
        RECT 57.045 128.505 57.710 128.675 ;
        RECT 57.995 128.630 58.165 129.430 ;
        RECT 58.350 129.195 58.615 129.555 ;
        RECT 58.985 129.445 59.925 129.615 ;
        RECT 59.755 129.195 59.925 129.445 ;
        RECT 58.350 128.945 59.025 129.195 ;
        RECT 59.245 128.945 59.585 129.195 ;
        RECT 59.755 128.865 60.045 129.195 ;
        RECT 59.755 128.775 59.925 128.865 ;
        RECT 57.045 128.125 57.215 128.505 ;
        RECT 57.395 127.955 57.725 128.335 ;
        RECT 57.905 128.125 58.165 128.630 ;
        RECT 58.535 128.585 59.925 128.775 ;
        RECT 58.535 128.225 58.865 128.585 ;
        RECT 60.215 128.415 60.465 129.785 ;
        RECT 61.555 129.340 61.845 130.505 ;
        RECT 62.475 129.415 64.145 130.505 ;
        RECT 62.475 128.895 63.225 129.415 ;
        RECT 64.375 129.365 64.585 130.505 ;
        RECT 64.755 129.355 65.085 130.335 ;
        RECT 65.255 129.365 65.485 130.505 ;
        RECT 65.695 129.415 69.205 130.505 ;
        RECT 69.380 130.070 74.725 130.505 ;
        RECT 63.395 128.725 64.145 129.245 ;
        RECT 59.485 127.955 59.735 128.415 ;
        RECT 59.905 128.125 60.465 128.415 ;
        RECT 61.555 127.955 61.845 128.680 ;
        RECT 62.475 127.955 64.145 128.725 ;
        RECT 64.375 127.955 64.585 128.775 ;
        RECT 64.755 128.755 65.005 129.355 ;
        RECT 65.175 128.945 65.505 129.195 ;
        RECT 65.695 128.895 67.385 129.415 ;
        RECT 64.755 128.125 65.085 128.755 ;
        RECT 65.255 127.955 65.485 128.775 ;
        RECT 67.555 128.725 69.205 129.245 ;
        RECT 70.970 128.820 71.320 130.070 ;
        RECT 74.985 129.575 75.155 130.335 ;
        RECT 75.335 129.745 75.665 130.505 ;
        RECT 74.985 129.405 75.650 129.575 ;
        RECT 75.835 129.430 76.105 130.335 ;
        RECT 65.695 127.955 69.205 128.725 ;
        RECT 72.800 128.500 73.140 129.330 ;
        RECT 75.480 129.260 75.650 129.405 ;
        RECT 74.915 128.855 75.245 129.225 ;
        RECT 75.480 128.930 75.765 129.260 ;
        RECT 75.480 128.675 75.650 128.930 ;
        RECT 74.985 128.505 75.650 128.675 ;
        RECT 75.935 128.630 76.105 129.430 ;
        RECT 76.365 129.575 76.535 130.335 ;
        RECT 76.715 129.745 77.045 130.505 ;
        RECT 76.365 129.405 77.030 129.575 ;
        RECT 77.215 129.430 77.485 130.335 ;
        RECT 76.860 129.260 77.030 129.405 ;
        RECT 76.295 128.855 76.625 129.225 ;
        RECT 76.860 128.930 77.145 129.260 ;
        RECT 76.860 128.675 77.030 128.930 ;
        RECT 69.380 127.955 74.725 128.500 ;
        RECT 74.985 128.125 75.155 128.505 ;
        RECT 75.335 127.955 75.665 128.335 ;
        RECT 75.845 128.125 76.105 128.630 ;
        RECT 76.365 128.505 77.030 128.675 ;
        RECT 77.315 128.630 77.485 129.430 ;
        RECT 76.365 128.125 76.535 128.505 ;
        RECT 76.715 127.955 77.045 128.335 ;
        RECT 77.225 128.125 77.485 128.630 ;
        RECT 77.655 129.430 77.925 130.335 ;
        RECT 78.095 129.745 78.425 130.505 ;
        RECT 78.605 129.575 78.775 130.335 ;
        RECT 77.655 128.630 77.825 129.430 ;
        RECT 78.110 129.405 78.775 129.575 ;
        RECT 79.045 129.525 79.375 130.335 ;
        RECT 79.545 129.705 79.785 130.505 ;
        RECT 78.110 129.260 78.280 129.405 ;
        RECT 79.045 129.355 79.760 129.525 ;
        RECT 77.995 128.930 78.280 129.260 ;
        RECT 78.110 128.675 78.280 128.930 ;
        RECT 78.515 128.855 78.845 129.225 ;
        RECT 79.040 128.945 79.420 129.185 ;
        RECT 79.590 129.115 79.760 129.355 ;
        RECT 79.965 129.485 80.135 130.335 ;
        RECT 80.305 129.705 80.635 130.505 ;
        RECT 80.805 129.485 80.975 130.335 ;
        RECT 79.965 129.315 80.975 129.485 ;
        RECT 81.145 129.355 81.475 130.505 ;
        RECT 81.795 129.415 85.305 130.505 ;
        RECT 79.590 128.945 80.090 129.115 ;
        RECT 79.590 128.775 79.760 128.945 ;
        RECT 80.480 128.805 80.975 129.315 ;
        RECT 81.795 128.895 83.485 129.415 ;
        RECT 85.515 129.365 85.745 130.505 ;
        RECT 85.915 129.355 86.245 130.335 ;
        RECT 86.415 129.365 86.625 130.505 ;
        RECT 80.475 128.775 80.975 128.805 ;
        RECT 77.655 128.125 77.915 128.630 ;
        RECT 78.110 128.505 78.775 128.675 ;
        RECT 78.095 127.955 78.425 128.335 ;
        RECT 78.605 128.125 78.775 128.505 ;
        RECT 79.125 128.605 79.760 128.775 ;
        RECT 79.965 128.605 80.975 128.775 ;
        RECT 79.125 128.125 79.295 128.605 ;
        RECT 79.475 127.955 79.715 128.435 ;
        RECT 79.965 128.125 80.135 128.605 ;
        RECT 80.305 127.955 80.635 128.435 ;
        RECT 80.805 128.125 80.975 128.605 ;
        RECT 81.145 127.955 81.475 128.755 ;
        RECT 83.655 128.725 85.305 129.245 ;
        RECT 85.495 128.945 85.825 129.195 ;
        RECT 81.795 127.955 85.305 128.725 ;
        RECT 85.515 127.955 85.745 128.775 ;
        RECT 85.995 128.755 86.245 129.355 ;
        RECT 87.315 129.340 87.605 130.505 ;
        RECT 88.785 129.575 88.955 130.335 ;
        RECT 89.135 129.745 89.465 130.505 ;
        RECT 88.785 129.405 89.450 129.575 ;
        RECT 89.635 129.430 89.905 130.335 ;
        RECT 89.280 129.260 89.450 129.405 ;
        RECT 88.715 128.855 89.045 129.225 ;
        RECT 89.280 128.930 89.565 129.260 ;
        RECT 85.915 128.125 86.245 128.755 ;
        RECT 86.415 127.955 86.625 128.775 ;
        RECT 87.315 127.955 87.605 128.680 ;
        RECT 89.280 128.675 89.450 128.930 ;
        RECT 88.785 128.505 89.450 128.675 ;
        RECT 89.735 128.630 89.905 129.430 ;
        RECT 90.115 129.365 90.345 130.505 ;
        RECT 90.515 129.355 90.845 130.335 ;
        RECT 91.015 129.365 91.225 130.505 ;
        RECT 91.975 129.365 92.185 130.505 ;
        RECT 90.095 128.945 90.425 129.195 ;
        RECT 88.785 128.125 88.955 128.505 ;
        RECT 89.135 127.955 89.465 128.335 ;
        RECT 89.645 128.125 89.905 128.630 ;
        RECT 90.115 127.955 90.345 128.775 ;
        RECT 90.595 128.755 90.845 129.355 ;
        RECT 92.355 129.355 92.685 130.335 ;
        RECT 92.855 129.365 93.085 130.505 ;
        RECT 93.385 129.575 93.555 130.335 ;
        RECT 93.735 129.745 94.065 130.505 ;
        RECT 93.385 129.405 94.050 129.575 ;
        RECT 94.235 129.430 94.505 130.335 ;
        RECT 90.515 128.125 90.845 128.755 ;
        RECT 91.015 127.955 91.225 128.775 ;
        RECT 91.975 127.955 92.185 128.775 ;
        RECT 92.355 128.755 92.605 129.355 ;
        RECT 93.880 129.260 94.050 129.405 ;
        RECT 92.775 128.945 93.105 129.195 ;
        RECT 93.315 128.855 93.645 129.225 ;
        RECT 93.880 128.930 94.165 129.260 ;
        RECT 92.355 128.125 92.685 128.755 ;
        RECT 92.855 127.955 93.085 128.775 ;
        RECT 93.880 128.675 94.050 128.930 ;
        RECT 93.385 128.505 94.050 128.675 ;
        RECT 94.335 128.630 94.505 129.430 ;
        RECT 94.765 129.575 94.935 130.335 ;
        RECT 95.115 129.745 95.445 130.505 ;
        RECT 94.765 129.405 95.430 129.575 ;
        RECT 95.615 129.430 95.885 130.335 ;
        RECT 95.260 129.260 95.430 129.405 ;
        RECT 94.695 128.855 95.025 129.225 ;
        RECT 95.260 128.930 95.545 129.260 ;
        RECT 95.260 128.675 95.430 128.930 ;
        RECT 93.385 128.125 93.555 128.505 ;
        RECT 93.735 127.955 94.065 128.335 ;
        RECT 94.245 128.125 94.505 128.630 ;
        RECT 94.765 128.505 95.430 128.675 ;
        RECT 95.715 128.630 95.885 129.430 ;
        RECT 96.115 129.365 96.325 130.505 ;
        RECT 96.495 129.355 96.825 130.335 ;
        RECT 96.995 129.365 97.225 130.505 ;
        RECT 98.445 129.575 98.615 130.335 ;
        RECT 98.795 129.745 99.125 130.505 ;
        RECT 98.445 129.405 99.110 129.575 ;
        RECT 99.295 129.430 99.565 130.335 ;
        RECT 94.765 128.125 94.935 128.505 ;
        RECT 95.115 127.955 95.445 128.335 ;
        RECT 95.625 128.125 95.885 128.630 ;
        RECT 96.115 127.955 96.325 128.775 ;
        RECT 96.495 128.755 96.745 129.355 ;
        RECT 98.940 129.260 99.110 129.405 ;
        RECT 96.915 128.945 97.245 129.195 ;
        RECT 98.375 128.855 98.705 129.225 ;
        RECT 98.940 128.930 99.225 129.260 ;
        RECT 96.495 128.125 96.825 128.755 ;
        RECT 96.995 127.955 97.225 128.775 ;
        RECT 98.940 128.675 99.110 128.930 ;
        RECT 98.445 128.505 99.110 128.675 ;
        RECT 99.395 128.630 99.565 129.430 ;
        RECT 100.235 129.365 100.465 130.505 ;
        RECT 100.635 129.355 100.965 130.335 ;
        RECT 101.135 129.365 101.345 130.505 ;
        RECT 101.580 129.835 101.835 130.335 ;
        RECT 102.005 130.005 102.335 130.505 ;
        RECT 101.580 129.665 102.330 129.835 ;
        RECT 100.215 128.945 100.545 129.195 ;
        RECT 98.445 128.125 98.615 128.505 ;
        RECT 98.795 127.955 99.125 128.335 ;
        RECT 99.305 128.125 99.565 128.630 ;
        RECT 100.235 127.955 100.465 128.775 ;
        RECT 100.715 128.755 100.965 129.355 ;
        RECT 101.580 128.845 101.930 129.495 ;
        RECT 100.635 128.125 100.965 128.755 ;
        RECT 101.135 127.955 101.345 128.775 ;
        RECT 102.100 128.675 102.330 129.665 ;
        RECT 101.580 128.505 102.330 128.675 ;
        RECT 101.580 128.215 101.835 128.505 ;
        RECT 102.005 127.955 102.335 128.335 ;
        RECT 102.505 128.215 102.675 130.335 ;
        RECT 102.845 129.535 103.170 130.320 ;
        RECT 103.340 130.045 103.590 130.505 ;
        RECT 103.760 130.005 104.010 130.335 ;
        RECT 104.225 130.005 104.905 130.335 ;
        RECT 103.760 129.875 103.930 130.005 ;
        RECT 103.535 129.705 103.930 129.875 ;
        RECT 102.905 128.485 103.365 129.535 ;
        RECT 103.535 128.345 103.705 129.705 ;
        RECT 104.100 129.445 104.565 129.835 ;
        RECT 103.875 128.635 104.225 129.255 ;
        RECT 104.395 128.855 104.565 129.445 ;
        RECT 104.735 129.225 104.905 130.005 ;
        RECT 105.075 129.905 105.245 130.245 ;
        RECT 105.480 130.075 105.810 130.505 ;
        RECT 105.980 129.905 106.150 130.245 ;
        RECT 106.445 130.045 106.815 130.505 ;
        RECT 105.075 129.735 106.150 129.905 ;
        RECT 106.985 129.875 107.155 130.335 ;
        RECT 107.390 129.995 108.260 130.335 ;
        RECT 108.430 130.045 108.680 130.505 ;
        RECT 106.595 129.705 107.155 129.875 ;
        RECT 106.595 129.565 106.765 129.705 ;
        RECT 105.265 129.395 106.765 129.565 ;
        RECT 107.460 129.535 107.920 129.825 ;
        RECT 104.735 129.055 106.425 129.225 ;
        RECT 104.395 128.635 104.750 128.855 ;
        RECT 104.920 128.345 105.090 129.055 ;
        RECT 105.295 128.635 106.085 128.885 ;
        RECT 106.255 128.875 106.425 129.055 ;
        RECT 106.595 128.705 106.765 129.395 ;
        RECT 103.035 127.955 103.365 128.315 ;
        RECT 103.535 128.175 104.030 128.345 ;
        RECT 104.235 128.175 105.090 128.345 ;
        RECT 105.965 127.955 106.295 128.415 ;
        RECT 106.505 128.315 106.765 128.705 ;
        RECT 106.955 129.525 107.920 129.535 ;
        RECT 108.090 129.615 108.260 129.995 ;
        RECT 108.850 129.955 109.020 130.245 ;
        RECT 109.200 130.125 109.530 130.505 ;
        RECT 108.850 129.785 109.650 129.955 ;
        RECT 106.955 129.365 107.630 129.525 ;
        RECT 108.090 129.445 109.310 129.615 ;
        RECT 106.955 128.575 107.165 129.365 ;
        RECT 108.090 129.355 108.260 129.445 ;
        RECT 107.335 128.575 107.685 129.195 ;
        RECT 107.855 129.185 108.260 129.355 ;
        RECT 107.855 128.405 108.025 129.185 ;
        RECT 108.195 128.735 108.415 129.015 ;
        RECT 108.595 128.905 109.135 129.275 ;
        RECT 109.480 129.165 109.650 129.785 ;
        RECT 109.825 129.445 109.995 130.505 ;
        RECT 110.205 129.495 110.495 130.335 ;
        RECT 110.665 129.665 110.835 130.505 ;
        RECT 111.045 129.495 111.295 130.335 ;
        RECT 111.505 129.665 111.675 130.505 ;
        RECT 110.205 129.325 111.930 129.495 ;
        RECT 108.195 128.565 108.725 128.735 ;
        RECT 106.505 128.145 106.855 128.315 ;
        RECT 107.075 128.125 108.025 128.405 ;
        RECT 108.195 127.955 108.385 128.395 ;
        RECT 108.555 128.335 108.725 128.565 ;
        RECT 108.895 128.505 109.135 128.905 ;
        RECT 109.305 129.155 109.650 129.165 ;
        RECT 109.305 128.945 111.335 129.155 ;
        RECT 109.305 128.690 109.630 128.945 ;
        RECT 111.520 128.775 111.930 129.325 ;
        RECT 112.155 129.415 113.365 130.505 ;
        RECT 112.155 128.875 112.675 129.415 ;
        RECT 109.305 128.335 109.625 128.690 ;
        RECT 108.555 128.165 109.625 128.335 ;
        RECT 109.825 127.955 109.995 128.765 ;
        RECT 110.165 128.605 111.930 128.775 ;
        RECT 112.845 128.705 113.365 129.245 ;
        RECT 110.165 128.125 110.495 128.605 ;
        RECT 110.665 127.955 110.835 128.425 ;
        RECT 111.005 128.125 111.335 128.605 ;
        RECT 111.505 127.955 111.675 128.425 ;
        RECT 112.155 127.955 113.365 128.705 ;
        RECT 26.970 127.785 113.450 127.955 ;
        RECT 27.055 127.035 28.265 127.785 ;
        RECT 27.055 126.495 27.575 127.035 ;
        RECT 28.955 126.965 29.165 127.785 ;
        RECT 29.335 126.985 29.665 127.615 ;
        RECT 27.745 126.325 28.265 126.865 ;
        RECT 29.335 126.385 29.585 126.985 ;
        RECT 29.835 126.965 30.065 127.785 ;
        RECT 30.365 127.235 30.535 127.615 ;
        RECT 30.715 127.405 31.045 127.785 ;
        RECT 30.365 127.065 31.030 127.235 ;
        RECT 31.225 127.110 31.485 127.615 ;
        RECT 29.755 126.545 30.085 126.795 ;
        RECT 30.295 126.515 30.625 126.885 ;
        RECT 30.860 126.810 31.030 127.065 ;
        RECT 30.860 126.480 31.145 126.810 ;
        RECT 27.055 125.235 28.265 126.325 ;
        RECT 28.955 125.235 29.165 126.375 ;
        RECT 29.335 125.405 29.665 126.385 ;
        RECT 29.835 125.235 30.065 126.375 ;
        RECT 30.860 126.335 31.030 126.480 ;
        RECT 30.365 126.165 31.030 126.335 ;
        RECT 31.315 126.310 31.485 127.110 ;
        RECT 31.655 127.035 32.865 127.785 ;
        RECT 33.125 127.235 33.295 127.615 ;
        RECT 33.475 127.405 33.805 127.785 ;
        RECT 33.125 127.065 33.790 127.235 ;
        RECT 33.985 127.110 34.245 127.615 ;
        RECT 30.365 125.405 30.535 126.165 ;
        RECT 30.715 125.235 31.045 125.995 ;
        RECT 31.215 125.405 31.485 126.310 ;
        RECT 31.655 126.325 32.175 126.865 ;
        RECT 32.345 126.495 32.865 127.035 ;
        RECT 33.055 126.515 33.385 126.885 ;
        RECT 33.620 126.810 33.790 127.065 ;
        RECT 33.620 126.480 33.905 126.810 ;
        RECT 33.620 126.335 33.790 126.480 ;
        RECT 31.655 125.235 32.865 126.325 ;
        RECT 33.125 126.165 33.790 126.335 ;
        RECT 34.075 126.310 34.245 127.110 ;
        RECT 34.505 127.235 34.675 127.615 ;
        RECT 34.855 127.405 35.185 127.785 ;
        RECT 34.505 127.065 35.170 127.235 ;
        RECT 35.365 127.110 35.625 127.615 ;
        RECT 34.435 126.515 34.765 126.885 ;
        RECT 35.000 126.810 35.170 127.065 ;
        RECT 35.000 126.480 35.285 126.810 ;
        RECT 35.000 126.335 35.170 126.480 ;
        RECT 33.125 125.405 33.295 126.165 ;
        RECT 33.475 125.235 33.805 125.995 ;
        RECT 33.975 125.405 34.245 126.310 ;
        RECT 34.505 126.165 35.170 126.335 ;
        RECT 35.455 126.310 35.625 127.110 ;
        RECT 35.885 127.235 36.055 127.615 ;
        RECT 36.235 127.405 36.565 127.785 ;
        RECT 35.885 127.065 36.550 127.235 ;
        RECT 36.745 127.110 37.005 127.615 ;
        RECT 35.815 126.515 36.145 126.885 ;
        RECT 36.380 126.810 36.550 127.065 ;
        RECT 36.380 126.480 36.665 126.810 ;
        RECT 36.380 126.335 36.550 126.480 ;
        RECT 34.505 125.405 34.675 126.165 ;
        RECT 34.855 125.235 35.185 125.995 ;
        RECT 35.355 125.405 35.625 126.310 ;
        RECT 35.885 126.165 36.550 126.335 ;
        RECT 36.835 126.310 37.005 127.110 ;
        RECT 37.180 127.235 37.435 127.525 ;
        RECT 37.605 127.405 37.935 127.785 ;
        RECT 37.180 127.065 37.930 127.235 ;
        RECT 35.885 125.405 36.055 126.165 ;
        RECT 36.235 125.235 36.565 125.995 ;
        RECT 36.735 125.405 37.005 126.310 ;
        RECT 37.180 126.245 37.530 126.895 ;
        RECT 37.700 126.075 37.930 127.065 ;
        RECT 37.180 125.905 37.930 126.075 ;
        RECT 37.180 125.405 37.435 125.905 ;
        RECT 37.605 125.235 37.935 125.735 ;
        RECT 38.105 125.405 38.275 127.525 ;
        RECT 38.635 127.425 38.965 127.785 ;
        RECT 39.135 127.395 39.630 127.565 ;
        RECT 39.835 127.395 40.690 127.565 ;
        RECT 38.505 126.205 38.965 127.255 ;
        RECT 38.445 125.420 38.770 126.205 ;
        RECT 39.135 126.035 39.305 127.395 ;
        RECT 39.475 126.485 39.825 127.105 ;
        RECT 39.995 126.885 40.350 127.105 ;
        RECT 39.995 126.295 40.165 126.885 ;
        RECT 40.520 126.685 40.690 127.395 ;
        RECT 41.565 127.325 41.895 127.785 ;
        RECT 42.105 127.425 42.455 127.595 ;
        RECT 40.895 126.855 41.685 127.105 ;
        RECT 42.105 127.035 42.365 127.425 ;
        RECT 42.675 127.335 43.625 127.615 ;
        RECT 43.795 127.345 43.985 127.785 ;
        RECT 44.155 127.405 45.225 127.575 ;
        RECT 41.855 126.685 42.025 126.865 ;
        RECT 39.135 125.865 39.530 126.035 ;
        RECT 39.700 125.905 40.165 126.295 ;
        RECT 40.335 126.515 42.025 126.685 ;
        RECT 39.360 125.735 39.530 125.865 ;
        RECT 40.335 125.735 40.505 126.515 ;
        RECT 42.195 126.345 42.365 127.035 ;
        RECT 40.865 126.175 42.365 126.345 ;
        RECT 42.555 126.375 42.765 127.165 ;
        RECT 42.935 126.545 43.285 127.165 ;
        RECT 43.455 126.555 43.625 127.335 ;
        RECT 44.155 127.175 44.325 127.405 ;
        RECT 43.795 127.005 44.325 127.175 ;
        RECT 43.795 126.725 44.015 127.005 ;
        RECT 44.495 126.835 44.735 127.235 ;
        RECT 43.455 126.385 43.860 126.555 ;
        RECT 44.195 126.465 44.735 126.835 ;
        RECT 44.905 127.050 45.225 127.405 ;
        RECT 44.905 126.795 45.230 127.050 ;
        RECT 45.425 126.975 45.595 127.785 ;
        RECT 45.765 127.135 46.095 127.615 ;
        RECT 46.265 127.315 46.435 127.785 ;
        RECT 46.605 127.135 46.935 127.615 ;
        RECT 47.105 127.315 47.275 127.785 ;
        RECT 45.765 126.965 47.530 127.135 ;
        RECT 48.675 127.060 48.965 127.785 ;
        RECT 49.745 126.985 50.075 127.785 ;
        RECT 50.245 127.135 50.415 127.615 ;
        RECT 50.585 127.305 50.915 127.785 ;
        RECT 51.085 127.135 51.255 127.615 ;
        RECT 51.505 127.305 51.745 127.785 ;
        RECT 51.925 127.135 52.095 127.615 ;
        RECT 44.905 126.585 46.935 126.795 ;
        RECT 44.905 126.575 45.250 126.585 ;
        RECT 42.555 126.215 43.230 126.375 ;
        RECT 43.690 126.295 43.860 126.385 ;
        RECT 42.555 126.205 43.520 126.215 ;
        RECT 42.195 126.035 42.365 126.175 ;
        RECT 38.940 125.235 39.190 125.695 ;
        RECT 39.360 125.405 39.610 125.735 ;
        RECT 39.825 125.405 40.505 125.735 ;
        RECT 40.675 125.835 41.750 126.005 ;
        RECT 42.195 125.865 42.755 126.035 ;
        RECT 43.060 125.915 43.520 126.205 ;
        RECT 43.690 126.125 44.910 126.295 ;
        RECT 40.675 125.495 40.845 125.835 ;
        RECT 41.080 125.235 41.410 125.665 ;
        RECT 41.580 125.495 41.750 125.835 ;
        RECT 42.045 125.235 42.415 125.695 ;
        RECT 42.585 125.405 42.755 125.865 ;
        RECT 43.690 125.745 43.860 126.125 ;
        RECT 45.080 125.955 45.250 126.575 ;
        RECT 47.120 126.415 47.530 126.965 ;
        RECT 42.990 125.405 43.860 125.745 ;
        RECT 44.450 125.785 45.250 125.955 ;
        RECT 44.030 125.235 44.280 125.695 ;
        RECT 44.450 125.495 44.620 125.785 ;
        RECT 44.800 125.235 45.130 125.615 ;
        RECT 45.425 125.235 45.595 126.295 ;
        RECT 45.805 126.245 47.530 126.415 ;
        RECT 50.245 126.965 51.255 127.135 ;
        RECT 51.460 126.965 52.095 127.135 ;
        RECT 53.335 126.965 53.545 127.785 ;
        RECT 53.715 126.985 54.045 127.615 ;
        RECT 50.245 126.425 50.740 126.965 ;
        RECT 51.460 126.795 51.630 126.965 ;
        RECT 51.130 126.625 51.630 126.795 ;
        RECT 45.805 125.405 46.095 126.245 ;
        RECT 46.265 125.235 46.435 126.075 ;
        RECT 46.645 125.405 46.895 126.245 ;
        RECT 47.105 125.235 47.275 126.075 ;
        RECT 48.675 125.235 48.965 126.400 ;
        RECT 49.745 125.235 50.075 126.385 ;
        RECT 50.245 126.255 51.255 126.425 ;
        RECT 50.245 125.405 50.415 126.255 ;
        RECT 50.585 125.235 50.915 126.035 ;
        RECT 51.085 125.405 51.255 126.255 ;
        RECT 51.460 126.385 51.630 126.625 ;
        RECT 51.800 126.555 52.180 126.795 ;
        RECT 53.715 126.385 53.965 126.985 ;
        RECT 54.215 126.965 54.445 127.785 ;
        RECT 54.745 127.235 54.915 127.615 ;
        RECT 55.095 127.405 55.425 127.785 ;
        RECT 54.745 127.065 55.410 127.235 ;
        RECT 55.605 127.110 55.865 127.615 ;
        RECT 54.135 126.545 54.465 126.795 ;
        RECT 54.675 126.515 55.005 126.885 ;
        RECT 55.240 126.810 55.410 127.065 ;
        RECT 55.240 126.480 55.525 126.810 ;
        RECT 51.460 126.215 52.175 126.385 ;
        RECT 51.435 125.235 51.675 126.035 ;
        RECT 51.845 125.405 52.175 126.215 ;
        RECT 53.335 125.235 53.545 126.375 ;
        RECT 53.715 125.405 54.045 126.385 ;
        RECT 54.215 125.235 54.445 126.375 ;
        RECT 55.240 126.335 55.410 126.480 ;
        RECT 54.745 126.165 55.410 126.335 ;
        RECT 55.695 126.310 55.865 127.110 ;
        RECT 56.040 127.235 56.295 127.525 ;
        RECT 56.465 127.405 56.795 127.785 ;
        RECT 56.040 127.065 56.790 127.235 ;
        RECT 54.745 125.405 54.915 126.165 ;
        RECT 55.095 125.235 55.425 125.995 ;
        RECT 55.595 125.405 55.865 126.310 ;
        RECT 56.040 126.245 56.390 126.895 ;
        RECT 56.560 126.075 56.790 127.065 ;
        RECT 56.040 125.905 56.790 126.075 ;
        RECT 56.040 125.405 56.295 125.905 ;
        RECT 56.465 125.235 56.795 125.735 ;
        RECT 56.965 125.405 57.135 127.525 ;
        RECT 57.495 127.425 57.825 127.785 ;
        RECT 57.995 127.395 58.490 127.565 ;
        RECT 58.695 127.395 59.550 127.565 ;
        RECT 57.365 126.205 57.825 127.255 ;
        RECT 57.305 125.420 57.630 126.205 ;
        RECT 57.995 126.035 58.165 127.395 ;
        RECT 58.335 126.485 58.685 127.105 ;
        RECT 58.855 126.885 59.210 127.105 ;
        RECT 58.855 126.295 59.025 126.885 ;
        RECT 59.380 126.685 59.550 127.395 ;
        RECT 60.425 127.325 60.755 127.785 ;
        RECT 60.965 127.425 61.315 127.595 ;
        RECT 59.755 126.855 60.545 127.105 ;
        RECT 60.965 127.035 61.225 127.425 ;
        RECT 61.535 127.335 62.485 127.615 ;
        RECT 62.655 127.345 62.845 127.785 ;
        RECT 63.015 127.405 64.085 127.575 ;
        RECT 60.715 126.685 60.885 126.865 ;
        RECT 57.995 125.865 58.390 126.035 ;
        RECT 58.560 125.905 59.025 126.295 ;
        RECT 59.195 126.515 60.885 126.685 ;
        RECT 58.220 125.735 58.390 125.865 ;
        RECT 59.195 125.735 59.365 126.515 ;
        RECT 61.055 126.345 61.225 127.035 ;
        RECT 59.725 126.175 61.225 126.345 ;
        RECT 61.415 126.375 61.625 127.165 ;
        RECT 61.795 126.545 62.145 127.165 ;
        RECT 62.315 126.555 62.485 127.335 ;
        RECT 63.015 127.175 63.185 127.405 ;
        RECT 62.655 127.005 63.185 127.175 ;
        RECT 62.655 126.725 62.875 127.005 ;
        RECT 63.355 126.835 63.595 127.235 ;
        RECT 62.315 126.385 62.720 126.555 ;
        RECT 63.055 126.465 63.595 126.835 ;
        RECT 63.765 127.050 64.085 127.405 ;
        RECT 63.765 126.795 64.090 127.050 ;
        RECT 64.285 126.975 64.455 127.785 ;
        RECT 64.625 127.135 64.955 127.615 ;
        RECT 65.125 127.315 65.295 127.785 ;
        RECT 65.465 127.135 65.795 127.615 ;
        RECT 65.965 127.315 66.135 127.785 ;
        RECT 66.705 127.235 66.875 127.615 ;
        RECT 67.055 127.405 67.385 127.785 ;
        RECT 64.625 126.965 66.390 127.135 ;
        RECT 66.705 127.065 67.370 127.235 ;
        RECT 67.565 127.110 67.825 127.615 ;
        RECT 63.765 126.585 65.795 126.795 ;
        RECT 63.765 126.575 64.110 126.585 ;
        RECT 61.415 126.215 62.090 126.375 ;
        RECT 62.550 126.295 62.720 126.385 ;
        RECT 61.415 126.205 62.380 126.215 ;
        RECT 61.055 126.035 61.225 126.175 ;
        RECT 57.800 125.235 58.050 125.695 ;
        RECT 58.220 125.405 58.470 125.735 ;
        RECT 58.685 125.405 59.365 125.735 ;
        RECT 59.535 125.835 60.610 126.005 ;
        RECT 61.055 125.865 61.615 126.035 ;
        RECT 61.920 125.915 62.380 126.205 ;
        RECT 62.550 126.125 63.770 126.295 ;
        RECT 59.535 125.495 59.705 125.835 ;
        RECT 59.940 125.235 60.270 125.665 ;
        RECT 60.440 125.495 60.610 125.835 ;
        RECT 60.905 125.235 61.275 125.695 ;
        RECT 61.445 125.405 61.615 125.865 ;
        RECT 62.550 125.745 62.720 126.125 ;
        RECT 63.940 125.955 64.110 126.575 ;
        RECT 65.980 126.415 66.390 126.965 ;
        RECT 66.635 126.515 66.965 126.885 ;
        RECT 67.200 126.810 67.370 127.065 ;
        RECT 61.850 125.405 62.720 125.745 ;
        RECT 63.310 125.785 64.110 125.955 ;
        RECT 62.890 125.235 63.140 125.695 ;
        RECT 63.310 125.495 63.480 125.785 ;
        RECT 63.660 125.235 63.990 125.615 ;
        RECT 64.285 125.235 64.455 126.295 ;
        RECT 64.665 126.245 66.390 126.415 ;
        RECT 67.200 126.480 67.485 126.810 ;
        RECT 67.200 126.335 67.370 126.480 ;
        RECT 64.665 125.405 64.955 126.245 ;
        RECT 65.125 125.235 65.295 126.075 ;
        RECT 65.505 125.405 65.755 126.245 ;
        RECT 66.705 126.165 67.370 126.335 ;
        RECT 67.655 126.310 67.825 127.110 ;
        RECT 68.035 126.965 68.265 127.785 ;
        RECT 68.435 126.985 68.765 127.615 ;
        RECT 68.015 126.545 68.345 126.795 ;
        RECT 68.515 126.385 68.765 126.985 ;
        RECT 68.935 126.965 69.145 127.785 ;
        RECT 69.465 127.235 69.635 127.615 ;
        RECT 69.815 127.405 70.145 127.785 ;
        RECT 69.465 127.065 70.130 127.235 ;
        RECT 70.325 127.110 70.585 127.615 ;
        RECT 69.395 126.515 69.725 126.885 ;
        RECT 69.960 126.810 70.130 127.065 ;
        RECT 65.965 125.235 66.135 126.075 ;
        RECT 66.705 125.405 66.875 126.165 ;
        RECT 67.055 125.235 67.385 125.995 ;
        RECT 67.555 125.405 67.825 126.310 ;
        RECT 68.035 125.235 68.265 126.375 ;
        RECT 68.435 125.405 68.765 126.385 ;
        RECT 69.960 126.480 70.245 126.810 ;
        RECT 68.935 125.235 69.145 126.375 ;
        RECT 69.960 126.335 70.130 126.480 ;
        RECT 69.465 126.165 70.130 126.335 ;
        RECT 70.415 126.310 70.585 127.110 ;
        RECT 71.215 127.015 72.885 127.785 ;
        RECT 73.145 127.235 73.315 127.615 ;
        RECT 73.495 127.405 73.825 127.785 ;
        RECT 73.145 127.065 73.810 127.235 ;
        RECT 74.005 127.110 74.265 127.615 ;
        RECT 69.465 125.405 69.635 126.165 ;
        RECT 69.815 125.235 70.145 125.995 ;
        RECT 70.315 125.405 70.585 126.310 ;
        RECT 71.215 126.325 71.965 126.845 ;
        RECT 72.135 126.495 72.885 127.015 ;
        RECT 73.075 126.515 73.405 126.885 ;
        RECT 73.640 126.810 73.810 127.065 ;
        RECT 73.640 126.480 73.925 126.810 ;
        RECT 73.640 126.335 73.810 126.480 ;
        RECT 71.215 125.235 72.885 126.325 ;
        RECT 73.145 126.165 73.810 126.335 ;
        RECT 74.095 126.310 74.265 127.110 ;
        RECT 74.435 127.060 74.725 127.785 ;
        RECT 74.900 127.235 75.155 127.525 ;
        RECT 75.325 127.405 75.655 127.785 ;
        RECT 74.900 127.065 75.650 127.235 ;
        RECT 73.145 125.405 73.315 126.165 ;
        RECT 73.495 125.235 73.825 125.995 ;
        RECT 73.995 125.405 74.265 126.310 ;
        RECT 74.435 125.235 74.725 126.400 ;
        RECT 74.900 126.245 75.250 126.895 ;
        RECT 75.420 126.075 75.650 127.065 ;
        RECT 74.900 125.905 75.650 126.075 ;
        RECT 74.900 125.405 75.155 125.905 ;
        RECT 75.325 125.235 75.655 125.735 ;
        RECT 75.825 125.405 75.995 127.525 ;
        RECT 76.355 127.425 76.685 127.785 ;
        RECT 76.855 127.395 77.350 127.565 ;
        RECT 77.555 127.395 78.410 127.565 ;
        RECT 76.225 126.205 76.685 127.255 ;
        RECT 76.165 125.420 76.490 126.205 ;
        RECT 76.855 126.035 77.025 127.395 ;
        RECT 77.195 126.485 77.545 127.105 ;
        RECT 77.715 126.885 78.070 127.105 ;
        RECT 77.715 126.295 77.885 126.885 ;
        RECT 78.240 126.685 78.410 127.395 ;
        RECT 79.285 127.325 79.615 127.785 ;
        RECT 79.825 127.425 80.175 127.595 ;
        RECT 78.615 126.855 79.405 127.105 ;
        RECT 79.825 127.035 80.085 127.425 ;
        RECT 80.395 127.335 81.345 127.615 ;
        RECT 81.515 127.345 81.705 127.785 ;
        RECT 81.875 127.405 82.945 127.575 ;
        RECT 79.575 126.685 79.745 126.865 ;
        RECT 76.855 125.865 77.250 126.035 ;
        RECT 77.420 125.905 77.885 126.295 ;
        RECT 78.055 126.515 79.745 126.685 ;
        RECT 77.080 125.735 77.250 125.865 ;
        RECT 78.055 125.735 78.225 126.515 ;
        RECT 79.915 126.345 80.085 127.035 ;
        RECT 78.585 126.175 80.085 126.345 ;
        RECT 80.275 126.375 80.485 127.165 ;
        RECT 80.655 126.545 81.005 127.165 ;
        RECT 81.175 126.555 81.345 127.335 ;
        RECT 81.875 127.175 82.045 127.405 ;
        RECT 81.515 127.005 82.045 127.175 ;
        RECT 81.515 126.725 81.735 127.005 ;
        RECT 82.215 126.835 82.455 127.235 ;
        RECT 81.175 126.385 81.580 126.555 ;
        RECT 81.915 126.465 82.455 126.835 ;
        RECT 82.625 127.050 82.945 127.405 ;
        RECT 82.625 126.795 82.950 127.050 ;
        RECT 83.145 126.975 83.315 127.785 ;
        RECT 83.485 127.135 83.815 127.615 ;
        RECT 83.985 127.315 84.155 127.785 ;
        RECT 84.325 127.135 84.655 127.615 ;
        RECT 84.825 127.315 84.995 127.785 ;
        RECT 86.485 127.235 86.655 127.615 ;
        RECT 86.835 127.405 87.165 127.785 ;
        RECT 83.485 126.965 85.250 127.135 ;
        RECT 86.485 127.065 87.150 127.235 ;
        RECT 87.345 127.110 87.605 127.615 ;
        RECT 88.085 127.315 88.255 127.785 ;
        RECT 88.425 127.135 88.755 127.615 ;
        RECT 88.925 127.315 89.095 127.785 ;
        RECT 89.265 127.135 89.595 127.615 ;
        RECT 82.625 126.585 84.655 126.795 ;
        RECT 82.625 126.575 82.970 126.585 ;
        RECT 80.275 126.215 80.950 126.375 ;
        RECT 81.410 126.295 81.580 126.385 ;
        RECT 80.275 126.205 81.240 126.215 ;
        RECT 79.915 126.035 80.085 126.175 ;
        RECT 76.660 125.235 76.910 125.695 ;
        RECT 77.080 125.405 77.330 125.735 ;
        RECT 77.545 125.405 78.225 125.735 ;
        RECT 78.395 125.835 79.470 126.005 ;
        RECT 79.915 125.865 80.475 126.035 ;
        RECT 80.780 125.915 81.240 126.205 ;
        RECT 81.410 126.125 82.630 126.295 ;
        RECT 78.395 125.495 78.565 125.835 ;
        RECT 78.800 125.235 79.130 125.665 ;
        RECT 79.300 125.495 79.470 125.835 ;
        RECT 79.765 125.235 80.135 125.695 ;
        RECT 80.305 125.405 80.475 125.865 ;
        RECT 81.410 125.745 81.580 126.125 ;
        RECT 82.800 125.955 82.970 126.575 ;
        RECT 84.840 126.415 85.250 126.965 ;
        RECT 86.415 126.515 86.745 126.885 ;
        RECT 86.980 126.810 87.150 127.065 ;
        RECT 80.710 125.405 81.580 125.745 ;
        RECT 82.170 125.785 82.970 125.955 ;
        RECT 81.750 125.235 82.000 125.695 ;
        RECT 82.170 125.495 82.340 125.785 ;
        RECT 82.520 125.235 82.850 125.615 ;
        RECT 83.145 125.235 83.315 126.295 ;
        RECT 83.525 126.245 85.250 126.415 ;
        RECT 86.980 126.480 87.265 126.810 ;
        RECT 86.980 126.335 87.150 126.480 ;
        RECT 83.525 125.405 83.815 126.245 ;
        RECT 83.985 125.235 84.155 126.075 ;
        RECT 84.365 125.405 84.615 126.245 ;
        RECT 86.485 126.165 87.150 126.335 ;
        RECT 87.435 126.310 87.605 127.110 ;
        RECT 84.825 125.235 84.995 126.075 ;
        RECT 86.485 125.405 86.655 126.165 ;
        RECT 86.835 125.235 87.165 125.995 ;
        RECT 87.335 125.405 87.605 126.310 ;
        RECT 87.830 126.965 89.595 127.135 ;
        RECT 89.765 126.975 89.935 127.785 ;
        RECT 90.135 127.405 91.205 127.575 ;
        RECT 90.135 127.050 90.455 127.405 ;
        RECT 87.830 126.415 88.240 126.965 ;
        RECT 90.130 126.795 90.455 127.050 ;
        RECT 88.425 126.585 90.455 126.795 ;
        RECT 90.110 126.575 90.455 126.585 ;
        RECT 90.625 126.835 90.865 127.235 ;
        RECT 91.035 127.175 91.205 127.405 ;
        RECT 91.375 127.345 91.565 127.785 ;
        RECT 91.735 127.335 92.685 127.615 ;
        RECT 92.905 127.425 93.255 127.595 ;
        RECT 91.035 127.005 91.565 127.175 ;
        RECT 87.830 126.245 89.555 126.415 ;
        RECT 88.085 125.235 88.255 126.075 ;
        RECT 88.465 125.405 88.715 126.245 ;
        RECT 88.925 125.235 89.095 126.075 ;
        RECT 89.265 125.405 89.555 126.245 ;
        RECT 89.765 125.235 89.935 126.295 ;
        RECT 90.110 125.955 90.280 126.575 ;
        RECT 90.625 126.465 91.165 126.835 ;
        RECT 91.345 126.725 91.565 127.005 ;
        RECT 91.735 126.555 91.905 127.335 ;
        RECT 91.500 126.385 91.905 126.555 ;
        RECT 92.075 126.545 92.425 127.165 ;
        RECT 91.500 126.295 91.670 126.385 ;
        RECT 92.595 126.375 92.805 127.165 ;
        RECT 90.450 126.125 91.670 126.295 ;
        RECT 92.130 126.215 92.805 126.375 ;
        RECT 90.110 125.785 90.910 125.955 ;
        RECT 90.230 125.235 90.560 125.615 ;
        RECT 90.740 125.495 90.910 125.785 ;
        RECT 91.500 125.745 91.670 126.125 ;
        RECT 91.840 126.205 92.805 126.215 ;
        RECT 92.995 127.035 93.255 127.425 ;
        RECT 93.465 127.325 93.795 127.785 ;
        RECT 94.670 127.395 95.525 127.565 ;
        RECT 95.730 127.395 96.225 127.565 ;
        RECT 96.395 127.425 96.725 127.785 ;
        RECT 92.995 126.345 93.165 127.035 ;
        RECT 93.335 126.685 93.505 126.865 ;
        RECT 93.675 126.855 94.465 127.105 ;
        RECT 94.670 126.685 94.840 127.395 ;
        RECT 95.010 126.885 95.365 127.105 ;
        RECT 93.335 126.515 95.025 126.685 ;
        RECT 91.840 125.915 92.300 126.205 ;
        RECT 92.995 126.175 94.495 126.345 ;
        RECT 92.995 126.035 93.165 126.175 ;
        RECT 92.605 125.865 93.165 126.035 ;
        RECT 91.080 125.235 91.330 125.695 ;
        RECT 91.500 125.405 92.370 125.745 ;
        RECT 92.605 125.405 92.775 125.865 ;
        RECT 93.610 125.835 94.685 126.005 ;
        RECT 92.945 125.235 93.315 125.695 ;
        RECT 93.610 125.495 93.780 125.835 ;
        RECT 93.950 125.235 94.280 125.665 ;
        RECT 94.515 125.495 94.685 125.835 ;
        RECT 94.855 125.735 95.025 126.515 ;
        RECT 95.195 126.295 95.365 126.885 ;
        RECT 95.535 126.485 95.885 127.105 ;
        RECT 95.195 125.905 95.660 126.295 ;
        RECT 96.055 126.035 96.225 127.395 ;
        RECT 96.395 126.205 96.855 127.255 ;
        RECT 95.830 125.865 96.225 126.035 ;
        RECT 95.830 125.735 96.000 125.865 ;
        RECT 94.855 125.405 95.535 125.735 ;
        RECT 95.750 125.405 96.000 125.735 ;
        RECT 96.170 125.235 96.420 125.695 ;
        RECT 96.590 125.420 96.915 126.205 ;
        RECT 97.085 125.405 97.255 127.525 ;
        RECT 97.425 127.405 97.755 127.785 ;
        RECT 97.925 127.235 98.180 127.525 ;
        RECT 97.430 127.065 98.180 127.235 ;
        RECT 98.355 127.110 98.615 127.615 ;
        RECT 98.795 127.405 99.125 127.785 ;
        RECT 99.305 127.235 99.475 127.615 ;
        RECT 97.430 126.075 97.660 127.065 ;
        RECT 97.830 126.245 98.180 126.895 ;
        RECT 98.355 126.310 98.525 127.110 ;
        RECT 98.810 127.065 99.475 127.235 ;
        RECT 98.810 126.810 98.980 127.065 ;
        RECT 100.195 127.060 100.485 127.785 ;
        RECT 101.580 127.235 101.835 127.525 ;
        RECT 102.005 127.405 102.335 127.785 ;
        RECT 101.580 127.065 102.330 127.235 ;
        RECT 98.695 126.480 98.980 126.810 ;
        RECT 99.215 126.515 99.545 126.885 ;
        RECT 98.810 126.335 98.980 126.480 ;
        RECT 97.430 125.905 98.180 126.075 ;
        RECT 97.425 125.235 97.755 125.735 ;
        RECT 97.925 125.405 98.180 125.905 ;
        RECT 98.355 125.405 98.625 126.310 ;
        RECT 98.810 126.165 99.475 126.335 ;
        RECT 98.795 125.235 99.125 125.995 ;
        RECT 99.305 125.405 99.475 126.165 ;
        RECT 100.195 125.235 100.485 126.400 ;
        RECT 101.580 126.245 101.930 126.895 ;
        RECT 102.100 126.075 102.330 127.065 ;
        RECT 101.580 125.905 102.330 126.075 ;
        RECT 101.580 125.405 101.835 125.905 ;
        RECT 102.005 125.235 102.335 125.735 ;
        RECT 102.505 125.405 102.675 127.525 ;
        RECT 103.035 127.425 103.365 127.785 ;
        RECT 103.535 127.395 104.030 127.565 ;
        RECT 104.235 127.395 105.090 127.565 ;
        RECT 102.905 126.205 103.365 127.255 ;
        RECT 102.845 125.420 103.170 126.205 ;
        RECT 103.535 126.035 103.705 127.395 ;
        RECT 103.875 126.485 104.225 127.105 ;
        RECT 104.395 126.885 104.750 127.105 ;
        RECT 104.395 126.295 104.565 126.885 ;
        RECT 104.920 126.685 105.090 127.395 ;
        RECT 105.965 127.325 106.295 127.785 ;
        RECT 106.505 127.425 106.855 127.595 ;
        RECT 105.295 126.855 106.085 127.105 ;
        RECT 106.505 127.035 106.765 127.425 ;
        RECT 107.075 127.335 108.025 127.615 ;
        RECT 108.195 127.345 108.385 127.785 ;
        RECT 108.555 127.405 109.625 127.575 ;
        RECT 106.255 126.685 106.425 126.865 ;
        RECT 103.535 125.865 103.930 126.035 ;
        RECT 104.100 125.905 104.565 126.295 ;
        RECT 104.735 126.515 106.425 126.685 ;
        RECT 103.760 125.735 103.930 125.865 ;
        RECT 104.735 125.735 104.905 126.515 ;
        RECT 106.595 126.345 106.765 127.035 ;
        RECT 105.265 126.175 106.765 126.345 ;
        RECT 106.955 126.375 107.165 127.165 ;
        RECT 107.335 126.545 107.685 127.165 ;
        RECT 107.855 126.555 108.025 127.335 ;
        RECT 108.555 127.175 108.725 127.405 ;
        RECT 108.195 127.005 108.725 127.175 ;
        RECT 108.195 126.725 108.415 127.005 ;
        RECT 108.895 126.835 109.135 127.235 ;
        RECT 107.855 126.385 108.260 126.555 ;
        RECT 108.595 126.465 109.135 126.835 ;
        RECT 109.305 127.050 109.625 127.405 ;
        RECT 109.305 126.795 109.630 127.050 ;
        RECT 109.825 126.975 109.995 127.785 ;
        RECT 110.165 127.135 110.495 127.615 ;
        RECT 110.665 127.315 110.835 127.785 ;
        RECT 111.005 127.135 111.335 127.615 ;
        RECT 111.505 127.315 111.675 127.785 ;
        RECT 110.165 126.965 111.930 127.135 ;
        RECT 112.155 127.035 113.365 127.785 ;
        RECT 109.305 126.585 111.335 126.795 ;
        RECT 109.305 126.575 109.650 126.585 ;
        RECT 106.955 126.215 107.630 126.375 ;
        RECT 108.090 126.295 108.260 126.385 ;
        RECT 106.955 126.205 107.920 126.215 ;
        RECT 106.595 126.035 106.765 126.175 ;
        RECT 103.340 125.235 103.590 125.695 ;
        RECT 103.760 125.405 104.010 125.735 ;
        RECT 104.225 125.405 104.905 125.735 ;
        RECT 105.075 125.835 106.150 126.005 ;
        RECT 106.595 125.865 107.155 126.035 ;
        RECT 107.460 125.915 107.920 126.205 ;
        RECT 108.090 126.125 109.310 126.295 ;
        RECT 105.075 125.495 105.245 125.835 ;
        RECT 105.480 125.235 105.810 125.665 ;
        RECT 105.980 125.495 106.150 125.835 ;
        RECT 106.445 125.235 106.815 125.695 ;
        RECT 106.985 125.405 107.155 125.865 ;
        RECT 108.090 125.745 108.260 126.125 ;
        RECT 109.480 125.955 109.650 126.575 ;
        RECT 111.520 126.415 111.930 126.965 ;
        RECT 107.390 125.405 108.260 125.745 ;
        RECT 108.850 125.785 109.650 125.955 ;
        RECT 108.430 125.235 108.680 125.695 ;
        RECT 108.850 125.495 109.020 125.785 ;
        RECT 109.200 125.235 109.530 125.615 ;
        RECT 109.825 125.235 109.995 126.295 ;
        RECT 110.205 126.245 111.930 126.415 ;
        RECT 112.155 126.325 112.675 126.865 ;
        RECT 112.845 126.495 113.365 127.035 ;
        RECT 110.205 125.405 110.495 126.245 ;
        RECT 110.665 125.235 110.835 126.075 ;
        RECT 111.045 125.405 111.295 126.245 ;
        RECT 111.505 125.235 111.675 126.075 ;
        RECT 112.155 125.235 113.365 126.325 ;
        RECT 26.970 125.065 113.450 125.235 ;
        RECT 27.055 123.975 28.265 125.065 ;
        RECT 27.055 123.265 27.575 123.805 ;
        RECT 27.745 123.435 28.265 123.975 ;
        RECT 28.495 123.925 28.705 125.065 ;
        RECT 28.875 123.915 29.205 124.895 ;
        RECT 29.375 123.925 29.605 125.065 ;
        RECT 29.815 123.975 31.485 125.065 ;
        RECT 27.055 122.515 28.265 123.265 ;
        RECT 28.495 122.515 28.705 123.335 ;
        RECT 28.875 123.315 29.125 123.915 ;
        RECT 29.295 123.505 29.625 123.755 ;
        RECT 29.815 123.455 30.565 123.975 ;
        RECT 31.715 123.925 31.925 125.065 ;
        RECT 32.095 123.915 32.425 124.895 ;
        RECT 32.595 123.925 32.825 125.065 ;
        RECT 33.075 123.925 33.305 125.065 ;
        RECT 33.475 123.915 33.805 124.895 ;
        RECT 33.975 123.925 34.185 125.065 ;
        RECT 34.455 123.925 34.685 125.065 ;
        RECT 34.855 123.915 35.185 124.895 ;
        RECT 35.355 123.925 35.565 125.065 ;
        RECT 28.875 122.685 29.205 123.315 ;
        RECT 29.375 122.515 29.605 123.335 ;
        RECT 30.735 123.285 31.485 123.805 ;
        RECT 29.815 122.515 31.485 123.285 ;
        RECT 31.715 122.515 31.925 123.335 ;
        RECT 32.095 123.315 32.345 123.915 ;
        RECT 32.515 123.505 32.845 123.755 ;
        RECT 33.055 123.505 33.385 123.755 ;
        RECT 32.095 122.685 32.425 123.315 ;
        RECT 32.595 122.515 32.825 123.335 ;
        RECT 33.075 122.515 33.305 123.335 ;
        RECT 33.555 123.315 33.805 123.915 ;
        RECT 34.435 123.505 34.765 123.755 ;
        RECT 33.475 122.685 33.805 123.315 ;
        RECT 33.975 122.515 34.185 123.335 ;
        RECT 34.455 122.515 34.685 123.335 ;
        RECT 34.935 123.315 35.185 123.915 ;
        RECT 35.795 123.900 36.085 125.065 ;
        RECT 36.295 123.925 36.525 125.065 ;
        RECT 36.695 123.915 37.025 124.895 ;
        RECT 37.195 123.925 37.405 125.065 ;
        RECT 37.725 124.135 37.895 124.895 ;
        RECT 38.075 124.305 38.405 125.065 ;
        RECT 37.725 123.965 38.390 124.135 ;
        RECT 38.575 123.990 38.845 124.895 ;
        RECT 36.275 123.505 36.605 123.755 ;
        RECT 34.855 122.685 35.185 123.315 ;
        RECT 35.355 122.515 35.565 123.335 ;
        RECT 35.795 122.515 36.085 123.240 ;
        RECT 36.295 122.515 36.525 123.335 ;
        RECT 36.775 123.315 37.025 123.915 ;
        RECT 38.220 123.820 38.390 123.965 ;
        RECT 37.655 123.415 37.985 123.785 ;
        RECT 38.220 123.490 38.505 123.820 ;
        RECT 36.695 122.685 37.025 123.315 ;
        RECT 37.195 122.515 37.405 123.335 ;
        RECT 38.220 123.235 38.390 123.490 ;
        RECT 37.725 123.065 38.390 123.235 ;
        RECT 38.675 123.190 38.845 123.990 ;
        RECT 39.055 123.925 39.285 125.065 ;
        RECT 39.455 123.915 39.785 124.895 ;
        RECT 39.955 123.925 40.165 125.065 ;
        RECT 40.400 124.395 40.655 124.895 ;
        RECT 40.825 124.565 41.155 125.065 ;
        RECT 40.400 124.225 41.150 124.395 ;
        RECT 39.035 123.505 39.365 123.755 ;
        RECT 37.725 122.685 37.895 123.065 ;
        RECT 38.075 122.515 38.405 122.895 ;
        RECT 38.585 122.685 38.845 123.190 ;
        RECT 39.055 122.515 39.285 123.335 ;
        RECT 39.535 123.315 39.785 123.915 ;
        RECT 40.400 123.405 40.750 124.055 ;
        RECT 39.455 122.685 39.785 123.315 ;
        RECT 39.955 122.515 40.165 123.335 ;
        RECT 40.920 123.235 41.150 124.225 ;
        RECT 40.400 123.065 41.150 123.235 ;
        RECT 40.400 122.775 40.655 123.065 ;
        RECT 40.825 122.515 41.155 122.895 ;
        RECT 41.325 122.775 41.495 124.895 ;
        RECT 41.665 124.095 41.990 124.880 ;
        RECT 42.160 124.605 42.410 125.065 ;
        RECT 42.580 124.565 42.830 124.895 ;
        RECT 43.045 124.565 43.725 124.895 ;
        RECT 42.580 124.435 42.750 124.565 ;
        RECT 42.355 124.265 42.750 124.435 ;
        RECT 41.725 123.045 42.185 124.095 ;
        RECT 42.355 122.905 42.525 124.265 ;
        RECT 42.920 124.005 43.385 124.395 ;
        RECT 42.695 123.195 43.045 123.815 ;
        RECT 43.215 123.415 43.385 124.005 ;
        RECT 43.555 123.785 43.725 124.565 ;
        RECT 43.895 124.465 44.065 124.805 ;
        RECT 44.300 124.635 44.630 125.065 ;
        RECT 44.800 124.465 44.970 124.805 ;
        RECT 45.265 124.605 45.635 125.065 ;
        RECT 43.895 124.295 44.970 124.465 ;
        RECT 45.805 124.435 45.975 124.895 ;
        RECT 46.210 124.555 47.080 124.895 ;
        RECT 47.250 124.605 47.500 125.065 ;
        RECT 45.415 124.265 45.975 124.435 ;
        RECT 45.415 124.125 45.585 124.265 ;
        RECT 44.085 123.955 45.585 124.125 ;
        RECT 46.280 124.095 46.740 124.385 ;
        RECT 43.555 123.615 45.245 123.785 ;
        RECT 43.215 123.195 43.570 123.415 ;
        RECT 43.740 122.905 43.910 123.615 ;
        RECT 44.115 123.195 44.905 123.445 ;
        RECT 45.075 123.435 45.245 123.615 ;
        RECT 45.415 123.265 45.585 123.955 ;
        RECT 41.855 122.515 42.185 122.875 ;
        RECT 42.355 122.735 42.850 122.905 ;
        RECT 43.055 122.735 43.910 122.905 ;
        RECT 44.785 122.515 45.115 122.975 ;
        RECT 45.325 122.875 45.585 123.265 ;
        RECT 45.775 124.085 46.740 124.095 ;
        RECT 46.910 124.175 47.080 124.555 ;
        RECT 47.670 124.515 47.840 124.805 ;
        RECT 48.020 124.685 48.350 125.065 ;
        RECT 47.670 124.345 48.470 124.515 ;
        RECT 45.775 123.925 46.450 124.085 ;
        RECT 46.910 124.005 48.130 124.175 ;
        RECT 45.775 123.135 45.985 123.925 ;
        RECT 46.910 123.915 47.080 124.005 ;
        RECT 46.155 123.135 46.505 123.755 ;
        RECT 46.675 123.745 47.080 123.915 ;
        RECT 46.675 122.965 46.845 123.745 ;
        RECT 47.015 123.295 47.235 123.575 ;
        RECT 47.415 123.465 47.955 123.835 ;
        RECT 48.300 123.725 48.470 124.345 ;
        RECT 48.645 124.005 48.815 125.065 ;
        RECT 49.025 124.055 49.315 124.895 ;
        RECT 49.485 124.225 49.655 125.065 ;
        RECT 49.865 124.055 50.115 124.895 ;
        RECT 50.325 124.225 50.495 125.065 ;
        RECT 51.285 124.225 51.455 125.065 ;
        RECT 51.665 124.055 51.915 124.895 ;
        RECT 52.125 124.225 52.295 125.065 ;
        RECT 52.465 124.055 52.755 124.895 ;
        RECT 49.025 123.885 50.750 124.055 ;
        RECT 47.015 123.125 47.545 123.295 ;
        RECT 45.325 122.705 45.675 122.875 ;
        RECT 45.895 122.685 46.845 122.965 ;
        RECT 47.015 122.515 47.205 122.955 ;
        RECT 47.375 122.895 47.545 123.125 ;
        RECT 47.715 123.065 47.955 123.465 ;
        RECT 48.125 123.715 48.470 123.725 ;
        RECT 48.125 123.505 50.155 123.715 ;
        RECT 48.125 123.250 48.450 123.505 ;
        RECT 50.340 123.335 50.750 123.885 ;
        RECT 48.125 122.895 48.445 123.250 ;
        RECT 47.375 122.725 48.445 122.895 ;
        RECT 48.645 122.515 48.815 123.325 ;
        RECT 48.985 123.165 50.750 123.335 ;
        RECT 51.030 123.885 52.755 124.055 ;
        RECT 52.965 124.005 53.135 125.065 ;
        RECT 53.430 124.685 53.760 125.065 ;
        RECT 53.940 124.515 54.110 124.805 ;
        RECT 54.280 124.605 54.530 125.065 ;
        RECT 53.310 124.345 54.110 124.515 ;
        RECT 54.700 124.555 55.570 124.895 ;
        RECT 51.030 123.335 51.440 123.885 ;
        RECT 53.310 123.725 53.480 124.345 ;
        RECT 54.700 124.175 54.870 124.555 ;
        RECT 55.805 124.435 55.975 124.895 ;
        RECT 56.145 124.605 56.515 125.065 ;
        RECT 56.810 124.465 56.980 124.805 ;
        RECT 57.150 124.635 57.480 125.065 ;
        RECT 57.715 124.465 57.885 124.805 ;
        RECT 53.650 124.005 54.870 124.175 ;
        RECT 55.040 124.095 55.500 124.385 ;
        RECT 55.805 124.265 56.365 124.435 ;
        RECT 56.810 124.295 57.885 124.465 ;
        RECT 58.055 124.565 58.735 124.895 ;
        RECT 58.950 124.565 59.200 124.895 ;
        RECT 59.370 124.605 59.620 125.065 ;
        RECT 56.195 124.125 56.365 124.265 ;
        RECT 55.040 124.085 56.005 124.095 ;
        RECT 54.700 123.915 54.870 124.005 ;
        RECT 55.330 123.925 56.005 124.085 ;
        RECT 53.310 123.715 53.655 123.725 ;
        RECT 51.625 123.505 53.655 123.715 ;
        RECT 51.030 123.165 52.795 123.335 ;
        RECT 48.985 122.685 49.315 123.165 ;
        RECT 49.485 122.515 49.655 122.985 ;
        RECT 49.825 122.685 50.155 123.165 ;
        RECT 50.325 122.515 50.495 122.985 ;
        RECT 51.285 122.515 51.455 122.985 ;
        RECT 51.625 122.685 51.955 123.165 ;
        RECT 52.125 122.515 52.295 122.985 ;
        RECT 52.465 122.685 52.795 123.165 ;
        RECT 52.965 122.515 53.135 123.325 ;
        RECT 53.330 123.250 53.655 123.505 ;
        RECT 53.335 122.895 53.655 123.250 ;
        RECT 53.825 123.465 54.365 123.835 ;
        RECT 54.700 123.745 55.105 123.915 ;
        RECT 53.825 123.065 54.065 123.465 ;
        RECT 54.545 123.295 54.765 123.575 ;
        RECT 54.235 123.125 54.765 123.295 ;
        RECT 54.235 122.895 54.405 123.125 ;
        RECT 54.935 122.965 55.105 123.745 ;
        RECT 55.275 123.135 55.625 123.755 ;
        RECT 55.795 123.135 56.005 123.925 ;
        RECT 56.195 123.955 57.695 124.125 ;
        RECT 56.195 123.265 56.365 123.955 ;
        RECT 58.055 123.785 58.225 124.565 ;
        RECT 59.030 124.435 59.200 124.565 ;
        RECT 56.535 123.615 58.225 123.785 ;
        RECT 58.395 124.005 58.860 124.395 ;
        RECT 59.030 124.265 59.425 124.435 ;
        RECT 56.535 123.435 56.705 123.615 ;
        RECT 53.335 122.725 54.405 122.895 ;
        RECT 54.575 122.515 54.765 122.955 ;
        RECT 54.935 122.685 55.885 122.965 ;
        RECT 56.195 122.875 56.455 123.265 ;
        RECT 56.875 123.195 57.665 123.445 ;
        RECT 56.105 122.705 56.455 122.875 ;
        RECT 56.665 122.515 56.995 122.975 ;
        RECT 57.870 122.905 58.040 123.615 ;
        RECT 58.395 123.415 58.565 124.005 ;
        RECT 58.210 123.195 58.565 123.415 ;
        RECT 58.735 123.195 59.085 123.815 ;
        RECT 59.255 122.905 59.425 124.265 ;
        RECT 59.790 124.095 60.115 124.880 ;
        RECT 59.595 123.045 60.055 124.095 ;
        RECT 57.870 122.735 58.725 122.905 ;
        RECT 58.930 122.735 59.425 122.905 ;
        RECT 59.595 122.515 59.925 122.875 ;
        RECT 60.285 122.775 60.455 124.895 ;
        RECT 60.625 124.565 60.955 125.065 ;
        RECT 61.125 124.395 61.380 124.895 ;
        RECT 60.630 124.225 61.380 124.395 ;
        RECT 60.630 123.235 60.860 124.225 ;
        RECT 61.030 123.405 61.380 124.055 ;
        RECT 61.555 123.900 61.845 125.065 ;
        RECT 62.325 124.225 62.495 125.065 ;
        RECT 62.705 124.055 62.955 124.895 ;
        RECT 63.165 124.225 63.335 125.065 ;
        RECT 63.505 124.055 63.795 124.895 ;
        RECT 62.070 123.885 63.795 124.055 ;
        RECT 64.005 124.005 64.175 125.065 ;
        RECT 64.470 124.685 64.800 125.065 ;
        RECT 64.980 124.515 65.150 124.805 ;
        RECT 65.320 124.605 65.570 125.065 ;
        RECT 64.350 124.345 65.150 124.515 ;
        RECT 65.740 124.555 66.610 124.895 ;
        RECT 62.070 123.335 62.480 123.885 ;
        RECT 64.350 123.725 64.520 124.345 ;
        RECT 65.740 124.175 65.910 124.555 ;
        RECT 66.845 124.435 67.015 124.895 ;
        RECT 67.185 124.605 67.555 125.065 ;
        RECT 67.850 124.465 68.020 124.805 ;
        RECT 68.190 124.635 68.520 125.065 ;
        RECT 68.755 124.465 68.925 124.805 ;
        RECT 64.690 124.005 65.910 124.175 ;
        RECT 66.080 124.095 66.540 124.385 ;
        RECT 66.845 124.265 67.405 124.435 ;
        RECT 67.850 124.295 68.925 124.465 ;
        RECT 69.095 124.565 69.775 124.895 ;
        RECT 69.990 124.565 70.240 124.895 ;
        RECT 70.410 124.605 70.660 125.065 ;
        RECT 67.235 124.125 67.405 124.265 ;
        RECT 66.080 124.085 67.045 124.095 ;
        RECT 65.740 123.915 65.910 124.005 ;
        RECT 66.370 123.925 67.045 124.085 ;
        RECT 64.350 123.715 64.695 123.725 ;
        RECT 62.665 123.505 64.695 123.715 ;
        RECT 60.630 123.065 61.380 123.235 ;
        RECT 60.625 122.515 60.955 122.895 ;
        RECT 61.125 122.775 61.380 123.065 ;
        RECT 61.555 122.515 61.845 123.240 ;
        RECT 62.070 123.165 63.835 123.335 ;
        RECT 62.325 122.515 62.495 122.985 ;
        RECT 62.665 122.685 62.995 123.165 ;
        RECT 63.165 122.515 63.335 122.985 ;
        RECT 63.505 122.685 63.835 123.165 ;
        RECT 64.005 122.515 64.175 123.325 ;
        RECT 64.370 123.250 64.695 123.505 ;
        RECT 64.375 122.895 64.695 123.250 ;
        RECT 64.865 123.465 65.405 123.835 ;
        RECT 65.740 123.745 66.145 123.915 ;
        RECT 64.865 123.065 65.105 123.465 ;
        RECT 65.585 123.295 65.805 123.575 ;
        RECT 65.275 123.125 65.805 123.295 ;
        RECT 65.275 122.895 65.445 123.125 ;
        RECT 65.975 122.965 66.145 123.745 ;
        RECT 66.315 123.135 66.665 123.755 ;
        RECT 66.835 123.135 67.045 123.925 ;
        RECT 67.235 123.955 68.735 124.125 ;
        RECT 67.235 123.265 67.405 123.955 ;
        RECT 69.095 123.785 69.265 124.565 ;
        RECT 70.070 124.435 70.240 124.565 ;
        RECT 67.575 123.615 69.265 123.785 ;
        RECT 69.435 124.005 69.900 124.395 ;
        RECT 70.070 124.265 70.465 124.435 ;
        RECT 67.575 123.435 67.745 123.615 ;
        RECT 64.375 122.725 65.445 122.895 ;
        RECT 65.615 122.515 65.805 122.955 ;
        RECT 65.975 122.685 66.925 122.965 ;
        RECT 67.235 122.875 67.495 123.265 ;
        RECT 67.915 123.195 68.705 123.445 ;
        RECT 67.145 122.705 67.495 122.875 ;
        RECT 67.705 122.515 68.035 122.975 ;
        RECT 68.910 122.905 69.080 123.615 ;
        RECT 69.435 123.415 69.605 124.005 ;
        RECT 69.250 123.195 69.605 123.415 ;
        RECT 69.775 123.195 70.125 123.815 ;
        RECT 70.295 122.905 70.465 124.265 ;
        RECT 70.830 124.095 71.155 124.880 ;
        RECT 70.635 123.045 71.095 124.095 ;
        RECT 68.910 122.735 69.765 122.905 ;
        RECT 69.970 122.735 70.465 122.905 ;
        RECT 70.635 122.515 70.965 122.875 ;
        RECT 71.325 122.775 71.495 124.895 ;
        RECT 71.665 124.565 71.995 125.065 ;
        RECT 72.165 124.395 72.420 124.895 ;
        RECT 71.670 124.225 72.420 124.395 ;
        RECT 72.905 124.225 73.075 125.065 ;
        RECT 71.670 123.235 71.900 124.225 ;
        RECT 73.285 124.055 73.535 124.895 ;
        RECT 73.745 124.225 73.915 125.065 ;
        RECT 74.085 124.055 74.375 124.895 ;
        RECT 72.070 123.405 72.420 124.055 ;
        RECT 72.650 123.885 74.375 124.055 ;
        RECT 74.585 124.005 74.755 125.065 ;
        RECT 75.050 124.685 75.380 125.065 ;
        RECT 75.560 124.515 75.730 124.805 ;
        RECT 75.900 124.605 76.150 125.065 ;
        RECT 74.930 124.345 75.730 124.515 ;
        RECT 76.320 124.555 77.190 124.895 ;
        RECT 72.650 123.335 73.060 123.885 ;
        RECT 74.930 123.725 75.100 124.345 ;
        RECT 76.320 124.175 76.490 124.555 ;
        RECT 77.425 124.435 77.595 124.895 ;
        RECT 77.765 124.605 78.135 125.065 ;
        RECT 78.430 124.465 78.600 124.805 ;
        RECT 78.770 124.635 79.100 125.065 ;
        RECT 79.335 124.465 79.505 124.805 ;
        RECT 75.270 124.005 76.490 124.175 ;
        RECT 76.660 124.095 77.120 124.385 ;
        RECT 77.425 124.265 77.985 124.435 ;
        RECT 78.430 124.295 79.505 124.465 ;
        RECT 79.675 124.565 80.355 124.895 ;
        RECT 80.570 124.565 80.820 124.895 ;
        RECT 80.990 124.605 81.240 125.065 ;
        RECT 77.815 124.125 77.985 124.265 ;
        RECT 76.660 124.085 77.625 124.095 ;
        RECT 76.320 123.915 76.490 124.005 ;
        RECT 76.950 123.925 77.625 124.085 ;
        RECT 74.930 123.715 75.275 123.725 ;
        RECT 73.245 123.505 75.275 123.715 ;
        RECT 71.670 123.065 72.420 123.235 ;
        RECT 72.650 123.165 74.415 123.335 ;
        RECT 71.665 122.515 71.995 122.895 ;
        RECT 72.165 122.775 72.420 123.065 ;
        RECT 72.905 122.515 73.075 122.985 ;
        RECT 73.245 122.685 73.575 123.165 ;
        RECT 73.745 122.515 73.915 122.985 ;
        RECT 74.085 122.685 74.415 123.165 ;
        RECT 74.585 122.515 74.755 123.325 ;
        RECT 74.950 123.250 75.275 123.505 ;
        RECT 74.955 122.895 75.275 123.250 ;
        RECT 75.445 123.465 75.985 123.835 ;
        RECT 76.320 123.745 76.725 123.915 ;
        RECT 75.445 123.065 75.685 123.465 ;
        RECT 76.165 123.295 76.385 123.575 ;
        RECT 75.855 123.125 76.385 123.295 ;
        RECT 75.855 122.895 76.025 123.125 ;
        RECT 76.555 122.965 76.725 123.745 ;
        RECT 76.895 123.135 77.245 123.755 ;
        RECT 77.415 123.135 77.625 123.925 ;
        RECT 77.815 123.955 79.315 124.125 ;
        RECT 77.815 123.265 77.985 123.955 ;
        RECT 79.675 123.785 79.845 124.565 ;
        RECT 80.650 124.435 80.820 124.565 ;
        RECT 78.155 123.615 79.845 123.785 ;
        RECT 80.015 124.005 80.480 124.395 ;
        RECT 80.650 124.265 81.045 124.435 ;
        RECT 78.155 123.435 78.325 123.615 ;
        RECT 74.955 122.725 76.025 122.895 ;
        RECT 76.195 122.515 76.385 122.955 ;
        RECT 76.555 122.685 77.505 122.965 ;
        RECT 77.815 122.875 78.075 123.265 ;
        RECT 78.495 123.195 79.285 123.445 ;
        RECT 77.725 122.705 78.075 122.875 ;
        RECT 78.285 122.515 78.615 122.975 ;
        RECT 79.490 122.905 79.660 123.615 ;
        RECT 80.015 123.415 80.185 124.005 ;
        RECT 79.830 123.195 80.185 123.415 ;
        RECT 80.355 123.195 80.705 123.815 ;
        RECT 80.875 122.905 81.045 124.265 ;
        RECT 81.410 124.095 81.735 124.880 ;
        RECT 81.215 123.045 81.675 124.095 ;
        RECT 79.490 122.735 80.345 122.905 ;
        RECT 80.550 122.735 81.045 122.905 ;
        RECT 81.215 122.515 81.545 122.875 ;
        RECT 81.905 122.775 82.075 124.895 ;
        RECT 82.245 124.565 82.575 125.065 ;
        RECT 82.745 124.395 83.000 124.895 ;
        RECT 82.250 124.225 83.000 124.395 ;
        RECT 82.250 123.235 82.480 124.225 ;
        RECT 82.650 123.405 83.000 124.055 ;
        RECT 83.235 123.925 83.445 125.065 ;
        RECT 83.615 123.915 83.945 124.895 ;
        RECT 84.115 123.925 84.345 125.065 ;
        RECT 84.615 123.925 84.825 125.065 ;
        RECT 84.995 123.915 85.325 124.895 ;
        RECT 85.495 123.925 85.725 125.065 ;
        RECT 85.995 123.925 86.205 125.065 ;
        RECT 86.375 123.915 86.705 124.895 ;
        RECT 86.875 123.925 87.105 125.065 ;
        RECT 82.250 123.065 83.000 123.235 ;
        RECT 82.245 122.515 82.575 122.895 ;
        RECT 82.745 122.775 83.000 123.065 ;
        RECT 83.235 122.515 83.445 123.335 ;
        RECT 83.615 123.315 83.865 123.915 ;
        RECT 84.035 123.505 84.365 123.755 ;
        RECT 83.615 122.685 83.945 123.315 ;
        RECT 84.115 122.515 84.345 123.335 ;
        RECT 84.615 122.515 84.825 123.335 ;
        RECT 84.995 123.315 85.245 123.915 ;
        RECT 85.415 123.505 85.745 123.755 ;
        RECT 84.995 122.685 85.325 123.315 ;
        RECT 85.495 122.515 85.725 123.335 ;
        RECT 85.995 122.515 86.205 123.335 ;
        RECT 86.375 123.315 86.625 123.915 ;
        RECT 87.315 123.900 87.605 125.065 ;
        RECT 88.085 124.225 88.255 125.065 ;
        RECT 88.465 124.055 88.715 124.895 ;
        RECT 88.925 124.225 89.095 125.065 ;
        RECT 89.265 124.055 89.555 124.895 ;
        RECT 87.830 123.885 89.555 124.055 ;
        RECT 89.765 124.005 89.935 125.065 ;
        RECT 90.230 124.685 90.560 125.065 ;
        RECT 90.740 124.515 90.910 124.805 ;
        RECT 91.080 124.605 91.330 125.065 ;
        RECT 90.110 124.345 90.910 124.515 ;
        RECT 91.500 124.555 92.370 124.895 ;
        RECT 86.795 123.505 87.125 123.755 ;
        RECT 87.830 123.335 88.240 123.885 ;
        RECT 90.110 123.725 90.280 124.345 ;
        RECT 91.500 124.175 91.670 124.555 ;
        RECT 92.605 124.435 92.775 124.895 ;
        RECT 92.945 124.605 93.315 125.065 ;
        RECT 93.610 124.465 93.780 124.805 ;
        RECT 93.950 124.635 94.280 125.065 ;
        RECT 94.515 124.465 94.685 124.805 ;
        RECT 90.450 124.005 91.670 124.175 ;
        RECT 91.840 124.095 92.300 124.385 ;
        RECT 92.605 124.265 93.165 124.435 ;
        RECT 93.610 124.295 94.685 124.465 ;
        RECT 94.855 124.565 95.535 124.895 ;
        RECT 95.750 124.565 96.000 124.895 ;
        RECT 96.170 124.605 96.420 125.065 ;
        RECT 92.995 124.125 93.165 124.265 ;
        RECT 91.840 124.085 92.805 124.095 ;
        RECT 91.500 123.915 91.670 124.005 ;
        RECT 92.130 123.925 92.805 124.085 ;
        RECT 90.110 123.715 90.455 123.725 ;
        RECT 88.425 123.505 90.455 123.715 ;
        RECT 86.375 122.685 86.705 123.315 ;
        RECT 86.875 122.515 87.105 123.335 ;
        RECT 87.315 122.515 87.605 123.240 ;
        RECT 87.830 123.165 89.595 123.335 ;
        RECT 88.085 122.515 88.255 122.985 ;
        RECT 88.425 122.685 88.755 123.165 ;
        RECT 88.925 122.515 89.095 122.985 ;
        RECT 89.265 122.685 89.595 123.165 ;
        RECT 89.765 122.515 89.935 123.325 ;
        RECT 90.130 123.250 90.455 123.505 ;
        RECT 90.135 122.895 90.455 123.250 ;
        RECT 90.625 123.465 91.165 123.835 ;
        RECT 91.500 123.745 91.905 123.915 ;
        RECT 90.625 123.065 90.865 123.465 ;
        RECT 91.345 123.295 91.565 123.575 ;
        RECT 91.035 123.125 91.565 123.295 ;
        RECT 91.035 122.895 91.205 123.125 ;
        RECT 91.735 122.965 91.905 123.745 ;
        RECT 92.075 123.135 92.425 123.755 ;
        RECT 92.595 123.135 92.805 123.925 ;
        RECT 92.995 123.955 94.495 124.125 ;
        RECT 92.995 123.265 93.165 123.955 ;
        RECT 94.855 123.785 95.025 124.565 ;
        RECT 95.830 124.435 96.000 124.565 ;
        RECT 93.335 123.615 95.025 123.785 ;
        RECT 95.195 124.005 95.660 124.395 ;
        RECT 95.830 124.265 96.225 124.435 ;
        RECT 93.335 123.435 93.505 123.615 ;
        RECT 90.135 122.725 91.205 122.895 ;
        RECT 91.375 122.515 91.565 122.955 ;
        RECT 91.735 122.685 92.685 122.965 ;
        RECT 92.995 122.875 93.255 123.265 ;
        RECT 93.675 123.195 94.465 123.445 ;
        RECT 92.905 122.705 93.255 122.875 ;
        RECT 93.465 122.515 93.795 122.975 ;
        RECT 94.670 122.905 94.840 123.615 ;
        RECT 95.195 123.415 95.365 124.005 ;
        RECT 95.010 123.195 95.365 123.415 ;
        RECT 95.535 123.195 95.885 123.815 ;
        RECT 96.055 122.905 96.225 124.265 ;
        RECT 96.590 124.095 96.915 124.880 ;
        RECT 96.395 123.045 96.855 124.095 ;
        RECT 94.670 122.735 95.525 122.905 ;
        RECT 95.730 122.735 96.225 122.905 ;
        RECT 96.395 122.515 96.725 122.875 ;
        RECT 97.085 122.775 97.255 124.895 ;
        RECT 97.425 124.565 97.755 125.065 ;
        RECT 97.925 124.395 98.180 124.895 ;
        RECT 97.430 124.225 98.180 124.395 ;
        RECT 98.665 124.225 98.835 125.065 ;
        RECT 97.430 123.235 97.660 124.225 ;
        RECT 99.045 124.055 99.295 124.895 ;
        RECT 99.505 124.225 99.675 125.065 ;
        RECT 99.845 124.055 100.135 124.895 ;
        RECT 97.830 123.405 98.180 124.055 ;
        RECT 98.410 123.885 100.135 124.055 ;
        RECT 100.345 124.005 100.515 125.065 ;
        RECT 100.810 124.685 101.140 125.065 ;
        RECT 101.320 124.515 101.490 124.805 ;
        RECT 101.660 124.605 101.910 125.065 ;
        RECT 100.690 124.345 101.490 124.515 ;
        RECT 102.080 124.555 102.950 124.895 ;
        RECT 98.410 123.335 98.820 123.885 ;
        RECT 100.690 123.725 100.860 124.345 ;
        RECT 102.080 124.175 102.250 124.555 ;
        RECT 103.185 124.435 103.355 124.895 ;
        RECT 103.525 124.605 103.895 125.065 ;
        RECT 104.190 124.465 104.360 124.805 ;
        RECT 104.530 124.635 104.860 125.065 ;
        RECT 105.095 124.465 105.265 124.805 ;
        RECT 101.030 124.005 102.250 124.175 ;
        RECT 102.420 124.095 102.880 124.385 ;
        RECT 103.185 124.265 103.745 124.435 ;
        RECT 104.190 124.295 105.265 124.465 ;
        RECT 105.435 124.565 106.115 124.895 ;
        RECT 106.330 124.565 106.580 124.895 ;
        RECT 106.750 124.605 107.000 125.065 ;
        RECT 103.575 124.125 103.745 124.265 ;
        RECT 102.420 124.085 103.385 124.095 ;
        RECT 102.080 123.915 102.250 124.005 ;
        RECT 102.710 123.925 103.385 124.085 ;
        RECT 100.690 123.715 101.035 123.725 ;
        RECT 99.005 123.505 101.035 123.715 ;
        RECT 97.430 123.065 98.180 123.235 ;
        RECT 98.410 123.165 100.175 123.335 ;
        RECT 97.425 122.515 97.755 122.895 ;
        RECT 97.925 122.775 98.180 123.065 ;
        RECT 98.665 122.515 98.835 122.985 ;
        RECT 99.005 122.685 99.335 123.165 ;
        RECT 99.505 122.515 99.675 122.985 ;
        RECT 99.845 122.685 100.175 123.165 ;
        RECT 100.345 122.515 100.515 123.325 ;
        RECT 100.710 123.250 101.035 123.505 ;
        RECT 100.715 122.895 101.035 123.250 ;
        RECT 101.205 123.465 101.745 123.835 ;
        RECT 102.080 123.745 102.485 123.915 ;
        RECT 101.205 123.065 101.445 123.465 ;
        RECT 101.925 123.295 102.145 123.575 ;
        RECT 101.615 123.125 102.145 123.295 ;
        RECT 101.615 122.895 101.785 123.125 ;
        RECT 102.315 122.965 102.485 123.745 ;
        RECT 102.655 123.135 103.005 123.755 ;
        RECT 103.175 123.135 103.385 123.925 ;
        RECT 103.575 123.955 105.075 124.125 ;
        RECT 103.575 123.265 103.745 123.955 ;
        RECT 105.435 123.785 105.605 124.565 ;
        RECT 106.410 124.435 106.580 124.565 ;
        RECT 103.915 123.615 105.605 123.785 ;
        RECT 105.775 124.005 106.240 124.395 ;
        RECT 106.410 124.265 106.805 124.435 ;
        RECT 103.915 123.435 104.085 123.615 ;
        RECT 100.715 122.725 101.785 122.895 ;
        RECT 101.955 122.515 102.145 122.955 ;
        RECT 102.315 122.685 103.265 122.965 ;
        RECT 103.575 122.875 103.835 123.265 ;
        RECT 104.255 123.195 105.045 123.445 ;
        RECT 103.485 122.705 103.835 122.875 ;
        RECT 104.045 122.515 104.375 122.975 ;
        RECT 105.250 122.905 105.420 123.615 ;
        RECT 105.775 123.415 105.945 124.005 ;
        RECT 105.590 123.195 105.945 123.415 ;
        RECT 106.115 123.195 106.465 123.815 ;
        RECT 106.635 122.905 106.805 124.265 ;
        RECT 107.170 124.095 107.495 124.880 ;
        RECT 106.975 123.045 107.435 124.095 ;
        RECT 105.250 122.735 106.105 122.905 ;
        RECT 106.310 122.735 106.805 122.905 ;
        RECT 106.975 122.515 107.305 122.875 ;
        RECT 107.665 122.775 107.835 124.895 ;
        RECT 108.005 124.565 108.335 125.065 ;
        RECT 108.505 124.395 108.760 124.895 ;
        RECT 108.010 124.225 108.760 124.395 ;
        RECT 108.010 123.235 108.240 124.225 ;
        RECT 108.410 123.405 108.760 124.055 ;
        RECT 108.995 123.925 109.205 125.065 ;
        RECT 109.375 123.915 109.705 124.895 ;
        RECT 109.875 123.925 110.105 125.065 ;
        RECT 110.315 123.990 110.585 124.895 ;
        RECT 110.755 124.305 111.085 125.065 ;
        RECT 111.265 124.135 111.435 124.895 ;
        RECT 108.010 123.065 108.760 123.235 ;
        RECT 108.005 122.515 108.335 122.895 ;
        RECT 108.505 122.775 108.760 123.065 ;
        RECT 108.995 122.515 109.205 123.335 ;
        RECT 109.375 123.315 109.625 123.915 ;
        RECT 109.795 123.505 110.125 123.755 ;
        RECT 109.375 122.685 109.705 123.315 ;
        RECT 109.875 122.515 110.105 123.335 ;
        RECT 110.315 123.190 110.485 123.990 ;
        RECT 110.770 123.965 111.435 124.135 ;
        RECT 112.155 123.975 113.365 125.065 ;
        RECT 110.770 123.820 110.940 123.965 ;
        RECT 110.655 123.490 110.940 123.820 ;
        RECT 110.770 123.235 110.940 123.490 ;
        RECT 111.175 123.415 111.505 123.785 ;
        RECT 112.155 123.435 112.675 123.975 ;
        RECT 112.845 123.265 113.365 123.805 ;
        RECT 110.315 122.685 110.575 123.190 ;
        RECT 110.770 123.065 111.435 123.235 ;
        RECT 110.755 122.515 111.085 122.895 ;
        RECT 111.265 122.685 111.435 123.065 ;
        RECT 112.155 122.515 113.365 123.265 ;
        RECT 26.970 122.345 113.450 122.515 ;
        RECT 27.055 121.595 28.265 122.345 ;
        RECT 27.055 121.055 27.575 121.595 ;
        RECT 28.435 121.575 30.105 122.345 ;
        RECT 30.280 121.800 35.625 122.345 ;
        RECT 27.745 120.885 28.265 121.425 ;
        RECT 27.055 119.795 28.265 120.885 ;
        RECT 28.435 120.885 29.185 121.405 ;
        RECT 29.355 121.055 30.105 121.575 ;
        RECT 28.435 119.795 30.105 120.885 ;
        RECT 31.870 120.230 32.220 121.480 ;
        RECT 33.700 120.970 34.040 121.800 ;
        RECT 35.795 121.620 36.085 122.345 ;
        RECT 36.565 121.875 36.735 122.345 ;
        RECT 36.905 121.695 37.235 122.175 ;
        RECT 37.405 121.875 37.575 122.345 ;
        RECT 37.745 121.695 38.075 122.175 ;
        RECT 36.310 121.525 38.075 121.695 ;
        RECT 38.245 121.535 38.415 122.345 ;
        RECT 38.615 121.965 39.685 122.135 ;
        RECT 38.615 121.610 38.935 121.965 ;
        RECT 36.310 120.975 36.720 121.525 ;
        RECT 38.610 121.355 38.935 121.610 ;
        RECT 36.905 121.145 38.935 121.355 ;
        RECT 38.590 121.135 38.935 121.145 ;
        RECT 39.105 121.395 39.345 121.795 ;
        RECT 39.515 121.735 39.685 121.965 ;
        RECT 39.855 121.905 40.045 122.345 ;
        RECT 40.215 121.895 41.165 122.175 ;
        RECT 41.385 121.985 41.735 122.155 ;
        RECT 39.515 121.565 40.045 121.735 ;
        RECT 30.280 119.795 35.625 120.230 ;
        RECT 35.795 119.795 36.085 120.960 ;
        RECT 36.310 120.805 38.035 120.975 ;
        RECT 36.565 119.795 36.735 120.635 ;
        RECT 36.945 119.965 37.195 120.805 ;
        RECT 37.405 119.795 37.575 120.635 ;
        RECT 37.745 119.965 38.035 120.805 ;
        RECT 38.245 119.795 38.415 120.855 ;
        RECT 38.590 120.515 38.760 121.135 ;
        RECT 39.105 121.025 39.645 121.395 ;
        RECT 39.825 121.285 40.045 121.565 ;
        RECT 40.215 121.115 40.385 121.895 ;
        RECT 39.980 120.945 40.385 121.115 ;
        RECT 40.555 121.105 40.905 121.725 ;
        RECT 39.980 120.855 40.150 120.945 ;
        RECT 41.075 120.935 41.285 121.725 ;
        RECT 38.930 120.685 40.150 120.855 ;
        RECT 40.610 120.775 41.285 120.935 ;
        RECT 38.590 120.345 39.390 120.515 ;
        RECT 38.710 119.795 39.040 120.175 ;
        RECT 39.220 120.055 39.390 120.345 ;
        RECT 39.980 120.305 40.150 120.685 ;
        RECT 40.320 120.765 41.285 120.775 ;
        RECT 41.475 121.595 41.735 121.985 ;
        RECT 41.945 121.885 42.275 122.345 ;
        RECT 43.150 121.955 44.005 122.125 ;
        RECT 44.210 121.955 44.705 122.125 ;
        RECT 44.875 121.985 45.205 122.345 ;
        RECT 41.475 120.905 41.645 121.595 ;
        RECT 41.815 121.245 41.985 121.425 ;
        RECT 42.155 121.415 42.945 121.665 ;
        RECT 43.150 121.245 43.320 121.955 ;
        RECT 43.490 121.445 43.845 121.665 ;
        RECT 41.815 121.075 43.505 121.245 ;
        RECT 40.320 120.475 40.780 120.765 ;
        RECT 41.475 120.735 42.975 120.905 ;
        RECT 41.475 120.595 41.645 120.735 ;
        RECT 41.085 120.425 41.645 120.595 ;
        RECT 39.560 119.795 39.810 120.255 ;
        RECT 39.980 119.965 40.850 120.305 ;
        RECT 41.085 119.965 41.255 120.425 ;
        RECT 42.090 120.395 43.165 120.565 ;
        RECT 41.425 119.795 41.795 120.255 ;
        RECT 42.090 120.055 42.260 120.395 ;
        RECT 42.430 119.795 42.760 120.225 ;
        RECT 42.995 120.055 43.165 120.395 ;
        RECT 43.335 120.295 43.505 121.075 ;
        RECT 43.675 120.855 43.845 121.445 ;
        RECT 44.015 121.045 44.365 121.665 ;
        RECT 43.675 120.465 44.140 120.855 ;
        RECT 44.535 120.595 44.705 121.955 ;
        RECT 44.875 120.765 45.335 121.815 ;
        RECT 44.310 120.425 44.705 120.595 ;
        RECT 44.310 120.295 44.480 120.425 ;
        RECT 43.335 119.965 44.015 120.295 ;
        RECT 44.230 119.965 44.480 120.295 ;
        RECT 44.650 119.795 44.900 120.255 ;
        RECT 45.070 119.980 45.395 120.765 ;
        RECT 45.565 119.965 45.735 122.085 ;
        RECT 45.905 121.965 46.235 122.345 ;
        RECT 46.405 121.795 46.660 122.085 ;
        RECT 45.910 121.625 46.660 121.795 ;
        RECT 45.910 120.635 46.140 121.625 ;
        RECT 47.355 121.525 47.565 122.345 ;
        RECT 47.735 121.545 48.065 122.175 ;
        RECT 46.310 120.805 46.660 121.455 ;
        RECT 47.735 120.945 47.985 121.545 ;
        RECT 48.235 121.525 48.465 122.345 ;
        RECT 48.675 121.620 48.965 122.345 ;
        RECT 50.145 121.795 50.315 122.175 ;
        RECT 50.495 121.965 50.825 122.345 ;
        RECT 50.145 121.625 50.810 121.795 ;
        RECT 51.005 121.670 51.265 122.175 ;
        RECT 48.155 121.105 48.485 121.355 ;
        RECT 50.075 121.075 50.405 121.445 ;
        RECT 50.640 121.370 50.810 121.625 ;
        RECT 50.640 121.040 50.925 121.370 ;
        RECT 45.910 120.465 46.660 120.635 ;
        RECT 45.905 119.795 46.235 120.295 ;
        RECT 46.405 119.965 46.660 120.465 ;
        RECT 47.355 119.795 47.565 120.935 ;
        RECT 47.735 119.965 48.065 120.945 ;
        RECT 48.235 119.795 48.465 120.935 ;
        RECT 48.675 119.795 48.965 120.960 ;
        RECT 50.640 120.895 50.810 121.040 ;
        RECT 50.145 120.725 50.810 120.895 ;
        RECT 51.095 120.870 51.265 121.670 ;
        RECT 51.435 121.575 53.105 122.345 ;
        RECT 50.145 119.965 50.315 120.725 ;
        RECT 50.495 119.795 50.825 120.555 ;
        RECT 50.995 119.965 51.265 120.870 ;
        RECT 51.435 120.885 52.185 121.405 ;
        RECT 52.355 121.055 53.105 121.575 ;
        RECT 53.275 121.670 53.535 122.175 ;
        RECT 53.715 121.965 54.045 122.345 ;
        RECT 54.225 121.795 54.395 122.175 ;
        RECT 51.435 119.795 53.105 120.885 ;
        RECT 53.275 120.870 53.445 121.670 ;
        RECT 53.730 121.625 54.395 121.795 ;
        RECT 53.730 121.370 53.900 121.625 ;
        RECT 55.635 121.525 55.845 122.345 ;
        RECT 56.015 121.545 56.345 122.175 ;
        RECT 53.615 121.040 53.900 121.370 ;
        RECT 54.135 121.075 54.465 121.445 ;
        RECT 53.730 120.895 53.900 121.040 ;
        RECT 56.015 120.945 56.265 121.545 ;
        RECT 56.515 121.525 56.745 122.345 ;
        RECT 57.415 121.575 60.005 122.345 ;
        RECT 56.435 121.105 56.765 121.355 ;
        RECT 53.275 119.965 53.545 120.870 ;
        RECT 53.730 120.725 54.395 120.895 ;
        RECT 53.715 119.795 54.045 120.555 ;
        RECT 54.225 119.965 54.395 120.725 ;
        RECT 55.635 119.795 55.845 120.935 ;
        RECT 56.015 119.965 56.345 120.945 ;
        RECT 56.515 119.795 56.745 120.935 ;
        RECT 57.415 120.885 58.625 121.405 ;
        RECT 58.795 121.055 60.005 121.575 ;
        RECT 60.215 121.525 60.445 122.345 ;
        RECT 60.615 121.545 60.945 122.175 ;
        RECT 60.195 121.105 60.525 121.355 ;
        RECT 60.695 120.945 60.945 121.545 ;
        RECT 61.115 121.525 61.325 122.345 ;
        RECT 61.555 121.620 61.845 122.345 ;
        RECT 62.515 121.525 62.745 122.345 ;
        RECT 62.915 121.545 63.245 122.175 ;
        RECT 62.495 121.105 62.825 121.355 ;
        RECT 57.415 119.795 60.005 120.885 ;
        RECT 60.215 119.795 60.445 120.935 ;
        RECT 60.615 119.965 60.945 120.945 ;
        RECT 61.115 119.795 61.325 120.935 ;
        RECT 61.555 119.795 61.845 120.960 ;
        RECT 62.995 120.945 63.245 121.545 ;
        RECT 63.415 121.525 63.625 122.345 ;
        RECT 64.165 121.875 64.335 122.345 ;
        RECT 64.505 121.695 64.835 122.175 ;
        RECT 65.005 121.875 65.175 122.345 ;
        RECT 65.345 121.695 65.675 122.175 ;
        RECT 63.910 121.525 65.675 121.695 ;
        RECT 65.845 121.535 66.015 122.345 ;
        RECT 66.215 121.965 67.285 122.135 ;
        RECT 66.215 121.610 66.535 121.965 ;
        RECT 62.515 119.795 62.745 120.935 ;
        RECT 62.915 119.965 63.245 120.945 ;
        RECT 63.910 120.975 64.320 121.525 ;
        RECT 66.210 121.355 66.535 121.610 ;
        RECT 64.505 121.145 66.535 121.355 ;
        RECT 66.190 121.135 66.535 121.145 ;
        RECT 66.705 121.395 66.945 121.795 ;
        RECT 67.115 121.735 67.285 121.965 ;
        RECT 67.455 121.905 67.645 122.345 ;
        RECT 67.815 121.895 68.765 122.175 ;
        RECT 68.985 121.985 69.335 122.155 ;
        RECT 67.115 121.565 67.645 121.735 ;
        RECT 63.415 119.795 63.625 120.935 ;
        RECT 63.910 120.805 65.635 120.975 ;
        RECT 64.165 119.795 64.335 120.635 ;
        RECT 64.545 119.965 64.795 120.805 ;
        RECT 65.005 119.795 65.175 120.635 ;
        RECT 65.345 119.965 65.635 120.805 ;
        RECT 65.845 119.795 66.015 120.855 ;
        RECT 66.190 120.515 66.360 121.135 ;
        RECT 66.705 121.025 67.245 121.395 ;
        RECT 67.425 121.285 67.645 121.565 ;
        RECT 67.815 121.115 67.985 121.895 ;
        RECT 67.580 120.945 67.985 121.115 ;
        RECT 68.155 121.105 68.505 121.725 ;
        RECT 67.580 120.855 67.750 120.945 ;
        RECT 68.675 120.935 68.885 121.725 ;
        RECT 66.530 120.685 67.750 120.855 ;
        RECT 68.210 120.775 68.885 120.935 ;
        RECT 66.190 120.345 66.990 120.515 ;
        RECT 66.310 119.795 66.640 120.175 ;
        RECT 66.820 120.055 66.990 120.345 ;
        RECT 67.580 120.305 67.750 120.685 ;
        RECT 67.920 120.765 68.885 120.775 ;
        RECT 69.075 121.595 69.335 121.985 ;
        RECT 69.545 121.885 69.875 122.345 ;
        RECT 70.750 121.955 71.605 122.125 ;
        RECT 71.810 121.955 72.305 122.125 ;
        RECT 72.475 121.985 72.805 122.345 ;
        RECT 69.075 120.905 69.245 121.595 ;
        RECT 69.415 121.245 69.585 121.425 ;
        RECT 69.755 121.415 70.545 121.665 ;
        RECT 70.750 121.245 70.920 121.955 ;
        RECT 71.090 121.445 71.445 121.665 ;
        RECT 69.415 121.075 71.105 121.245 ;
        RECT 67.920 120.475 68.380 120.765 ;
        RECT 69.075 120.735 70.575 120.905 ;
        RECT 69.075 120.595 69.245 120.735 ;
        RECT 68.685 120.425 69.245 120.595 ;
        RECT 67.160 119.795 67.410 120.255 ;
        RECT 67.580 119.965 68.450 120.305 ;
        RECT 68.685 119.965 68.855 120.425 ;
        RECT 69.690 120.395 70.765 120.565 ;
        RECT 69.025 119.795 69.395 120.255 ;
        RECT 69.690 120.055 69.860 120.395 ;
        RECT 70.030 119.795 70.360 120.225 ;
        RECT 70.595 120.055 70.765 120.395 ;
        RECT 70.935 120.295 71.105 121.075 ;
        RECT 71.275 120.855 71.445 121.445 ;
        RECT 71.615 121.045 71.965 121.665 ;
        RECT 71.275 120.465 71.740 120.855 ;
        RECT 72.135 120.595 72.305 121.955 ;
        RECT 72.475 120.765 72.935 121.815 ;
        RECT 71.910 120.425 72.305 120.595 ;
        RECT 71.910 120.295 72.080 120.425 ;
        RECT 70.935 119.965 71.615 120.295 ;
        RECT 71.830 119.965 72.080 120.295 ;
        RECT 72.250 119.795 72.500 120.255 ;
        RECT 72.670 119.980 72.995 120.765 ;
        RECT 73.165 119.965 73.335 122.085 ;
        RECT 73.505 121.965 73.835 122.345 ;
        RECT 74.005 121.795 74.260 122.085 ;
        RECT 73.510 121.625 74.260 121.795 ;
        RECT 73.510 120.635 73.740 121.625 ;
        RECT 74.435 121.620 74.725 122.345 ;
        RECT 75.415 121.525 75.625 122.345 ;
        RECT 75.795 121.545 76.125 122.175 ;
        RECT 73.910 120.805 74.260 121.455 ;
        RECT 73.510 120.465 74.260 120.635 ;
        RECT 73.505 119.795 73.835 120.295 ;
        RECT 74.005 119.965 74.260 120.465 ;
        RECT 74.435 119.795 74.725 120.960 ;
        RECT 75.795 120.945 76.045 121.545 ;
        RECT 76.295 121.525 76.525 122.345 ;
        RECT 76.740 121.795 76.995 122.085 ;
        RECT 77.165 121.965 77.495 122.345 ;
        RECT 76.740 121.625 77.490 121.795 ;
        RECT 76.215 121.105 76.545 121.355 ;
        RECT 75.415 119.795 75.625 120.935 ;
        RECT 75.795 119.965 76.125 120.945 ;
        RECT 76.295 119.795 76.525 120.935 ;
        RECT 76.740 120.805 77.090 121.455 ;
        RECT 77.260 120.635 77.490 121.625 ;
        RECT 76.740 120.465 77.490 120.635 ;
        RECT 76.740 119.965 76.995 120.465 ;
        RECT 77.165 119.795 77.495 120.295 ;
        RECT 77.665 119.965 77.835 122.085 ;
        RECT 78.195 121.985 78.525 122.345 ;
        RECT 78.695 121.955 79.190 122.125 ;
        RECT 79.395 121.955 80.250 122.125 ;
        RECT 78.065 120.765 78.525 121.815 ;
        RECT 78.005 119.980 78.330 120.765 ;
        RECT 78.695 120.595 78.865 121.955 ;
        RECT 79.035 121.045 79.385 121.665 ;
        RECT 79.555 121.445 79.910 121.665 ;
        RECT 79.555 120.855 79.725 121.445 ;
        RECT 80.080 121.245 80.250 121.955 ;
        RECT 81.125 121.885 81.455 122.345 ;
        RECT 81.665 121.985 82.015 122.155 ;
        RECT 80.455 121.415 81.245 121.665 ;
        RECT 81.665 121.595 81.925 121.985 ;
        RECT 82.235 121.895 83.185 122.175 ;
        RECT 83.355 121.905 83.545 122.345 ;
        RECT 83.715 121.965 84.785 122.135 ;
        RECT 81.415 121.245 81.585 121.425 ;
        RECT 78.695 120.425 79.090 120.595 ;
        RECT 79.260 120.465 79.725 120.855 ;
        RECT 79.895 121.075 81.585 121.245 ;
        RECT 78.920 120.295 79.090 120.425 ;
        RECT 79.895 120.295 80.065 121.075 ;
        RECT 81.755 120.905 81.925 121.595 ;
        RECT 80.425 120.735 81.925 120.905 ;
        RECT 82.115 120.935 82.325 121.725 ;
        RECT 82.495 121.105 82.845 121.725 ;
        RECT 83.015 121.115 83.185 121.895 ;
        RECT 83.715 121.735 83.885 121.965 ;
        RECT 83.355 121.565 83.885 121.735 ;
        RECT 83.355 121.285 83.575 121.565 ;
        RECT 84.055 121.395 84.295 121.795 ;
        RECT 83.015 120.945 83.420 121.115 ;
        RECT 83.755 121.025 84.295 121.395 ;
        RECT 84.465 121.610 84.785 121.965 ;
        RECT 84.465 121.355 84.790 121.610 ;
        RECT 84.985 121.535 85.155 122.345 ;
        RECT 85.325 121.695 85.655 122.175 ;
        RECT 85.825 121.875 85.995 122.345 ;
        RECT 86.165 121.695 86.495 122.175 ;
        RECT 86.665 121.875 86.835 122.345 ;
        RECT 85.325 121.525 87.090 121.695 ;
        RECT 87.315 121.620 87.605 122.345 ;
        RECT 87.815 121.525 88.045 122.345 ;
        RECT 88.215 121.545 88.545 122.175 ;
        RECT 84.465 121.145 86.495 121.355 ;
        RECT 84.465 121.135 84.810 121.145 ;
        RECT 82.115 120.775 82.790 120.935 ;
        RECT 83.250 120.855 83.420 120.945 ;
        RECT 82.115 120.765 83.080 120.775 ;
        RECT 81.755 120.595 81.925 120.735 ;
        RECT 78.500 119.795 78.750 120.255 ;
        RECT 78.920 119.965 79.170 120.295 ;
        RECT 79.385 119.965 80.065 120.295 ;
        RECT 80.235 120.395 81.310 120.565 ;
        RECT 81.755 120.425 82.315 120.595 ;
        RECT 82.620 120.475 83.080 120.765 ;
        RECT 83.250 120.685 84.470 120.855 ;
        RECT 80.235 120.055 80.405 120.395 ;
        RECT 80.640 119.795 80.970 120.225 ;
        RECT 81.140 120.055 81.310 120.395 ;
        RECT 81.605 119.795 81.975 120.255 ;
        RECT 82.145 119.965 82.315 120.425 ;
        RECT 83.250 120.305 83.420 120.685 ;
        RECT 84.640 120.515 84.810 121.135 ;
        RECT 86.680 120.975 87.090 121.525 ;
        RECT 87.795 121.105 88.125 121.355 ;
        RECT 82.550 119.965 83.420 120.305 ;
        RECT 84.010 120.345 84.810 120.515 ;
        RECT 83.590 119.795 83.840 120.255 ;
        RECT 84.010 120.055 84.180 120.345 ;
        RECT 84.360 119.795 84.690 120.175 ;
        RECT 84.985 119.795 85.155 120.855 ;
        RECT 85.365 120.805 87.090 120.975 ;
        RECT 85.365 119.965 85.655 120.805 ;
        RECT 85.825 119.795 85.995 120.635 ;
        RECT 86.205 119.965 86.455 120.805 ;
        RECT 86.665 119.795 86.835 120.635 ;
        RECT 87.315 119.795 87.605 120.960 ;
        RECT 88.295 120.945 88.545 121.545 ;
        RECT 88.715 121.525 88.925 122.345 ;
        RECT 89.925 121.875 90.095 122.345 ;
        RECT 90.265 121.695 90.595 122.175 ;
        RECT 90.765 121.875 90.935 122.345 ;
        RECT 91.105 121.695 91.435 122.175 ;
        RECT 89.670 121.525 91.435 121.695 ;
        RECT 91.605 121.535 91.775 122.345 ;
        RECT 91.975 121.965 93.045 122.135 ;
        RECT 91.975 121.610 92.295 121.965 ;
        RECT 87.815 119.795 88.045 120.935 ;
        RECT 88.215 119.965 88.545 120.945 ;
        RECT 89.670 120.975 90.080 121.525 ;
        RECT 91.970 121.355 92.295 121.610 ;
        RECT 90.265 121.145 92.295 121.355 ;
        RECT 91.950 121.135 92.295 121.145 ;
        RECT 92.465 121.395 92.705 121.795 ;
        RECT 92.875 121.735 93.045 121.965 ;
        RECT 93.215 121.905 93.405 122.345 ;
        RECT 93.575 121.895 94.525 122.175 ;
        RECT 94.745 121.985 95.095 122.155 ;
        RECT 92.875 121.565 93.405 121.735 ;
        RECT 88.715 119.795 88.925 120.935 ;
        RECT 89.670 120.805 91.395 120.975 ;
        RECT 89.925 119.795 90.095 120.635 ;
        RECT 90.305 119.965 90.555 120.805 ;
        RECT 90.765 119.795 90.935 120.635 ;
        RECT 91.105 119.965 91.395 120.805 ;
        RECT 91.605 119.795 91.775 120.855 ;
        RECT 91.950 120.515 92.120 121.135 ;
        RECT 92.465 121.025 93.005 121.395 ;
        RECT 93.185 121.285 93.405 121.565 ;
        RECT 93.575 121.115 93.745 121.895 ;
        RECT 93.340 120.945 93.745 121.115 ;
        RECT 93.915 121.105 94.265 121.725 ;
        RECT 93.340 120.855 93.510 120.945 ;
        RECT 94.435 120.935 94.645 121.725 ;
        RECT 92.290 120.685 93.510 120.855 ;
        RECT 93.970 120.775 94.645 120.935 ;
        RECT 91.950 120.345 92.750 120.515 ;
        RECT 92.070 119.795 92.400 120.175 ;
        RECT 92.580 120.055 92.750 120.345 ;
        RECT 93.340 120.305 93.510 120.685 ;
        RECT 93.680 120.765 94.645 120.775 ;
        RECT 94.835 121.595 95.095 121.985 ;
        RECT 95.305 121.885 95.635 122.345 ;
        RECT 96.510 121.955 97.365 122.125 ;
        RECT 97.570 121.955 98.065 122.125 ;
        RECT 98.235 121.985 98.565 122.345 ;
        RECT 94.835 120.905 95.005 121.595 ;
        RECT 95.175 121.245 95.345 121.425 ;
        RECT 95.515 121.415 96.305 121.665 ;
        RECT 96.510 121.245 96.680 121.955 ;
        RECT 96.850 121.445 97.205 121.665 ;
        RECT 95.175 121.075 96.865 121.245 ;
        RECT 93.680 120.475 94.140 120.765 ;
        RECT 94.835 120.735 96.335 120.905 ;
        RECT 94.835 120.595 95.005 120.735 ;
        RECT 94.445 120.425 95.005 120.595 ;
        RECT 92.920 119.795 93.170 120.255 ;
        RECT 93.340 119.965 94.210 120.305 ;
        RECT 94.445 119.965 94.615 120.425 ;
        RECT 95.450 120.395 96.525 120.565 ;
        RECT 94.785 119.795 95.155 120.255 ;
        RECT 95.450 120.055 95.620 120.395 ;
        RECT 95.790 119.795 96.120 120.225 ;
        RECT 96.355 120.055 96.525 120.395 ;
        RECT 96.695 120.295 96.865 121.075 ;
        RECT 97.035 120.855 97.205 121.445 ;
        RECT 97.375 121.045 97.725 121.665 ;
        RECT 97.035 120.465 97.500 120.855 ;
        RECT 97.895 120.595 98.065 121.955 ;
        RECT 98.235 120.765 98.695 121.815 ;
        RECT 97.670 120.425 98.065 120.595 ;
        RECT 97.670 120.295 97.840 120.425 ;
        RECT 96.695 119.965 97.375 120.295 ;
        RECT 97.590 119.965 97.840 120.295 ;
        RECT 98.010 119.795 98.260 120.255 ;
        RECT 98.430 119.980 98.755 120.765 ;
        RECT 98.925 119.965 99.095 122.085 ;
        RECT 99.265 121.965 99.595 122.345 ;
        RECT 99.765 121.795 100.020 122.085 ;
        RECT 99.270 121.625 100.020 121.795 ;
        RECT 99.270 120.635 99.500 121.625 ;
        RECT 100.195 121.620 100.485 122.345 ;
        RECT 101.885 121.875 102.055 122.345 ;
        RECT 102.225 121.695 102.555 122.175 ;
        RECT 102.725 121.875 102.895 122.345 ;
        RECT 103.065 121.695 103.395 122.175 ;
        RECT 101.630 121.525 103.395 121.695 ;
        RECT 103.565 121.535 103.735 122.345 ;
        RECT 103.935 121.965 105.005 122.135 ;
        RECT 103.935 121.610 104.255 121.965 ;
        RECT 99.670 120.805 100.020 121.455 ;
        RECT 101.630 120.975 102.040 121.525 ;
        RECT 103.930 121.355 104.255 121.610 ;
        RECT 102.225 121.145 104.255 121.355 ;
        RECT 103.910 121.135 104.255 121.145 ;
        RECT 104.425 121.395 104.665 121.795 ;
        RECT 104.835 121.735 105.005 121.965 ;
        RECT 105.175 121.905 105.365 122.345 ;
        RECT 105.535 121.895 106.485 122.175 ;
        RECT 106.705 121.985 107.055 122.155 ;
        RECT 104.835 121.565 105.365 121.735 ;
        RECT 99.270 120.465 100.020 120.635 ;
        RECT 99.265 119.795 99.595 120.295 ;
        RECT 99.765 119.965 100.020 120.465 ;
        RECT 100.195 119.795 100.485 120.960 ;
        RECT 101.630 120.805 103.355 120.975 ;
        RECT 101.885 119.795 102.055 120.635 ;
        RECT 102.265 119.965 102.515 120.805 ;
        RECT 102.725 119.795 102.895 120.635 ;
        RECT 103.065 119.965 103.355 120.805 ;
        RECT 103.565 119.795 103.735 120.855 ;
        RECT 103.910 120.515 104.080 121.135 ;
        RECT 104.425 121.025 104.965 121.395 ;
        RECT 105.145 121.285 105.365 121.565 ;
        RECT 105.535 121.115 105.705 121.895 ;
        RECT 105.300 120.945 105.705 121.115 ;
        RECT 105.875 121.105 106.225 121.725 ;
        RECT 105.300 120.855 105.470 120.945 ;
        RECT 106.395 120.935 106.605 121.725 ;
        RECT 104.250 120.685 105.470 120.855 ;
        RECT 105.930 120.775 106.605 120.935 ;
        RECT 103.910 120.345 104.710 120.515 ;
        RECT 104.030 119.795 104.360 120.175 ;
        RECT 104.540 120.055 104.710 120.345 ;
        RECT 105.300 120.305 105.470 120.685 ;
        RECT 105.640 120.765 106.605 120.775 ;
        RECT 106.795 121.595 107.055 121.985 ;
        RECT 107.265 121.885 107.595 122.345 ;
        RECT 108.470 121.955 109.325 122.125 ;
        RECT 109.530 121.955 110.025 122.125 ;
        RECT 110.195 121.985 110.525 122.345 ;
        RECT 106.795 120.905 106.965 121.595 ;
        RECT 107.135 121.245 107.305 121.425 ;
        RECT 107.475 121.415 108.265 121.665 ;
        RECT 108.470 121.245 108.640 121.955 ;
        RECT 108.810 121.445 109.165 121.665 ;
        RECT 107.135 121.075 108.825 121.245 ;
        RECT 105.640 120.475 106.100 120.765 ;
        RECT 106.795 120.735 108.295 120.905 ;
        RECT 106.795 120.595 106.965 120.735 ;
        RECT 106.405 120.425 106.965 120.595 ;
        RECT 104.880 119.795 105.130 120.255 ;
        RECT 105.300 119.965 106.170 120.305 ;
        RECT 106.405 119.965 106.575 120.425 ;
        RECT 107.410 120.395 108.485 120.565 ;
        RECT 106.745 119.795 107.115 120.255 ;
        RECT 107.410 120.055 107.580 120.395 ;
        RECT 107.750 119.795 108.080 120.225 ;
        RECT 108.315 120.055 108.485 120.395 ;
        RECT 108.655 120.295 108.825 121.075 ;
        RECT 108.995 120.855 109.165 121.445 ;
        RECT 109.335 121.045 109.685 121.665 ;
        RECT 108.995 120.465 109.460 120.855 ;
        RECT 109.855 120.595 110.025 121.955 ;
        RECT 110.195 120.765 110.655 121.815 ;
        RECT 109.630 120.425 110.025 120.595 ;
        RECT 109.630 120.295 109.800 120.425 ;
        RECT 108.655 119.965 109.335 120.295 ;
        RECT 109.550 119.965 109.800 120.295 ;
        RECT 109.970 119.795 110.220 120.255 ;
        RECT 110.390 119.980 110.715 120.765 ;
        RECT 110.885 119.965 111.055 122.085 ;
        RECT 111.225 121.965 111.555 122.345 ;
        RECT 111.725 121.795 111.980 122.085 ;
        RECT 111.230 121.625 111.980 121.795 ;
        RECT 111.230 120.635 111.460 121.625 ;
        RECT 112.155 121.595 113.365 122.345 ;
        RECT 111.630 120.805 111.980 121.455 ;
        RECT 112.155 120.885 112.675 121.425 ;
        RECT 112.845 121.055 113.365 121.595 ;
        RECT 111.230 120.465 111.980 120.635 ;
        RECT 111.225 119.795 111.555 120.295 ;
        RECT 111.725 119.965 111.980 120.465 ;
        RECT 112.155 119.795 113.365 120.885 ;
        RECT 26.970 119.625 113.450 119.795 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 46.820 206.990 47.140 207.050 ;
        RECT 99.720 206.990 100.040 207.050 ;
        RECT 46.820 206.850 100.040 206.990 ;
        RECT 46.820 206.790 47.140 206.850 ;
        RECT 99.720 206.790 100.040 206.850 ;
        RECT 54.180 205.970 54.500 206.030 ;
        RECT 84.080 205.970 84.400 206.030 ;
        RECT 54.180 205.830 84.400 205.970 ;
        RECT 54.180 205.770 54.500 205.830 ;
        RECT 84.080 205.770 84.400 205.830 ;
        RECT 88.680 205.970 89.000 206.030 ;
        RECT 111.220 205.970 111.540 206.030 ;
        RECT 88.680 205.830 111.540 205.970 ;
        RECT 88.680 205.770 89.000 205.830 ;
        RECT 111.220 205.770 111.540 205.830 ;
        RECT 45.900 205.630 46.220 205.690 ;
        RECT 94.660 205.630 94.980 205.690 ;
        RECT 45.900 205.490 94.980 205.630 ;
        RECT 45.900 205.430 46.220 205.490 ;
        RECT 94.660 205.430 94.980 205.490 ;
        RECT 40.840 205.290 41.160 205.350 ;
        RECT 95.120 205.290 95.440 205.350 ;
        RECT 40.840 205.150 95.440 205.290 ;
        RECT 40.840 205.090 41.160 205.150 ;
        RECT 95.120 205.090 95.440 205.150 ;
        RECT 56.940 204.950 57.260 205.010 ;
        RECT 68.900 204.950 69.220 205.010 ;
        RECT 56.940 204.810 69.220 204.950 ;
        RECT 56.940 204.750 57.260 204.810 ;
        RECT 68.900 204.750 69.220 204.810 ;
        RECT 81.780 204.950 82.100 205.010 ;
        RECT 88.680 204.950 89.000 205.010 ;
        RECT 81.780 204.810 89.000 204.950 ;
        RECT 81.780 204.750 82.100 204.810 ;
        RECT 88.680 204.750 89.000 204.810 ;
        RECT 89.140 204.950 89.460 205.010 ;
        RECT 107.080 204.950 107.400 205.010 ;
        RECT 89.140 204.810 107.400 204.950 ;
        RECT 89.140 204.750 89.460 204.810 ;
        RECT 107.080 204.750 107.400 204.810 ;
        RECT 39.000 204.610 39.320 204.670 ;
        RECT 96.040 204.610 96.360 204.670 ;
        RECT 39.000 204.470 96.360 204.610 ;
        RECT 39.000 204.410 39.320 204.470 ;
        RECT 96.040 204.410 96.360 204.470 ;
        RECT 26.970 203.790 113.450 204.270 ;
        RECT 39.920 203.390 40.240 203.650 ;
        RECT 40.840 203.390 41.160 203.650 ;
        RECT 44.980 203.390 45.300 203.650 ;
        RECT 46.820 203.390 47.140 203.650 ;
        RECT 61.540 203.590 61.860 203.650 ;
        RECT 62.475 203.590 62.765 203.635 ;
        RECT 63.380 203.590 63.700 203.650 ;
        RECT 69.360 203.590 69.680 203.650 ;
        RECT 47.370 203.450 59.010 203.590 ;
        RECT 47.370 203.250 47.510 203.450 ;
        RECT 41.850 203.110 47.510 203.250 ;
        RECT 29.815 202.910 30.105 202.955 ;
        RECT 30.275 202.910 30.565 202.955 ;
        RECT 31.655 202.910 31.945 202.955 ;
        RECT 32.560 202.910 32.880 202.970 ;
        RECT 29.815 202.770 32.880 202.910 ;
        RECT 29.815 202.725 30.105 202.770 ;
        RECT 30.275 202.725 30.565 202.770 ;
        RECT 31.655 202.725 31.945 202.770 ;
        RECT 32.560 202.710 32.880 202.770 ;
        RECT 39.000 202.710 39.320 202.970 ;
        RECT 41.850 202.955 41.990 203.110 ;
        RECT 41.315 202.910 41.605 202.955 ;
        RECT 41.775 202.910 42.065 202.955 ;
        RECT 41.315 202.770 42.065 202.910 ;
        RECT 41.315 202.725 41.605 202.770 ;
        RECT 41.775 202.725 42.065 202.770 ;
        RECT 43.140 202.710 43.460 202.970 ;
        RECT 44.610 202.955 44.750 203.110 ;
        RECT 44.535 202.725 44.825 202.955 ;
        RECT 45.900 202.710 46.220 202.970 ;
        RECT 47.295 202.910 47.585 202.955 ;
        RECT 49.580 202.910 49.900 202.970 ;
        RECT 50.130 202.955 50.270 203.450 ;
        RECT 50.500 203.250 50.820 203.310 ;
        RECT 57.860 203.250 58.180 203.310 ;
        RECT 50.500 203.110 58.180 203.250 ;
        RECT 50.500 203.050 50.820 203.110 ;
        RECT 57.860 203.050 58.180 203.110 ;
        RECT 58.870 203.250 59.010 203.450 ;
        RECT 61.540 203.450 62.765 203.590 ;
        RECT 61.540 203.390 61.860 203.450 ;
        RECT 62.475 203.405 62.765 203.450 ;
        RECT 63.010 203.450 63.700 203.590 ;
        RECT 63.010 203.295 63.150 203.450 ;
        RECT 63.380 203.390 63.700 203.450 ;
        RECT 64.390 203.450 69.680 203.590 ;
        RECT 58.870 203.110 61.770 203.250 ;
        RECT 47.295 202.770 49.900 202.910 ;
        RECT 47.295 202.725 47.585 202.770 ;
        RECT 49.580 202.710 49.900 202.770 ;
        RECT 50.055 202.725 50.345 202.955 ;
        RECT 51.420 202.910 51.740 202.970 ;
        RECT 52.355 202.910 52.645 202.955 ;
        RECT 51.420 202.770 52.645 202.910 ;
        RECT 51.420 202.710 51.740 202.770 ;
        RECT 52.355 202.725 52.645 202.770 ;
        RECT 53.275 202.725 53.565 202.955 ;
        RECT 42.220 202.370 42.540 202.630 ;
        RECT 29.355 202.230 29.645 202.275 ;
        RECT 43.600 202.230 43.920 202.290 ;
        RECT 29.355 202.090 43.920 202.230 ;
        RECT 29.355 202.045 29.645 202.090 ;
        RECT 43.600 202.030 43.920 202.090 ;
        RECT 44.075 202.230 44.365 202.275 ;
        RECT 52.800 202.230 53.120 202.290 ;
        RECT 44.075 202.090 53.120 202.230 ;
        RECT 44.075 202.045 44.365 202.090 ;
        RECT 52.800 202.030 53.120 202.090 ;
        RECT 27.500 201.890 27.820 201.950 ;
        RECT 30.735 201.890 31.025 201.935 ;
        RECT 27.500 201.750 31.025 201.890 ;
        RECT 27.500 201.690 27.820 201.750 ;
        RECT 30.735 201.705 31.025 201.750 ;
        RECT 32.100 201.690 32.420 201.950 ;
        RECT 48.215 201.890 48.505 201.935 ;
        RECT 50.040 201.890 50.360 201.950 ;
        RECT 48.215 201.750 50.360 201.890 ;
        RECT 48.215 201.705 48.505 201.750 ;
        RECT 50.040 201.690 50.360 201.750 ;
        RECT 50.500 201.690 50.820 201.950 ;
        RECT 50.960 201.890 51.280 201.950 ;
        RECT 51.895 201.890 52.185 201.935 ;
        RECT 50.960 201.750 52.185 201.890 ;
        RECT 53.350 201.890 53.490 202.725 ;
        RECT 54.640 202.710 54.960 202.970 ;
        RECT 56.020 202.710 56.340 202.970 ;
        RECT 56.940 202.710 57.260 202.970 ;
        RECT 58.870 202.955 59.010 203.110 ;
        RECT 58.335 202.910 58.625 202.955 ;
        RECT 58.795 202.910 59.085 202.955 ;
        RECT 58.335 202.770 59.085 202.910 ;
        RECT 58.335 202.725 58.625 202.770 ;
        RECT 58.795 202.725 59.085 202.770 ;
        RECT 61.080 202.710 61.400 202.970 ;
        RECT 61.630 202.910 61.770 203.110 ;
        RECT 62.935 203.065 63.225 203.295 ;
        RECT 63.380 202.910 63.700 202.970 ;
        RECT 61.630 202.770 63.700 202.910 ;
        RECT 63.380 202.710 63.700 202.770 ;
        RECT 63.855 202.910 64.145 202.955 ;
        RECT 64.390 202.910 64.530 203.450 ;
        RECT 69.360 203.390 69.680 203.450 ;
        RECT 69.820 203.590 70.140 203.650 ;
        RECT 75.815 203.590 76.105 203.635 ;
        RECT 91.900 203.590 92.220 203.650 ;
        RECT 69.820 203.450 92.220 203.590 ;
        RECT 69.820 203.390 70.140 203.450 ;
        RECT 75.815 203.405 76.105 203.450 ;
        RECT 91.900 203.390 92.220 203.450 ;
        RECT 96.040 203.390 96.360 203.650 ;
        RECT 100.180 203.590 100.500 203.650 ;
        RECT 100.180 203.450 110.070 203.590 ;
        RECT 100.180 203.390 100.500 203.450 ;
        RECT 81.780 203.295 82.100 203.310 ;
        RECT 70.755 203.250 71.045 203.295 ;
        RECT 64.850 203.110 71.045 203.250 ;
        RECT 64.850 202.970 64.990 203.110 ;
        RECT 70.755 203.065 71.045 203.110 ;
        RECT 78.215 203.250 78.505 203.295 ;
        RECT 81.455 203.250 82.105 203.295 ;
        RECT 78.215 203.110 82.105 203.250 ;
        RECT 78.215 203.065 78.805 203.110 ;
        RECT 81.455 203.065 82.105 203.110 ;
        RECT 84.540 203.250 84.860 203.310 ;
        RECT 91.440 203.250 91.760 203.310 ;
        RECT 92.375 203.250 92.665 203.295 ;
        RECT 84.540 203.110 85.690 203.250 ;
        RECT 63.855 202.770 64.530 202.910 ;
        RECT 63.855 202.725 64.145 202.770 ;
        RECT 64.760 202.710 65.080 202.970 ;
        RECT 65.680 202.910 66.000 202.970 ;
        RECT 67.995 202.910 68.285 202.955 ;
        RECT 65.680 202.770 68.285 202.910 ;
        RECT 65.680 202.710 66.000 202.770 ;
        RECT 67.995 202.725 68.285 202.770 ;
        RECT 68.900 202.710 69.220 202.970 ;
        RECT 69.360 202.710 69.680 202.970 ;
        RECT 71.200 202.910 71.520 202.970 ;
        RECT 75.340 202.910 75.660 202.970 ;
        RECT 71.200 202.770 75.660 202.910 ;
        RECT 71.200 202.710 71.520 202.770 ;
        RECT 75.340 202.710 75.660 202.770 ;
        RECT 78.515 202.750 78.805 203.065 ;
        RECT 81.780 203.050 82.100 203.065 ;
        RECT 84.540 203.050 84.860 203.110 ;
        RECT 85.550 202.955 85.690 203.110 ;
        RECT 91.440 203.110 92.665 203.250 ;
        RECT 91.440 203.050 91.760 203.110 ;
        RECT 92.375 203.065 92.665 203.110 ;
        RECT 95.120 203.250 95.440 203.310 ;
        RECT 102.135 203.250 102.425 203.295 ;
        RECT 105.375 203.250 106.025 203.295 ;
        RECT 95.120 203.110 106.025 203.250 ;
        RECT 95.120 203.050 95.440 203.110 ;
        RECT 102.135 203.065 102.725 203.110 ;
        RECT 105.375 203.065 106.025 203.110 ;
        RECT 79.595 202.910 79.885 202.955 ;
        RECT 83.175 202.910 83.465 202.955 ;
        RECT 85.010 202.910 85.300 202.955 ;
        RECT 79.595 202.770 85.300 202.910 ;
        RECT 79.595 202.725 79.885 202.770 ;
        RECT 83.175 202.725 83.465 202.770 ;
        RECT 85.010 202.725 85.300 202.770 ;
        RECT 85.475 202.725 85.765 202.955 ;
        RECT 86.840 202.710 87.160 202.970 ;
        RECT 89.140 202.710 89.460 202.970 ;
        RECT 91.915 202.910 92.205 202.955 ;
        RECT 97.420 202.910 97.740 202.970 ;
        RECT 97.895 202.910 98.185 202.955 ;
        RECT 91.915 202.770 98.185 202.910 ;
        RECT 91.915 202.725 92.205 202.770 ;
        RECT 97.420 202.710 97.740 202.770 ;
        RECT 97.895 202.725 98.185 202.770 ;
        RECT 102.435 202.750 102.725 203.065 ;
        RECT 108.000 203.050 108.320 203.310 ;
        RECT 109.930 202.955 110.070 203.450 ;
        RECT 103.515 202.910 103.805 202.955 ;
        RECT 107.095 202.910 107.385 202.955 ;
        RECT 108.930 202.910 109.220 202.955 ;
        RECT 103.515 202.770 109.220 202.910 ;
        RECT 103.515 202.725 103.805 202.770 ;
        RECT 107.095 202.725 107.385 202.770 ;
        RECT 108.930 202.725 109.220 202.770 ;
        RECT 109.855 202.725 110.145 202.955 ;
        RECT 64.300 202.570 64.620 202.630 ;
        RECT 55.650 202.430 64.620 202.570 ;
        RECT 54.180 202.030 54.500 202.290 ;
        RECT 55.650 202.275 55.790 202.430 ;
        RECT 64.300 202.370 64.620 202.430 ;
        RECT 65.220 202.370 65.540 202.630 ;
        RECT 68.455 202.570 68.745 202.615 ;
        RECT 73.040 202.570 73.360 202.630 ;
        RECT 73.515 202.570 73.805 202.615 ;
        RECT 76.735 202.570 77.025 202.615 ;
        RECT 65.770 202.430 70.740 202.570 ;
        RECT 55.575 202.045 55.865 202.275 ;
        RECT 56.480 202.030 56.800 202.290 ;
        RECT 58.780 202.230 59.100 202.290 ;
        RECT 57.030 202.090 59.100 202.230 ;
        RECT 57.030 201.890 57.170 202.090 ;
        RECT 58.780 202.030 59.100 202.090 ;
        RECT 59.255 202.230 59.545 202.275 ;
        RECT 64.760 202.230 65.080 202.290 ;
        RECT 65.770 202.230 65.910 202.430 ;
        RECT 68.455 202.385 68.745 202.430 ;
        RECT 70.600 202.290 70.740 202.430 ;
        RECT 73.040 202.430 77.025 202.570 ;
        RECT 73.040 202.370 73.360 202.430 ;
        RECT 73.515 202.385 73.805 202.430 ;
        RECT 76.735 202.385 77.025 202.430 ;
        RECT 84.095 202.570 84.385 202.615 ;
        RECT 95.595 202.570 95.885 202.615 ;
        RECT 96.500 202.570 96.820 202.630 ;
        RECT 84.095 202.430 95.350 202.570 ;
        RECT 84.095 202.385 84.385 202.430 ;
        RECT 59.255 202.090 65.080 202.230 ;
        RECT 59.255 202.045 59.545 202.090 ;
        RECT 64.760 202.030 65.080 202.090 ;
        RECT 65.310 202.090 65.910 202.230 ;
        RECT 66.615 202.230 66.905 202.275 ;
        RECT 67.520 202.230 67.840 202.290 ;
        RECT 66.615 202.090 67.840 202.230 ;
        RECT 70.600 202.230 71.060 202.290 ;
        RECT 75.800 202.230 76.120 202.290 ;
        RECT 70.600 202.090 76.120 202.230 ;
        RECT 53.350 201.750 57.170 201.890 ;
        RECT 57.400 201.890 57.720 201.950 ;
        RECT 57.875 201.890 58.165 201.935 ;
        RECT 57.400 201.750 58.165 201.890 ;
        RECT 50.960 201.690 51.280 201.750 ;
        RECT 51.895 201.705 52.185 201.750 ;
        RECT 57.400 201.690 57.720 201.750 ;
        RECT 57.875 201.705 58.165 201.750 ;
        RECT 58.320 201.890 58.640 201.950 ;
        RECT 60.175 201.890 60.465 201.935 ;
        RECT 58.320 201.750 60.465 201.890 ;
        RECT 58.320 201.690 58.640 201.750 ;
        RECT 60.175 201.705 60.465 201.750 ;
        RECT 61.540 201.890 61.860 201.950 ;
        RECT 65.310 201.890 65.450 202.090 ;
        RECT 66.615 202.045 66.905 202.090 ;
        RECT 67.520 202.030 67.840 202.090 ;
        RECT 70.740 202.030 71.060 202.090 ;
        RECT 75.800 202.030 76.120 202.090 ;
        RECT 79.595 202.230 79.885 202.275 ;
        RECT 82.715 202.230 83.005 202.275 ;
        RECT 84.605 202.230 84.895 202.275 ;
        RECT 79.595 202.090 84.895 202.230 ;
        RECT 79.595 202.045 79.885 202.090 ;
        RECT 82.715 202.045 83.005 202.090 ;
        RECT 84.605 202.045 84.895 202.090 ;
        RECT 61.540 201.750 65.450 201.890 ;
        RECT 61.540 201.690 61.860 201.750 ;
        RECT 65.680 201.690 66.000 201.950 ;
        RECT 67.060 201.690 67.380 201.950 ;
        RECT 80.860 201.890 81.180 201.950 ;
        RECT 86.395 201.890 86.685 201.935 ;
        RECT 80.860 201.750 86.685 201.890 ;
        RECT 95.210 201.890 95.350 202.430 ;
        RECT 95.595 202.430 96.820 202.570 ;
        RECT 95.595 202.385 95.885 202.430 ;
        RECT 96.500 202.370 96.820 202.430 ;
        RECT 96.960 202.570 97.280 202.630 ;
        RECT 98.355 202.570 98.645 202.615 ;
        RECT 96.960 202.430 98.645 202.570 ;
        RECT 96.960 202.370 97.280 202.430 ;
        RECT 98.355 202.385 98.645 202.430 ;
        RECT 99.260 202.370 99.580 202.630 ;
        RECT 109.395 202.570 109.685 202.615 ;
        RECT 110.300 202.570 110.620 202.630 ;
        RECT 109.395 202.430 110.620 202.570 ;
        RECT 109.395 202.385 109.685 202.430 ;
        RECT 110.300 202.370 110.620 202.430 ;
        RECT 100.640 202.030 100.960 202.290 ;
        RECT 103.515 202.230 103.805 202.275 ;
        RECT 106.635 202.230 106.925 202.275 ;
        RECT 108.525 202.230 108.815 202.275 ;
        RECT 103.515 202.090 108.815 202.230 ;
        RECT 103.515 202.045 103.805 202.090 ;
        RECT 106.635 202.045 106.925 202.090 ;
        RECT 108.525 202.045 108.815 202.090 ;
        RECT 110.315 201.890 110.605 201.935 ;
        RECT 95.210 201.750 110.605 201.890 ;
        RECT 80.860 201.690 81.180 201.750 ;
        RECT 86.395 201.705 86.685 201.750 ;
        RECT 110.315 201.705 110.605 201.750 ;
        RECT 26.970 201.070 113.450 201.550 ;
        RECT 56.940 200.870 57.260 200.930 ;
        RECT 74.880 200.870 75.200 200.930 ;
        RECT 52.430 200.730 57.260 200.870 ;
        RECT 26.580 200.530 26.900 200.590 ;
        RECT 39.475 200.530 39.765 200.575 ;
        RECT 47.280 200.530 47.600 200.590 ;
        RECT 26.580 200.390 39.765 200.530 ;
        RECT 26.580 200.330 26.900 200.390 ;
        RECT 39.475 200.345 39.765 200.390 ;
        RECT 45.530 200.390 47.600 200.530 ;
        RECT 25.200 200.190 25.520 200.250 ;
        RECT 30.735 200.190 31.025 200.235 ;
        RECT 25.200 200.050 31.025 200.190 ;
        RECT 25.200 199.990 25.520 200.050 ;
        RECT 30.735 200.005 31.025 200.050 ;
        RECT 28.420 199.850 28.740 199.910 ;
        RECT 28.895 199.850 29.185 199.895 ;
        RECT 28.420 199.710 29.185 199.850 ;
        RECT 28.420 199.650 28.740 199.710 ;
        RECT 28.895 199.665 29.185 199.710 ;
        RECT 29.340 199.850 29.660 199.910 ;
        RECT 30.275 199.850 30.565 199.895 ;
        RECT 31.655 199.850 31.945 199.895 ;
        RECT 29.340 199.710 31.945 199.850 ;
        RECT 29.340 199.650 29.660 199.710 ;
        RECT 30.275 199.665 30.565 199.710 ;
        RECT 31.655 199.665 31.945 199.710 ;
        RECT 32.560 199.850 32.880 199.910 ;
        RECT 33.955 199.850 34.245 199.895 ;
        RECT 32.560 199.710 34.245 199.850 ;
        RECT 32.560 199.650 32.880 199.710 ;
        RECT 33.955 199.665 34.245 199.710 ;
        RECT 34.415 199.850 34.705 199.895 ;
        RECT 34.860 199.850 35.180 199.910 ;
        RECT 34.415 199.710 35.180 199.850 ;
        RECT 34.415 199.665 34.705 199.710 ;
        RECT 34.860 199.650 35.180 199.710 ;
        RECT 36.240 199.850 36.560 199.910 ;
        RECT 36.715 199.850 37.005 199.895 ;
        RECT 36.240 199.710 37.005 199.850 ;
        RECT 36.240 199.650 36.560 199.710 ;
        RECT 36.715 199.665 37.005 199.710 ;
        RECT 38.080 199.650 38.400 199.910 ;
        RECT 40.840 199.650 41.160 199.910 ;
        RECT 41.315 199.665 41.605 199.895 ;
        RECT 32.115 199.510 32.405 199.555 ;
        RECT 30.350 199.370 32.405 199.510 ;
        RECT 30.350 199.230 30.490 199.370 ;
        RECT 32.115 199.325 32.405 199.370 ;
        RECT 39.920 199.510 40.240 199.570 ;
        RECT 41.390 199.510 41.530 199.665 ;
        RECT 41.760 199.650 42.080 199.910 ;
        RECT 42.680 199.650 43.000 199.910 ;
        RECT 44.060 199.650 44.380 199.910 ;
        RECT 45.530 199.895 45.670 200.390 ;
        RECT 47.280 200.330 47.600 200.390 ;
        RECT 47.755 200.530 48.045 200.575 ;
        RECT 52.430 200.530 52.570 200.730 ;
        RECT 56.940 200.670 57.260 200.730 ;
        RECT 60.710 200.730 69.590 200.870 ;
        RECT 47.755 200.390 52.570 200.530 ;
        RECT 53.225 200.530 53.515 200.575 ;
        RECT 55.115 200.530 55.405 200.575 ;
        RECT 58.235 200.530 58.525 200.575 ;
        RECT 53.225 200.390 58.525 200.530 ;
        RECT 47.755 200.345 48.045 200.390 ;
        RECT 53.225 200.345 53.515 200.390 ;
        RECT 55.115 200.345 55.405 200.390 ;
        RECT 58.235 200.345 58.525 200.390 ;
        RECT 48.675 200.190 48.965 200.235 ;
        RECT 45.990 200.050 48.965 200.190 ;
        RECT 45.990 199.895 46.130 200.050 ;
        RECT 48.675 200.005 48.965 200.050 ;
        RECT 53.735 200.190 54.025 200.235 ;
        RECT 55.560 200.190 55.880 200.250 ;
        RECT 53.735 200.050 55.880 200.190 ;
        RECT 53.735 200.005 54.025 200.050 ;
        RECT 55.560 199.990 55.880 200.050 ;
        RECT 56.480 200.190 56.800 200.250 ;
        RECT 60.710 200.190 60.850 200.730 ;
        RECT 64.300 200.530 64.620 200.590 ;
        RECT 69.450 200.530 69.590 200.730 ;
        RECT 71.290 200.730 75.200 200.870 ;
        RECT 71.290 200.530 71.430 200.730 ;
        RECT 74.880 200.670 75.200 200.730 ;
        RECT 75.340 200.870 75.660 200.930 ;
        RECT 79.495 200.870 79.785 200.915 ;
        RECT 96.960 200.870 97.280 200.930 ;
        RECT 75.340 200.730 79.785 200.870 ;
        RECT 75.340 200.670 75.660 200.730 ;
        RECT 79.495 200.685 79.785 200.730 ;
        RECT 89.690 200.730 97.280 200.870 ;
        RECT 64.300 200.390 68.670 200.530 ;
        RECT 69.450 200.390 71.430 200.530 ;
        RECT 71.625 200.530 71.915 200.575 ;
        RECT 73.515 200.530 73.805 200.575 ;
        RECT 76.635 200.530 76.925 200.575 ;
        RECT 71.625 200.390 76.925 200.530 ;
        RECT 64.300 200.330 64.620 200.390 ;
        RECT 56.480 200.050 60.850 200.190 ;
        RECT 61.095 200.190 61.385 200.235 ;
        RECT 62.475 200.190 62.765 200.235 ;
        RECT 66.140 200.190 66.460 200.250 ;
        RECT 61.095 200.050 66.460 200.190 ;
        RECT 56.480 199.990 56.800 200.050 ;
        RECT 61.095 200.005 61.385 200.050 ;
        RECT 62.475 200.005 62.765 200.050 ;
        RECT 66.140 199.990 66.460 200.050 ;
        RECT 67.980 199.990 68.300 200.250 ;
        RECT 68.530 200.190 68.670 200.390 ;
        RECT 71.625 200.345 71.915 200.390 ;
        RECT 73.515 200.345 73.805 200.390 ;
        RECT 76.635 200.345 76.925 200.390 ;
        RECT 83.175 200.530 83.465 200.575 ;
        RECT 89.690 200.530 89.830 200.730 ;
        RECT 96.960 200.670 97.280 200.730 ;
        RECT 83.175 200.390 89.830 200.530 ;
        RECT 90.025 200.530 90.315 200.575 ;
        RECT 91.915 200.530 92.205 200.575 ;
        RECT 95.035 200.530 95.325 200.575 ;
        RECT 90.025 200.390 95.325 200.530 ;
        RECT 83.175 200.345 83.465 200.390 ;
        RECT 90.025 200.345 90.315 200.390 ;
        RECT 91.915 200.345 92.205 200.390 ;
        RECT 95.035 200.345 95.325 200.390 ;
        RECT 96.040 200.330 96.360 200.590 ;
        RECT 99.225 200.530 99.515 200.575 ;
        RECT 101.115 200.530 101.405 200.575 ;
        RECT 104.235 200.530 104.525 200.575 ;
        RECT 99.225 200.390 104.525 200.530 ;
        RECT 99.225 200.345 99.515 200.390 ;
        RECT 101.115 200.345 101.405 200.390 ;
        RECT 104.235 200.345 104.525 200.390 ;
        RECT 72.135 200.190 72.425 200.235 ;
        RECT 68.530 200.050 72.425 200.190 ;
        RECT 72.135 200.005 72.425 200.050 ;
        RECT 83.620 199.990 83.940 200.250 ;
        RECT 84.080 200.190 84.400 200.250 ;
        RECT 90.535 200.190 90.825 200.235 ;
        RECT 84.080 200.050 90.825 200.190 ;
        RECT 84.080 199.990 84.400 200.050 ;
        RECT 90.535 200.005 90.825 200.050 ;
        RECT 90.980 200.190 91.300 200.250 ;
        RECT 96.130 200.190 96.270 200.330 ;
        RECT 97.895 200.190 98.185 200.235 ;
        RECT 90.980 200.050 98.185 200.190 ;
        RECT 90.980 199.990 91.300 200.050 ;
        RECT 97.895 200.005 98.185 200.050 ;
        RECT 99.720 199.990 100.040 200.250 ;
        RECT 45.455 199.665 45.745 199.895 ;
        RECT 45.915 199.665 46.205 199.895 ;
        RECT 47.280 199.850 47.600 199.910 ;
        RECT 49.120 199.850 49.440 199.910 ;
        RECT 51.420 199.850 51.740 199.910 ;
        RECT 47.280 199.710 51.740 199.850 ;
        RECT 47.280 199.650 47.600 199.710 ;
        RECT 49.120 199.650 49.440 199.710 ;
        RECT 51.420 199.650 51.740 199.710 ;
        RECT 51.880 199.650 52.200 199.910 ;
        RECT 52.355 199.665 52.645 199.895 ;
        RECT 52.820 199.850 53.110 199.895 ;
        RECT 54.655 199.850 54.945 199.895 ;
        RECT 58.235 199.850 58.525 199.895 ;
        RECT 52.820 199.710 58.525 199.850 ;
        RECT 52.820 199.665 53.110 199.710 ;
        RECT 54.655 199.665 54.945 199.710 ;
        RECT 58.235 199.665 58.525 199.710 ;
        RECT 39.920 199.370 41.530 199.510 ;
        RECT 43.615 199.510 43.905 199.555 ;
        RECT 50.040 199.510 50.360 199.570 ;
        RECT 43.615 199.370 50.360 199.510 ;
        RECT 52.430 199.510 52.570 199.665 ;
        RECT 53.720 199.510 54.040 199.570 ;
        RECT 52.430 199.370 54.040 199.510 ;
        RECT 39.920 199.310 40.240 199.370 ;
        RECT 43.615 199.325 43.905 199.370 ;
        RECT 50.040 199.310 50.360 199.370 ;
        RECT 53.720 199.310 54.040 199.370 ;
        RECT 56.015 199.510 56.665 199.555 ;
        RECT 57.400 199.510 57.720 199.570 ;
        RECT 59.315 199.555 59.605 199.870 ;
        RECT 65.235 199.850 65.525 199.895 ;
        RECT 67.535 199.850 67.825 199.895 ;
        RECT 65.235 199.710 67.825 199.850 ;
        RECT 65.235 199.665 65.525 199.710 ;
        RECT 67.535 199.665 67.825 199.710 ;
        RECT 68.915 199.665 69.205 199.895 ;
        RECT 70.755 199.665 71.045 199.895 ;
        RECT 71.220 199.850 71.510 199.895 ;
        RECT 73.055 199.850 73.345 199.895 ;
        RECT 76.635 199.850 76.925 199.895 ;
        RECT 71.220 199.710 76.925 199.850 ;
        RECT 71.220 199.665 71.510 199.710 ;
        RECT 73.055 199.665 73.345 199.710 ;
        RECT 76.635 199.665 76.925 199.710 ;
        RECT 59.315 199.510 59.905 199.555 ;
        RECT 56.015 199.370 59.905 199.510 ;
        RECT 56.015 199.325 56.665 199.370 ;
        RECT 57.400 199.310 57.720 199.370 ;
        RECT 59.615 199.325 59.905 199.370 ;
        RECT 63.840 199.510 64.160 199.570 ;
        RECT 66.600 199.510 66.920 199.570 ;
        RECT 68.990 199.510 69.130 199.665 ;
        RECT 63.840 199.370 66.370 199.510 ;
        RECT 63.840 199.310 64.160 199.370 ;
        RECT 29.800 198.970 30.120 199.230 ;
        RECT 30.260 198.970 30.580 199.230 ;
        RECT 31.180 199.170 31.500 199.230 ;
        RECT 33.495 199.170 33.785 199.215 ;
        RECT 31.180 199.030 33.785 199.170 ;
        RECT 31.180 198.970 31.500 199.030 ;
        RECT 33.495 198.985 33.785 199.030 ;
        RECT 35.320 198.970 35.640 199.230 ;
        RECT 37.635 199.170 37.925 199.215 ;
        RECT 38.540 199.170 38.860 199.230 ;
        RECT 37.635 199.030 38.860 199.170 ;
        RECT 37.635 198.985 37.925 199.030 ;
        RECT 38.540 198.970 38.860 199.030 ;
        RECT 39.000 198.970 39.320 199.230 ;
        RECT 44.980 198.970 45.300 199.230 ;
        RECT 46.835 199.170 47.125 199.215 ;
        RECT 52.800 199.170 53.120 199.230 ;
        RECT 46.835 199.030 53.120 199.170 ;
        RECT 46.835 198.985 47.125 199.030 ;
        RECT 52.800 198.970 53.120 199.030 ;
        RECT 55.560 199.170 55.880 199.230 ;
        RECT 65.695 199.170 65.985 199.215 ;
        RECT 55.560 199.030 65.985 199.170 ;
        RECT 66.230 199.170 66.370 199.370 ;
        RECT 66.600 199.370 69.130 199.510 ;
        RECT 66.600 199.310 66.920 199.370 ;
        RECT 69.360 199.170 69.680 199.230 ;
        RECT 66.230 199.030 69.680 199.170 ;
        RECT 55.560 198.970 55.880 199.030 ;
        RECT 65.695 198.985 65.985 199.030 ;
        RECT 69.360 198.970 69.680 199.030 ;
        RECT 69.820 198.970 70.140 199.230 ;
        RECT 70.830 199.170 70.970 199.665 ;
        RECT 77.715 199.555 78.005 199.870 ;
        RECT 80.415 199.850 80.705 199.895 ;
        RECT 88.220 199.850 88.540 199.910 ;
        RECT 80.415 199.710 88.540 199.850 ;
        RECT 80.415 199.665 80.705 199.710 ;
        RECT 88.220 199.650 88.540 199.710 ;
        RECT 88.695 199.665 88.985 199.895 ;
        RECT 89.155 199.665 89.445 199.895 ;
        RECT 89.620 199.850 89.910 199.895 ;
        RECT 91.455 199.850 91.745 199.895 ;
        RECT 95.035 199.850 95.325 199.895 ;
        RECT 89.620 199.710 95.325 199.850 ;
        RECT 89.620 199.665 89.910 199.710 ;
        RECT 91.455 199.665 91.745 199.710 ;
        RECT 95.035 199.665 95.325 199.710 ;
        RECT 74.415 199.510 75.065 199.555 ;
        RECT 77.715 199.510 78.305 199.555 ;
        RECT 80.860 199.510 81.180 199.570 ;
        RECT 74.415 199.370 81.180 199.510 ;
        RECT 74.415 199.325 75.065 199.370 ;
        RECT 78.015 199.325 78.305 199.370 ;
        RECT 80.860 199.310 81.180 199.370 ;
        RECT 82.700 199.510 83.020 199.570 ;
        RECT 88.770 199.510 88.910 199.665 ;
        RECT 82.700 199.370 88.910 199.510 ;
        RECT 82.700 199.310 83.020 199.370 ;
        RECT 87.850 199.230 87.990 199.370 ;
        RECT 84.540 199.170 84.860 199.230 ;
        RECT 70.830 199.030 84.860 199.170 ;
        RECT 84.540 198.970 84.860 199.030 ;
        RECT 86.840 198.970 87.160 199.230 ;
        RECT 87.760 198.970 88.080 199.230 ;
        RECT 88.235 199.170 88.525 199.215 ;
        RECT 88.680 199.170 89.000 199.230 ;
        RECT 88.235 199.030 89.000 199.170 ;
        RECT 89.230 199.170 89.370 199.665 ;
        RECT 96.115 199.555 96.405 199.870 ;
        RECT 98.355 199.665 98.645 199.895 ;
        RECT 98.820 199.850 99.110 199.895 ;
        RECT 100.655 199.850 100.945 199.895 ;
        RECT 104.235 199.850 104.525 199.895 ;
        RECT 98.820 199.710 104.525 199.850 ;
        RECT 98.820 199.665 99.110 199.710 ;
        RECT 100.655 199.665 100.945 199.710 ;
        RECT 104.235 199.665 104.525 199.710 ;
        RECT 105.240 199.870 105.560 199.910 ;
        RECT 92.815 199.510 93.465 199.555 ;
        RECT 96.115 199.510 96.705 199.555 ;
        RECT 97.880 199.510 98.200 199.570 ;
        RECT 92.815 199.370 98.200 199.510 ;
        RECT 92.815 199.325 93.465 199.370 ;
        RECT 96.415 199.325 96.705 199.370 ;
        RECT 97.880 199.310 98.200 199.370 ;
        RECT 98.430 199.230 98.570 199.665 ;
        RECT 105.240 199.650 105.605 199.870 ;
        RECT 106.620 199.850 106.940 199.910 ;
        RECT 107.555 199.850 107.845 199.895 ;
        RECT 106.620 199.710 107.845 199.850 ;
        RECT 106.620 199.650 106.940 199.710 ;
        RECT 107.555 199.665 107.845 199.710 ;
        RECT 105.315 199.555 105.605 199.650 ;
        RECT 102.015 199.510 102.665 199.555 ;
        RECT 105.315 199.510 105.905 199.555 ;
        RECT 102.015 199.370 105.905 199.510 ;
        RECT 102.015 199.325 102.665 199.370 ;
        RECT 105.615 199.325 105.905 199.370 ;
        RECT 98.340 199.170 98.660 199.230 ;
        RECT 89.230 199.030 98.660 199.170 ;
        RECT 88.235 198.985 88.525 199.030 ;
        RECT 88.680 198.970 89.000 199.030 ;
        RECT 98.340 198.970 98.660 199.030 ;
        RECT 107.080 198.970 107.400 199.230 ;
        RECT 110.760 198.970 111.080 199.230 ;
        RECT 26.970 198.350 113.450 198.830 ;
        RECT 51.420 198.150 51.740 198.210 ;
        RECT 55.100 198.150 55.420 198.210 ;
        RECT 58.780 198.150 59.100 198.210 ;
        RECT 42.310 198.010 55.420 198.150 ;
        RECT 32.100 197.810 32.420 197.870 ;
        RECT 41.760 197.810 42.080 197.870 ;
        RECT 32.100 197.670 33.710 197.810 ;
        RECT 32.100 197.610 32.420 197.670 ;
        RECT 33.570 197.530 33.710 197.670 ;
        RECT 35.410 197.670 42.080 197.810 ;
        RECT 29.340 197.470 29.660 197.530 ;
        RECT 33.035 197.470 33.325 197.515 ;
        RECT 29.340 197.330 33.325 197.470 ;
        RECT 29.340 197.270 29.660 197.330 ;
        RECT 33.035 197.285 33.325 197.330 ;
        RECT 33.480 197.270 33.800 197.530 ;
        RECT 35.410 197.515 35.550 197.670 ;
        RECT 41.760 197.610 42.080 197.670 ;
        RECT 35.335 197.285 35.625 197.515 ;
        RECT 39.475 197.285 39.765 197.515 ;
        RECT 39.935 197.470 40.225 197.515 ;
        RECT 40.380 197.470 40.700 197.530 ;
        RECT 42.310 197.515 42.450 198.010 ;
        RECT 51.420 197.950 51.740 198.010 ;
        RECT 55.100 197.950 55.420 198.010 ;
        RECT 56.570 198.010 59.100 198.150 ;
        RECT 55.560 197.810 55.880 197.870 ;
        RECT 43.230 197.670 55.880 197.810 ;
        RECT 43.230 197.530 43.370 197.670 ;
        RECT 55.560 197.610 55.880 197.670 ;
        RECT 39.935 197.330 40.700 197.470 ;
        RECT 39.935 197.285 40.225 197.330 ;
        RECT 26.120 197.130 26.440 197.190 ;
        RECT 28.435 197.130 28.725 197.175 ;
        RECT 26.120 196.990 28.725 197.130 ;
        RECT 26.120 196.930 26.440 196.990 ;
        RECT 28.435 196.945 28.725 196.990 ;
        RECT 31.640 197.130 31.960 197.190 ;
        RECT 39.550 197.130 39.690 197.285 ;
        RECT 40.380 197.270 40.700 197.330 ;
        RECT 41.315 197.285 41.605 197.515 ;
        RECT 42.235 197.285 42.525 197.515 ;
        RECT 31.640 196.990 39.690 197.130 ;
        RECT 31.640 196.930 31.960 196.990 ;
        RECT 27.960 196.790 28.280 196.850 ;
        RECT 32.575 196.790 32.865 196.835 ;
        RECT 27.960 196.650 32.865 196.790 ;
        RECT 27.960 196.590 28.280 196.650 ;
        RECT 32.575 196.605 32.865 196.650 ;
        RECT 38.095 196.790 38.385 196.835 ;
        RECT 39.000 196.790 39.320 196.850 ;
        RECT 41.390 196.790 41.530 197.285 ;
        RECT 42.680 197.270 43.000 197.530 ;
        RECT 43.140 197.270 43.460 197.530 ;
        RECT 45.455 197.470 45.745 197.515 ;
        RECT 46.360 197.470 46.680 197.530 ;
        RECT 56.570 197.515 56.710 198.010 ;
        RECT 58.780 197.950 59.100 198.010 ;
        RECT 59.240 198.150 59.560 198.210 ;
        RECT 59.240 198.010 67.750 198.150 ;
        RECT 59.240 197.950 59.560 198.010 ;
        RECT 58.320 197.610 58.640 197.870 ;
        RECT 60.615 197.810 61.265 197.855 ;
        RECT 64.215 197.810 64.505 197.855 ;
        RECT 64.760 197.810 65.080 197.870 ;
        RECT 60.615 197.670 65.080 197.810 ;
        RECT 67.610 197.810 67.750 198.010 ;
        RECT 67.980 197.950 68.300 198.210 ;
        RECT 68.455 198.150 68.745 198.195 ;
        RECT 70.740 198.150 71.060 198.210 ;
        RECT 68.455 198.010 71.060 198.150 ;
        RECT 68.455 197.965 68.745 198.010 ;
        RECT 70.740 197.950 71.060 198.010 ;
        RECT 73.500 198.150 73.820 198.210 ;
        RECT 82.700 198.150 83.020 198.210 ;
        RECT 73.500 198.010 83.020 198.150 ;
        RECT 73.500 197.950 73.820 198.010 ;
        RECT 82.700 197.950 83.020 198.010 ;
        RECT 83.620 198.150 83.940 198.210 ;
        RECT 91.440 198.150 91.760 198.210 ;
        RECT 83.620 198.010 91.760 198.150 ;
        RECT 83.620 197.950 83.940 198.010 ;
        RECT 91.440 197.950 91.760 198.010 ;
        RECT 95.120 197.950 95.440 198.210 ;
        RECT 96.960 197.950 97.280 198.210 ;
        RECT 97.420 197.950 97.740 198.210 ;
        RECT 97.970 198.010 110.990 198.150 ;
        RECT 84.100 197.810 84.390 197.855 ;
        RECT 85.960 197.810 86.250 197.855 ;
        RECT 67.610 197.670 78.330 197.810 ;
        RECT 60.615 197.625 61.265 197.670 ;
        RECT 63.915 197.625 64.505 197.670 ;
        RECT 45.455 197.330 46.680 197.470 ;
        RECT 45.455 197.285 45.745 197.330 ;
        RECT 46.360 197.270 46.680 197.330 ;
        RECT 56.495 197.285 56.785 197.515 ;
        RECT 57.420 197.470 57.710 197.515 ;
        RECT 59.255 197.470 59.545 197.515 ;
        RECT 62.835 197.470 63.125 197.515 ;
        RECT 57.420 197.330 63.125 197.470 ;
        RECT 57.420 197.285 57.710 197.330 ;
        RECT 59.255 197.285 59.545 197.330 ;
        RECT 62.835 197.285 63.125 197.330 ;
        RECT 63.915 197.310 64.205 197.625 ;
        RECT 64.760 197.610 65.080 197.670 ;
        RECT 67.535 197.470 67.825 197.515 ;
        RECT 68.440 197.470 68.760 197.530 ;
        RECT 64.850 197.330 68.760 197.470 ;
        RECT 64.850 197.190 64.990 197.330 ;
        RECT 67.535 197.285 67.825 197.330 ;
        RECT 68.440 197.270 68.760 197.330 ;
        RECT 68.900 197.270 69.220 197.530 ;
        RECT 69.375 197.470 69.665 197.515 ;
        RECT 69.835 197.470 70.125 197.515 ;
        RECT 70.280 197.470 70.600 197.530 ;
        RECT 69.375 197.330 70.600 197.470 ;
        RECT 69.375 197.285 69.665 197.330 ;
        RECT 69.835 197.285 70.125 197.330 ;
        RECT 44.520 196.930 44.840 197.190 ;
        RECT 45.900 197.130 46.220 197.190 ;
        RECT 48.215 197.130 48.505 197.175 ;
        RECT 45.900 196.990 48.505 197.130 ;
        RECT 45.900 196.930 46.220 196.990 ;
        RECT 48.215 196.945 48.505 196.990 ;
        RECT 52.340 196.930 52.660 197.190 ;
        RECT 53.720 197.130 54.040 197.190 ;
        RECT 56.955 197.130 57.245 197.175 ;
        RECT 53.720 196.990 57.245 197.130 ;
        RECT 53.720 196.930 54.040 196.990 ;
        RECT 56.955 196.945 57.245 196.990 ;
        RECT 64.760 196.930 65.080 197.190 ;
        RECT 66.600 197.130 66.920 197.190 ;
        RECT 65.310 196.990 66.920 197.130 ;
        RECT 38.095 196.650 39.320 196.790 ;
        RECT 38.095 196.605 38.385 196.650 ;
        RECT 39.000 196.590 39.320 196.650 ;
        RECT 40.010 196.650 41.530 196.790 ;
        RECT 44.060 196.790 44.380 196.850 ;
        RECT 57.825 196.790 58.115 196.835 ;
        RECT 59.715 196.790 60.005 196.835 ;
        RECT 62.835 196.790 63.125 196.835 ;
        RECT 44.060 196.650 56.940 196.790 ;
        RECT 40.010 196.510 40.150 196.650 ;
        RECT 44.060 196.590 44.380 196.650 ;
        RECT 31.655 196.450 31.945 196.495 ;
        RECT 32.100 196.450 32.420 196.510 ;
        RECT 31.655 196.310 32.420 196.450 ;
        RECT 31.655 196.265 31.945 196.310 ;
        RECT 32.100 196.250 32.420 196.310 ;
        RECT 33.940 196.250 34.260 196.510 ;
        RECT 37.620 196.450 37.940 196.510 ;
        RECT 38.555 196.450 38.845 196.495 ;
        RECT 37.620 196.310 38.845 196.450 ;
        RECT 37.620 196.250 37.940 196.310 ;
        RECT 38.555 196.265 38.845 196.310 ;
        RECT 39.920 196.250 40.240 196.510 ;
        RECT 40.855 196.450 41.145 196.495 ;
        RECT 45.440 196.450 45.760 196.510 ;
        RECT 40.855 196.310 45.760 196.450 ;
        RECT 40.855 196.265 41.145 196.310 ;
        RECT 45.440 196.250 45.760 196.310 ;
        RECT 46.820 196.450 47.140 196.510 ;
        RECT 49.135 196.450 49.425 196.495 ;
        RECT 46.820 196.310 49.425 196.450 ;
        RECT 46.820 196.250 47.140 196.310 ;
        RECT 49.135 196.265 49.425 196.310 ;
        RECT 53.275 196.450 53.565 196.495 ;
        RECT 54.180 196.450 54.500 196.510 ;
        RECT 53.275 196.310 54.500 196.450 ;
        RECT 56.800 196.450 56.940 196.650 ;
        RECT 57.825 196.650 63.125 196.790 ;
        RECT 57.825 196.605 58.115 196.650 ;
        RECT 59.715 196.605 60.005 196.650 ;
        RECT 62.835 196.605 63.125 196.650 ;
        RECT 63.840 196.790 64.160 196.850 ;
        RECT 65.310 196.790 65.450 196.990 ;
        RECT 66.600 196.930 66.920 196.990 ;
        RECT 67.075 197.130 67.365 197.175 ;
        RECT 69.450 197.130 69.590 197.285 ;
        RECT 70.280 197.270 70.600 197.330 ;
        RECT 71.675 197.470 71.965 197.515 ;
        RECT 73.040 197.470 73.360 197.530 ;
        RECT 71.675 197.330 73.360 197.470 ;
        RECT 71.675 197.285 71.965 197.330 ;
        RECT 73.040 197.270 73.360 197.330 ;
        RECT 74.895 197.285 75.185 197.515 ;
        RECT 75.800 197.470 76.120 197.530 ;
        RECT 77.195 197.470 77.485 197.515 ;
        RECT 75.800 197.330 77.485 197.470 ;
        RECT 67.075 196.990 69.590 197.130 ;
        RECT 67.075 196.945 67.365 196.990 ;
        RECT 71.200 196.930 71.520 197.190 ;
        RECT 72.120 197.175 72.440 197.190 ;
        RECT 72.120 196.945 72.550 197.175 ;
        RECT 72.120 196.930 72.440 196.945 ;
        RECT 63.840 196.650 65.450 196.790 ;
        RECT 66.140 196.790 66.460 196.850 ;
        RECT 74.970 196.790 75.110 197.285 ;
        RECT 75.800 197.270 76.120 197.330 ;
        RECT 77.195 197.285 77.485 197.330 ;
        RECT 75.340 197.130 75.660 197.190 ;
        RECT 76.720 197.130 77.040 197.190 ;
        RECT 75.340 196.990 77.040 197.130 ;
        RECT 78.190 197.130 78.330 197.670 ;
        RECT 84.100 197.670 86.250 197.810 ;
        RECT 84.100 197.625 84.390 197.670 ;
        RECT 85.960 197.625 86.250 197.670 ;
        RECT 86.880 197.810 87.170 197.855 ;
        RECT 88.680 197.810 89.000 197.870 ;
        RECT 90.140 197.810 90.430 197.855 ;
        RECT 86.880 197.670 90.430 197.810 ;
        RECT 86.880 197.625 87.170 197.670 ;
        RECT 79.940 197.270 80.260 197.530 ;
        RECT 83.175 197.470 83.465 197.515 ;
        RECT 84.540 197.470 84.860 197.530 ;
        RECT 83.175 197.330 84.860 197.470 ;
        RECT 83.175 197.285 83.465 197.330 ;
        RECT 84.540 197.270 84.860 197.330 ;
        RECT 85.000 197.270 85.320 197.530 ;
        RECT 86.035 197.470 86.250 197.625 ;
        RECT 88.680 197.610 89.000 197.670 ;
        RECT 90.140 197.625 90.430 197.670 ;
        RECT 90.980 197.810 91.300 197.870 ;
        RECT 94.675 197.810 94.965 197.855 ;
        RECT 90.980 197.670 94.965 197.810 ;
        RECT 90.980 197.610 91.300 197.670 ;
        RECT 94.675 197.625 94.965 197.670 ;
        RECT 95.580 197.810 95.900 197.870 ;
        RECT 97.970 197.810 98.110 198.010 ;
        RECT 95.580 197.670 98.110 197.810 ;
        RECT 98.800 197.810 99.120 197.870 ;
        RECT 103.055 197.810 103.345 197.855 ;
        RECT 106.295 197.810 106.945 197.855 ;
        RECT 98.800 197.670 106.945 197.810 ;
        RECT 88.280 197.470 88.570 197.515 ;
        RECT 86.035 197.330 88.570 197.470 ;
        RECT 88.280 197.285 88.570 197.330 ;
        RECT 91.900 197.470 92.220 197.530 ;
        RECT 93.755 197.470 94.045 197.515 ;
        RECT 91.900 197.330 94.045 197.470 ;
        RECT 94.750 197.470 94.890 197.625 ;
        RECT 95.580 197.610 95.900 197.670 ;
        RECT 98.800 197.610 99.120 197.670 ;
        RECT 103.055 197.625 103.645 197.670 ;
        RECT 106.295 197.625 106.945 197.670 ;
        RECT 100.180 197.470 100.500 197.530 ;
        RECT 94.750 197.330 100.500 197.470 ;
        RECT 91.900 197.270 92.220 197.330 ;
        RECT 93.755 197.285 94.045 197.330 ;
        RECT 100.180 197.270 100.500 197.330 ;
        RECT 103.355 197.310 103.645 197.625 ;
        RECT 108.920 197.610 109.240 197.870 ;
        RECT 104.435 197.470 104.725 197.515 ;
        RECT 108.015 197.470 108.305 197.515 ;
        RECT 109.850 197.470 110.140 197.515 ;
        RECT 104.435 197.330 110.140 197.470 ;
        RECT 104.435 197.285 104.725 197.330 ;
        RECT 108.015 197.285 108.305 197.330 ;
        RECT 109.850 197.285 110.140 197.330 ;
        RECT 110.300 197.270 110.620 197.530 ;
        RECT 110.850 197.470 110.990 198.010 ;
        RECT 111.220 197.950 111.540 198.210 ;
        RECT 111.680 197.470 112.000 197.530 ;
        RECT 110.850 197.330 112.000 197.470 ;
        RECT 111.680 197.270 112.000 197.330 ;
        RECT 84.080 197.130 84.400 197.190 ;
        RECT 78.190 196.990 84.400 197.130 ;
        RECT 75.340 196.930 75.660 196.990 ;
        RECT 76.720 196.930 77.040 196.990 ;
        RECT 84.080 196.930 84.400 196.990 ;
        RECT 86.840 197.130 87.160 197.190 ;
        RECT 96.960 197.130 97.280 197.190 ;
        RECT 86.840 196.990 97.280 197.130 ;
        RECT 86.840 196.930 87.160 196.990 ;
        RECT 96.960 196.930 97.280 196.990 ;
        RECT 98.355 197.130 98.645 197.175 ;
        RECT 98.800 197.130 99.120 197.190 ;
        RECT 99.720 197.130 100.040 197.190 ;
        RECT 98.355 196.990 100.040 197.130 ;
        RECT 98.355 196.945 98.645 196.990 ;
        RECT 98.800 196.930 99.120 196.990 ;
        RECT 99.720 196.930 100.040 196.990 ;
        RECT 105.240 197.130 105.560 197.190 ;
        RECT 111.220 197.130 111.540 197.190 ;
        RECT 105.240 196.990 111.540 197.130 ;
        RECT 105.240 196.930 105.560 196.990 ;
        RECT 111.220 196.930 111.540 196.990 ;
        RECT 66.140 196.650 75.110 196.790 ;
        RECT 83.640 196.790 83.930 196.835 ;
        RECT 85.500 196.790 85.790 196.835 ;
        RECT 88.280 196.790 88.570 196.835 ;
        RECT 83.640 196.650 88.570 196.790 ;
        RECT 63.840 196.590 64.160 196.650 ;
        RECT 66.140 196.590 66.460 196.650 ;
        RECT 83.640 196.605 83.930 196.650 ;
        RECT 85.500 196.605 85.790 196.650 ;
        RECT 88.280 196.605 88.570 196.650 ;
        RECT 91.440 196.790 91.760 196.850 ;
        RECT 92.145 196.790 92.435 196.835 ;
        RECT 91.440 196.650 92.435 196.790 ;
        RECT 91.440 196.590 91.760 196.650 ;
        RECT 92.145 196.605 92.435 196.650 ;
        RECT 92.835 196.790 93.125 196.835 ;
        RECT 94.660 196.790 94.980 196.850 ;
        RECT 92.835 196.650 94.980 196.790 ;
        RECT 92.835 196.605 93.125 196.650 ;
        RECT 94.660 196.590 94.980 196.650 ;
        RECT 104.435 196.790 104.725 196.835 ;
        RECT 107.555 196.790 107.845 196.835 ;
        RECT 109.445 196.790 109.735 196.835 ;
        RECT 104.435 196.650 109.735 196.790 ;
        RECT 104.435 196.605 104.725 196.650 ;
        RECT 107.555 196.605 107.845 196.650 ;
        RECT 109.445 196.605 109.735 196.650 ;
        RECT 64.300 196.450 64.620 196.510 ;
        RECT 56.800 196.310 64.620 196.450 ;
        RECT 53.275 196.265 53.565 196.310 ;
        RECT 54.180 196.250 54.500 196.310 ;
        RECT 64.300 196.250 64.620 196.310 ;
        RECT 73.055 196.450 73.345 196.495 ;
        RECT 74.420 196.450 74.740 196.510 ;
        RECT 73.055 196.310 74.740 196.450 ;
        RECT 73.055 196.265 73.345 196.310 ;
        RECT 74.420 196.250 74.740 196.310 ;
        RECT 75.355 196.450 75.645 196.495 ;
        RECT 76.260 196.450 76.580 196.510 ;
        RECT 75.355 196.310 76.580 196.450 ;
        RECT 75.355 196.265 75.645 196.310 ;
        RECT 76.260 196.250 76.580 196.310 ;
        RECT 78.575 196.450 78.865 196.495 ;
        RECT 79.480 196.450 79.800 196.510 ;
        RECT 78.575 196.310 79.800 196.450 ;
        RECT 78.575 196.265 78.865 196.310 ;
        RECT 79.480 196.250 79.800 196.310 ;
        RECT 82.715 196.450 83.005 196.495 ;
        RECT 99.720 196.450 100.040 196.510 ;
        RECT 82.715 196.310 100.040 196.450 ;
        RECT 82.715 196.265 83.005 196.310 ;
        RECT 99.720 196.250 100.040 196.310 ;
        RECT 101.560 196.250 101.880 196.510 ;
        RECT 26.970 195.630 113.450 196.110 ;
        RECT 31.640 195.230 31.960 195.490 ;
        RECT 51.420 195.430 51.740 195.490 ;
        RECT 51.895 195.430 52.185 195.475 ;
        RECT 43.690 195.290 49.810 195.430 ;
        RECT 39.460 194.890 39.780 195.150 ;
        RECT 32.575 194.750 32.865 194.795 ;
        RECT 33.020 194.750 33.340 194.810 ;
        RECT 32.575 194.610 33.340 194.750 ;
        RECT 32.575 194.565 32.865 194.610 ;
        RECT 33.020 194.550 33.340 194.610 ;
        RECT 33.480 194.750 33.800 194.810 ;
        RECT 40.380 194.750 40.700 194.810 ;
        RECT 43.155 194.750 43.445 194.795 ;
        RECT 43.690 194.750 43.830 195.290 ;
        RECT 44.025 195.090 44.315 195.135 ;
        RECT 45.915 195.090 46.205 195.135 ;
        RECT 49.035 195.090 49.325 195.135 ;
        RECT 44.025 194.950 49.325 195.090 ;
        RECT 49.670 195.090 49.810 195.290 ;
        RECT 51.420 195.290 52.185 195.430 ;
        RECT 51.420 195.230 51.740 195.290 ;
        RECT 51.895 195.245 52.185 195.290 ;
        RECT 52.800 195.230 53.120 195.490 ;
        RECT 62.920 195.230 63.240 195.490 ;
        RECT 64.315 195.430 64.605 195.475 ;
        RECT 65.220 195.430 65.540 195.490 ;
        RECT 64.315 195.290 65.540 195.430 ;
        RECT 64.315 195.245 64.605 195.290 ;
        RECT 65.220 195.230 65.540 195.290 ;
        RECT 66.140 195.230 66.460 195.490 ;
        RECT 69.360 195.430 69.680 195.490 ;
        RECT 67.150 195.290 68.670 195.430 ;
        RECT 49.670 194.950 52.570 195.090 ;
        RECT 44.025 194.905 44.315 194.950 ;
        RECT 45.915 194.905 46.205 194.950 ;
        RECT 49.035 194.905 49.325 194.950 ;
        RECT 33.480 194.610 36.930 194.750 ;
        RECT 33.480 194.550 33.800 194.610 ;
        RECT 36.790 194.470 36.930 194.610 ;
        RECT 40.380 194.610 41.530 194.750 ;
        RECT 40.380 194.550 40.700 194.610 ;
        RECT 28.880 194.210 29.200 194.470 ;
        RECT 35.335 194.410 35.625 194.455 ;
        RECT 35.780 194.410 36.100 194.470 ;
        RECT 35.335 194.270 36.100 194.410 ;
        RECT 35.335 194.225 35.625 194.270 ;
        RECT 35.780 194.210 36.100 194.270 ;
        RECT 36.700 194.210 37.020 194.470 ;
        RECT 38.095 194.410 38.385 194.455 ;
        RECT 38.095 194.270 40.610 194.410 ;
        RECT 38.095 194.225 38.385 194.270 ;
        RECT 37.160 193.530 37.480 193.790 ;
        RECT 38.080 193.730 38.400 193.790 ;
        RECT 39.015 193.730 39.305 193.775 ;
        RECT 38.080 193.590 39.305 193.730 ;
        RECT 40.470 193.730 40.610 194.270 ;
        RECT 40.840 194.210 41.160 194.470 ;
        RECT 41.390 194.455 41.530 194.610 ;
        RECT 43.155 194.610 43.830 194.750 ;
        RECT 43.155 194.565 43.445 194.610 ;
        RECT 41.315 194.225 41.605 194.455 ;
        RECT 41.760 194.210 42.080 194.470 ;
        RECT 52.430 194.455 52.570 194.950 ;
        RECT 52.890 194.750 53.030 195.230 ;
        RECT 53.225 195.090 53.515 195.135 ;
        RECT 55.115 195.090 55.405 195.135 ;
        RECT 58.235 195.090 58.525 195.135 ;
        RECT 67.150 195.090 67.290 195.290 ;
        RECT 53.225 194.950 58.525 195.090 ;
        RECT 53.225 194.905 53.515 194.950 ;
        RECT 55.115 194.905 55.405 194.950 ;
        RECT 58.235 194.905 58.525 194.950 ;
        RECT 65.310 194.950 67.290 195.090 ;
        RECT 53.735 194.750 54.025 194.795 ;
        RECT 52.890 194.610 54.025 194.750 ;
        RECT 53.735 194.565 54.025 194.610 ;
        RECT 57.400 194.750 57.720 194.810 ;
        RECT 65.310 194.750 65.450 194.950 ;
        RECT 67.995 194.905 68.285 195.135 ;
        RECT 68.530 195.090 68.670 195.290 ;
        RECT 69.360 195.290 80.630 195.430 ;
        RECT 69.360 195.230 69.680 195.290 ;
        RECT 71.200 195.090 71.520 195.150 ;
        RECT 72.135 195.090 72.425 195.135 ;
        RECT 68.530 194.950 72.425 195.090 ;
        RECT 57.400 194.610 65.450 194.750 ;
        RECT 68.070 194.750 68.210 194.905 ;
        RECT 71.200 194.890 71.520 194.950 ;
        RECT 72.135 194.905 72.425 194.950 ;
        RECT 74.995 195.090 75.285 195.135 ;
        RECT 78.115 195.090 78.405 195.135 ;
        RECT 80.005 195.090 80.295 195.135 ;
        RECT 74.995 194.950 80.295 195.090 ;
        RECT 80.490 195.090 80.630 195.290 ;
        RECT 83.160 195.230 83.480 195.490 ;
        RECT 84.080 195.430 84.400 195.490 ;
        RECT 89.615 195.430 89.905 195.475 ;
        RECT 84.080 195.290 89.905 195.430 ;
        RECT 84.080 195.230 84.400 195.290 ;
        RECT 89.615 195.245 89.905 195.290 ;
        RECT 90.060 195.430 90.380 195.490 ;
        RECT 100.640 195.430 100.960 195.490 ;
        RECT 90.060 195.290 100.960 195.430 ;
        RECT 90.060 195.230 90.380 195.290 ;
        RECT 83.620 195.090 83.940 195.150 ;
        RECT 90.980 195.090 91.300 195.150 ;
        RECT 80.490 194.950 83.940 195.090 ;
        RECT 74.995 194.905 75.285 194.950 ;
        RECT 78.115 194.905 78.405 194.950 ;
        RECT 80.005 194.905 80.295 194.950 ;
        RECT 83.620 194.890 83.940 194.950 ;
        RECT 84.630 194.950 91.300 195.090 ;
        RECT 84.630 194.810 84.770 194.950 ;
        RECT 90.980 194.890 91.300 194.950 ;
        RECT 93.755 195.090 94.045 195.135 ;
        RECT 95.120 195.090 95.440 195.150 ;
        RECT 93.755 194.950 95.440 195.090 ;
        RECT 93.755 194.905 94.045 194.950 ;
        RECT 95.120 194.890 95.440 194.950 ;
        RECT 68.440 194.750 68.760 194.810 ;
        RECT 70.755 194.750 71.045 194.795 ;
        RECT 73.040 194.750 73.360 194.810 ;
        RECT 68.070 194.610 69.130 194.750 ;
        RECT 57.400 194.550 57.720 194.610 ;
        RECT 68.440 194.550 68.760 194.610 ;
        RECT 42.695 194.410 42.985 194.455 ;
        RECT 43.620 194.410 43.910 194.455 ;
        RECT 45.455 194.410 45.745 194.455 ;
        RECT 49.035 194.410 49.325 194.455 ;
        RECT 42.695 194.270 43.370 194.410 ;
        RECT 42.695 194.225 42.985 194.270 ;
        RECT 43.230 194.070 43.370 194.270 ;
        RECT 43.620 194.270 49.325 194.410 ;
        RECT 43.620 194.225 43.910 194.270 ;
        RECT 45.455 194.225 45.745 194.270 ;
        RECT 49.035 194.225 49.325 194.270 ;
        RECT 44.060 194.070 44.380 194.130 ;
        RECT 43.230 193.930 44.380 194.070 ;
        RECT 44.060 193.870 44.380 193.930 ;
        RECT 44.520 193.870 44.840 194.130 ;
        RECT 50.115 194.115 50.405 194.430 ;
        RECT 52.355 194.225 52.645 194.455 ;
        RECT 52.820 194.410 53.110 194.455 ;
        RECT 54.655 194.410 54.945 194.455 ;
        RECT 58.235 194.410 58.525 194.455 ;
        RECT 52.820 194.270 58.525 194.410 ;
        RECT 52.820 194.225 53.110 194.270 ;
        RECT 54.655 194.225 54.945 194.270 ;
        RECT 58.235 194.225 58.525 194.270 ;
        RECT 46.815 194.070 47.465 194.115 ;
        RECT 50.115 194.070 50.705 194.115 ;
        RECT 50.960 194.070 51.280 194.130 ;
        RECT 46.815 193.930 51.280 194.070 ;
        RECT 52.430 194.070 52.570 194.225 ;
        RECT 53.720 194.070 54.040 194.130 ;
        RECT 52.430 193.930 54.040 194.070 ;
        RECT 46.815 193.885 47.465 193.930 ;
        RECT 50.415 193.885 50.705 193.930 ;
        RECT 50.960 193.870 51.280 193.930 ;
        RECT 53.720 193.870 54.040 193.930 ;
        RECT 56.015 194.070 56.665 194.115 ;
        RECT 56.940 194.070 57.260 194.130 ;
        RECT 59.315 194.115 59.605 194.430 ;
        RECT 63.840 194.210 64.160 194.470 ;
        RECT 64.760 194.410 65.080 194.470 ;
        RECT 65.235 194.410 65.525 194.455 ;
        RECT 64.760 194.270 65.525 194.410 ;
        RECT 64.760 194.210 65.080 194.270 ;
        RECT 65.235 194.225 65.525 194.270 ;
        RECT 67.075 194.225 67.365 194.455 ;
        RECT 59.315 194.070 59.905 194.115 ;
        RECT 56.015 193.930 59.905 194.070 ;
        RECT 56.015 193.885 56.665 193.930 ;
        RECT 56.940 193.870 57.260 193.930 ;
        RECT 59.615 193.885 59.905 193.930 ;
        RECT 43.140 193.730 43.460 193.790 ;
        RECT 40.470 193.590 43.460 193.730 ;
        RECT 38.080 193.530 38.400 193.590 ;
        RECT 39.015 193.545 39.305 193.590 ;
        RECT 43.140 193.530 43.460 193.590 ;
        RECT 58.780 193.730 59.100 193.790 ;
        RECT 61.095 193.730 61.385 193.775 ;
        RECT 58.780 193.590 61.385 193.730 ;
        RECT 58.780 193.530 59.100 193.590 ;
        RECT 61.095 193.545 61.385 193.590 ;
        RECT 65.220 193.730 65.540 193.790 ;
        RECT 67.150 193.730 67.290 194.225 ;
        RECT 67.995 193.885 68.285 194.115 ;
        RECT 68.990 194.070 69.130 194.610 ;
        RECT 70.755 194.610 73.360 194.750 ;
        RECT 70.755 194.565 71.045 194.610 ;
        RECT 73.040 194.550 73.360 194.610 ;
        RECT 79.480 194.550 79.800 194.810 ;
        RECT 80.875 194.750 81.165 194.795 ;
        RECT 84.540 194.750 84.860 194.810 ;
        RECT 80.875 194.610 84.860 194.750 ;
        RECT 80.875 194.565 81.165 194.610 ;
        RECT 84.540 194.550 84.860 194.610 ;
        RECT 85.920 194.550 86.240 194.810 ;
        RECT 86.840 194.750 87.160 194.810 ;
        RECT 91.915 194.750 92.205 194.795 ;
        RECT 86.840 194.610 92.205 194.750 ;
        RECT 86.840 194.550 87.160 194.610 ;
        RECT 91.915 194.565 92.205 194.610 ;
        RECT 92.375 194.565 92.665 194.795 ;
        RECT 95.670 194.750 95.810 195.290 ;
        RECT 100.640 195.230 100.960 195.290 ;
        RECT 101.100 195.430 101.420 195.490 ;
        RECT 101.575 195.430 101.865 195.475 ;
        RECT 101.100 195.290 101.865 195.430 ;
        RECT 101.100 195.230 101.420 195.290 ;
        RECT 101.575 195.245 101.865 195.290 ;
        RECT 111.220 195.230 111.540 195.490 ;
        RECT 97.880 195.090 98.200 195.150 ;
        RECT 105.240 195.090 105.560 195.150 ;
        RECT 97.880 194.950 105.560 195.090 ;
        RECT 97.880 194.890 98.200 194.950 ;
        RECT 105.240 194.890 105.560 194.950 ;
        RECT 95.670 194.610 99.490 194.750 ;
        RECT 70.295 194.410 70.585 194.455 ;
        RECT 72.120 194.410 72.440 194.470 ;
        RECT 70.295 194.270 72.440 194.410 ;
        RECT 70.295 194.225 70.585 194.270 ;
        RECT 72.120 194.210 72.440 194.270 ;
        RECT 73.915 194.115 74.205 194.430 ;
        RECT 74.995 194.410 75.285 194.455 ;
        RECT 78.575 194.410 78.865 194.455 ;
        RECT 80.410 194.410 80.700 194.455 ;
        RECT 74.995 194.270 80.700 194.410 ;
        RECT 74.995 194.225 75.285 194.270 ;
        RECT 78.575 194.225 78.865 194.270 ;
        RECT 80.410 194.225 80.700 194.270 ;
        RECT 81.795 194.225 82.085 194.455 ;
        RECT 82.255 194.410 82.545 194.455 ;
        RECT 83.620 194.410 83.940 194.470 ;
        RECT 82.255 194.270 83.940 194.410 ;
        RECT 82.255 194.225 82.545 194.270 ;
        RECT 73.615 194.070 74.205 194.115 ;
        RECT 76.855 194.070 77.505 194.115 ;
        RECT 81.870 194.070 82.010 194.225 ;
        RECT 83.620 194.210 83.940 194.270 ;
        RECT 84.080 194.410 84.400 194.470 ;
        RECT 85.475 194.410 85.765 194.455 ;
        RECT 87.760 194.410 88.080 194.470 ;
        RECT 88.235 194.410 88.525 194.455 ;
        RECT 84.080 194.270 87.530 194.410 ;
        RECT 84.080 194.210 84.400 194.270 ;
        RECT 85.475 194.225 85.765 194.270 ;
        RECT 68.990 193.930 72.810 194.070 ;
        RECT 65.220 193.590 67.290 193.730 ;
        RECT 68.070 193.730 68.210 193.885 ;
        RECT 70.280 193.730 70.600 193.790 ;
        RECT 68.070 193.590 70.600 193.730 ;
        RECT 65.220 193.530 65.540 193.590 ;
        RECT 70.280 193.530 70.600 193.590 ;
        RECT 71.675 193.730 71.965 193.775 ;
        RECT 72.120 193.730 72.440 193.790 ;
        RECT 71.675 193.590 72.440 193.730 ;
        RECT 72.670 193.730 72.810 193.930 ;
        RECT 73.615 193.930 82.010 194.070 ;
        RECT 87.390 194.070 87.530 194.270 ;
        RECT 87.760 194.270 88.525 194.410 ;
        RECT 87.760 194.210 88.080 194.270 ;
        RECT 88.235 194.225 88.525 194.270 ;
        RECT 88.680 194.210 89.000 194.470 ;
        RECT 91.440 194.410 91.760 194.470 ;
        RECT 89.230 194.270 91.760 194.410 ;
        RECT 89.230 194.070 89.370 194.270 ;
        RECT 91.440 194.210 91.760 194.270 ;
        RECT 92.450 194.070 92.590 194.565 ;
        RECT 94.200 194.410 94.520 194.470 ;
        RECT 95.135 194.410 95.425 194.455 ;
        RECT 94.200 194.270 95.425 194.410 ;
        RECT 94.200 194.210 94.520 194.270 ;
        RECT 95.135 194.225 95.425 194.270 ;
        RECT 95.580 194.210 95.900 194.470 ;
        RECT 96.130 194.455 96.270 194.610 ;
        RECT 96.055 194.225 96.345 194.455 ;
        RECT 96.500 194.410 96.820 194.470 ;
        RECT 99.350 194.455 99.490 194.610 ;
        RECT 99.720 194.550 100.040 194.810 ;
        RECT 100.195 194.565 100.485 194.795 ;
        RECT 104.335 194.750 104.625 194.795 ;
        RECT 102.570 194.610 104.625 194.750 ;
        RECT 96.975 194.410 97.265 194.455 ;
        RECT 96.500 194.270 97.265 194.410 ;
        RECT 96.500 194.210 96.820 194.270 ;
        RECT 96.975 194.225 97.265 194.270 ;
        RECT 99.275 194.225 99.565 194.455 ;
        RECT 100.270 194.410 100.410 194.565 ;
        RECT 102.570 194.470 102.710 194.610 ;
        RECT 104.335 194.565 104.625 194.610 ;
        RECT 104.780 194.750 105.100 194.810 ;
        RECT 104.780 194.610 109.150 194.750 ;
        RECT 104.780 194.550 105.100 194.610 ;
        RECT 102.480 194.410 102.800 194.470 ;
        RECT 99.810 194.270 102.800 194.410 ;
        RECT 98.800 194.070 99.120 194.130 ;
        RECT 99.810 194.070 99.950 194.270 ;
        RECT 102.480 194.210 102.800 194.270 ;
        RECT 103.875 194.225 104.165 194.455 ;
        RECT 106.160 194.410 106.480 194.470 ;
        RECT 107.095 194.410 107.385 194.455 ;
        RECT 106.160 194.270 107.385 194.410 ;
        RECT 87.390 193.930 89.370 194.070 ;
        RECT 91.530 193.930 99.950 194.070 ;
        RECT 100.180 194.070 100.500 194.130 ;
        RECT 103.950 194.070 104.090 194.225 ;
        RECT 106.160 194.210 106.480 194.270 ;
        RECT 107.095 194.225 107.385 194.270 ;
        RECT 107.555 194.225 107.845 194.455 ;
        RECT 107.630 194.070 107.770 194.225 ;
        RECT 108.000 194.210 108.320 194.470 ;
        RECT 109.010 194.455 109.150 194.610 ;
        RECT 108.935 194.225 109.225 194.455 ;
        RECT 109.380 194.410 109.700 194.470 ;
        RECT 110.315 194.410 110.605 194.455 ;
        RECT 109.380 194.270 110.605 194.410 ;
        RECT 109.380 194.210 109.700 194.270 ;
        RECT 110.315 194.225 110.605 194.270 ;
        RECT 111.680 194.210 112.000 194.470 ;
        RECT 100.180 193.930 104.090 194.070 ;
        RECT 107.170 193.930 107.770 194.070 ;
        RECT 73.615 193.885 73.905 193.930 ;
        RECT 76.855 193.885 77.505 193.930 ;
        RECT 91.530 193.790 91.670 193.930 ;
        RECT 98.800 193.870 99.120 193.930 ;
        RECT 100.180 193.870 100.500 193.930 ;
        RECT 107.170 193.790 107.310 193.930 ;
        RECT 74.880 193.730 75.200 193.790 ;
        RECT 75.800 193.730 76.120 193.790 ;
        RECT 72.670 193.590 76.120 193.730 ;
        RECT 71.675 193.545 71.965 193.590 ;
        RECT 72.120 193.530 72.440 193.590 ;
        RECT 74.880 193.530 75.200 193.590 ;
        RECT 75.800 193.530 76.120 193.590 ;
        RECT 80.400 193.730 80.720 193.790 ;
        RECT 85.015 193.730 85.305 193.775 ;
        RECT 80.400 193.590 85.305 193.730 ;
        RECT 80.400 193.530 80.720 193.590 ;
        RECT 85.015 193.545 85.305 193.590 ;
        RECT 85.920 193.730 86.240 193.790 ;
        RECT 91.440 193.730 91.760 193.790 ;
        RECT 85.920 193.590 91.760 193.730 ;
        RECT 85.920 193.530 86.240 193.590 ;
        RECT 91.440 193.530 91.760 193.590 ;
        RECT 96.960 193.730 97.280 193.790 ;
        RECT 97.435 193.730 97.725 193.775 ;
        RECT 96.960 193.590 97.725 193.730 ;
        RECT 96.960 193.530 97.280 193.590 ;
        RECT 97.435 193.545 97.725 193.590 ;
        RECT 99.720 193.730 100.040 193.790 ;
        RECT 103.415 193.730 103.705 193.775 ;
        RECT 99.720 193.590 103.705 193.730 ;
        RECT 99.720 193.530 100.040 193.590 ;
        RECT 103.415 193.545 103.705 193.590 ;
        RECT 105.240 193.730 105.560 193.790 ;
        RECT 105.715 193.730 106.005 193.775 ;
        RECT 105.240 193.590 106.005 193.730 ;
        RECT 105.240 193.530 105.560 193.590 ;
        RECT 105.715 193.545 106.005 193.590 ;
        RECT 107.080 193.530 107.400 193.790 ;
        RECT 108.920 193.730 109.240 193.790 ;
        RECT 109.395 193.730 109.685 193.775 ;
        RECT 108.920 193.590 109.685 193.730 ;
        RECT 108.920 193.530 109.240 193.590 ;
        RECT 109.395 193.545 109.685 193.590 ;
        RECT 26.970 192.910 113.450 193.390 ;
        RECT 40.840 192.710 41.160 192.770 ;
        RECT 42.220 192.710 42.540 192.770 ;
        RECT 40.840 192.570 42.540 192.710 ;
        RECT 40.840 192.510 41.160 192.570 ;
        RECT 42.220 192.510 42.540 192.570 ;
        RECT 43.140 192.710 43.460 192.770 ;
        RECT 43.615 192.710 43.905 192.755 ;
        RECT 43.140 192.570 43.905 192.710 ;
        RECT 43.140 192.510 43.460 192.570 ;
        RECT 43.615 192.525 43.905 192.570 ;
        RECT 51.420 192.510 51.740 192.770 ;
        RECT 52.340 192.510 52.660 192.770 ;
        RECT 54.180 192.510 54.500 192.770 ;
        RECT 54.655 192.710 54.945 192.755 ;
        RECT 55.100 192.710 55.420 192.770 ;
        RECT 67.060 192.755 67.380 192.770 ;
        RECT 54.655 192.570 55.420 192.710 ;
        RECT 54.655 192.525 54.945 192.570 ;
        RECT 55.100 192.510 55.420 192.570 ;
        RECT 57.030 192.570 60.390 192.710 ;
        RECT 30.720 192.370 31.040 192.430 ;
        RECT 33.430 192.370 33.720 192.415 ;
        RECT 36.690 192.370 36.980 192.415 ;
        RECT 30.720 192.230 36.980 192.370 ;
        RECT 30.720 192.170 31.040 192.230 ;
        RECT 33.430 192.185 33.720 192.230 ;
        RECT 36.690 192.185 36.980 192.230 ;
        RECT 37.610 192.370 37.900 192.415 ;
        RECT 39.470 192.370 39.760 192.415 ;
        RECT 46.820 192.370 47.140 192.430 ;
        RECT 50.040 192.370 50.360 192.430 ;
        RECT 37.610 192.230 39.760 192.370 ;
        RECT 37.610 192.185 37.900 192.230 ;
        RECT 39.470 192.185 39.760 192.230 ;
        RECT 40.930 192.230 47.140 192.370 ;
        RECT 27.500 192.030 27.820 192.090 ;
        RECT 28.895 192.030 29.185 192.075 ;
        RECT 27.500 191.890 29.185 192.030 ;
        RECT 27.500 191.830 27.820 191.890 ;
        RECT 28.895 191.845 29.185 191.890 ;
        RECT 35.290 192.030 35.580 192.075 ;
        RECT 37.610 192.030 37.825 192.185 ;
        RECT 35.290 191.890 37.825 192.030 ;
        RECT 35.290 191.845 35.580 191.890 ;
        RECT 38.080 191.830 38.400 192.090 ;
        RECT 38.540 191.830 38.860 192.090 ;
        RECT 40.930 192.075 41.070 192.230 ;
        RECT 46.820 192.170 47.140 192.230 ;
        RECT 49.210 192.230 50.360 192.370 ;
        RECT 40.855 191.845 41.145 192.075 ;
        RECT 42.220 191.830 42.540 192.090 ;
        RECT 49.210 192.075 49.350 192.230 ;
        RECT 50.040 192.170 50.360 192.230 ;
        RECT 50.975 192.370 51.265 192.415 ;
        RECT 56.480 192.370 56.800 192.430 ;
        RECT 50.975 192.230 56.800 192.370 ;
        RECT 50.975 192.185 51.265 192.230 ;
        RECT 56.480 192.170 56.800 192.230 ;
        RECT 45.455 191.845 45.745 192.075 ;
        RECT 49.135 191.845 49.425 192.075 ;
        RECT 49.595 192.030 49.885 192.075 ;
        RECT 57.030 192.030 57.170 192.570 ;
        RECT 60.250 192.370 60.390 192.570 ;
        RECT 66.995 192.525 67.380 192.755 ;
        RECT 70.740 192.710 71.060 192.770 ;
        RECT 96.960 192.710 97.280 192.770 ;
        RECT 108.920 192.710 109.240 192.770 ;
        RECT 67.060 192.510 67.380 192.525 ;
        RECT 67.610 192.570 71.060 192.710 ;
        RECT 60.615 192.370 61.265 192.415 ;
        RECT 64.215 192.370 64.505 192.415 ;
        RECT 60.250 192.230 64.505 192.370 ;
        RECT 60.615 192.185 61.265 192.230 ;
        RECT 63.915 192.185 64.505 192.230 ;
        RECT 65.220 192.370 65.540 192.430 ;
        RECT 67.610 192.370 67.750 192.570 ;
        RECT 70.740 192.510 71.060 192.570 ;
        RECT 78.190 192.570 97.280 192.710 ;
        RECT 65.220 192.230 67.750 192.370 ;
        RECT 67.995 192.370 68.285 192.415 ;
        RECT 68.900 192.370 69.220 192.430 ;
        RECT 67.995 192.230 69.220 192.370 ;
        RECT 49.595 191.890 57.170 192.030 ;
        RECT 57.420 192.030 57.710 192.075 ;
        RECT 59.255 192.030 59.545 192.075 ;
        RECT 62.835 192.030 63.125 192.075 ;
        RECT 57.420 191.890 63.125 192.030 ;
        RECT 49.595 191.845 49.885 191.890 ;
        RECT 57.420 191.845 57.710 191.890 ;
        RECT 59.255 191.845 59.545 191.890 ;
        RECT 62.835 191.845 63.125 191.890 ;
        RECT 63.915 191.870 64.205 192.185 ;
        RECT 65.220 192.170 65.540 192.230 ;
        RECT 67.995 192.185 68.285 192.230 ;
        RECT 67.520 192.030 67.840 192.090 ;
        RECT 68.070 192.030 68.210 192.185 ;
        RECT 68.900 192.170 69.220 192.230 ;
        RECT 69.360 192.370 69.680 192.430 ;
        RECT 69.835 192.370 70.125 192.415 ;
        RECT 69.360 192.230 70.125 192.370 ;
        RECT 69.360 192.170 69.680 192.230 ;
        RECT 69.835 192.185 70.125 192.230 ;
        RECT 67.520 191.890 68.210 192.030 ;
        RECT 68.455 192.030 68.745 192.075 ;
        RECT 68.455 191.980 70.740 192.030 ;
        RECT 71.200 191.980 71.520 192.090 ;
        RECT 68.455 191.890 71.520 191.980 ;
        RECT 38.170 191.690 38.310 191.830 ;
        RECT 40.395 191.690 40.685 191.735 ;
        RECT 38.170 191.550 40.685 191.690 ;
        RECT 40.395 191.505 40.685 191.550 ;
        RECT 41.300 191.690 41.620 191.750 ;
        RECT 45.530 191.690 45.670 191.845 ;
        RECT 67.520 191.830 67.840 191.890 ;
        RECT 68.455 191.845 68.745 191.890 ;
        RECT 70.600 191.840 71.520 191.890 ;
        RECT 71.200 191.830 71.520 191.840 ;
        RECT 71.660 192.050 71.980 192.090 ;
        RECT 71.660 192.030 72.350 192.050 ;
        RECT 72.580 192.030 72.900 192.090 ;
        RECT 71.660 191.910 72.900 192.030 ;
        RECT 71.660 191.830 71.980 191.910 ;
        RECT 72.210 191.890 72.900 191.910 ;
        RECT 72.580 191.830 72.900 191.890 ;
        RECT 73.040 191.830 73.360 192.090 ;
        RECT 73.500 191.830 73.820 192.090 ;
        RECT 78.190 192.075 78.330 192.570 ;
        RECT 96.960 192.510 97.280 192.570 ;
        RECT 97.510 192.570 109.240 192.710 ;
        RECT 87.760 192.415 88.080 192.430 ;
        RECT 84.490 192.370 84.780 192.415 ;
        RECT 87.750 192.370 88.080 192.415 ;
        RECT 84.490 192.230 88.080 192.370 ;
        RECT 84.490 192.185 84.780 192.230 ;
        RECT 87.750 192.185 88.080 192.230 ;
        RECT 87.760 192.170 88.080 192.185 ;
        RECT 88.670 192.370 88.960 192.415 ;
        RECT 90.530 192.370 90.820 192.415 ;
        RECT 97.510 192.370 97.650 192.570 ;
        RECT 108.920 192.510 109.240 192.570 ;
        RECT 88.670 192.230 90.820 192.370 ;
        RECT 88.670 192.185 88.960 192.230 ;
        RECT 90.530 192.185 90.820 192.230 ;
        RECT 91.070 192.230 97.650 192.370 ;
        RECT 78.115 191.845 78.405 192.075 ;
        RECT 79.035 192.030 79.325 192.075 ;
        RECT 85.460 192.030 85.780 192.090 ;
        RECT 79.035 191.890 85.780 192.030 ;
        RECT 79.035 191.845 79.325 191.890 ;
        RECT 85.460 191.830 85.780 191.890 ;
        RECT 86.350 192.030 86.640 192.075 ;
        RECT 88.670 192.030 88.885 192.185 ;
        RECT 86.350 191.890 88.885 192.030 ;
        RECT 89.615 192.030 89.905 192.075 ;
        RECT 91.070 192.030 91.210 192.230 ;
        RECT 89.615 191.890 91.210 192.030 ;
        RECT 86.350 191.845 86.640 191.890 ;
        RECT 89.615 191.845 89.905 191.890 ;
        RECT 91.440 191.830 91.760 192.090 ;
        RECT 94.675 192.030 94.965 192.075 ;
        RECT 91.990 191.890 94.965 192.030 ;
        RECT 97.895 191.965 98.185 192.195 ;
        RECT 103.860 192.170 104.180 192.430 ;
        RECT 104.320 192.370 104.640 192.430 ;
        RECT 106.155 192.370 106.805 192.415 ;
        RECT 109.755 192.370 110.045 192.415 ;
        RECT 104.320 192.230 110.045 192.370 ;
        RECT 104.320 192.170 104.640 192.230 ;
        RECT 106.155 192.185 106.805 192.230 ;
        RECT 109.455 192.185 110.045 192.230 ;
        RECT 98.800 192.030 99.120 192.090 ;
        RECT 99.735 192.030 100.025 192.075 ;
        RECT 41.300 191.550 45.670 191.690 ;
        RECT 41.300 191.490 41.620 191.550 ;
        RECT 45.915 191.505 46.205 191.735 ;
        RECT 46.820 191.690 47.140 191.750 ;
        RECT 55.115 191.690 55.405 191.735 ;
        RECT 56.480 191.690 56.800 191.750 ;
        RECT 46.820 191.550 56.800 191.690 ;
        RECT 35.290 191.350 35.580 191.395 ;
        RECT 38.070 191.350 38.360 191.395 ;
        RECT 39.930 191.350 40.220 191.395 ;
        RECT 35.290 191.210 40.220 191.350 ;
        RECT 35.290 191.165 35.580 191.210 ;
        RECT 38.070 191.165 38.360 191.210 ;
        RECT 39.930 191.165 40.220 191.210 ;
        RECT 29.815 191.010 30.105 191.055 ;
        RECT 30.260 191.010 30.580 191.070 ;
        RECT 29.815 190.870 30.580 191.010 ;
        RECT 29.815 190.825 30.105 190.870 ;
        RECT 30.260 190.810 30.580 190.870 ;
        RECT 31.425 191.010 31.715 191.055 ;
        RECT 33.020 191.010 33.340 191.070 ;
        RECT 41.390 191.010 41.530 191.490 ;
        RECT 41.775 191.350 42.065 191.395 ;
        RECT 44.520 191.350 44.840 191.410 ;
        RECT 41.775 191.210 44.840 191.350 ;
        RECT 45.990 191.350 46.130 191.505 ;
        RECT 46.820 191.490 47.140 191.550 ;
        RECT 55.115 191.505 55.405 191.550 ;
        RECT 56.480 191.490 56.800 191.550 ;
        RECT 56.955 191.505 57.245 191.735 ;
        RECT 52.340 191.350 52.660 191.410 ;
        RECT 45.990 191.210 52.660 191.350 ;
        RECT 41.775 191.165 42.065 191.210 ;
        RECT 44.520 191.150 44.840 191.210 ;
        RECT 52.340 191.150 52.660 191.210 ;
        RECT 53.720 191.350 54.040 191.410 ;
        RECT 57.030 191.350 57.170 191.505 ;
        RECT 58.320 191.490 58.640 191.750 ;
        RECT 61.540 191.690 61.860 191.750 ;
        RECT 72.135 191.690 72.425 191.735 ;
        RECT 74.880 191.690 75.200 191.750 ;
        RECT 61.540 191.550 70.740 191.690 ;
        RECT 61.540 191.490 61.860 191.550 ;
        RECT 53.720 191.210 57.170 191.350 ;
        RECT 57.825 191.350 58.115 191.395 ;
        RECT 59.715 191.350 60.005 191.395 ;
        RECT 62.835 191.350 63.125 191.395 ;
        RECT 57.825 191.210 63.125 191.350 ;
        RECT 53.720 191.150 54.040 191.210 ;
        RECT 57.825 191.165 58.115 191.210 ;
        RECT 59.715 191.165 60.005 191.210 ;
        RECT 62.835 191.165 63.125 191.210 ;
        RECT 63.380 191.350 63.700 191.410 ;
        RECT 65.695 191.350 65.985 191.395 ;
        RECT 63.380 191.210 65.985 191.350 ;
        RECT 70.600 191.350 70.740 191.550 ;
        RECT 72.135 191.550 75.200 191.690 ;
        RECT 72.135 191.505 72.425 191.550 ;
        RECT 74.880 191.490 75.200 191.550 ;
        RECT 81.795 191.690 82.085 191.735 ;
        RECT 91.990 191.690 92.130 191.890 ;
        RECT 94.675 191.845 94.965 191.890 ;
        RECT 97.970 191.750 98.110 191.965 ;
        RECT 98.800 191.890 100.025 192.030 ;
        RECT 98.800 191.830 99.120 191.890 ;
        RECT 99.735 191.845 100.025 191.890 ;
        RECT 101.560 191.830 101.880 192.090 ;
        RECT 102.960 192.030 103.250 192.075 ;
        RECT 104.795 192.030 105.085 192.075 ;
        RECT 108.375 192.030 108.665 192.075 ;
        RECT 102.960 191.890 108.665 192.030 ;
        RECT 102.960 191.845 103.250 191.890 ;
        RECT 104.795 191.845 105.085 191.890 ;
        RECT 108.375 191.845 108.665 191.890 ;
        RECT 109.455 191.870 109.745 192.185 ;
        RECT 81.795 191.550 92.130 191.690 ;
        RECT 92.360 191.690 92.680 191.750 ;
        RECT 93.295 191.690 93.585 191.735 ;
        RECT 92.360 191.550 93.585 191.690 ;
        RECT 81.795 191.505 82.085 191.550 ;
        RECT 92.360 191.490 92.680 191.550 ;
        RECT 93.295 191.505 93.585 191.550 ;
        RECT 94.215 191.505 94.505 191.735 ;
        RECT 97.420 191.690 97.740 191.750 ;
        RECT 96.590 191.550 97.740 191.690 ;
        RECT 86.350 191.350 86.640 191.395 ;
        RECT 89.130 191.350 89.420 191.395 ;
        RECT 90.990 191.350 91.280 191.395 ;
        RECT 70.600 191.210 75.110 191.350 ;
        RECT 63.380 191.150 63.700 191.210 ;
        RECT 65.695 191.165 65.985 191.210 ;
        RECT 31.425 190.870 41.530 191.010 ;
        RECT 43.155 191.010 43.445 191.055 ;
        RECT 45.440 191.010 45.760 191.070 ;
        RECT 43.155 190.870 45.760 191.010 ;
        RECT 31.425 190.825 31.715 190.870 ;
        RECT 33.020 190.810 33.340 190.870 ;
        RECT 43.155 190.825 43.445 190.870 ;
        RECT 45.440 190.810 45.760 190.870 ;
        RECT 51.420 191.010 51.740 191.070 ;
        RECT 55.100 191.010 55.420 191.070 ;
        RECT 51.420 190.870 55.420 191.010 ;
        RECT 51.420 190.810 51.740 190.870 ;
        RECT 55.100 190.810 55.420 190.870 ;
        RECT 61.080 191.010 61.400 191.070 ;
        RECT 66.155 191.010 66.445 191.055 ;
        RECT 61.080 190.870 66.445 191.010 ;
        RECT 61.080 190.810 61.400 190.870 ;
        RECT 66.155 190.825 66.445 190.870 ;
        RECT 67.075 191.010 67.365 191.055 ;
        RECT 67.980 191.010 68.300 191.070 ;
        RECT 67.075 190.870 68.300 191.010 ;
        RECT 67.075 190.825 67.365 190.870 ;
        RECT 67.980 190.810 68.300 190.870 ;
        RECT 68.440 191.010 68.760 191.070 ;
        RECT 74.970 191.055 75.110 191.210 ;
        RECT 86.350 191.210 91.280 191.350 ;
        RECT 86.350 191.165 86.640 191.210 ;
        RECT 89.130 191.165 89.420 191.210 ;
        RECT 90.990 191.165 91.280 191.210 ;
        RECT 91.900 191.350 92.220 191.410 ;
        RECT 94.290 191.350 94.430 191.505 ;
        RECT 96.590 191.395 96.730 191.550 ;
        RECT 97.420 191.490 97.740 191.550 ;
        RECT 97.880 191.490 98.200 191.750 ;
        RECT 98.340 191.690 98.660 191.750 ;
        RECT 102.495 191.690 102.785 191.735 ;
        RECT 98.340 191.550 102.785 191.690 ;
        RECT 98.340 191.490 98.660 191.550 ;
        RECT 102.495 191.505 102.785 191.550 ;
        RECT 91.900 191.210 94.430 191.350 ;
        RECT 91.900 191.150 92.220 191.210 ;
        RECT 96.515 191.165 96.805 191.395 ;
        RECT 98.815 191.350 99.105 191.395 ;
        RECT 99.260 191.350 99.580 191.410 ;
        RECT 98.815 191.210 99.580 191.350 ;
        RECT 98.815 191.165 99.105 191.210 ;
        RECT 99.260 191.150 99.580 191.210 ;
        RECT 103.365 191.350 103.655 191.395 ;
        RECT 105.255 191.350 105.545 191.395 ;
        RECT 108.375 191.350 108.665 191.395 ;
        RECT 103.365 191.210 108.665 191.350 ;
        RECT 103.365 191.165 103.655 191.210 ;
        RECT 105.255 191.165 105.545 191.210 ;
        RECT 108.375 191.165 108.665 191.210 ;
        RECT 71.215 191.010 71.505 191.055 ;
        RECT 68.440 190.870 71.505 191.010 ;
        RECT 68.440 190.810 68.760 190.870 ;
        RECT 71.215 190.825 71.505 190.870 ;
        RECT 74.895 190.825 75.185 191.055 ;
        RECT 80.400 191.010 80.720 191.070 ;
        RECT 82.485 191.010 82.775 191.055 ;
        RECT 80.400 190.870 82.775 191.010 ;
        RECT 80.400 190.810 80.720 190.870 ;
        RECT 82.485 190.825 82.775 190.870 ;
        RECT 86.840 191.010 87.160 191.070 ;
        RECT 90.060 191.010 90.380 191.070 ;
        RECT 86.840 190.870 90.380 191.010 ;
        RECT 86.840 190.810 87.160 190.870 ;
        RECT 90.060 190.810 90.380 190.870 ;
        RECT 90.520 191.010 90.840 191.070 ;
        RECT 96.975 191.010 97.265 191.055 ;
        RECT 90.520 190.870 97.265 191.010 ;
        RECT 90.520 190.810 90.840 190.870 ;
        RECT 96.975 190.825 97.265 190.870 ;
        RECT 97.420 191.010 97.740 191.070 ;
        RECT 101.115 191.010 101.405 191.055 ;
        RECT 97.420 190.870 101.405 191.010 ;
        RECT 97.420 190.810 97.740 190.870 ;
        RECT 101.115 190.825 101.405 190.870 ;
        RECT 109.840 191.010 110.160 191.070 ;
        RECT 111.235 191.010 111.525 191.055 ;
        RECT 109.840 190.870 111.525 191.010 ;
        RECT 109.840 190.810 110.160 190.870 ;
        RECT 111.235 190.825 111.525 190.870 ;
        RECT 26.970 190.190 113.450 190.670 ;
        RECT 35.335 189.990 35.625 190.035 ;
        RECT 36.240 189.990 36.560 190.050 ;
        RECT 35.335 189.850 36.560 189.990 ;
        RECT 35.335 189.805 35.625 189.850 ;
        RECT 36.240 189.790 36.560 189.850 ;
        RECT 36.700 189.990 37.020 190.050 ;
        RECT 39.460 189.990 39.780 190.050 ;
        RECT 41.300 189.990 41.620 190.050 ;
        RECT 51.880 189.990 52.200 190.050 ;
        RECT 56.035 189.990 56.325 190.035 ;
        RECT 36.700 189.850 38.310 189.990 ;
        RECT 36.700 189.790 37.020 189.850 ;
        RECT 29.340 189.110 29.660 189.370 ;
        RECT 32.560 189.110 32.880 189.370 ;
        RECT 33.020 189.110 33.340 189.370 ;
        RECT 29.430 188.970 29.570 189.110 ;
        RECT 29.815 188.970 30.105 189.015 ;
        RECT 29.430 188.830 30.105 188.970 ;
        RECT 29.815 188.785 30.105 188.830 ;
        RECT 30.275 188.970 30.565 189.015 ;
        RECT 31.640 188.970 31.960 189.030 ;
        RECT 30.275 188.830 31.960 188.970 ;
        RECT 30.275 188.785 30.565 188.830 ;
        RECT 31.640 188.770 31.960 188.830 ;
        RECT 32.100 188.970 32.420 189.030 ;
        RECT 33.495 188.970 33.785 189.015 ;
        RECT 32.100 188.830 33.785 188.970 ;
        RECT 32.100 188.770 32.420 188.830 ;
        RECT 33.495 188.785 33.785 188.830 ;
        RECT 36.700 188.770 37.020 189.030 ;
        RECT 38.170 189.015 38.310 189.850 ;
        RECT 39.460 189.850 51.650 189.990 ;
        RECT 39.460 189.790 39.780 189.850 ;
        RECT 41.300 189.790 41.620 189.850 ;
        RECT 38.095 188.970 38.385 189.015 ;
        RECT 38.540 188.970 38.860 189.030 ;
        RECT 39.550 189.015 39.690 189.790 ;
        RECT 42.695 189.650 42.985 189.695 ;
        RECT 44.060 189.650 44.380 189.710 ;
        RECT 42.695 189.510 44.380 189.650 ;
        RECT 42.695 189.465 42.985 189.510 ;
        RECT 44.060 189.450 44.380 189.510 ;
        RECT 46.015 189.650 46.305 189.695 ;
        RECT 49.135 189.650 49.425 189.695 ;
        RECT 51.025 189.650 51.315 189.695 ;
        RECT 46.015 189.510 51.315 189.650 ;
        RECT 46.015 189.465 46.305 189.510 ;
        RECT 49.135 189.465 49.425 189.510 ;
        RECT 51.025 189.465 51.315 189.510 ;
        RECT 48.660 189.310 48.980 189.370 ;
        RECT 40.930 189.170 48.980 189.310 ;
        RECT 40.930 189.030 41.070 189.170 ;
        RECT 48.660 189.110 48.980 189.170 ;
        RECT 50.500 189.110 50.820 189.370 ;
        RECT 51.510 189.310 51.650 189.850 ;
        RECT 51.880 189.850 56.325 189.990 ;
        RECT 51.880 189.790 52.200 189.850 ;
        RECT 56.035 189.805 56.325 189.850 ;
        RECT 67.535 189.990 67.825 190.035 ;
        RECT 82.715 189.990 83.005 190.035 ;
        RECT 89.140 189.990 89.460 190.050 ;
        RECT 67.535 189.850 74.650 189.990 ;
        RECT 67.535 189.805 67.825 189.850 ;
        RECT 64.760 189.650 65.080 189.710 ;
        RECT 69.820 189.650 70.140 189.710 ;
        RECT 73.040 189.650 73.360 189.710 ;
        RECT 64.760 189.510 73.360 189.650 ;
        RECT 64.760 189.450 65.080 189.510 ;
        RECT 69.820 189.450 70.140 189.510 ;
        RECT 56.020 189.310 56.340 189.370 ;
        RECT 51.510 189.170 52.570 189.310 ;
        RECT 38.095 188.830 38.860 188.970 ;
        RECT 38.095 188.785 38.385 188.830 ;
        RECT 38.540 188.770 38.860 188.830 ;
        RECT 39.475 188.785 39.765 189.015 ;
        RECT 40.395 188.785 40.685 189.015 ;
        RECT 29.355 188.630 29.645 188.675 ;
        RECT 40.470 188.630 40.610 188.785 ;
        RECT 40.840 188.770 41.160 189.030 ;
        RECT 41.315 188.950 41.605 189.015 ;
        RECT 42.680 188.950 43.000 189.030 ;
        RECT 44.980 188.990 45.300 189.030 ;
        RECT 52.430 189.015 52.570 189.170 ;
        RECT 53.350 189.170 56.340 189.310 ;
        RECT 41.315 188.810 43.000 188.950 ;
        RECT 41.315 188.785 41.605 188.810 ;
        RECT 42.680 188.770 43.000 188.810 ;
        RECT 44.935 188.770 45.300 188.990 ;
        RECT 46.015 188.970 46.305 189.015 ;
        RECT 49.595 188.970 49.885 189.015 ;
        RECT 51.430 188.970 51.720 189.015 ;
        RECT 46.015 188.830 51.720 188.970 ;
        RECT 46.015 188.785 46.305 188.830 ;
        RECT 49.595 188.785 49.885 188.830 ;
        RECT 51.430 188.785 51.720 188.830 ;
        RECT 51.895 188.785 52.185 189.015 ;
        RECT 52.355 188.785 52.645 189.015 ;
        RECT 44.935 188.675 45.225 188.770 ;
        RECT 44.635 188.630 45.225 188.675 ;
        RECT 47.875 188.630 48.525 188.675 ;
        RECT 29.355 188.490 36.930 188.630 ;
        RECT 40.470 188.490 41.990 188.630 ;
        RECT 29.355 188.445 29.645 188.490 ;
        RECT 36.790 188.350 36.930 188.490 ;
        RECT 31.195 188.290 31.485 188.335 ;
        RECT 36.240 188.290 36.560 188.350 ;
        RECT 31.195 188.150 36.560 188.290 ;
        RECT 31.195 188.105 31.485 188.150 ;
        RECT 36.240 188.090 36.560 188.150 ;
        RECT 36.700 188.090 37.020 188.350 ;
        RECT 37.160 188.290 37.480 188.350 ;
        RECT 37.635 188.290 37.925 188.335 ;
        RECT 37.160 188.150 37.925 188.290 ;
        RECT 37.160 188.090 37.480 188.150 ;
        RECT 37.635 188.105 37.925 188.150 ;
        RECT 38.555 188.290 38.845 188.335 ;
        RECT 40.380 188.290 40.700 188.350 ;
        RECT 38.555 188.150 40.700 188.290 ;
        RECT 41.850 188.290 41.990 188.490 ;
        RECT 44.635 188.490 48.525 188.630 ;
        RECT 44.635 188.445 44.925 188.490 ;
        RECT 47.875 188.445 48.525 188.490 ;
        RECT 49.120 188.630 49.440 188.690 ;
        RECT 50.500 188.630 50.820 188.690 ;
        RECT 51.970 188.630 52.110 188.785 ;
        RECT 52.800 188.770 53.120 189.030 ;
        RECT 53.350 189.015 53.490 189.170 ;
        RECT 56.020 189.110 56.340 189.170 ;
        RECT 56.480 189.310 56.800 189.370 ;
        RECT 58.795 189.310 59.085 189.355 ;
        RECT 56.480 189.170 59.085 189.310 ;
        RECT 56.480 189.110 56.800 189.170 ;
        RECT 58.795 189.125 59.085 189.170 ;
        RECT 66.140 189.310 66.460 189.370 ;
        RECT 70.370 189.355 70.510 189.510 ;
        RECT 73.040 189.450 73.360 189.510 ;
        RECT 69.375 189.310 69.665 189.355 ;
        RECT 70.295 189.310 70.585 189.355 ;
        RECT 66.140 189.170 69.665 189.310 ;
        RECT 70.185 189.170 70.585 189.310 ;
        RECT 66.140 189.110 66.460 189.170 ;
        RECT 69.375 189.125 69.665 189.170 ;
        RECT 70.295 189.125 70.585 189.170 ;
        RECT 70.755 189.310 71.045 189.355 ;
        RECT 74.510 189.310 74.650 189.850 ;
        RECT 82.715 189.850 89.460 189.990 ;
        RECT 82.715 189.805 83.005 189.850 ;
        RECT 89.140 189.790 89.460 189.850 ;
        RECT 90.060 189.990 90.380 190.050 ;
        RECT 98.815 189.990 99.105 190.035 ;
        RECT 90.060 189.850 99.105 189.990 ;
        RECT 90.060 189.790 90.380 189.850 ;
        RECT 98.815 189.805 99.105 189.850 ;
        RECT 106.160 189.990 106.480 190.050 ;
        RECT 110.760 189.990 111.080 190.050 ;
        RECT 106.160 189.850 111.080 189.990 ;
        RECT 106.160 189.790 106.480 189.850 ;
        RECT 110.760 189.790 111.080 189.850 ;
        RECT 74.895 189.650 75.185 189.695 ;
        RECT 74.895 189.510 87.530 189.650 ;
        RECT 74.895 189.465 75.185 189.510 ;
        RECT 79.495 189.310 79.785 189.355 ;
        RECT 83.635 189.310 83.925 189.355 ;
        RECT 85.920 189.310 86.240 189.370 ;
        RECT 70.755 189.170 72.810 189.310 ;
        RECT 74.510 189.170 86.240 189.310 ;
        RECT 87.390 189.310 87.530 189.510 ;
        RECT 87.760 189.450 88.080 189.710 ;
        RECT 89.600 189.650 89.920 189.710 ;
        RECT 91.900 189.650 92.220 189.710 ;
        RECT 89.600 189.510 92.220 189.650 ;
        RECT 89.600 189.450 89.920 189.510 ;
        RECT 91.900 189.450 92.220 189.510 ;
        RECT 92.475 189.650 92.765 189.695 ;
        RECT 95.595 189.650 95.885 189.695 ;
        RECT 97.485 189.650 97.775 189.695 ;
        RECT 92.475 189.510 97.775 189.650 ;
        RECT 92.475 189.465 92.765 189.510 ;
        RECT 95.595 189.465 95.885 189.510 ;
        RECT 97.485 189.465 97.775 189.510 ;
        RECT 103.515 189.650 103.805 189.695 ;
        RECT 106.635 189.650 106.925 189.695 ;
        RECT 108.525 189.650 108.815 189.695 ;
        RECT 103.515 189.510 108.815 189.650 ;
        RECT 103.515 189.465 103.805 189.510 ;
        RECT 106.635 189.465 106.925 189.510 ;
        RECT 108.525 189.465 108.815 189.510 ;
        RECT 87.390 189.170 90.750 189.310 ;
        RECT 70.755 189.125 71.045 189.170 ;
        RECT 71.290 189.030 71.430 189.170 ;
        RECT 53.275 188.785 53.565 189.015 ;
        RECT 53.735 188.785 54.025 189.015 ;
        RECT 54.195 188.970 54.485 189.015 ;
        RECT 55.560 188.970 55.880 189.030 ;
        RECT 54.195 188.830 55.880 188.970 ;
        RECT 54.195 188.785 54.485 188.830 ;
        RECT 52.890 188.630 53.030 188.770 ;
        RECT 49.120 188.490 51.650 188.630 ;
        RECT 51.970 188.490 53.030 188.630 ;
        RECT 49.120 188.430 49.440 188.490 ;
        RECT 50.500 188.430 50.820 188.490 ;
        RECT 43.155 188.290 43.445 188.335 ;
        RECT 50.960 188.290 51.280 188.350 ;
        RECT 41.850 188.150 51.280 188.290 ;
        RECT 51.510 188.290 51.650 188.490 ;
        RECT 53.810 188.290 53.950 188.785 ;
        RECT 55.560 188.770 55.880 188.830 ;
        RECT 60.160 188.770 60.480 189.030 ;
        RECT 61.080 188.970 61.400 189.030 ;
        RECT 63.380 188.970 63.700 189.030 ;
        RECT 64.775 188.970 65.065 189.015 ;
        RECT 61.080 188.830 65.065 188.970 ;
        RECT 61.080 188.770 61.400 188.830 ;
        RECT 63.380 188.770 63.700 188.830 ;
        RECT 64.775 188.785 65.065 188.830 ;
        RECT 69.835 188.785 70.125 189.015 ;
        RECT 57.875 188.630 58.165 188.675 ;
        RECT 62.015 188.630 62.305 188.675 ;
        RECT 57.875 188.490 62.305 188.630 ;
        RECT 57.875 188.445 58.165 188.490 ;
        RECT 62.015 188.445 62.305 188.490 ;
        RECT 66.140 188.430 66.460 188.690 ;
        RECT 66.600 188.630 66.920 188.690 ;
        RECT 68.455 188.630 68.745 188.675 ;
        RECT 66.600 188.490 68.745 188.630 ;
        RECT 69.910 188.630 70.050 188.785 ;
        RECT 71.200 188.770 71.520 189.030 ;
        RECT 72.135 188.785 72.425 189.015 ;
        RECT 72.670 188.970 72.810 189.170 ;
        RECT 79.495 189.125 79.785 189.170 ;
        RECT 83.635 189.125 83.925 189.170 ;
        RECT 85.920 189.110 86.240 189.170 ;
        RECT 74.880 188.970 75.200 189.030 ;
        RECT 72.670 188.830 75.200 188.970 ;
        RECT 70.280 188.630 70.600 188.690 ;
        RECT 69.910 188.490 70.600 188.630 ;
        RECT 72.210 188.630 72.350 188.785 ;
        RECT 74.880 188.770 75.200 188.830 ;
        RECT 75.815 188.970 76.105 189.015 ;
        RECT 78.100 188.970 78.420 189.030 ;
        RECT 75.815 188.830 78.420 188.970 ;
        RECT 75.815 188.785 76.105 188.830 ;
        RECT 78.100 188.770 78.420 188.830 ;
        RECT 78.575 188.970 78.865 189.015 ;
        RECT 80.875 188.970 81.165 189.015 ;
        RECT 84.555 188.970 84.845 189.015 ;
        RECT 78.575 188.830 84.845 188.970 ;
        RECT 78.575 188.785 78.865 188.830 ;
        RECT 80.875 188.785 81.165 188.830 ;
        RECT 84.555 188.785 84.845 188.830 ;
        RECT 88.220 188.970 88.540 189.030 ;
        RECT 88.695 188.970 88.985 189.015 ;
        RECT 88.220 188.830 88.985 188.970 ;
        RECT 88.220 188.770 88.540 188.830 ;
        RECT 88.695 188.785 88.985 188.830 ;
        RECT 89.140 188.630 89.460 188.690 ;
        RECT 72.210 188.490 89.460 188.630 ;
        RECT 66.600 188.430 66.920 188.490 ;
        RECT 68.455 188.445 68.745 188.490 ;
        RECT 70.280 188.430 70.600 188.490 ;
        RECT 89.140 188.430 89.460 188.490 ;
        RECT 51.510 188.150 53.950 188.290 ;
        RECT 55.100 188.290 55.420 188.350 ;
        RECT 55.575 188.290 55.865 188.335 ;
        RECT 55.100 188.150 55.865 188.290 ;
        RECT 38.555 188.105 38.845 188.150 ;
        RECT 40.380 188.090 40.700 188.150 ;
        RECT 43.155 188.105 43.445 188.150 ;
        RECT 50.960 188.090 51.280 188.150 ;
        RECT 55.100 188.090 55.420 188.150 ;
        RECT 55.575 188.105 55.865 188.150 ;
        RECT 58.335 188.290 58.625 188.335 ;
        RECT 58.780 188.290 59.100 188.350 ;
        RECT 58.335 188.150 59.100 188.290 ;
        RECT 58.335 188.105 58.625 188.150 ;
        RECT 58.780 188.090 59.100 188.150 ;
        RECT 61.095 188.290 61.385 188.335 ;
        RECT 65.680 188.290 66.000 188.350 ;
        RECT 61.095 188.150 66.000 188.290 ;
        RECT 61.095 188.105 61.385 188.150 ;
        RECT 65.680 188.090 66.000 188.150 ;
        RECT 67.980 188.290 68.300 188.350 ;
        RECT 69.360 188.290 69.680 188.350 ;
        RECT 67.980 188.150 69.680 188.290 ;
        RECT 70.370 188.290 70.510 188.430 ;
        RECT 73.500 188.290 73.820 188.350 ;
        RECT 70.370 188.150 73.820 188.290 ;
        RECT 67.980 188.090 68.300 188.150 ;
        RECT 69.360 188.090 69.680 188.150 ;
        RECT 73.500 188.090 73.820 188.150 ;
        RECT 80.400 188.090 80.720 188.350 ;
        RECT 85.000 188.090 85.320 188.350 ;
        RECT 86.855 188.290 87.145 188.335 ;
        RECT 90.060 188.290 90.380 188.350 ;
        RECT 86.855 188.150 90.380 188.290 ;
        RECT 90.610 188.290 90.750 189.170 ;
        RECT 96.960 189.110 97.280 189.370 ;
        RECT 98.340 189.310 98.660 189.370 ;
        RECT 105.700 189.310 106.020 189.370 ;
        RECT 109.395 189.310 109.685 189.355 ;
        RECT 110.300 189.310 110.620 189.370 ;
        RECT 98.340 189.170 110.620 189.310 ;
        RECT 98.340 189.110 98.660 189.170 ;
        RECT 105.700 189.110 106.020 189.170 ;
        RECT 109.395 189.125 109.685 189.170 ;
        RECT 110.300 189.110 110.620 189.170 ;
        RECT 91.440 188.990 91.760 189.030 ;
        RECT 91.395 188.770 91.760 188.990 ;
        RECT 92.475 188.970 92.765 189.015 ;
        RECT 96.055 188.970 96.345 189.015 ;
        RECT 97.890 188.970 98.180 189.015 ;
        RECT 92.475 188.830 98.180 188.970 ;
        RECT 92.475 188.785 92.765 188.830 ;
        RECT 96.055 188.785 96.345 188.830 ;
        RECT 97.890 188.785 98.180 188.830 ;
        RECT 99.720 188.770 100.040 189.030 ;
        RECT 91.395 188.675 91.685 188.770 ;
        RECT 91.095 188.630 91.685 188.675 ;
        RECT 94.335 188.630 94.985 188.675 ;
        RECT 91.095 188.490 94.985 188.630 ;
        RECT 91.095 188.445 91.385 188.490 ;
        RECT 94.335 188.445 94.985 188.490 ;
        RECT 101.100 188.630 101.420 188.690 ;
        RECT 102.435 188.675 102.725 188.990 ;
        RECT 103.515 188.970 103.805 189.015 ;
        RECT 107.095 188.970 107.385 189.015 ;
        RECT 108.930 188.970 109.220 189.015 ;
        RECT 103.515 188.830 109.220 188.970 ;
        RECT 103.515 188.785 103.805 188.830 ;
        RECT 107.095 188.785 107.385 188.830 ;
        RECT 108.930 188.785 109.220 188.830 ;
        RECT 109.840 188.970 110.160 189.030 ;
        RECT 110.775 188.970 111.065 189.015 ;
        RECT 109.840 188.830 111.065 188.970 ;
        RECT 109.840 188.770 110.160 188.830 ;
        RECT 110.775 188.785 111.065 188.830 ;
        RECT 102.135 188.630 102.725 188.675 ;
        RECT 105.375 188.630 106.025 188.675 ;
        RECT 101.100 188.490 106.025 188.630 ;
        RECT 101.100 188.430 101.420 188.490 ;
        RECT 102.135 188.445 102.425 188.490 ;
        RECT 105.375 188.445 106.025 188.490 ;
        RECT 108.000 188.430 108.320 188.690 ;
        RECT 100.180 188.290 100.500 188.350 ;
        RECT 90.610 188.150 100.500 188.290 ;
        RECT 86.855 188.105 87.145 188.150 ;
        RECT 90.060 188.090 90.380 188.150 ;
        RECT 100.180 188.090 100.500 188.150 ;
        RECT 100.640 188.090 100.960 188.350 ;
        RECT 109.855 188.290 110.145 188.335 ;
        RECT 110.300 188.290 110.620 188.350 ;
        RECT 109.855 188.150 110.620 188.290 ;
        RECT 109.855 188.105 110.145 188.150 ;
        RECT 110.300 188.090 110.620 188.150 ;
        RECT 26.970 187.470 113.450 187.950 ;
        RECT 38.095 187.270 38.385 187.315 ;
        RECT 41.760 187.270 42.080 187.330 ;
        RECT 38.095 187.130 42.080 187.270 ;
        RECT 38.095 187.085 38.385 187.130 ;
        RECT 41.760 187.070 42.080 187.130 ;
        RECT 51.420 187.070 51.740 187.330 ;
        RECT 54.655 187.085 54.945 187.315 ;
        RECT 58.320 187.270 58.640 187.330 ;
        RECT 55.650 187.130 58.640 187.270 ;
        RECT 30.375 186.930 30.665 186.975 ;
        RECT 31.180 186.930 31.500 186.990 ;
        RECT 33.615 186.930 34.265 186.975 ;
        RECT 30.375 186.790 34.265 186.930 ;
        RECT 30.375 186.745 30.965 186.790 ;
        RECT 30.675 186.430 30.965 186.745 ;
        RECT 31.180 186.730 31.500 186.790 ;
        RECT 33.615 186.745 34.265 186.790 ;
        RECT 36.255 186.930 36.545 186.975 ;
        RECT 37.620 186.930 37.940 186.990 ;
        RECT 36.255 186.790 37.940 186.930 ;
        RECT 36.255 186.745 36.545 186.790 ;
        RECT 37.620 186.730 37.940 186.790 ;
        RECT 39.575 186.930 39.865 186.975 ;
        RECT 42.815 186.930 43.465 186.975 ;
        RECT 39.575 186.790 43.465 186.930 ;
        RECT 39.575 186.745 40.165 186.790 ;
        RECT 42.815 186.745 43.465 186.790 ;
        RECT 31.755 186.590 32.045 186.635 ;
        RECT 35.335 186.590 35.625 186.635 ;
        RECT 37.170 186.590 37.460 186.635 ;
        RECT 31.755 186.450 37.460 186.590 ;
        RECT 31.755 186.405 32.045 186.450 ;
        RECT 35.335 186.405 35.625 186.450 ;
        RECT 37.170 186.405 37.460 186.450 ;
        RECT 39.875 186.430 40.165 186.745 ;
        RECT 45.440 186.730 45.760 186.990 ;
        RECT 45.900 186.930 46.220 186.990 ;
        RECT 51.895 186.930 52.185 186.975 ;
        RECT 45.900 186.790 52.185 186.930 ;
        RECT 54.730 186.930 54.870 187.085 ;
        RECT 55.650 186.930 55.790 187.130 ;
        RECT 58.320 187.070 58.640 187.130 ;
        RECT 59.700 187.270 60.020 187.330 ;
        RECT 64.300 187.270 64.620 187.330 ;
        RECT 68.440 187.270 68.760 187.330 ;
        RECT 59.700 187.130 64.620 187.270 ;
        RECT 59.700 187.070 60.020 187.130 ;
        RECT 64.300 187.070 64.620 187.130 ;
        RECT 65.310 187.130 68.760 187.270 ;
        RECT 54.730 186.790 55.790 186.930 ;
        RECT 45.900 186.730 46.220 186.790 ;
        RECT 51.895 186.745 52.185 186.790 ;
        RECT 65.310 186.650 65.450 187.130 ;
        RECT 68.440 187.070 68.760 187.130 ;
        RECT 68.915 187.270 69.205 187.315 ;
        RECT 69.360 187.270 69.680 187.330 ;
        RECT 68.915 187.130 69.680 187.270 ;
        RECT 68.915 187.085 69.205 187.130 ;
        RECT 69.360 187.070 69.680 187.130 ;
        RECT 69.820 187.070 70.140 187.330 ;
        RECT 70.295 187.270 70.585 187.315 ;
        RECT 71.200 187.270 71.520 187.330 ;
        RECT 70.295 187.130 71.520 187.270 ;
        RECT 70.295 187.085 70.585 187.130 ;
        RECT 71.200 187.070 71.520 187.130 ;
        RECT 74.880 187.070 75.200 187.330 ;
        RECT 77.180 187.270 77.500 187.330 ;
        RECT 85.000 187.270 85.320 187.330 ;
        RECT 89.600 187.270 89.920 187.330 ;
        RECT 77.180 187.130 89.920 187.270 ;
        RECT 77.180 187.070 77.500 187.130 ;
        RECT 85.000 187.070 85.320 187.130 ;
        RECT 89.600 187.070 89.920 187.130 ;
        RECT 91.900 187.270 92.220 187.330 ;
        RECT 100.640 187.270 100.960 187.330 ;
        RECT 102.035 187.270 102.325 187.315 ;
        RECT 91.900 187.130 98.570 187.270 ;
        RECT 91.900 187.070 92.220 187.130 ;
        RECT 69.910 186.930 70.050 187.070 ;
        RECT 66.230 186.790 70.050 186.930 ;
        RECT 70.740 186.930 71.060 186.990 ;
        RECT 72.595 186.930 72.885 186.975 ;
        RECT 75.655 186.930 75.945 186.975 ;
        RECT 70.740 186.790 72.885 186.930 ;
        RECT 40.955 186.590 41.245 186.635 ;
        RECT 44.535 186.590 44.825 186.635 ;
        RECT 46.370 186.590 46.660 186.635 ;
        RECT 40.955 186.450 46.660 186.590 ;
        RECT 37.635 186.250 37.925 186.295 ;
        RECT 38.080 186.250 38.400 186.310 ;
        RECT 37.635 186.110 38.400 186.250 ;
        RECT 37.635 186.065 37.925 186.110 ;
        RECT 38.080 186.050 38.400 186.110 ;
        RECT 39.460 186.250 39.780 186.310 ;
        RECT 40.010 186.250 40.150 186.430 ;
        RECT 40.955 186.405 41.245 186.450 ;
        RECT 44.535 186.405 44.825 186.450 ;
        RECT 46.370 186.405 46.660 186.450 ;
        RECT 47.295 186.405 47.585 186.635 ;
        RECT 53.735 186.590 54.025 186.635 ;
        RECT 55.115 186.590 55.405 186.635 ;
        RECT 53.735 186.450 55.405 186.590 ;
        RECT 53.735 186.405 54.025 186.450 ;
        RECT 55.115 186.405 55.405 186.450 ;
        RECT 57.950 186.450 59.010 186.590 ;
        RECT 39.460 186.110 40.150 186.250 ;
        RECT 43.600 186.250 43.920 186.310 ;
        RECT 46.835 186.250 47.125 186.295 ;
        RECT 43.600 186.110 47.125 186.250 ;
        RECT 39.460 186.050 39.780 186.110 ;
        RECT 43.600 186.050 43.920 186.110 ;
        RECT 46.835 186.065 47.125 186.110 ;
        RECT 31.755 185.910 32.045 185.955 ;
        RECT 34.875 185.910 35.165 185.955 ;
        RECT 36.765 185.910 37.055 185.955 ;
        RECT 31.755 185.770 37.055 185.910 ;
        RECT 31.755 185.725 32.045 185.770 ;
        RECT 34.875 185.725 35.165 185.770 ;
        RECT 36.765 185.725 37.055 185.770 ;
        RECT 40.955 185.910 41.245 185.955 ;
        RECT 44.075 185.910 44.365 185.955 ;
        RECT 45.965 185.910 46.255 185.955 ;
        RECT 40.955 185.770 46.255 185.910 ;
        RECT 40.955 185.725 41.245 185.770 ;
        RECT 44.075 185.725 44.365 185.770 ;
        RECT 45.965 185.725 46.255 185.770 ;
        RECT 26.120 185.570 26.440 185.630 ;
        RECT 28.895 185.570 29.185 185.615 ;
        RECT 33.940 185.570 34.260 185.630 ;
        RECT 26.120 185.430 34.260 185.570 ;
        RECT 26.120 185.370 26.440 185.430 ;
        RECT 28.895 185.385 29.185 185.430 ;
        RECT 33.940 185.370 34.260 185.430 ;
        RECT 44.520 185.570 44.840 185.630 ;
        RECT 47.370 185.570 47.510 186.405 ;
        RECT 47.740 186.250 48.060 186.310 ;
        RECT 52.355 186.250 52.645 186.295 ;
        RECT 54.640 186.250 54.960 186.310 ;
        RECT 57.950 186.250 58.090 186.450 ;
        RECT 47.740 186.110 58.090 186.250 ;
        RECT 47.740 186.050 48.060 186.110 ;
        RECT 52.355 186.065 52.645 186.110 ;
        RECT 54.640 186.050 54.960 186.110 ;
        RECT 58.335 186.065 58.625 186.295 ;
        RECT 58.870 186.250 59.010 186.450 ;
        RECT 60.620 186.390 60.940 186.650 ;
        RECT 61.080 186.390 61.400 186.650 ;
        RECT 65.220 186.390 65.540 186.650 ;
        RECT 66.230 186.635 66.370 186.790 ;
        RECT 70.740 186.730 71.060 186.790 ;
        RECT 72.595 186.745 72.885 186.790 ;
        RECT 73.130 186.790 75.945 186.930 ;
        RECT 66.155 186.405 66.445 186.635 ;
        RECT 68.440 186.390 68.760 186.650 ;
        RECT 68.900 186.590 69.220 186.650 ;
        RECT 73.130 186.590 73.270 186.790 ;
        RECT 75.655 186.745 75.945 186.790 ;
        RECT 76.720 186.730 77.040 186.990 ;
        RECT 85.920 186.975 86.240 186.990 ;
        RECT 82.355 186.930 82.645 186.975 ;
        RECT 85.595 186.930 86.245 186.975 ;
        RECT 82.355 186.790 86.245 186.930 ;
        RECT 82.355 186.745 82.945 186.790 ;
        RECT 85.595 186.745 86.245 186.790 ;
        RECT 88.235 186.930 88.525 186.975 ;
        RECT 90.520 186.930 90.840 186.990 ;
        RECT 88.235 186.790 90.840 186.930 ;
        RECT 88.235 186.745 88.525 186.790 ;
        RECT 78.575 186.590 78.865 186.635 ;
        RECT 68.900 186.450 73.270 186.590 ;
        RECT 75.430 186.450 78.865 186.590 ;
        RECT 68.900 186.390 69.220 186.450 ;
        RECT 75.430 186.310 75.570 186.450 ;
        RECT 78.575 186.405 78.865 186.450 ;
        RECT 79.035 186.405 79.325 186.635 ;
        RECT 79.495 186.590 79.785 186.635 ;
        RECT 79.940 186.590 80.260 186.650 ;
        RECT 79.495 186.450 80.260 186.590 ;
        RECT 79.495 186.405 79.785 186.450 ;
        RECT 61.555 186.250 61.845 186.295 ;
        RECT 58.870 186.110 61.845 186.250 ;
        RECT 61.555 186.065 61.845 186.110 ;
        RECT 66.615 186.065 66.905 186.295 ;
        RECT 67.075 186.065 67.365 186.295 ;
        RECT 67.535 186.250 67.825 186.295 ;
        RECT 70.280 186.250 70.600 186.310 ;
        RECT 67.535 186.110 70.600 186.250 ;
        RECT 67.535 186.065 67.825 186.110 ;
        RECT 49.580 185.710 49.900 185.970 ;
        RECT 50.040 185.910 50.360 185.970 ;
        RECT 54.180 185.910 54.500 185.970 ;
        RECT 50.040 185.770 54.500 185.910 ;
        RECT 58.410 185.910 58.550 186.065 ;
        RECT 58.795 185.910 59.085 185.955 ;
        RECT 58.410 185.770 59.085 185.910 ;
        RECT 50.040 185.710 50.360 185.770 ;
        RECT 54.180 185.710 54.500 185.770 ;
        RECT 58.795 185.725 59.085 185.770 ;
        RECT 44.520 185.430 47.510 185.570 ;
        RECT 48.215 185.570 48.505 185.615 ;
        RECT 52.800 185.570 53.120 185.630 ;
        RECT 48.215 185.430 53.120 185.570 ;
        RECT 66.690 185.570 66.830 186.065 ;
        RECT 67.150 185.910 67.290 186.065 ;
        RECT 70.280 186.050 70.600 186.110 ;
        RECT 75.340 186.050 75.660 186.310 ;
        RECT 75.800 186.250 76.120 186.310 ;
        RECT 79.110 186.250 79.250 186.405 ;
        RECT 79.940 186.390 80.260 186.450 ;
        RECT 80.400 186.390 80.720 186.650 ;
        RECT 82.655 186.430 82.945 186.745 ;
        RECT 85.920 186.730 86.240 186.745 ;
        RECT 90.520 186.730 90.840 186.790 ;
        RECT 93.295 186.930 93.585 186.975 ;
        RECT 97.880 186.930 98.200 186.990 ;
        RECT 93.295 186.790 98.200 186.930 ;
        RECT 93.295 186.745 93.585 186.790 ;
        RECT 97.880 186.730 98.200 186.790 ;
        RECT 83.735 186.590 84.025 186.635 ;
        RECT 87.315 186.590 87.605 186.635 ;
        RECT 89.150 186.590 89.440 186.635 ;
        RECT 83.735 186.450 89.440 186.590 ;
        RECT 83.735 186.405 84.025 186.450 ;
        RECT 87.315 186.405 87.605 186.450 ;
        RECT 89.150 186.405 89.440 186.450 ;
        RECT 90.060 186.390 90.380 186.650 ;
        RECT 93.740 186.590 94.060 186.650 ;
        RECT 95.135 186.590 95.425 186.635 ;
        RECT 93.740 186.450 95.425 186.590 ;
        RECT 93.740 186.390 94.060 186.450 ;
        RECT 95.135 186.405 95.425 186.450 ;
        RECT 95.580 186.390 95.900 186.650 ;
        RECT 96.040 186.390 96.360 186.650 ;
        RECT 96.500 186.590 96.820 186.650 ;
        RECT 96.975 186.590 97.265 186.635 ;
        RECT 96.500 186.450 97.265 186.590 ;
        RECT 96.500 186.390 96.820 186.450 ;
        RECT 96.975 186.405 97.265 186.450 ;
        RECT 97.435 186.590 97.725 186.635 ;
        RECT 98.430 186.590 98.570 187.130 ;
        RECT 100.640 187.130 102.325 187.270 ;
        RECT 100.640 187.070 100.960 187.130 ;
        RECT 102.035 187.085 102.325 187.130 ;
        RECT 107.080 187.270 107.400 187.330 ;
        RECT 107.080 187.130 110.070 187.270 ;
        RECT 107.080 187.070 107.400 187.130 ;
        RECT 98.800 186.730 99.120 186.990 ;
        RECT 100.180 186.930 100.500 186.990 ;
        RECT 102.495 186.930 102.785 186.975 ;
        RECT 100.180 186.790 102.785 186.930 ;
        RECT 100.180 186.730 100.500 186.790 ;
        RECT 102.495 186.745 102.785 186.790 ;
        RECT 107.170 186.790 108.690 186.930 ;
        RECT 97.435 186.450 98.570 186.590 ;
        RECT 98.890 186.590 99.030 186.730 ;
        RECT 104.780 186.590 105.100 186.650 ;
        RECT 107.170 186.590 107.310 186.790 ;
        RECT 98.890 186.450 107.310 186.590 ;
        RECT 97.435 186.405 97.725 186.450 ;
        RECT 104.780 186.390 105.100 186.450 ;
        RECT 107.540 186.390 107.860 186.650 ;
        RECT 108.550 186.635 108.690 186.790 ;
        RECT 108.475 186.405 108.765 186.635 ;
        RECT 109.380 186.390 109.700 186.650 ;
        RECT 109.930 186.635 110.070 187.130 ;
        RECT 109.855 186.405 110.145 186.635 ;
        RECT 110.315 186.590 110.605 186.635 ;
        RECT 110.760 186.590 111.080 186.650 ;
        RECT 110.315 186.450 111.080 186.590 ;
        RECT 110.315 186.405 110.605 186.450 ;
        RECT 110.760 186.390 111.080 186.450 ;
        RECT 75.800 186.110 79.250 186.250 ;
        RECT 85.000 186.250 85.320 186.310 ;
        RECT 89.615 186.250 89.905 186.295 ;
        RECT 90.980 186.250 91.300 186.310 ;
        RECT 85.000 186.110 91.300 186.250 ;
        RECT 75.800 186.050 76.120 186.110 ;
        RECT 85.000 186.050 85.320 186.110 ;
        RECT 89.615 186.065 89.905 186.110 ;
        RECT 90.980 186.050 91.300 186.110 ;
        RECT 94.200 186.250 94.520 186.310 ;
        RECT 95.670 186.250 95.810 186.390 ;
        RECT 94.200 186.110 95.810 186.250 ;
        RECT 98.815 186.250 99.105 186.295 ;
        RECT 100.180 186.250 100.500 186.310 ;
        RECT 101.100 186.250 101.420 186.310 ;
        RECT 98.815 186.110 101.420 186.250 ;
        RECT 94.200 186.050 94.520 186.110 ;
        RECT 98.815 186.065 99.105 186.110 ;
        RECT 100.180 186.050 100.500 186.110 ;
        RECT 101.100 186.050 101.420 186.110 ;
        RECT 101.575 186.250 101.865 186.295 ;
        RECT 102.480 186.250 102.800 186.310 ;
        RECT 101.575 186.110 102.800 186.250 ;
        RECT 101.575 186.065 101.865 186.110 ;
        RECT 102.480 186.050 102.800 186.110 ;
        RECT 102.940 186.250 103.260 186.310 ;
        RECT 111.695 186.250 111.985 186.295 ;
        RECT 102.940 186.110 111.985 186.250 ;
        RECT 102.940 186.050 103.260 186.110 ;
        RECT 111.695 186.065 111.985 186.110 ;
        RECT 71.200 185.910 71.520 185.970 ;
        RECT 67.150 185.770 71.520 185.910 ;
        RECT 71.200 185.710 71.520 185.770 ;
        RECT 72.580 185.710 72.900 185.970 ;
        RECT 73.500 185.910 73.820 185.970 ;
        RECT 77.195 185.910 77.485 185.955 ;
        RECT 83.735 185.910 84.025 185.955 ;
        RECT 86.855 185.910 87.145 185.955 ;
        RECT 88.745 185.910 89.035 185.955 ;
        RECT 94.660 185.910 94.980 185.970 ;
        RECT 73.500 185.770 77.485 185.910 ;
        RECT 73.500 185.710 73.820 185.770 ;
        RECT 77.195 185.725 77.485 185.770 ;
        RECT 77.730 185.770 83.390 185.910 ;
        RECT 72.670 185.570 72.810 185.710 ;
        RECT 66.690 185.430 72.810 185.570 ;
        RECT 75.815 185.570 76.105 185.615 ;
        RECT 77.730 185.570 77.870 185.770 ;
        RECT 75.815 185.430 77.870 185.570 ;
        RECT 78.100 185.570 78.420 185.630 ;
        RECT 80.875 185.570 81.165 185.615 ;
        RECT 81.320 185.570 81.640 185.630 ;
        RECT 78.100 185.430 81.640 185.570 ;
        RECT 83.250 185.570 83.390 185.770 ;
        RECT 83.735 185.770 89.035 185.910 ;
        RECT 83.735 185.725 84.025 185.770 ;
        RECT 86.855 185.725 87.145 185.770 ;
        RECT 88.745 185.725 89.035 185.770 ;
        RECT 89.690 185.770 94.980 185.910 ;
        RECT 89.690 185.570 89.830 185.770 ;
        RECT 94.660 185.710 94.980 185.770 ;
        RECT 104.335 185.910 104.625 185.955 ;
        RECT 106.620 185.910 106.940 185.970 ;
        RECT 104.335 185.770 106.940 185.910 ;
        RECT 104.335 185.725 104.625 185.770 ;
        RECT 106.620 185.710 106.940 185.770 ;
        RECT 83.250 185.430 89.830 185.570 ;
        RECT 90.060 185.570 90.380 185.630 ;
        RECT 93.755 185.570 94.045 185.615 ;
        RECT 90.060 185.430 94.045 185.570 ;
        RECT 44.520 185.370 44.840 185.430 ;
        RECT 48.215 185.385 48.505 185.430 ;
        RECT 52.800 185.370 53.120 185.430 ;
        RECT 75.815 185.385 76.105 185.430 ;
        RECT 78.100 185.370 78.420 185.430 ;
        RECT 80.875 185.385 81.165 185.430 ;
        RECT 81.320 185.370 81.640 185.430 ;
        RECT 90.060 185.370 90.380 185.430 ;
        RECT 93.755 185.385 94.045 185.430 ;
        RECT 104.795 185.570 105.085 185.615 ;
        RECT 107.080 185.570 107.400 185.630 ;
        RECT 104.795 185.430 107.400 185.570 ;
        RECT 104.795 185.385 105.085 185.430 ;
        RECT 107.080 185.370 107.400 185.430 ;
        RECT 26.970 184.750 113.450 185.230 ;
        RECT 34.860 184.550 35.180 184.610 ;
        RECT 36.715 184.550 37.005 184.595 ;
        RECT 40.840 184.550 41.160 184.610 ;
        RECT 34.860 184.410 37.005 184.550 ;
        RECT 34.860 184.350 35.180 184.410 ;
        RECT 36.715 184.365 37.005 184.410 ;
        RECT 39.550 184.410 41.160 184.550 ;
        RECT 28.880 184.210 29.200 184.270 ;
        RECT 31.655 184.210 31.945 184.255 ;
        RECT 39.550 184.210 39.690 184.410 ;
        RECT 40.840 184.350 41.160 184.410 ;
        RECT 41.315 184.550 41.605 184.595 ;
        RECT 42.220 184.550 42.540 184.610 ;
        RECT 41.315 184.410 42.540 184.550 ;
        RECT 41.315 184.365 41.605 184.410 ;
        RECT 42.220 184.350 42.540 184.410 ;
        RECT 45.455 184.550 45.745 184.595 ;
        RECT 46.360 184.550 46.680 184.610 ;
        RECT 45.455 184.410 46.680 184.550 ;
        RECT 45.455 184.365 45.745 184.410 ;
        RECT 46.360 184.350 46.680 184.410 ;
        RECT 54.640 184.550 54.960 184.610 ;
        RECT 55.115 184.550 55.405 184.595 ;
        RECT 60.160 184.550 60.480 184.610 ;
        RECT 61.095 184.550 61.385 184.595 ;
        RECT 54.640 184.410 58.090 184.550 ;
        RECT 54.640 184.350 54.960 184.410 ;
        RECT 55.115 184.365 55.405 184.410 ;
        RECT 28.880 184.070 31.945 184.210 ;
        RECT 28.880 184.010 29.200 184.070 ;
        RECT 31.655 184.025 31.945 184.070 ;
        RECT 34.490 184.070 39.690 184.210 ;
        RECT 29.355 183.870 29.645 183.915 ;
        RECT 31.180 183.870 31.500 183.930 ;
        RECT 29.355 183.730 31.500 183.870 ;
        RECT 29.355 183.685 29.645 183.730 ;
        RECT 31.180 183.670 31.500 183.730 ;
        RECT 32.100 183.870 32.420 183.930 ;
        RECT 34.490 183.915 34.630 184.070 ;
        RECT 39.550 183.915 39.690 184.070 ;
        RECT 40.380 184.210 40.700 184.270 ;
        RECT 48.315 184.210 48.605 184.255 ;
        RECT 51.435 184.210 51.725 184.255 ;
        RECT 53.325 184.210 53.615 184.255 ;
        RECT 40.380 184.070 47.510 184.210 ;
        RECT 40.380 184.010 40.700 184.070 ;
        RECT 34.415 183.870 34.705 183.915 ;
        RECT 39.015 183.870 39.305 183.915 ;
        RECT 32.100 183.730 34.705 183.870 ;
        RECT 32.100 183.670 32.420 183.730 ;
        RECT 34.415 183.685 34.705 183.730 ;
        RECT 35.870 183.730 39.305 183.870 ;
        RECT 35.870 183.590 36.010 183.730 ;
        RECT 39.015 183.685 39.305 183.730 ;
        RECT 39.475 183.685 39.765 183.915 ;
        RECT 40.840 183.870 41.160 183.930 ;
        RECT 44.075 183.870 44.365 183.915 ;
        RECT 46.820 183.870 47.140 183.930 ;
        RECT 40.840 183.730 47.140 183.870 ;
        RECT 40.840 183.670 41.160 183.730 ;
        RECT 44.075 183.685 44.365 183.730 ;
        RECT 46.820 183.670 47.140 183.730 ;
        RECT 26.120 183.530 26.440 183.590 ;
        RECT 29.815 183.530 30.105 183.575 ;
        RECT 30.275 183.530 30.565 183.575 ;
        RECT 26.120 183.390 30.565 183.530 ;
        RECT 26.120 183.330 26.440 183.390 ;
        RECT 29.815 183.345 30.105 183.390 ;
        RECT 30.275 183.345 30.565 183.390 ;
        RECT 33.495 183.530 33.785 183.575 ;
        RECT 35.780 183.530 36.100 183.590 ;
        RECT 33.495 183.390 36.100 183.530 ;
        RECT 33.495 183.345 33.785 183.390 ;
        RECT 35.780 183.330 36.100 183.390 ;
        RECT 43.155 183.530 43.445 183.575 ;
        RECT 45.900 183.530 46.220 183.590 ;
        RECT 47.370 183.550 47.510 184.070 ;
        RECT 48.315 184.070 53.615 184.210 ;
        RECT 48.315 184.025 48.605 184.070 ;
        RECT 51.435 184.025 51.725 184.070 ;
        RECT 53.325 184.025 53.615 184.070 ;
        RECT 52.800 183.670 53.120 183.930 ;
        RECT 57.950 183.915 58.090 184.410 ;
        RECT 60.160 184.410 61.385 184.550 ;
        RECT 60.160 184.350 60.480 184.410 ;
        RECT 61.095 184.365 61.385 184.410 ;
        RECT 73.975 184.550 74.265 184.595 ;
        RECT 74.880 184.550 75.200 184.610 ;
        RECT 79.480 184.550 79.800 184.610 ;
        RECT 73.975 184.410 75.200 184.550 ;
        RECT 73.975 184.365 74.265 184.410 ;
        RECT 74.880 184.350 75.200 184.410 ;
        RECT 75.890 184.410 79.800 184.550 ;
        RECT 68.440 184.210 68.760 184.270 ;
        RECT 70.740 184.210 71.060 184.270 ;
        RECT 75.890 184.210 76.030 184.410 ;
        RECT 79.480 184.350 79.800 184.410 ;
        RECT 106.175 184.550 106.465 184.595 ;
        RECT 109.840 184.550 110.160 184.610 ;
        RECT 106.175 184.410 110.160 184.550 ;
        RECT 106.175 184.365 106.465 184.410 ;
        RECT 109.840 184.350 110.160 184.410 ;
        RECT 76.720 184.210 77.040 184.270 ;
        RECT 68.440 184.070 71.060 184.210 ;
        RECT 68.440 184.010 68.760 184.070 ;
        RECT 70.740 184.010 71.060 184.070 ;
        RECT 71.290 184.070 76.030 184.210 ;
        RECT 76.350 184.070 77.040 184.210 ;
        RECT 57.875 183.685 58.165 183.915 ;
        RECT 58.795 183.870 59.085 183.915 ;
        RECT 60.620 183.870 60.940 183.930 ;
        RECT 62.015 183.870 62.305 183.915 ;
        RECT 58.795 183.730 62.305 183.870 ;
        RECT 58.795 183.685 59.085 183.730 ;
        RECT 60.620 183.670 60.940 183.730 ;
        RECT 62.015 183.685 62.305 183.730 ;
        RECT 64.760 183.670 65.080 183.930 ;
        RECT 67.520 183.870 67.840 183.930 ;
        RECT 67.520 183.730 69.130 183.870 ;
        RECT 67.520 183.670 67.840 183.730 ;
        RECT 43.155 183.390 46.220 183.530 ;
        RECT 43.155 183.345 43.445 183.390 ;
        RECT 45.900 183.330 46.220 183.390 ;
        RECT 38.555 183.190 38.845 183.235 ;
        RECT 39.000 183.190 39.320 183.250 ;
        RECT 47.235 183.235 47.525 183.550 ;
        RECT 48.315 183.530 48.605 183.575 ;
        RECT 51.895 183.530 52.185 183.575 ;
        RECT 53.730 183.530 54.020 183.575 ;
        RECT 48.315 183.390 54.020 183.530 ;
        RECT 48.315 183.345 48.605 183.390 ;
        RECT 51.895 183.345 52.185 183.390 ;
        RECT 53.730 183.345 54.020 183.390 ;
        RECT 54.180 183.330 54.500 183.590 ;
        RECT 56.480 183.330 56.800 183.590 ;
        RECT 65.695 183.530 65.985 183.575 ;
        RECT 59.330 183.390 65.985 183.530 ;
        RECT 43.615 183.190 43.905 183.235 ;
        RECT 38.555 183.050 43.905 183.190 ;
        RECT 38.555 183.005 38.845 183.050 ;
        RECT 39.000 182.990 39.320 183.050 ;
        RECT 43.615 183.005 43.905 183.050 ;
        RECT 46.935 183.190 47.525 183.235 ;
        RECT 50.175 183.190 50.825 183.235 ;
        RECT 46.935 183.050 50.825 183.190 ;
        RECT 46.935 183.005 47.225 183.050 ;
        RECT 50.175 183.005 50.825 183.050 ;
        RECT 52.340 183.190 52.660 183.250 ;
        RECT 59.330 183.235 59.470 183.390 ;
        RECT 65.695 183.345 65.985 183.390 ;
        RECT 68.455 183.345 68.745 183.575 ;
        RECT 59.255 183.190 59.545 183.235 ;
        RECT 68.530 183.190 68.670 183.345 ;
        RECT 52.340 183.050 59.545 183.190 ;
        RECT 52.340 182.990 52.660 183.050 ;
        RECT 59.255 183.005 59.545 183.050 ;
        RECT 59.790 183.050 68.670 183.190 ;
        RECT 68.990 183.190 69.130 183.730 ;
        RECT 70.295 183.530 70.585 183.575 ;
        RECT 70.830 183.530 70.970 184.010 ;
        RECT 71.290 183.575 71.430 184.070 ;
        RECT 73.515 183.870 73.805 183.915 ;
        RECT 74.880 183.870 75.200 183.930 ;
        RECT 73.515 183.730 75.200 183.870 ;
        RECT 73.515 183.685 73.805 183.730 ;
        RECT 74.880 183.670 75.200 183.730 ;
        RECT 70.295 183.390 70.970 183.530 ;
        RECT 70.295 183.345 70.585 183.390 ;
        RECT 71.215 183.345 71.505 183.575 ;
        RECT 71.675 183.345 71.965 183.575 ;
        RECT 72.135 183.345 72.425 183.575 ;
        RECT 75.340 183.530 75.660 183.590 ;
        RECT 74.050 183.390 75.660 183.530 ;
        RECT 70.740 183.190 71.060 183.250 ;
        RECT 71.750 183.190 71.890 183.345 ;
        RECT 68.990 183.050 71.890 183.190 ;
        RECT 72.210 183.190 72.350 183.345 ;
        RECT 73.040 183.190 73.360 183.250 ;
        RECT 72.210 183.050 73.360 183.190 ;
        RECT 29.340 182.850 29.660 182.910 ;
        RECT 30.735 182.850 31.025 182.895 ;
        RECT 29.340 182.710 31.025 182.850 ;
        RECT 29.340 182.650 29.660 182.710 ;
        RECT 30.735 182.665 31.025 182.710 ;
        RECT 33.940 182.850 34.260 182.910 ;
        RECT 47.740 182.850 48.060 182.910 ;
        RECT 33.940 182.710 48.060 182.850 ;
        RECT 33.940 182.650 34.260 182.710 ;
        RECT 47.740 182.650 48.060 182.710 ;
        RECT 50.960 182.850 51.280 182.910 ;
        RECT 59.790 182.850 59.930 183.050 ;
        RECT 70.740 182.990 71.060 183.050 ;
        RECT 73.040 182.990 73.360 183.050 ;
        RECT 50.960 182.710 59.930 182.850 ;
        RECT 64.300 182.850 64.620 182.910 ;
        RECT 67.520 182.850 67.840 182.910 ;
        RECT 64.300 182.710 67.840 182.850 ;
        RECT 50.960 182.650 51.280 182.710 ;
        RECT 64.300 182.650 64.620 182.710 ;
        RECT 67.520 182.650 67.840 182.710 ;
        RECT 67.980 182.850 68.300 182.910 ;
        RECT 74.050 182.850 74.190 183.390 ;
        RECT 75.340 183.330 75.660 183.390 ;
        RECT 75.800 183.330 76.120 183.590 ;
        RECT 76.350 183.575 76.490 184.070 ;
        RECT 76.720 184.010 77.040 184.070 ;
        RECT 77.180 184.210 77.500 184.270 ;
        RECT 80.400 184.210 80.720 184.270 ;
        RECT 77.180 184.070 80.720 184.210 ;
        RECT 77.180 184.010 77.500 184.070 ;
        RECT 80.400 184.010 80.720 184.070 ;
        RECT 85.920 184.210 86.240 184.270 ;
        RECT 96.515 184.210 96.805 184.255 ;
        RECT 85.920 184.070 96.805 184.210 ;
        RECT 85.920 184.010 86.240 184.070 ;
        RECT 96.515 184.025 96.805 184.070 ;
        RECT 96.960 184.210 97.280 184.270 ;
        RECT 102.940 184.210 103.260 184.270 ;
        RECT 96.960 184.070 103.260 184.210 ;
        RECT 96.960 184.010 97.280 184.070 ;
        RECT 102.940 184.010 103.260 184.070 ;
        RECT 85.460 183.870 85.780 183.930 ;
        RECT 100.640 183.870 100.960 183.930 ;
        RECT 85.460 183.730 100.960 183.870 ;
        RECT 85.460 183.670 85.780 183.730 ;
        RECT 76.275 183.345 76.565 183.575 ;
        RECT 77.180 183.330 77.500 183.590 ;
        RECT 78.100 183.530 78.420 183.590 ;
        RECT 79.035 183.530 79.325 183.575 ;
        RECT 78.100 183.390 79.325 183.530 ;
        RECT 78.100 183.330 78.420 183.390 ;
        RECT 79.035 183.345 79.325 183.390 ;
        RECT 79.495 183.345 79.785 183.575 ;
        RECT 79.955 183.345 80.245 183.575 ;
        RECT 80.400 183.530 80.720 183.590 ;
        RECT 80.875 183.530 81.165 183.575 ;
        RECT 84.540 183.530 84.860 183.590 ;
        RECT 80.400 183.390 84.860 183.530 ;
        RECT 67.980 182.710 74.190 182.850 ;
        RECT 75.430 182.850 75.570 183.330 ;
        RECT 75.890 183.190 76.030 183.330 ;
        RECT 79.570 183.190 79.710 183.345 ;
        RECT 75.890 183.050 79.710 183.190 ;
        RECT 80.030 183.190 80.170 183.345 ;
        RECT 80.400 183.330 80.720 183.390 ;
        RECT 80.875 183.345 81.165 183.390 ;
        RECT 84.540 183.330 84.860 183.390 ;
        RECT 85.015 183.345 85.305 183.575 ;
        RECT 85.935 183.530 86.225 183.575 ;
        RECT 87.300 183.530 87.620 183.590 ;
        RECT 85.935 183.390 87.620 183.530 ;
        RECT 85.935 183.345 86.225 183.390 ;
        RECT 84.080 183.190 84.400 183.250 ;
        RECT 80.030 183.050 84.400 183.190 ;
        RECT 84.080 182.990 84.400 183.050 ;
        RECT 85.090 182.910 85.230 183.345 ;
        RECT 87.300 183.330 87.620 183.390 ;
        RECT 88.680 183.330 89.000 183.590 ;
        RECT 89.690 183.575 89.830 183.730 ;
        RECT 100.640 183.670 100.960 183.730 ;
        RECT 89.615 183.345 89.905 183.575 ;
        RECT 90.075 183.345 90.365 183.575 ;
        RECT 89.140 183.190 89.460 183.250 ;
        RECT 90.150 183.190 90.290 183.345 ;
        RECT 90.520 183.330 90.840 183.590 ;
        RECT 92.835 183.530 93.125 183.575 ;
        RECT 96.040 183.530 96.360 183.590 ;
        RECT 92.835 183.390 96.360 183.530 ;
        RECT 92.835 183.345 93.125 183.390 ;
        RECT 96.040 183.330 96.360 183.390 ;
        RECT 96.975 183.530 97.265 183.575 ;
        RECT 97.420 183.530 97.740 183.590 ;
        RECT 98.355 183.530 98.645 183.575 ;
        RECT 96.975 183.390 98.645 183.530 ;
        RECT 96.975 183.345 97.265 183.390 ;
        RECT 97.420 183.330 97.740 183.390 ;
        RECT 98.355 183.345 98.645 183.390 ;
        RECT 99.735 183.530 100.025 183.575 ;
        RECT 100.180 183.530 100.500 183.590 ;
        RECT 99.735 183.390 100.500 183.530 ;
        RECT 99.735 183.345 100.025 183.390 ;
        RECT 100.180 183.330 100.500 183.390 ;
        RECT 102.940 183.330 103.260 183.590 ;
        RECT 106.160 183.530 106.480 183.590 ;
        RECT 106.635 183.530 106.925 183.575 ;
        RECT 106.160 183.390 106.925 183.530 ;
        RECT 106.160 183.330 106.480 183.390 ;
        RECT 106.635 183.345 106.925 183.390 ;
        RECT 109.855 183.530 110.145 183.575 ;
        RECT 111.695 183.530 111.985 183.575 ;
        RECT 109.855 183.390 111.985 183.530 ;
        RECT 109.855 183.345 110.145 183.390 ;
        RECT 111.695 183.345 111.985 183.390 ;
        RECT 94.200 183.190 94.520 183.250 ;
        RECT 89.140 183.050 94.520 183.190 ;
        RECT 89.140 182.990 89.460 183.050 ;
        RECT 94.200 182.990 94.520 183.050 ;
        RECT 94.660 183.190 94.980 183.250 ;
        RECT 94.660 183.050 98.110 183.190 ;
        RECT 94.660 182.990 94.980 183.050 ;
        RECT 77.180 182.850 77.500 182.910 ;
        RECT 75.430 182.710 77.500 182.850 ;
        RECT 67.980 182.650 68.300 182.710 ;
        RECT 77.180 182.650 77.500 182.710 ;
        RECT 77.655 182.850 77.945 182.895 ;
        RECT 79.940 182.850 80.260 182.910 ;
        RECT 77.655 182.710 80.260 182.850 ;
        RECT 77.655 182.665 77.945 182.710 ;
        RECT 79.940 182.650 80.260 182.710 ;
        RECT 85.000 182.650 85.320 182.910 ;
        RECT 86.380 182.650 86.700 182.910 ;
        RECT 90.520 182.850 90.840 182.910 ;
        RECT 91.915 182.850 92.205 182.895 ;
        RECT 90.520 182.710 92.205 182.850 ;
        RECT 90.520 182.650 90.840 182.710 ;
        RECT 91.915 182.665 92.205 182.710 ;
        RECT 95.595 182.850 95.885 182.895 ;
        RECT 96.500 182.850 96.820 182.910 ;
        RECT 97.970 182.895 98.110 183.050 ;
        RECT 95.595 182.710 96.820 182.850 ;
        RECT 95.595 182.665 95.885 182.710 ;
        RECT 96.500 182.650 96.820 182.710 ;
        RECT 97.895 182.665 98.185 182.895 ;
        RECT 102.480 182.650 102.800 182.910 ;
        RECT 110.760 182.650 111.080 182.910 ;
        RECT 26.970 182.030 113.450 182.510 ;
        RECT 30.735 181.830 31.025 181.875 ;
        RECT 33.020 181.830 33.340 181.890 ;
        RECT 30.735 181.690 33.340 181.830 ;
        RECT 30.735 181.645 31.025 181.690 ;
        RECT 33.020 181.630 33.340 181.690 ;
        RECT 37.620 181.830 37.940 181.890 ;
        RECT 41.760 181.830 42.080 181.890 ;
        RECT 37.620 181.690 42.080 181.830 ;
        RECT 37.620 181.630 37.940 181.690 ;
        RECT 41.760 181.630 42.080 181.690 ;
        RECT 44.520 181.630 44.840 181.890 ;
        RECT 49.580 181.830 49.900 181.890 ;
        RECT 49.210 181.690 49.900 181.830 ;
        RECT 27.040 181.490 27.360 181.550 ;
        RECT 32.215 181.490 32.505 181.535 ;
        RECT 35.455 181.490 36.105 181.535 ;
        RECT 27.040 181.350 36.105 181.490 ;
        RECT 27.040 181.290 27.360 181.350 ;
        RECT 32.215 181.305 32.805 181.350 ;
        RECT 35.455 181.305 36.105 181.350 ;
        RECT 38.540 181.490 38.860 181.550 ;
        RECT 38.540 181.350 40.150 181.490 ;
        RECT 28.880 181.150 29.200 181.210 ;
        RECT 30.275 181.150 30.565 181.195 ;
        RECT 28.880 181.010 30.565 181.150 ;
        RECT 28.880 180.950 29.200 181.010 ;
        RECT 30.275 180.965 30.565 181.010 ;
        RECT 32.515 180.990 32.805 181.305 ;
        RECT 38.540 181.290 38.860 181.350 ;
        RECT 40.010 181.210 40.150 181.350 ;
        RECT 40.380 181.290 40.700 181.550 ;
        RECT 49.210 181.490 49.350 181.690 ;
        RECT 49.580 181.630 49.900 181.690 ;
        RECT 56.020 181.830 56.340 181.890 ;
        RECT 58.335 181.830 58.625 181.875 ;
        RECT 64.760 181.830 65.080 181.890 ;
        RECT 56.020 181.690 65.080 181.830 ;
        RECT 56.020 181.630 56.340 181.690 ;
        RECT 58.335 181.645 58.625 181.690 ;
        RECT 64.760 181.630 65.080 181.690 ;
        RECT 66.140 181.830 66.460 181.890 ;
        RECT 69.835 181.830 70.125 181.875 ;
        RECT 66.140 181.690 70.125 181.830 ;
        RECT 66.140 181.630 66.460 181.690 ;
        RECT 69.835 181.645 70.125 181.690 ;
        RECT 75.340 181.830 75.660 181.890 ;
        RECT 75.815 181.830 76.105 181.875 ;
        RECT 75.340 181.690 76.105 181.830 ;
        RECT 75.340 181.630 75.660 181.690 ;
        RECT 75.815 181.645 76.105 181.690 ;
        RECT 80.875 181.830 81.165 181.875 ;
        RECT 88.220 181.830 88.540 181.890 ;
        RECT 80.875 181.690 88.540 181.830 ;
        RECT 80.875 181.645 81.165 181.690 ;
        RECT 88.220 181.630 88.540 181.690 ;
        RECT 94.675 181.645 94.965 181.875 ;
        RECT 107.080 181.830 107.400 181.890 ;
        RECT 102.110 181.690 107.400 181.830 ;
        RECT 41.850 181.350 49.350 181.490 ;
        RECT 59.815 181.490 60.105 181.535 ;
        RECT 63.055 181.490 63.705 181.535 ;
        RECT 59.815 181.350 63.705 181.490 ;
        RECT 33.595 181.150 33.885 181.195 ;
        RECT 37.175 181.150 37.465 181.195 ;
        RECT 39.010 181.150 39.300 181.195 ;
        RECT 33.595 181.010 39.300 181.150 ;
        RECT 33.595 180.965 33.885 181.010 ;
        RECT 37.175 180.965 37.465 181.010 ;
        RECT 39.010 180.965 39.300 181.010 ;
        RECT 39.920 180.950 40.240 181.210 ;
        RECT 41.850 181.195 41.990 181.350 ;
        RECT 59.815 181.305 60.405 181.350 ;
        RECT 63.055 181.305 63.705 181.350 ;
        RECT 41.775 180.965 42.065 181.195 ;
        RECT 46.375 180.965 46.665 181.195 ;
        RECT 46.835 180.965 47.125 181.195 ;
        RECT 29.815 180.810 30.105 180.855 ;
        RECT 37.620 180.810 37.940 180.870 ;
        RECT 29.815 180.670 37.940 180.810 ;
        RECT 29.815 180.625 30.105 180.670 ;
        RECT 37.620 180.610 37.940 180.670 ;
        RECT 38.080 180.810 38.400 180.870 ;
        RECT 39.475 180.810 39.765 180.855 ;
        RECT 43.600 180.810 43.920 180.870 ;
        RECT 38.080 180.670 43.920 180.810 ;
        RECT 38.080 180.610 38.400 180.670 ;
        RECT 39.475 180.625 39.765 180.670 ;
        RECT 43.600 180.610 43.920 180.670 ;
        RECT 44.980 180.610 45.300 180.870 ;
        RECT 33.595 180.470 33.885 180.515 ;
        RECT 36.715 180.470 37.005 180.515 ;
        RECT 38.605 180.470 38.895 180.515 ;
        RECT 33.595 180.330 38.895 180.470 ;
        RECT 33.595 180.285 33.885 180.330 ;
        RECT 36.715 180.285 37.005 180.330 ;
        RECT 38.605 180.285 38.895 180.330 ;
        RECT 35.320 180.130 35.640 180.190 ;
        RECT 38.160 180.130 38.450 180.175 ;
        RECT 35.320 179.990 38.450 180.130 ;
        RECT 46.450 180.130 46.590 180.965 ;
        RECT 46.910 180.810 47.050 180.965 ;
        RECT 47.280 180.950 47.600 181.210 ;
        RECT 48.200 180.950 48.520 181.210 ;
        RECT 49.135 181.150 49.425 181.195 ;
        RECT 49.580 181.150 49.900 181.210 ;
        RECT 60.115 181.150 60.405 181.305 ;
        RECT 65.680 181.290 66.000 181.550 ;
        RECT 67.060 181.490 67.380 181.550 ;
        RECT 70.755 181.490 71.045 181.535 ;
        RECT 67.060 181.350 71.045 181.490 ;
        RECT 67.060 181.290 67.380 181.350 ;
        RECT 68.070 181.195 68.210 181.350 ;
        RECT 70.755 181.305 71.045 181.350 ;
        RECT 71.200 181.490 71.520 181.550 ;
        RECT 72.580 181.490 72.900 181.550 ;
        RECT 81.320 181.490 81.640 181.550 ;
        RECT 86.395 181.490 86.685 181.535 ;
        RECT 86.840 181.490 87.160 181.550 ;
        RECT 71.200 181.350 72.350 181.490 ;
        RECT 71.200 181.290 71.520 181.350 ;
        RECT 49.135 181.010 49.900 181.150 ;
        RECT 49.135 180.965 49.425 181.010 ;
        RECT 49.580 180.950 49.900 181.010 ;
        RECT 56.800 181.010 60.405 181.150 ;
        RECT 50.500 180.810 50.820 180.870 ;
        RECT 46.910 180.670 50.820 180.810 ;
        RECT 50.500 180.610 50.820 180.670 ;
        RECT 52.340 180.810 52.660 180.870 ;
        RECT 56.800 180.810 56.940 181.010 ;
        RECT 60.115 180.990 60.405 181.010 ;
        RECT 61.195 181.150 61.485 181.195 ;
        RECT 64.775 181.150 65.065 181.195 ;
        RECT 66.610 181.150 66.900 181.195 ;
        RECT 61.195 181.010 66.900 181.150 ;
        RECT 61.195 180.965 61.485 181.010 ;
        RECT 64.775 180.965 65.065 181.010 ;
        RECT 66.610 180.965 66.900 181.010 ;
        RECT 67.995 180.965 68.285 181.195 ;
        RECT 69.835 180.965 70.125 181.195 ;
        RECT 70.280 181.150 70.600 181.210 ;
        RECT 72.210 181.195 72.350 181.350 ;
        RECT 72.580 181.350 73.270 181.490 ;
        RECT 72.580 181.290 72.900 181.350 ;
        RECT 73.130 181.195 73.270 181.350 ;
        RECT 75.890 181.350 80.170 181.490 ;
        RECT 75.890 181.210 76.030 181.350 ;
        RECT 71.675 181.150 71.965 181.195 ;
        RECT 70.280 181.010 71.965 181.150 ;
        RECT 52.340 180.670 56.940 180.810 ;
        RECT 57.400 180.810 57.720 180.870 ;
        RECT 65.220 180.810 65.540 180.870 ;
        RECT 57.400 180.670 66.830 180.810 ;
        RECT 52.340 180.610 52.660 180.670 ;
        RECT 57.400 180.610 57.720 180.670 ;
        RECT 65.220 180.610 65.540 180.670 ;
        RECT 56.020 180.470 56.340 180.530 ;
        RECT 52.430 180.330 56.340 180.470 ;
        RECT 52.430 180.130 52.570 180.330 ;
        RECT 56.020 180.270 56.340 180.330 ;
        RECT 61.195 180.470 61.485 180.515 ;
        RECT 64.315 180.470 64.605 180.515 ;
        RECT 66.205 180.470 66.495 180.515 ;
        RECT 61.195 180.330 66.495 180.470 ;
        RECT 66.690 180.470 66.830 180.670 ;
        RECT 67.060 180.610 67.380 180.870 ;
        RECT 68.455 180.810 68.745 180.855 ;
        RECT 67.610 180.670 68.745 180.810 ;
        RECT 67.610 180.470 67.750 180.670 ;
        RECT 68.455 180.625 68.745 180.670 ;
        RECT 69.375 180.625 69.665 180.855 ;
        RECT 69.910 180.810 70.050 180.965 ;
        RECT 70.280 180.950 70.600 181.010 ;
        RECT 71.675 180.965 71.965 181.010 ;
        RECT 72.135 180.965 72.425 181.195 ;
        RECT 73.055 180.965 73.345 181.195 ;
        RECT 74.420 181.150 74.740 181.210 ;
        RECT 74.895 181.150 75.185 181.195 ;
        RECT 74.420 181.010 75.185 181.150 ;
        RECT 74.420 180.950 74.740 181.010 ;
        RECT 74.895 180.965 75.185 181.010 ;
        RECT 75.800 180.950 76.120 181.210 ;
        RECT 79.035 181.150 79.325 181.195 ;
        RECT 79.480 181.150 79.800 181.210 ;
        RECT 79.035 181.010 79.800 181.150 ;
        RECT 80.030 181.150 80.170 181.350 ;
        RECT 81.320 181.350 83.850 181.490 ;
        RECT 81.320 181.290 81.640 181.350 ;
        RECT 80.030 181.010 82.470 181.150 ;
        RECT 79.035 180.965 79.325 181.010 ;
        RECT 79.480 180.950 79.800 181.010 ;
        RECT 70.740 180.810 71.060 180.870 ;
        RECT 72.595 180.810 72.885 180.855 ;
        RECT 69.910 180.670 70.510 180.810 ;
        RECT 66.690 180.330 67.750 180.470 ;
        RECT 61.195 180.285 61.485 180.330 ;
        RECT 64.315 180.285 64.605 180.330 ;
        RECT 66.205 180.285 66.495 180.330 ;
        RECT 46.450 179.990 52.570 180.130 ;
        RECT 53.720 180.130 54.040 180.190 ;
        RECT 55.575 180.130 55.865 180.175 ;
        RECT 67.060 180.130 67.380 180.190 ;
        RECT 53.720 179.990 67.380 180.130 ;
        RECT 69.450 180.130 69.590 180.625 ;
        RECT 70.370 180.470 70.510 180.670 ;
        RECT 70.740 180.670 72.885 180.810 ;
        RECT 70.740 180.610 71.060 180.670 ;
        RECT 72.595 180.625 72.885 180.670 ;
        RECT 76.720 180.810 77.040 180.870 ;
        RECT 77.655 180.810 77.945 180.855 ;
        RECT 76.720 180.670 77.945 180.810 ;
        RECT 76.720 180.610 77.040 180.670 ;
        RECT 77.655 180.625 77.945 180.670 ;
        RECT 78.575 180.625 78.865 180.855 ;
        RECT 73.040 180.470 73.360 180.530 ;
        RECT 76.810 180.470 76.950 180.610 ;
        RECT 70.370 180.330 71.890 180.470 ;
        RECT 71.200 180.130 71.520 180.190 ;
        RECT 69.450 179.990 71.520 180.130 ;
        RECT 71.750 180.130 71.890 180.330 ;
        RECT 73.040 180.330 76.950 180.470 ;
        RECT 78.650 180.470 78.790 180.625 ;
        RECT 81.320 180.610 81.640 180.870 ;
        RECT 82.330 180.810 82.470 181.010 ;
        RECT 82.700 180.950 83.020 181.210 ;
        RECT 83.710 181.195 83.850 181.350 ;
        RECT 86.395 181.350 87.160 181.490 ;
        RECT 86.395 181.305 86.685 181.350 ;
        RECT 86.840 181.290 87.160 181.350 ;
        RECT 88.675 181.490 89.325 181.535 ;
        RECT 92.275 181.490 92.565 181.535 ;
        RECT 94.200 181.490 94.520 181.550 ;
        RECT 88.675 181.350 94.520 181.490 ;
        RECT 88.675 181.305 89.325 181.350 ;
        RECT 91.975 181.305 92.565 181.350 ;
        RECT 83.175 180.965 83.465 181.195 ;
        RECT 83.635 180.965 83.925 181.195 ;
        RECT 83.250 180.810 83.390 180.965 ;
        RECT 84.540 180.950 84.860 181.210 ;
        RECT 85.000 180.950 85.320 181.210 ;
        RECT 85.480 181.150 85.770 181.195 ;
        RECT 87.315 181.150 87.605 181.195 ;
        RECT 90.895 181.150 91.185 181.195 ;
        RECT 85.480 181.010 91.185 181.150 ;
        RECT 85.480 180.965 85.770 181.010 ;
        RECT 87.315 180.965 87.605 181.010 ;
        RECT 90.895 180.965 91.185 181.010 ;
        RECT 91.975 180.990 92.265 181.305 ;
        RECT 94.200 181.290 94.520 181.350 ;
        RECT 94.750 181.150 94.890 181.645 ;
        RECT 101.560 181.290 101.880 181.550 ;
        RECT 92.450 181.010 94.890 181.150 ;
        RECT 82.330 180.670 83.390 180.810 ;
        RECT 84.630 180.810 84.770 180.950 ;
        RECT 92.450 180.810 92.590 181.010 ;
        RECT 95.580 180.950 95.900 181.210 ;
        RECT 96.500 181.150 96.820 181.210 ;
        RECT 97.895 181.150 98.185 181.195 ;
        RECT 96.500 181.010 98.185 181.150 ;
        RECT 96.500 180.950 96.820 181.010 ;
        RECT 97.895 180.965 98.185 181.010 ;
        RECT 98.355 181.150 98.645 181.195 ;
        RECT 102.110 181.150 102.250 181.690 ;
        RECT 107.080 181.630 107.400 181.690 ;
        RECT 106.620 181.535 106.940 181.550 ;
        RECT 106.155 181.490 106.940 181.535 ;
        RECT 109.755 181.490 110.045 181.535 ;
        RECT 106.155 181.350 110.045 181.490 ;
        RECT 106.155 181.305 106.940 181.350 ;
        RECT 106.620 181.290 106.940 181.305 ;
        RECT 109.455 181.305 110.045 181.350 ;
        RECT 98.355 181.010 102.250 181.150 ;
        RECT 102.960 181.150 103.250 181.195 ;
        RECT 104.795 181.150 105.085 181.195 ;
        RECT 108.375 181.150 108.665 181.195 ;
        RECT 102.960 181.010 108.665 181.150 ;
        RECT 98.355 180.965 98.645 181.010 ;
        RECT 102.960 180.965 103.250 181.010 ;
        RECT 104.795 180.965 105.085 181.010 ;
        RECT 108.375 180.965 108.665 181.010 ;
        RECT 109.455 180.990 109.745 181.305 ;
        RECT 84.630 180.670 92.590 180.810 ;
        RECT 93.755 180.810 94.045 180.855 ;
        RECT 96.040 180.810 96.360 180.870 ;
        RECT 93.755 180.670 96.360 180.810 ;
        RECT 93.755 180.625 94.045 180.670 ;
        RECT 96.040 180.610 96.360 180.670 ;
        RECT 97.420 180.810 97.740 180.870 ;
        RECT 98.815 180.810 99.105 180.855 ;
        RECT 102.495 180.810 102.785 180.855 ;
        RECT 105.700 180.810 106.020 180.870 ;
        RECT 111.220 180.810 111.540 180.870 ;
        RECT 97.420 180.670 99.105 180.810 ;
        RECT 97.420 180.610 97.740 180.670 ;
        RECT 98.815 180.625 99.105 180.670 ;
        RECT 99.350 180.670 111.540 180.810 ;
        RECT 81.780 180.470 82.100 180.530 ;
        RECT 78.650 180.330 82.100 180.470 ;
        RECT 73.040 180.270 73.360 180.330 ;
        RECT 81.780 180.270 82.100 180.330 ;
        RECT 85.885 180.470 86.175 180.515 ;
        RECT 87.775 180.470 88.065 180.515 ;
        RECT 90.895 180.470 91.185 180.515 ;
        RECT 85.885 180.330 91.185 180.470 ;
        RECT 85.885 180.285 86.175 180.330 ;
        RECT 87.775 180.285 88.065 180.330 ;
        RECT 90.895 180.285 91.185 180.330 ;
        RECT 94.660 180.470 94.980 180.530 ;
        RECT 99.350 180.470 99.490 180.670 ;
        RECT 102.495 180.625 102.785 180.670 ;
        RECT 105.700 180.610 106.020 180.670 ;
        RECT 111.220 180.610 111.540 180.670 ;
        RECT 94.660 180.330 99.490 180.470 ;
        RECT 94.660 180.270 94.980 180.330 ;
        RECT 100.640 180.270 100.960 180.530 ;
        RECT 103.365 180.470 103.655 180.515 ;
        RECT 105.255 180.470 105.545 180.515 ;
        RECT 108.375 180.470 108.665 180.515 ;
        RECT 103.365 180.330 108.665 180.470 ;
        RECT 103.365 180.285 103.655 180.330 ;
        RECT 105.255 180.285 105.545 180.330 ;
        RECT 108.375 180.285 108.665 180.330 ;
        RECT 73.960 180.130 74.280 180.190 ;
        RECT 71.750 179.990 74.280 180.130 ;
        RECT 35.320 179.930 35.640 179.990 ;
        RECT 38.160 179.945 38.450 179.990 ;
        RECT 53.720 179.930 54.040 179.990 ;
        RECT 55.575 179.945 55.865 179.990 ;
        RECT 67.060 179.930 67.380 179.990 ;
        RECT 71.200 179.930 71.520 179.990 ;
        RECT 73.960 179.930 74.280 179.990 ;
        RECT 74.880 180.130 75.200 180.190 ;
        RECT 82.700 180.130 83.020 180.190 ;
        RECT 74.880 179.990 83.020 180.130 ;
        RECT 74.880 179.930 75.200 179.990 ;
        RECT 82.700 179.930 83.020 179.990 ;
        RECT 88.220 180.130 88.540 180.190 ;
        RECT 96.055 180.130 96.345 180.175 ;
        RECT 88.220 179.990 96.345 180.130 ;
        RECT 88.220 179.930 88.540 179.990 ;
        RECT 96.055 179.945 96.345 179.990 ;
        RECT 101.100 180.130 101.420 180.190 ;
        RECT 103.785 180.130 104.075 180.175 ;
        RECT 101.100 179.990 104.075 180.130 ;
        RECT 101.100 179.930 101.420 179.990 ;
        RECT 103.785 179.945 104.075 179.990 ;
        RECT 104.320 180.130 104.640 180.190 ;
        RECT 111.235 180.130 111.525 180.175 ;
        RECT 104.320 179.990 111.525 180.130 ;
        RECT 104.320 179.930 104.640 179.990 ;
        RECT 111.235 179.945 111.525 179.990 ;
        RECT 26.970 179.310 113.450 179.790 ;
        RECT 30.735 179.110 31.025 179.155 ;
        RECT 39.460 179.110 39.780 179.170 ;
        RECT 30.735 178.970 39.780 179.110 ;
        RECT 30.735 178.925 31.025 178.970 ;
        RECT 39.460 178.910 39.780 178.970 ;
        RECT 40.380 179.110 40.700 179.170 ;
        RECT 46.360 179.110 46.680 179.170 ;
        RECT 40.380 178.970 46.680 179.110 ;
        RECT 40.380 178.910 40.700 178.970 ;
        RECT 46.360 178.910 46.680 178.970 ;
        RECT 50.500 179.110 50.820 179.170 ;
        RECT 51.895 179.110 52.185 179.155 ;
        RECT 50.500 178.970 52.185 179.110 ;
        RECT 50.500 178.910 50.820 178.970 ;
        RECT 51.895 178.925 52.185 178.970 ;
        RECT 55.560 179.110 55.880 179.170 ;
        RECT 63.380 179.110 63.700 179.170 ;
        RECT 55.560 178.970 63.700 179.110 ;
        RECT 28.420 178.770 28.740 178.830 ;
        RECT 31.655 178.770 31.945 178.815 ;
        RECT 28.420 178.630 31.945 178.770 ;
        RECT 28.420 178.570 28.740 178.630 ;
        RECT 31.655 178.585 31.945 178.630 ;
        RECT 36.700 178.770 37.020 178.830 ;
        RECT 46.835 178.770 47.125 178.815 ;
        RECT 36.700 178.630 47.125 178.770 ;
        RECT 36.700 178.570 37.020 178.630 ;
        RECT 46.835 178.585 47.125 178.630 ;
        RECT 32.100 178.430 32.420 178.490 ;
        RECT 34.415 178.430 34.705 178.475 ;
        RECT 32.100 178.290 34.705 178.430 ;
        RECT 32.100 178.230 32.420 178.290 ;
        RECT 34.415 178.245 34.705 178.290 ;
        RECT 38.555 178.430 38.845 178.475 ;
        RECT 45.900 178.430 46.220 178.490 ;
        RECT 38.555 178.290 46.220 178.430 ;
        RECT 51.970 178.430 52.110 178.925 ;
        RECT 55.560 178.910 55.880 178.970 ;
        RECT 51.970 178.290 58.090 178.430 ;
        RECT 38.555 178.245 38.845 178.290 ;
        RECT 45.900 178.230 46.220 178.290 ;
        RECT 28.880 177.890 29.200 178.150 ;
        RECT 30.275 177.905 30.565 178.135 ;
        RECT 35.320 178.090 35.640 178.150 ;
        RECT 32.650 177.950 35.640 178.090 ;
        RECT 26.120 177.750 26.440 177.810 ;
        RECT 27.040 177.750 27.360 177.810 ;
        RECT 30.350 177.750 30.490 177.905 ;
        RECT 26.120 177.610 30.490 177.750 ;
        RECT 26.120 177.550 26.440 177.610 ;
        RECT 27.040 177.550 27.360 177.610 ;
        RECT 29.815 177.410 30.105 177.455 ;
        RECT 32.650 177.410 32.790 177.950 ;
        RECT 35.320 177.890 35.640 177.950 ;
        RECT 36.715 177.905 37.005 178.135 ;
        RECT 37.620 178.090 37.940 178.150 ;
        RECT 38.095 178.090 38.385 178.135 ;
        RECT 37.620 177.950 38.385 178.090 ;
        RECT 33.955 177.750 34.245 177.795 ;
        RECT 35.780 177.750 36.100 177.810 ;
        RECT 33.955 177.610 36.100 177.750 ;
        RECT 36.790 177.750 36.930 177.905 ;
        RECT 37.620 177.890 37.940 177.950 ;
        RECT 38.095 177.905 38.385 177.950 ;
        RECT 39.475 177.905 39.765 178.135 ;
        RECT 38.540 177.750 38.860 177.810 ;
        RECT 36.790 177.610 38.860 177.750 ;
        RECT 33.955 177.565 34.245 177.610 ;
        RECT 35.780 177.550 36.100 177.610 ;
        RECT 38.540 177.550 38.860 177.610 ;
        RECT 29.815 177.270 32.790 177.410 ;
        RECT 33.495 177.410 33.785 177.455 ;
        RECT 34.860 177.410 35.180 177.470 ;
        RECT 33.495 177.270 35.180 177.410 ;
        RECT 29.815 177.225 30.105 177.270 ;
        RECT 33.495 177.225 33.785 177.270 ;
        RECT 34.860 177.210 35.180 177.270 ;
        RECT 37.620 177.210 37.940 177.470 ;
        RECT 39.550 177.410 39.690 177.905 ;
        RECT 40.380 177.890 40.700 178.150 ;
        RECT 40.840 177.890 41.160 178.150 ;
        RECT 41.315 177.905 41.605 178.135 ;
        RECT 42.220 178.090 42.540 178.150 ;
        RECT 43.155 178.090 43.445 178.135 ;
        RECT 42.220 177.950 43.445 178.090 ;
        RECT 39.920 177.750 40.240 177.810 ;
        RECT 41.390 177.750 41.530 177.905 ;
        RECT 42.220 177.890 42.540 177.950 ;
        RECT 43.155 177.905 43.445 177.950 ;
        RECT 43.600 178.090 43.920 178.150 ;
        RECT 44.075 178.090 44.365 178.135 ;
        RECT 43.600 177.950 44.365 178.090 ;
        RECT 43.600 177.890 43.920 177.950 ;
        RECT 44.075 177.905 44.365 177.950 ;
        RECT 44.520 177.890 44.840 178.150 ;
        RECT 44.995 177.905 45.285 178.135 ;
        RECT 50.055 178.090 50.345 178.135 ;
        RECT 50.055 177.950 51.650 178.090 ;
        RECT 50.055 177.905 50.345 177.950 ;
        RECT 45.070 177.750 45.210 177.905 ;
        RECT 39.920 177.610 41.530 177.750 ;
        RECT 44.610 177.610 45.210 177.750 ;
        RECT 39.920 177.550 40.240 177.610 ;
        RECT 44.610 177.470 44.750 177.610 ;
        RECT 41.300 177.410 41.620 177.470 ;
        RECT 39.550 177.270 41.620 177.410 ;
        RECT 41.300 177.210 41.620 177.270 ;
        RECT 42.680 177.210 43.000 177.470 ;
        RECT 44.520 177.210 44.840 177.470 ;
        RECT 46.375 177.410 46.665 177.455 ;
        RECT 46.820 177.410 47.140 177.470 ;
        RECT 46.375 177.270 47.140 177.410 ;
        RECT 51.510 177.410 51.650 177.950 ;
        RECT 52.815 177.905 53.105 178.135 ;
        RECT 52.890 177.750 53.030 177.905 ;
        RECT 53.720 177.890 54.040 178.150 ;
        RECT 57.400 177.750 57.720 177.810 ;
        RECT 52.890 177.610 57.720 177.750 ;
        RECT 57.950 177.750 58.090 178.290 ;
        RECT 58.410 178.090 58.550 178.970 ;
        RECT 63.380 178.910 63.700 178.970 ;
        RECT 63.840 179.110 64.160 179.170 ;
        RECT 71.660 179.110 71.980 179.170 ;
        RECT 63.840 178.970 71.980 179.110 ;
        RECT 63.840 178.910 64.160 178.970 ;
        RECT 71.660 178.910 71.980 178.970 ;
        RECT 73.040 178.910 73.360 179.170 ;
        RECT 74.435 179.110 74.725 179.155 ;
        RECT 74.880 179.110 75.200 179.170 ;
        RECT 74.435 178.970 75.200 179.110 ;
        RECT 74.435 178.925 74.725 178.970 ;
        RECT 74.880 178.910 75.200 178.970 ;
        RECT 79.035 179.110 79.325 179.155 ;
        RECT 85.000 179.110 85.320 179.170 ;
        RECT 94.660 179.110 94.980 179.170 ;
        RECT 79.035 178.970 85.320 179.110 ;
        RECT 79.035 178.925 79.325 178.970 ;
        RECT 85.000 178.910 85.320 178.970 ;
        RECT 91.070 178.970 94.980 179.110 ;
        RECT 61.080 178.770 61.400 178.830 ;
        RECT 80.400 178.770 80.720 178.830 ;
        RECT 61.080 178.630 80.720 178.770 ;
        RECT 61.080 178.570 61.400 178.630 ;
        RECT 58.780 178.430 59.100 178.490 ;
        RECT 58.780 178.290 64.530 178.430 ;
        RECT 58.780 178.230 59.100 178.290 ;
        RECT 59.255 178.090 59.545 178.135 ;
        RECT 58.410 177.950 59.545 178.090 ;
        RECT 59.255 177.905 59.545 177.950 ;
        RECT 59.715 177.905 60.005 178.135 ;
        RECT 60.175 178.090 60.465 178.135 ;
        RECT 60.620 178.090 60.940 178.150 ;
        RECT 60.175 177.950 60.940 178.090 ;
        RECT 60.175 177.905 60.465 177.950 ;
        RECT 59.790 177.750 59.930 177.905 ;
        RECT 60.620 177.890 60.940 177.950 ;
        RECT 61.080 177.890 61.400 178.150 ;
        RECT 63.380 177.890 63.700 178.150 ;
        RECT 63.840 177.890 64.160 178.150 ;
        RECT 64.390 178.135 64.530 178.290 ;
        RECT 64.315 177.905 64.605 178.135 ;
        RECT 64.850 178.090 64.990 178.630 ;
        RECT 80.400 178.570 80.720 178.630 ;
        RECT 71.660 178.430 71.980 178.490 ;
        RECT 75.800 178.430 76.120 178.490 ;
        RECT 91.070 178.475 91.210 178.970 ;
        RECT 94.660 178.910 94.980 178.970 ;
        RECT 98.800 179.110 99.120 179.170 ;
        RECT 101.115 179.110 101.405 179.155 ;
        RECT 98.800 178.970 101.405 179.110 ;
        RECT 98.800 178.910 99.120 178.970 ;
        RECT 101.115 178.925 101.405 178.970 ;
        RECT 91.865 178.770 92.155 178.815 ;
        RECT 93.755 178.770 94.045 178.815 ;
        RECT 96.875 178.770 97.165 178.815 ;
        RECT 91.865 178.630 97.165 178.770 ;
        RECT 91.865 178.585 92.155 178.630 ;
        RECT 93.755 178.585 94.045 178.630 ;
        RECT 96.875 178.585 97.165 178.630 ;
        RECT 99.735 178.770 100.025 178.815 ;
        RECT 103.400 178.770 103.720 178.830 ;
        RECT 99.735 178.630 103.720 178.770 ;
        RECT 99.735 178.585 100.025 178.630 ;
        RECT 103.400 178.570 103.720 178.630 ;
        RECT 105.355 178.770 105.645 178.815 ;
        RECT 108.475 178.770 108.765 178.815 ;
        RECT 110.365 178.770 110.655 178.815 ;
        RECT 105.355 178.630 110.655 178.770 ;
        RECT 105.355 178.585 105.645 178.630 ;
        RECT 108.475 178.585 108.765 178.630 ;
        RECT 110.365 178.585 110.655 178.630 ;
        RECT 71.660 178.290 76.120 178.430 ;
        RECT 71.660 178.230 71.980 178.290 ;
        RECT 75.800 178.230 76.120 178.290 ;
        RECT 90.995 178.245 91.285 178.475 ;
        RECT 92.375 178.430 92.665 178.475 ;
        RECT 109.380 178.430 109.700 178.490 ;
        RECT 92.375 178.290 109.700 178.430 ;
        RECT 92.375 178.245 92.665 178.290 ;
        RECT 65.235 178.090 65.525 178.135 ;
        RECT 64.850 177.950 65.525 178.090 ;
        RECT 65.235 177.905 65.525 177.950 ;
        RECT 67.075 177.905 67.365 178.135 ;
        RECT 63.930 177.750 64.070 177.890 ;
        RECT 67.150 177.750 67.290 177.905 ;
        RECT 67.520 177.890 67.840 178.150 ;
        RECT 67.980 177.890 68.300 178.150 ;
        RECT 68.440 178.090 68.760 178.150 ;
        RECT 68.915 178.090 69.205 178.135 ;
        RECT 68.440 177.950 69.205 178.090 ;
        RECT 68.440 177.890 68.760 177.950 ;
        RECT 68.915 177.905 69.205 177.950 ;
        RECT 70.755 178.090 71.045 178.135 ;
        RECT 72.580 178.090 72.900 178.150 ;
        RECT 74.420 178.090 74.740 178.150 ;
        RECT 70.755 177.950 74.740 178.090 ;
        RECT 70.755 177.905 71.045 177.950 ;
        RECT 72.580 177.890 72.900 177.950 ;
        RECT 74.420 177.890 74.740 177.950 ;
        RECT 75.355 178.090 75.645 178.135 ;
        RECT 76.260 178.090 76.580 178.150 ;
        RECT 75.355 177.950 86.610 178.090 ;
        RECT 75.355 177.905 75.645 177.950 ;
        RECT 57.950 177.610 64.070 177.750 ;
        RECT 65.310 177.610 67.290 177.750 ;
        RECT 57.400 177.550 57.720 177.610 ;
        RECT 52.800 177.410 53.120 177.470 ;
        RECT 51.510 177.270 53.120 177.410 ;
        RECT 46.375 177.225 46.665 177.270 ;
        RECT 46.820 177.210 47.140 177.270 ;
        RECT 52.800 177.210 53.120 177.270 ;
        RECT 57.860 177.210 58.180 177.470 ;
        RECT 60.160 177.410 60.480 177.470 ;
        RECT 62.015 177.410 62.305 177.455 ;
        RECT 60.160 177.270 62.305 177.410 ;
        RECT 60.160 177.210 60.480 177.270 ;
        RECT 62.015 177.225 62.305 177.270 ;
        RECT 62.460 177.410 62.780 177.470 ;
        RECT 65.310 177.410 65.450 177.610 ;
        RECT 71.660 177.550 71.980 177.810 ;
        RECT 73.960 177.750 74.280 177.810 ;
        RECT 75.430 177.750 75.570 177.905 ;
        RECT 76.260 177.890 76.580 177.950 ;
        RECT 73.960 177.610 75.570 177.750 ;
        RECT 85.475 177.750 85.765 177.795 ;
        RECT 85.920 177.750 86.240 177.810 ;
        RECT 85.475 177.610 86.240 177.750 ;
        RECT 86.470 177.750 86.610 177.950 ;
        RECT 86.840 177.890 87.160 178.150 ;
        RECT 90.075 178.090 90.365 178.135 ;
        RECT 91.070 178.090 91.210 178.245 ;
        RECT 109.380 178.230 109.700 178.290 ;
        RECT 111.220 178.230 111.540 178.490 ;
        RECT 90.075 177.950 91.210 178.090 ;
        RECT 91.460 178.090 91.750 178.135 ;
        RECT 93.295 178.090 93.585 178.135 ;
        RECT 96.875 178.090 97.165 178.135 ;
        RECT 91.460 177.950 97.165 178.090 ;
        RECT 90.075 177.905 90.365 177.950 ;
        RECT 91.460 177.905 91.750 177.950 ;
        RECT 93.295 177.905 93.585 177.950 ;
        RECT 96.875 177.905 97.165 177.950 ;
        RECT 97.880 178.110 98.200 178.150 ;
        RECT 97.880 177.890 98.245 178.110 ;
        RECT 100.195 178.090 100.485 178.135 ;
        RECT 104.320 178.110 104.640 178.150 ;
        RECT 97.955 177.795 98.245 177.890 ;
        RECT 98.890 177.950 100.485 178.090 ;
        RECT 94.655 177.750 95.305 177.795 ;
        RECT 97.955 177.750 98.545 177.795 ;
        RECT 86.470 177.610 94.430 177.750 ;
        RECT 73.960 177.550 74.280 177.610 ;
        RECT 85.475 177.565 85.765 177.610 ;
        RECT 85.920 177.550 86.240 177.610 ;
        RECT 62.460 177.270 65.450 177.410 ;
        RECT 62.460 177.210 62.780 177.270 ;
        RECT 65.680 177.210 66.000 177.470 ;
        RECT 69.820 177.210 70.140 177.470 ;
        RECT 70.740 177.410 71.060 177.470 ;
        RECT 74.050 177.410 74.190 177.550 ;
        RECT 70.740 177.270 74.190 177.410 ;
        RECT 80.400 177.410 80.720 177.470 ;
        RECT 86.395 177.410 86.685 177.455 ;
        RECT 80.400 177.270 86.685 177.410 ;
        RECT 94.290 177.410 94.430 177.610 ;
        RECT 94.655 177.610 98.545 177.750 ;
        RECT 94.655 177.565 95.305 177.610 ;
        RECT 98.255 177.565 98.545 177.610 ;
        RECT 95.580 177.410 95.900 177.470 ;
        RECT 98.890 177.410 99.030 177.950 ;
        RECT 100.195 177.905 100.485 177.950 ;
        RECT 104.275 177.890 104.640 178.110 ;
        RECT 105.355 178.090 105.645 178.135 ;
        RECT 108.935 178.090 109.225 178.135 ;
        RECT 110.770 178.090 111.060 178.135 ;
        RECT 105.355 177.950 111.060 178.090 ;
        RECT 105.355 177.905 105.645 177.950 ;
        RECT 108.935 177.905 109.225 177.950 ;
        RECT 110.770 177.905 111.060 177.950 ;
        RECT 104.275 177.795 104.565 177.890 ;
        RECT 103.975 177.750 104.565 177.795 ;
        RECT 107.215 177.750 107.865 177.795 ;
        RECT 103.975 177.610 107.865 177.750 ;
        RECT 103.975 177.565 104.265 177.610 ;
        RECT 107.215 177.565 107.865 177.610 ;
        RECT 109.840 177.550 110.160 177.810 ;
        RECT 94.290 177.270 99.030 177.410 ;
        RECT 100.180 177.410 100.500 177.470 ;
        RECT 102.495 177.410 102.785 177.455 ;
        RECT 104.780 177.410 105.100 177.470 ;
        RECT 100.180 177.270 105.100 177.410 ;
        RECT 70.740 177.210 71.060 177.270 ;
        RECT 80.400 177.210 80.720 177.270 ;
        RECT 86.395 177.225 86.685 177.270 ;
        RECT 95.580 177.210 95.900 177.270 ;
        RECT 100.180 177.210 100.500 177.270 ;
        RECT 102.495 177.225 102.785 177.270 ;
        RECT 104.780 177.210 105.100 177.270 ;
        RECT 26.970 176.590 113.450 177.070 ;
        RECT 30.720 176.390 31.040 176.450 ;
        RECT 47.755 176.390 48.045 176.435 ;
        RECT 52.340 176.390 52.660 176.450 ;
        RECT 71.660 176.390 71.980 176.450 ;
        RECT 30.720 176.250 31.870 176.390 ;
        RECT 30.720 176.190 31.040 176.250 ;
        RECT 29.360 176.050 29.650 176.095 ;
        RECT 31.220 176.050 31.510 176.095 ;
        RECT 29.360 175.910 31.510 176.050 ;
        RECT 31.730 176.050 31.870 176.250 ;
        RECT 47.755 176.250 52.660 176.390 ;
        RECT 47.755 176.205 48.045 176.250 ;
        RECT 52.340 176.190 52.660 176.250 ;
        RECT 70.830 176.250 71.980 176.390 ;
        RECT 32.140 176.050 32.430 176.095 ;
        RECT 35.400 176.050 35.690 176.095 ;
        RECT 31.730 175.910 35.690 176.050 ;
        RECT 29.360 175.865 29.650 175.910 ;
        RECT 31.220 175.865 31.510 175.910 ;
        RECT 32.140 175.865 32.430 175.910 ;
        RECT 35.400 175.865 35.690 175.910 ;
        RECT 36.240 176.050 36.560 176.110 ;
        RECT 39.475 176.050 39.765 176.095 ;
        RECT 36.240 175.910 39.765 176.050 ;
        RECT 29.800 175.710 30.120 175.770 ;
        RECT 30.275 175.710 30.565 175.755 ;
        RECT 29.800 175.570 30.565 175.710 ;
        RECT 31.295 175.710 31.510 175.865 ;
        RECT 36.240 175.850 36.560 175.910 ;
        RECT 39.475 175.865 39.765 175.910 ;
        RECT 41.755 176.050 42.405 176.095 ;
        RECT 43.140 176.050 43.460 176.110 ;
        RECT 45.355 176.050 45.645 176.095 ;
        RECT 41.755 175.910 45.645 176.050 ;
        RECT 41.755 175.865 42.405 175.910 ;
        RECT 43.140 175.850 43.460 175.910 ;
        RECT 45.055 175.865 45.645 175.910 ;
        RECT 45.900 176.050 46.220 176.110 ;
        RECT 58.435 176.050 58.725 176.095 ;
        RECT 61.675 176.050 62.325 176.095 ;
        RECT 45.900 175.910 62.325 176.050 ;
        RECT 33.540 175.710 33.830 175.755 ;
        RECT 31.295 175.570 33.830 175.710 ;
        RECT 29.800 175.510 30.120 175.570 ;
        RECT 30.275 175.525 30.565 175.570 ;
        RECT 33.540 175.525 33.830 175.570 ;
        RECT 38.560 175.710 38.850 175.755 ;
        RECT 40.395 175.710 40.685 175.755 ;
        RECT 43.975 175.710 44.265 175.755 ;
        RECT 38.560 175.570 44.265 175.710 ;
        RECT 38.560 175.525 38.850 175.570 ;
        RECT 40.395 175.525 40.685 175.570 ;
        RECT 43.975 175.525 44.265 175.570 ;
        RECT 45.055 175.550 45.345 175.865 ;
        RECT 45.900 175.850 46.220 175.910 ;
        RECT 58.435 175.865 59.025 175.910 ;
        RECT 61.675 175.865 62.325 175.910 ;
        RECT 64.315 176.050 64.605 176.095 ;
        RECT 64.760 176.050 65.080 176.110 ;
        RECT 70.830 176.095 70.970 176.250 ;
        RECT 71.660 176.190 71.980 176.250 ;
        RECT 82.240 176.390 82.560 176.450 ;
        RECT 82.240 176.250 95.350 176.390 ;
        RECT 82.240 176.190 82.560 176.250 ;
        RECT 64.315 175.910 65.080 176.050 ;
        RECT 64.315 175.865 64.605 175.910 ;
        RECT 47.295 175.710 47.585 175.755 ;
        RECT 54.640 175.710 54.960 175.770 ;
        RECT 56.480 175.710 56.800 175.770 ;
        RECT 47.295 175.570 56.800 175.710 ;
        RECT 47.295 175.525 47.585 175.570 ;
        RECT 54.640 175.510 54.960 175.570 ;
        RECT 56.480 175.510 56.800 175.570 ;
        RECT 58.735 175.550 59.025 175.865 ;
        RECT 64.760 175.850 65.080 175.910 ;
        RECT 67.995 176.050 68.285 176.095 ;
        RECT 70.755 176.050 71.045 176.095 ;
        RECT 74.420 176.050 74.740 176.110 ;
        RECT 67.995 175.910 71.045 176.050 ;
        RECT 67.995 175.865 68.285 175.910 ;
        RECT 70.755 175.865 71.045 175.910 ;
        RECT 71.750 175.910 74.740 176.050 ;
        RECT 71.750 175.770 71.890 175.910 ;
        RECT 74.420 175.850 74.740 175.910 ;
        RECT 78.510 176.050 78.800 176.095 ;
        RECT 80.860 176.050 81.180 176.110 ;
        RECT 81.770 176.050 82.060 176.095 ;
        RECT 78.510 175.910 82.060 176.050 ;
        RECT 78.510 175.865 78.800 175.910 ;
        RECT 80.860 175.850 81.180 175.910 ;
        RECT 81.770 175.865 82.060 175.910 ;
        RECT 82.690 176.050 82.980 176.095 ;
        RECT 84.550 176.050 84.840 176.095 ;
        RECT 82.690 175.910 84.840 176.050 ;
        RECT 82.690 175.865 82.980 175.910 ;
        RECT 84.550 175.865 84.840 175.910 ;
        RECT 59.815 175.710 60.105 175.755 ;
        RECT 63.395 175.710 63.685 175.755 ;
        RECT 65.230 175.710 65.520 175.755 ;
        RECT 59.815 175.570 65.520 175.710 ;
        RECT 59.815 175.525 60.105 175.570 ;
        RECT 63.395 175.525 63.685 175.570 ;
        RECT 65.230 175.525 65.520 175.570 ;
        RECT 68.900 175.510 69.220 175.770 ;
        RECT 70.280 175.710 70.600 175.770 ;
        RECT 71.215 175.710 71.505 175.755 ;
        RECT 70.280 175.570 71.505 175.710 ;
        RECT 70.280 175.510 70.600 175.570 ;
        RECT 71.215 175.525 71.505 175.570 ;
        RECT 71.660 175.510 71.980 175.770 ;
        RECT 72.580 175.510 72.900 175.770 ;
        RECT 73.055 175.710 73.345 175.755 ;
        RECT 73.960 175.710 74.280 175.770 ;
        RECT 73.055 175.570 74.280 175.710 ;
        RECT 73.055 175.525 73.345 175.570 ;
        RECT 28.420 175.370 28.740 175.430 ;
        RECT 38.080 175.370 38.400 175.430 ;
        RECT 28.420 175.230 38.400 175.370 ;
        RECT 28.420 175.170 28.740 175.230 ;
        RECT 38.080 175.170 38.400 175.230 ;
        RECT 49.595 175.185 49.885 175.415 ;
        RECT 50.500 175.370 50.820 175.430 ;
        RECT 53.275 175.370 53.565 175.415 ;
        RECT 61.540 175.370 61.860 175.430 ;
        RECT 50.500 175.230 61.860 175.370 ;
        RECT 28.900 175.030 29.190 175.075 ;
        RECT 30.760 175.030 31.050 175.075 ;
        RECT 33.540 175.030 33.830 175.075 ;
        RECT 28.900 174.890 33.830 175.030 ;
        RECT 28.900 174.845 29.190 174.890 ;
        RECT 30.760 174.845 31.050 174.890 ;
        RECT 33.540 174.845 33.830 174.890 ;
        RECT 38.965 175.030 39.255 175.075 ;
        RECT 40.855 175.030 41.145 175.075 ;
        RECT 43.975 175.030 44.265 175.075 ;
        RECT 38.965 174.890 44.265 175.030 ;
        RECT 49.670 175.030 49.810 175.185 ;
        RECT 50.500 175.170 50.820 175.230 ;
        RECT 53.275 175.185 53.565 175.230 ;
        RECT 61.540 175.170 61.860 175.230 ;
        RECT 65.695 175.370 65.985 175.415 ;
        RECT 67.060 175.370 67.380 175.430 ;
        RECT 68.440 175.370 68.760 175.430 ;
        RECT 65.695 175.230 68.760 175.370 ;
        RECT 68.990 175.370 69.130 175.510 ;
        RECT 73.130 175.370 73.270 175.525 ;
        RECT 73.960 175.510 74.280 175.570 ;
        RECT 74.895 175.525 75.185 175.755 ;
        RECT 80.370 175.710 80.660 175.755 ;
        RECT 82.690 175.710 82.905 175.865 ;
        RECT 85.920 175.850 86.240 176.110 ;
        RECT 94.660 175.850 94.980 176.110 ;
        RECT 95.210 176.050 95.350 176.250 ;
        RECT 96.500 176.190 96.820 176.450 ;
        RECT 98.815 176.390 99.105 176.435 ;
        RECT 99.720 176.390 100.040 176.450 ;
        RECT 98.815 176.250 100.040 176.390 ;
        RECT 98.815 176.205 99.105 176.250 ;
        RECT 99.720 176.190 100.040 176.250 ;
        RECT 102.020 176.390 102.340 176.450 ;
        RECT 102.495 176.390 102.785 176.435 ;
        RECT 102.020 176.250 102.785 176.390 ;
        RECT 102.020 176.190 102.340 176.250 ;
        RECT 102.495 176.205 102.785 176.250 ;
        RECT 104.795 176.390 105.085 176.435 ;
        RECT 106.160 176.390 106.480 176.450 ;
        RECT 104.795 176.250 106.480 176.390 ;
        RECT 104.795 176.205 105.085 176.250 ;
        RECT 106.160 176.190 106.480 176.250 ;
        RECT 107.080 176.190 107.400 176.450 ;
        RECT 96.975 176.050 97.265 176.095 ;
        RECT 95.210 175.910 97.265 176.050 ;
        RECT 96.975 175.865 97.265 175.910 ;
        RECT 80.370 175.570 82.905 175.710 ;
        RECT 85.000 175.710 85.320 175.770 ;
        RECT 85.475 175.710 85.765 175.755 ;
        RECT 85.000 175.570 85.765 175.710 ;
        RECT 80.370 175.525 80.660 175.570 ;
        RECT 68.990 175.230 73.270 175.370 ;
        RECT 65.695 175.185 65.985 175.230 ;
        RECT 67.060 175.170 67.380 175.230 ;
        RECT 68.440 175.170 68.760 175.230 ;
        RECT 54.180 175.030 54.500 175.090 ;
        RECT 56.955 175.030 57.245 175.075 ;
        RECT 49.670 174.890 57.245 175.030 ;
        RECT 38.965 174.845 39.255 174.890 ;
        RECT 40.855 174.845 41.145 174.890 ;
        RECT 43.975 174.845 44.265 174.890 ;
        RECT 54.180 174.830 54.500 174.890 ;
        RECT 56.955 174.845 57.245 174.890 ;
        RECT 59.815 175.030 60.105 175.075 ;
        RECT 62.935 175.030 63.225 175.075 ;
        RECT 64.825 175.030 65.115 175.075 ;
        RECT 74.970 175.030 75.110 175.525 ;
        RECT 85.000 175.510 85.320 175.570 ;
        RECT 85.475 175.525 85.765 175.570 ;
        RECT 88.680 175.710 89.000 175.770 ;
        RECT 101.100 175.710 101.420 175.770 ;
        RECT 88.680 175.570 101.420 175.710 ;
        RECT 88.680 175.510 89.000 175.570 ;
        RECT 101.100 175.510 101.420 175.570 ;
        RECT 102.480 175.710 102.800 175.770 ;
        RECT 102.955 175.710 103.245 175.755 ;
        RECT 106.635 175.710 106.925 175.755 ;
        RECT 102.480 175.570 106.925 175.710 ;
        RECT 102.480 175.510 102.800 175.570 ;
        RECT 102.955 175.525 103.245 175.570 ;
        RECT 106.635 175.525 106.925 175.570 ;
        RECT 109.395 175.525 109.685 175.755 ;
        RECT 76.505 175.370 76.795 175.415 ;
        RECT 81.780 175.370 82.100 175.430 ;
        RECT 76.505 175.230 82.100 175.370 ;
        RECT 76.505 175.185 76.795 175.230 ;
        RECT 81.780 175.170 82.100 175.230 ;
        RECT 83.635 175.370 83.925 175.415 ;
        RECT 87.760 175.370 88.080 175.430 ;
        RECT 83.635 175.230 88.080 175.370 ;
        RECT 83.635 175.185 83.925 175.230 ;
        RECT 87.760 175.170 88.080 175.230 ;
        RECT 95.580 175.370 95.900 175.430 ;
        RECT 97.420 175.370 97.740 175.430 ;
        RECT 101.575 175.370 101.865 175.415 ;
        RECT 105.715 175.370 106.005 175.415 ;
        RECT 95.580 175.230 106.005 175.370 ;
        RECT 95.580 175.170 95.900 175.230 ;
        RECT 97.420 175.170 97.740 175.230 ;
        RECT 101.575 175.185 101.865 175.230 ;
        RECT 105.715 175.185 106.005 175.230 ;
        RECT 59.815 174.890 65.115 175.030 ;
        RECT 59.815 174.845 60.105 174.890 ;
        RECT 62.935 174.845 63.225 174.890 ;
        RECT 64.825 174.845 65.115 174.890 ;
        RECT 65.310 174.890 75.110 175.030 ;
        RECT 80.370 175.030 80.660 175.075 ;
        RECT 83.150 175.030 83.440 175.075 ;
        RECT 85.010 175.030 85.300 175.075 ;
        RECT 80.370 174.890 85.300 175.030 ;
        RECT 27.040 174.690 27.360 174.750 ;
        RECT 31.180 174.690 31.500 174.750 ;
        RECT 27.040 174.550 31.500 174.690 ;
        RECT 27.040 174.490 27.360 174.550 ;
        RECT 31.180 174.490 31.500 174.550 ;
        RECT 36.240 174.690 36.560 174.750 ;
        RECT 37.405 174.690 37.695 174.735 ;
        RECT 39.920 174.690 40.240 174.750 ;
        RECT 36.240 174.550 40.240 174.690 ;
        RECT 36.240 174.490 36.560 174.550 ;
        RECT 37.405 174.505 37.695 174.550 ;
        RECT 39.920 174.490 40.240 174.550 ;
        RECT 43.140 174.690 43.460 174.750 ;
        RECT 46.835 174.690 47.125 174.735 ;
        RECT 43.140 174.550 47.125 174.690 ;
        RECT 43.140 174.490 43.460 174.550 ;
        RECT 46.835 174.505 47.125 174.550 ;
        RECT 52.355 174.690 52.645 174.735 ;
        RECT 54.640 174.690 54.960 174.750 ;
        RECT 52.355 174.550 54.960 174.690 ;
        RECT 52.355 174.505 52.645 174.550 ;
        RECT 54.640 174.490 54.960 174.550 ;
        RECT 56.020 174.490 56.340 174.750 ;
        RECT 60.620 174.690 60.940 174.750 ;
        RECT 65.310 174.690 65.450 174.890 ;
        RECT 80.370 174.845 80.660 174.890 ;
        RECT 83.150 174.845 83.440 174.890 ;
        RECT 85.010 174.845 85.300 174.890 ;
        RECT 86.840 175.030 87.160 175.090 ;
        RECT 100.640 175.030 100.960 175.090 ;
        RECT 109.470 175.030 109.610 175.525 ;
        RECT 110.300 175.170 110.620 175.430 ;
        RECT 86.840 174.890 92.130 175.030 ;
        RECT 86.840 174.830 87.160 174.890 ;
        RECT 60.620 174.550 65.450 174.690 ;
        RECT 65.680 174.690 66.000 174.750 ;
        RECT 66.615 174.690 66.905 174.735 ;
        RECT 65.680 174.550 66.905 174.690 ;
        RECT 60.620 174.490 60.940 174.550 ;
        RECT 65.680 174.490 66.000 174.550 ;
        RECT 66.615 174.505 66.905 174.550 ;
        RECT 67.980 174.690 68.300 174.750 ;
        RECT 69.835 174.690 70.125 174.735 ;
        RECT 67.980 174.550 70.125 174.690 ;
        RECT 67.980 174.490 68.300 174.550 ;
        RECT 69.835 174.505 70.125 174.550 ;
        RECT 75.340 174.490 75.660 174.750 ;
        RECT 84.540 174.690 84.860 174.750 ;
        RECT 91.440 174.690 91.760 174.750 ;
        RECT 84.540 174.550 91.760 174.690 ;
        RECT 91.990 174.690 92.130 174.890 ;
        RECT 100.640 174.890 109.610 175.030 ;
        RECT 100.640 174.830 100.960 174.890 ;
        RECT 105.700 174.690 106.020 174.750 ;
        RECT 91.990 174.550 106.020 174.690 ;
        RECT 84.540 174.490 84.860 174.550 ;
        RECT 91.440 174.490 91.760 174.550 ;
        RECT 105.700 174.490 106.020 174.550 ;
        RECT 107.080 174.690 107.400 174.750 ;
        RECT 108.935 174.690 109.225 174.735 ;
        RECT 107.080 174.550 109.225 174.690 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 107.080 174.490 107.400 174.550 ;
        RECT 108.935 174.505 109.225 174.550 ;
        RECT 26.970 173.870 113.450 174.350 ;
        RECT 42.220 173.670 42.540 173.730 ;
        RECT 52.800 173.670 53.120 173.730 ;
        RECT 32.650 173.530 35.090 173.670 ;
        RECT 31.640 173.130 31.960 173.390 ;
        RECT 28.435 172.990 28.725 173.035 ;
        RECT 32.650 172.990 32.790 173.530 ;
        RECT 34.400 172.990 34.720 173.050 ;
        RECT 28.435 172.850 32.790 172.990 ;
        RECT 33.110 172.850 34.720 172.990 ;
        RECT 34.950 172.990 35.090 173.530 ;
        RECT 42.220 173.530 53.120 173.670 ;
        RECT 42.220 173.470 42.540 173.530 ;
        RECT 52.800 173.470 53.120 173.530 ;
        RECT 56.480 173.670 56.800 173.730 ;
        RECT 68.900 173.670 69.220 173.730 ;
        RECT 56.480 173.530 69.220 173.670 ;
        RECT 56.480 173.470 56.800 173.530 ;
        RECT 68.900 173.470 69.220 173.530 ;
        RECT 72.595 173.670 72.885 173.715 ;
        RECT 73.040 173.670 73.360 173.730 ;
        RECT 72.595 173.530 73.360 173.670 ;
        RECT 72.595 173.485 72.885 173.530 ;
        RECT 73.040 173.470 73.360 173.530 ;
        RECT 83.160 173.670 83.480 173.730 ;
        RECT 86.840 173.670 87.160 173.730 ;
        RECT 103.400 173.670 103.720 173.730 ;
        RECT 83.160 173.530 87.160 173.670 ;
        RECT 83.160 173.470 83.480 173.530 ;
        RECT 86.840 173.470 87.160 173.530 ;
        RECT 99.810 173.530 103.720 173.670 ;
        RECT 41.265 173.330 41.555 173.375 ;
        RECT 43.155 173.330 43.445 173.375 ;
        RECT 46.275 173.330 46.565 173.375 ;
        RECT 41.265 173.190 46.565 173.330 ;
        RECT 41.265 173.145 41.555 173.190 ;
        RECT 43.155 173.145 43.445 173.190 ;
        RECT 46.275 173.145 46.565 173.190 ;
        RECT 50.465 173.330 50.755 173.375 ;
        RECT 52.355 173.330 52.645 173.375 ;
        RECT 55.475 173.330 55.765 173.375 ;
        RECT 50.465 173.190 55.765 173.330 ;
        RECT 50.465 173.145 50.755 173.190 ;
        RECT 52.355 173.145 52.645 173.190 ;
        RECT 55.475 173.145 55.765 173.190 ;
        RECT 64.875 173.330 65.165 173.375 ;
        RECT 67.995 173.330 68.285 173.375 ;
        RECT 69.885 173.330 70.175 173.375 ;
        RECT 64.875 173.190 70.175 173.330 ;
        RECT 64.875 173.145 65.165 173.190 ;
        RECT 67.995 173.145 68.285 173.190 ;
        RECT 69.885 173.145 70.175 173.190 ;
        RECT 75.125 173.330 75.415 173.375 ;
        RECT 77.640 173.330 77.960 173.390 ;
        RECT 75.125 173.190 77.960 173.330 ;
        RECT 75.125 173.145 75.415 173.190 ;
        RECT 77.640 173.130 77.960 173.190 ;
        RECT 78.990 173.330 79.280 173.375 ;
        RECT 81.770 173.330 82.060 173.375 ;
        RECT 83.630 173.330 83.920 173.375 ;
        RECT 78.990 173.190 83.920 173.330 ;
        RECT 78.990 173.145 79.280 173.190 ;
        RECT 81.770 173.145 82.060 173.190 ;
        RECT 83.630 173.145 83.920 173.190 ;
        RECT 91.870 173.330 92.160 173.375 ;
        RECT 94.650 173.330 94.940 173.375 ;
        RECT 96.510 173.330 96.800 173.375 ;
        RECT 99.260 173.330 99.580 173.390 ;
        RECT 91.870 173.190 96.800 173.330 ;
        RECT 91.870 173.145 92.160 173.190 ;
        RECT 94.650 173.145 94.940 173.190 ;
        RECT 96.510 173.145 96.800 173.190 ;
        RECT 97.970 173.190 99.580 173.330 ;
        RECT 37.160 172.990 37.480 173.050 ;
        RECT 41.775 172.990 42.065 173.035 ;
        RECT 34.950 172.850 36.930 172.990 ;
        RECT 28.435 172.805 28.725 172.850 ;
        RECT 29.355 172.650 29.645 172.695 ;
        RECT 29.800 172.650 30.120 172.710 ;
        RECT 29.355 172.510 30.120 172.650 ;
        RECT 29.355 172.465 29.645 172.510 ;
        RECT 29.800 172.450 30.120 172.510 ;
        RECT 32.100 172.650 32.420 172.710 ;
        RECT 33.110 172.650 33.250 172.850 ;
        RECT 34.400 172.790 34.720 172.850 ;
        RECT 32.100 172.510 33.250 172.650 ;
        RECT 33.955 172.650 34.245 172.695 ;
        RECT 35.780 172.650 36.100 172.710 ;
        RECT 33.955 172.510 36.100 172.650 ;
        RECT 36.790 172.650 36.930 172.850 ;
        RECT 37.160 172.850 42.065 172.990 ;
        RECT 37.160 172.790 37.480 172.850 ;
        RECT 41.775 172.805 42.065 172.850 ;
        RECT 49.135 172.805 49.425 173.035 ;
        RECT 49.595 172.990 49.885 173.035 ;
        RECT 53.720 172.990 54.040 173.050 ;
        RECT 49.595 172.850 54.040 172.990 ;
        RECT 49.595 172.805 49.885 172.850 ;
        RECT 38.080 172.650 38.400 172.710 ;
        RECT 39.475 172.650 39.765 172.695 ;
        RECT 40.380 172.650 40.700 172.710 ;
        RECT 36.790 172.510 37.850 172.650 ;
        RECT 32.100 172.450 32.420 172.510 ;
        RECT 33.955 172.465 34.245 172.510 ;
        RECT 35.780 172.450 36.100 172.510 ;
        RECT 30.275 172.310 30.565 172.355 ;
        RECT 37.160 172.310 37.480 172.370 ;
        RECT 30.275 172.170 37.480 172.310 ;
        RECT 37.710 172.310 37.850 172.510 ;
        RECT 38.080 172.510 40.700 172.650 ;
        RECT 38.080 172.450 38.400 172.510 ;
        RECT 39.475 172.465 39.765 172.510 ;
        RECT 40.380 172.450 40.700 172.510 ;
        RECT 40.860 172.650 41.150 172.695 ;
        RECT 42.695 172.650 42.985 172.695 ;
        RECT 46.275 172.650 46.565 172.695 ;
        RECT 40.860 172.510 46.565 172.650 ;
        RECT 40.860 172.465 41.150 172.510 ;
        RECT 42.695 172.465 42.985 172.510 ;
        RECT 46.275 172.465 46.565 172.510 ;
        RECT 47.280 172.670 47.600 172.710 ;
        RECT 47.280 172.450 47.645 172.670 ;
        RECT 42.220 172.310 42.540 172.370 ;
        RECT 47.355 172.355 47.645 172.450 ;
        RECT 37.710 172.170 42.540 172.310 ;
        RECT 30.275 172.125 30.565 172.170 ;
        RECT 37.160 172.110 37.480 172.170 ;
        RECT 42.220 172.110 42.540 172.170 ;
        RECT 44.055 172.310 44.705 172.355 ;
        RECT 47.355 172.310 47.945 172.355 ;
        RECT 44.055 172.170 47.945 172.310 ;
        RECT 49.210 172.310 49.350 172.805 ;
        RECT 53.720 172.790 54.040 172.850 ;
        RECT 60.175 172.990 60.465 173.035 ;
        RECT 60.620 172.990 60.940 173.050 ;
        RECT 67.060 172.990 67.380 173.050 ;
        RECT 60.175 172.850 60.940 172.990 ;
        RECT 60.175 172.805 60.465 172.850 ;
        RECT 60.620 172.790 60.940 172.850 ;
        RECT 61.170 172.850 67.380 172.990 ;
        RECT 61.170 172.695 61.310 172.850 ;
        RECT 67.060 172.790 67.380 172.850 ;
        RECT 70.755 172.990 71.045 173.035 ;
        RECT 70.755 172.850 82.010 172.990 ;
        RECT 70.755 172.805 71.045 172.850 ;
        RECT 50.060 172.650 50.350 172.695 ;
        RECT 51.895 172.650 52.185 172.695 ;
        RECT 55.475 172.650 55.765 172.695 ;
        RECT 50.060 172.510 55.765 172.650 ;
        RECT 50.060 172.465 50.350 172.510 ;
        RECT 51.895 172.465 52.185 172.510 ;
        RECT 55.475 172.465 55.765 172.510 ;
        RECT 50.500 172.310 50.820 172.370 ;
        RECT 49.210 172.170 50.820 172.310 ;
        RECT 44.055 172.125 44.705 172.170 ;
        RECT 47.655 172.125 47.945 172.170 ;
        RECT 50.500 172.110 50.820 172.170 ;
        RECT 50.975 172.125 51.265 172.355 ;
        RECT 51.420 172.310 51.740 172.370 ;
        RECT 56.555 172.355 56.845 172.670 ;
        RECT 61.095 172.465 61.385 172.695 ;
        RECT 63.795 172.355 64.085 172.670 ;
        RECT 64.875 172.650 65.165 172.695 ;
        RECT 68.455 172.650 68.745 172.695 ;
        RECT 70.290 172.650 70.580 172.695 ;
        RECT 64.875 172.510 70.580 172.650 ;
        RECT 64.875 172.465 65.165 172.510 ;
        RECT 68.455 172.465 68.745 172.510 ;
        RECT 70.290 172.465 70.580 172.510 ;
        RECT 73.040 172.450 73.360 172.710 ;
        RECT 73.960 172.650 74.280 172.710 ;
        RECT 78.990 172.650 79.280 172.695 ;
        RECT 81.870 172.650 82.010 172.850 ;
        RECT 82.240 172.790 82.560 173.050 ;
        RECT 84.095 172.990 84.385 173.035 ;
        RECT 85.000 172.990 85.320 173.050 ;
        RECT 84.095 172.850 85.320 172.990 ;
        RECT 84.095 172.805 84.385 172.850 ;
        RECT 84.170 172.650 84.310 172.805 ;
        RECT 85.000 172.790 85.320 172.850 ;
        RECT 95.135 172.990 95.425 173.035 ;
        RECT 97.970 172.990 98.110 173.190 ;
        RECT 99.260 173.130 99.580 173.190 ;
        RECT 95.135 172.850 98.110 172.990 ;
        RECT 95.135 172.805 95.425 172.850 ;
        RECT 98.355 172.805 98.645 173.035 ;
        RECT 98.800 172.990 99.120 173.050 ;
        RECT 99.810 172.990 99.950 173.530 ;
        RECT 103.400 173.470 103.720 173.530 ;
        RECT 105.700 173.670 106.020 173.730 ;
        RECT 110.300 173.670 110.620 173.730 ;
        RECT 105.700 173.530 112.370 173.670 ;
        RECT 105.700 173.470 106.020 173.530 ;
        RECT 110.300 173.470 110.620 173.530 ;
        RECT 101.115 173.330 101.405 173.375 ;
        RECT 102.940 173.330 103.260 173.390 ;
        RECT 101.115 173.190 103.260 173.330 ;
        RECT 101.115 173.145 101.405 173.190 ;
        RECT 102.940 173.130 103.260 173.190 ;
        RECT 104.435 173.330 104.725 173.375 ;
        RECT 107.555 173.330 107.845 173.375 ;
        RECT 109.445 173.330 109.735 173.375 ;
        RECT 104.435 173.190 109.735 173.330 ;
        RECT 104.435 173.145 104.725 173.190 ;
        RECT 107.555 173.145 107.845 173.190 ;
        RECT 109.445 173.145 109.735 173.190 ;
        RECT 98.800 172.850 99.950 172.990 ;
        RECT 73.960 172.510 76.030 172.650 ;
        RECT 73.960 172.450 74.280 172.510 ;
        RECT 53.255 172.310 53.905 172.355 ;
        RECT 56.555 172.310 57.145 172.355 ;
        RECT 51.420 172.170 57.145 172.310 ;
        RECT 33.495 171.970 33.785 172.015 ;
        RECT 39.920 171.970 40.240 172.030 ;
        RECT 33.495 171.830 40.240 171.970 ;
        RECT 33.495 171.785 33.785 171.830 ;
        RECT 39.920 171.770 40.240 171.830 ;
        RECT 41.300 171.970 41.620 172.030 ;
        RECT 51.050 171.970 51.190 172.125 ;
        RECT 51.420 172.110 51.740 172.170 ;
        RECT 53.255 172.125 53.905 172.170 ;
        RECT 56.855 172.125 57.145 172.170 ;
        RECT 63.495 172.310 64.085 172.355 ;
        RECT 66.735 172.310 67.385 172.355 ;
        RECT 69.375 172.310 69.665 172.355 ;
        RECT 74.880 172.310 75.200 172.370 ;
        RECT 63.495 172.170 69.130 172.310 ;
        RECT 63.495 172.125 63.785 172.170 ;
        RECT 66.735 172.125 67.385 172.170 ;
        RECT 41.300 171.830 51.190 171.970 ;
        RECT 55.560 171.970 55.880 172.030 ;
        RECT 58.335 171.970 58.625 172.015 ;
        RECT 55.560 171.830 58.625 171.970 ;
        RECT 41.300 171.770 41.620 171.830 ;
        RECT 55.560 171.770 55.880 171.830 ;
        RECT 58.335 171.785 58.625 171.830 ;
        RECT 60.620 171.970 60.940 172.030 ;
        RECT 62.015 171.970 62.305 172.015 ;
        RECT 60.620 171.830 62.305 171.970 ;
        RECT 68.990 171.970 69.130 172.170 ;
        RECT 69.375 172.170 75.200 172.310 ;
        RECT 69.375 172.125 69.665 172.170 ;
        RECT 74.880 172.110 75.200 172.170 ;
        RECT 75.340 171.970 75.660 172.030 ;
        RECT 68.990 171.830 75.660 171.970 ;
        RECT 75.890 171.970 76.030 172.510 ;
        RECT 78.990 172.510 81.525 172.650 ;
        RECT 81.870 172.510 84.310 172.650 ;
        RECT 78.990 172.465 79.280 172.510 ;
        RECT 80.400 172.355 80.720 172.370 ;
        RECT 77.130 172.310 77.420 172.355 ;
        RECT 80.390 172.310 80.720 172.355 ;
        RECT 77.130 172.170 80.720 172.310 ;
        RECT 77.130 172.125 77.420 172.170 ;
        RECT 80.390 172.125 80.720 172.170 ;
        RECT 81.310 172.355 81.525 172.510 ;
        RECT 84.555 172.465 84.845 172.695 ;
        RECT 91.870 172.650 92.160 172.695 ;
        RECT 94.660 172.650 94.980 172.710 ;
        RECT 96.975 172.650 97.265 172.695 ;
        RECT 91.870 172.510 94.405 172.650 ;
        RECT 91.870 172.465 92.160 172.510 ;
        RECT 81.310 172.310 81.600 172.355 ;
        RECT 83.170 172.310 83.460 172.355 ;
        RECT 81.310 172.170 83.460 172.310 ;
        RECT 81.310 172.125 81.600 172.170 ;
        RECT 83.170 172.125 83.460 172.170 ;
        RECT 80.400 172.110 80.720 172.125 ;
        RECT 84.630 171.970 84.770 172.465 ;
        RECT 86.380 172.310 86.700 172.370 ;
        RECT 94.190 172.355 94.405 172.510 ;
        RECT 94.660 172.510 97.265 172.650 ;
        RECT 94.660 172.450 94.980 172.510 ;
        RECT 96.975 172.465 97.265 172.510 ;
        RECT 90.010 172.310 90.300 172.355 ;
        RECT 93.270 172.310 93.560 172.355 ;
        RECT 86.380 172.170 93.560 172.310 ;
        RECT 86.380 172.110 86.700 172.170 ;
        RECT 90.010 172.125 90.300 172.170 ;
        RECT 93.270 172.125 93.560 172.170 ;
        RECT 94.190 172.310 94.480 172.355 ;
        RECT 96.050 172.310 96.340 172.355 ;
        RECT 98.430 172.310 98.570 172.805 ;
        RECT 98.800 172.790 99.120 172.850 ;
        RECT 101.560 172.790 101.880 173.050 ;
        RECT 103.860 172.990 104.180 173.050 ;
        RECT 103.030 172.850 104.180 172.990 ;
        RECT 99.260 172.650 99.580 172.710 ;
        RECT 103.030 172.650 103.170 172.850 ;
        RECT 103.860 172.790 104.180 172.850 ;
        RECT 110.315 172.990 110.605 173.035 ;
        RECT 111.220 172.990 111.540 173.050 ;
        RECT 112.230 172.990 112.370 173.530 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 110.315 172.850 111.540 172.990 ;
        RECT 110.315 172.805 110.605 172.850 ;
        RECT 111.220 172.790 111.540 172.850 ;
        RECT 111.770 172.850 112.370 172.990 ;
        RECT 111.770 172.710 111.910 172.850 ;
        RECT 99.260 172.510 103.170 172.650 ;
        RECT 99.260 172.450 99.580 172.510 ;
        RECT 94.190 172.170 96.340 172.310 ;
        RECT 94.190 172.125 94.480 172.170 ;
        RECT 96.050 172.125 96.340 172.170 ;
        RECT 97.970 172.170 98.570 172.310 ;
        RECT 100.640 172.310 100.960 172.370 ;
        RECT 103.355 172.355 103.645 172.670 ;
        RECT 104.435 172.650 104.725 172.695 ;
        RECT 108.015 172.650 108.305 172.695 ;
        RECT 109.850 172.650 110.140 172.695 ;
        RECT 104.435 172.510 110.140 172.650 ;
        RECT 104.435 172.465 104.725 172.510 ;
        RECT 108.015 172.465 108.305 172.510 ;
        RECT 109.850 172.465 110.140 172.510 ;
        RECT 111.680 172.450 112.000 172.710 ;
        RECT 103.055 172.310 103.645 172.355 ;
        RECT 106.295 172.310 106.945 172.355 ;
        RECT 100.640 172.170 106.945 172.310 ;
        RECT 75.890 171.830 84.770 171.970 ;
        RECT 85.475 171.970 85.765 172.015 ;
        RECT 85.920 171.970 86.240 172.030 ;
        RECT 85.475 171.830 86.240 171.970 ;
        RECT 60.620 171.770 60.940 171.830 ;
        RECT 62.015 171.785 62.305 171.830 ;
        RECT 75.340 171.770 75.660 171.830 ;
        RECT 85.475 171.785 85.765 171.830 ;
        RECT 85.920 171.770 86.240 171.830 ;
        RECT 88.005 171.970 88.295 172.015 ;
        RECT 91.900 171.970 92.220 172.030 ;
        RECT 88.005 171.830 92.220 171.970 ;
        RECT 88.005 171.785 88.295 171.830 ;
        RECT 91.900 171.770 92.220 171.830 ;
        RECT 92.360 171.970 92.680 172.030 ;
        RECT 95.580 171.970 95.900 172.030 ;
        RECT 97.970 171.970 98.110 172.170 ;
        RECT 100.640 172.110 100.960 172.170 ;
        RECT 103.055 172.125 103.345 172.170 ;
        RECT 106.295 172.125 106.945 172.170 ;
        RECT 108.935 172.310 109.225 172.355 ;
        RECT 110.760 172.310 111.080 172.370 ;
        RECT 108.935 172.170 111.080 172.310 ;
        RECT 108.935 172.125 109.225 172.170 ;
        RECT 110.760 172.110 111.080 172.170 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 92.360 171.830 98.110 171.970 ;
        RECT 99.275 171.970 99.565 172.015 ;
        RECT 104.320 171.970 104.640 172.030 ;
        RECT 99.275 171.830 104.640 171.970 ;
        RECT 92.360 171.770 92.680 171.830 ;
        RECT 95.580 171.770 95.900 171.830 ;
        RECT 99.275 171.785 99.565 171.830 ;
        RECT 104.320 171.770 104.640 171.830 ;
        RECT 104.780 171.970 105.100 172.030 ;
        RECT 108.460 171.970 108.780 172.030 ;
        RECT 104.780 171.830 108.780 171.970 ;
        RECT 104.780 171.770 105.100 171.830 ;
        RECT 108.460 171.770 108.780 171.830 ;
        RECT 110.300 171.970 110.620 172.030 ;
        RECT 111.235 171.970 111.525 172.015 ;
        RECT 110.300 171.830 111.525 171.970 ;
        RECT 110.300 171.770 110.620 171.830 ;
        RECT 111.235 171.785 111.525 171.830 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 26.970 171.150 113.450 171.630 ;
        RECT 25.200 170.950 25.520 171.010 ;
        RECT 34.860 170.950 35.180 171.010 ;
        RECT 37.405 170.950 37.695 170.995 ;
        RECT 25.200 170.810 31.870 170.950 ;
        RECT 25.200 170.750 25.520 170.810 ;
        RECT 29.360 170.610 29.650 170.655 ;
        RECT 31.220 170.610 31.510 170.655 ;
        RECT 29.360 170.470 31.510 170.610 ;
        RECT 31.730 170.610 31.870 170.810 ;
        RECT 34.860 170.810 37.695 170.950 ;
        RECT 34.860 170.750 35.180 170.810 ;
        RECT 37.405 170.765 37.695 170.810 ;
        RECT 38.080 170.950 38.400 171.010 ;
        RECT 40.840 170.950 41.160 171.010 ;
        RECT 38.080 170.810 41.160 170.950 ;
        RECT 38.080 170.750 38.400 170.810 ;
        RECT 40.840 170.750 41.160 170.810 ;
        RECT 42.680 170.950 43.000 171.010 ;
        RECT 46.360 170.950 46.680 171.010 ;
        RECT 42.680 170.810 46.680 170.950 ;
        RECT 42.680 170.750 43.000 170.810 ;
        RECT 46.360 170.750 46.680 170.810 ;
        RECT 51.435 170.950 51.725 170.995 ;
        RECT 51.435 170.810 52.570 170.950 ;
        RECT 51.435 170.765 51.725 170.810 ;
        RECT 32.140 170.610 32.430 170.655 ;
        RECT 35.400 170.610 35.690 170.655 ;
        RECT 50.975 170.610 51.265 170.655 ;
        RECT 31.730 170.470 35.690 170.610 ;
        RECT 29.360 170.425 29.650 170.470 ;
        RECT 31.220 170.425 31.510 170.470 ;
        RECT 32.140 170.425 32.430 170.470 ;
        RECT 35.400 170.425 35.690 170.470 ;
        RECT 35.870 170.470 51.265 170.610 ;
        RECT 52.430 170.610 52.570 170.810 ;
        RECT 53.260 170.750 53.580 171.010 ;
        RECT 54.640 170.950 54.960 171.010 ;
        RECT 55.115 170.950 55.405 170.995 ;
        RECT 63.395 170.950 63.685 170.995 ;
        RECT 54.640 170.810 55.405 170.950 ;
        RECT 54.640 170.750 54.960 170.810 ;
        RECT 55.115 170.765 55.405 170.810 ;
        RECT 58.870 170.810 63.685 170.950 ;
        RECT 56.020 170.610 56.340 170.670 ;
        RECT 58.870 170.610 59.010 170.810 ;
        RECT 63.395 170.765 63.685 170.810 ;
        RECT 74.880 170.750 75.200 171.010 ;
        RECT 77.640 170.950 77.960 171.010 ;
        RECT 79.480 170.950 79.800 171.010 ;
        RECT 77.640 170.810 79.800 170.950 ;
        RECT 77.640 170.750 77.960 170.810 ;
        RECT 79.480 170.750 79.800 170.810 ;
        RECT 80.860 170.750 81.180 171.010 ;
        RECT 85.920 170.950 86.240 171.010 ;
        RECT 81.410 170.810 86.240 170.950 ;
        RECT 52.430 170.470 59.010 170.610 ;
        RECT 59.255 170.610 59.545 170.655 ;
        RECT 62.935 170.610 63.225 170.655 ;
        RECT 65.695 170.610 65.985 170.655 ;
        RECT 59.255 170.470 65.985 170.610 ;
        RECT 28.420 170.070 28.740 170.330 ;
        RECT 30.260 170.070 30.580 170.330 ;
        RECT 31.295 170.270 31.510 170.425 ;
        RECT 33.540 170.270 33.830 170.315 ;
        RECT 31.295 170.130 33.830 170.270 ;
        RECT 33.540 170.085 33.830 170.130 ;
        RECT 35.870 169.990 36.010 170.470 ;
        RECT 50.975 170.425 51.265 170.470 ;
        RECT 56.020 170.410 56.340 170.470 ;
        RECT 59.255 170.425 59.545 170.470 ;
        RECT 62.935 170.425 63.225 170.470 ;
        RECT 65.695 170.425 65.985 170.470 ;
        RECT 70.740 170.610 71.060 170.670 ;
        RECT 73.960 170.610 74.280 170.670 ;
        RECT 81.410 170.610 81.550 170.810 ;
        RECT 85.920 170.750 86.240 170.810 ;
        RECT 91.900 170.950 92.220 171.010 ;
        RECT 92.835 170.950 93.125 170.995 ;
        RECT 91.900 170.810 93.125 170.950 ;
        RECT 91.900 170.750 92.220 170.810 ;
        RECT 92.835 170.765 93.125 170.810 ;
        RECT 95.135 170.950 95.425 170.995 ;
        RECT 98.340 170.950 98.660 171.010 ;
        RECT 102.020 170.950 102.340 171.010 ;
        RECT 95.135 170.810 98.660 170.950 ;
        RECT 95.135 170.765 95.425 170.810 ;
        RECT 98.340 170.750 98.660 170.810 ;
        RECT 98.890 170.810 102.340 170.950 ;
        RECT 70.740 170.470 73.730 170.610 ;
        RECT 70.740 170.410 71.060 170.470 ;
        RECT 46.820 170.070 47.140 170.330 ;
        RECT 47.295 170.270 47.585 170.315 ;
        RECT 51.420 170.270 51.740 170.330 ;
        RECT 47.295 170.130 51.740 170.270 ;
        RECT 47.295 170.085 47.585 170.130 ;
        RECT 51.420 170.070 51.740 170.130 ;
        RECT 54.640 170.270 54.960 170.330 ;
        RECT 59.715 170.270 60.005 170.315 ;
        RECT 54.640 170.130 60.005 170.270 ;
        RECT 54.640 170.070 54.960 170.130 ;
        RECT 59.715 170.085 60.005 170.130 ;
        RECT 61.080 170.270 61.400 170.330 ;
        RECT 68.455 170.270 68.745 170.315 ;
        RECT 61.080 170.130 68.745 170.270 ;
        RECT 61.080 170.070 61.400 170.130 ;
        RECT 68.455 170.085 68.745 170.130 ;
        RECT 68.900 170.270 69.220 170.330 ;
        RECT 70.295 170.270 70.585 170.315 ;
        RECT 68.900 170.130 70.585 170.270 ;
        RECT 68.900 170.070 69.220 170.130 ;
        RECT 70.295 170.085 70.585 170.130 ;
        RECT 71.675 170.270 71.965 170.315 ;
        RECT 73.040 170.270 73.360 170.330 ;
        RECT 73.590 170.315 73.730 170.470 ;
        RECT 73.960 170.470 81.550 170.610 ;
        RECT 84.030 170.610 84.320 170.655 ;
        RECT 85.460 170.610 85.780 170.670 ;
        RECT 87.290 170.610 87.580 170.655 ;
        RECT 84.030 170.470 87.580 170.610 ;
        RECT 73.960 170.410 74.280 170.470 ;
        RECT 84.030 170.425 84.320 170.470 ;
        RECT 85.460 170.410 85.780 170.470 ;
        RECT 87.290 170.425 87.580 170.470 ;
        RECT 88.210 170.610 88.500 170.655 ;
        RECT 90.070 170.610 90.360 170.655 ;
        RECT 88.210 170.470 90.360 170.610 ;
        RECT 88.210 170.425 88.500 170.470 ;
        RECT 90.070 170.425 90.360 170.470 ;
        RECT 71.675 170.130 73.360 170.270 ;
        RECT 71.675 170.085 71.965 170.130 ;
        RECT 73.040 170.070 73.360 170.130 ;
        RECT 73.515 170.270 73.805 170.315 ;
        RECT 75.340 170.270 75.660 170.330 ;
        RECT 73.515 170.130 75.660 170.270 ;
        RECT 73.515 170.085 73.805 170.130 ;
        RECT 75.340 170.070 75.660 170.130 ;
        RECT 75.815 170.085 76.105 170.315 ;
        RECT 78.115 170.270 78.405 170.315 ;
        RECT 79.480 170.270 79.800 170.330 ;
        RECT 78.115 170.130 79.800 170.270 ;
        RECT 78.115 170.085 78.405 170.130 ;
        RECT 35.780 169.730 36.100 169.990 ;
        RECT 36.240 169.930 36.560 169.990 ;
        RECT 52.355 169.930 52.645 169.975 ;
        RECT 36.240 169.790 52.645 169.930 ;
        RECT 36.240 169.730 36.560 169.790 ;
        RECT 52.355 169.745 52.645 169.790 ;
        RECT 53.720 169.930 54.040 169.990 ;
        RECT 55.560 169.930 55.880 169.990 ;
        RECT 53.720 169.790 55.880 169.930 ;
        RECT 28.900 169.590 29.190 169.635 ;
        RECT 30.760 169.590 31.050 169.635 ;
        RECT 33.540 169.590 33.830 169.635 ;
        RECT 28.900 169.450 33.830 169.590 ;
        RECT 28.900 169.405 29.190 169.450 ;
        RECT 30.760 169.405 31.050 169.450 ;
        RECT 33.540 169.405 33.830 169.450 ;
        RECT 45.440 169.590 45.760 169.650 ;
        RECT 49.135 169.590 49.425 169.635 ;
        RECT 45.440 169.450 49.425 169.590 ;
        RECT 52.430 169.590 52.570 169.745 ;
        RECT 53.720 169.730 54.040 169.790 ;
        RECT 55.560 169.730 55.880 169.790 ;
        RECT 56.495 169.745 56.785 169.975 ;
        RECT 60.635 169.930 60.925 169.975 ;
        RECT 62.475 169.930 62.765 169.975 ;
        RECT 75.890 169.930 76.030 170.085 ;
        RECT 79.480 170.070 79.800 170.130 ;
        RECT 81.335 170.270 81.625 170.315 ;
        RECT 83.160 170.270 83.480 170.330 ;
        RECT 81.335 170.130 83.480 170.270 ;
        RECT 81.335 170.085 81.625 170.130 ;
        RECT 83.160 170.070 83.480 170.130 ;
        RECT 85.890 170.270 86.180 170.315 ;
        RECT 88.210 170.270 88.425 170.425 ;
        RECT 93.280 170.410 93.600 170.670 ;
        RECT 98.890 170.610 99.030 170.810 ;
        RECT 102.020 170.750 102.340 170.810 ;
        RECT 104.320 170.750 104.640 171.010 ;
        RECT 110.760 170.950 111.080 171.010 ;
        RECT 111.680 170.950 112.000 171.010 ;
        RECT 105.330 170.810 106.850 170.950 ;
        RECT 105.330 170.610 105.470 170.810 ;
        RECT 97.970 170.470 99.030 170.610 ;
        RECT 104.870 170.470 105.470 170.610 ;
        RECT 106.710 170.610 106.850 170.810 ;
        RECT 110.760 170.810 112.000 170.950 ;
        RECT 110.760 170.750 111.080 170.810 ;
        RECT 111.680 170.750 112.000 170.810 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 106.710 170.470 108.230 170.610 ;
        RECT 90.995 170.270 91.285 170.315 ;
        RECT 94.660 170.270 94.980 170.330 ;
        RECT 85.890 170.130 88.425 170.270 ;
        RECT 88.770 170.130 89.830 170.270 ;
        RECT 85.890 170.085 86.180 170.130 ;
        RECT 60.635 169.790 63.150 169.930 ;
        RECT 60.635 169.745 60.925 169.790 ;
        RECT 62.475 169.745 62.765 169.790 ;
        RECT 54.640 169.590 54.960 169.650 ;
        RECT 56.570 169.590 56.710 169.745 ;
        RECT 60.710 169.590 60.850 169.745 ;
        RECT 52.430 169.450 60.850 169.590 ;
        RECT 45.440 169.390 45.760 169.450 ;
        RECT 49.135 169.405 49.425 169.450 ;
        RECT 54.640 169.390 54.960 169.450 ;
        RECT 40.380 169.250 40.700 169.310 ;
        RECT 42.680 169.250 43.000 169.310 ;
        RECT 40.380 169.110 43.000 169.250 ;
        RECT 40.380 169.050 40.700 169.110 ;
        RECT 42.680 169.050 43.000 169.110 ;
        RECT 48.215 169.250 48.505 169.295 ;
        RECT 49.580 169.250 49.900 169.310 ;
        RECT 48.215 169.110 49.900 169.250 ;
        RECT 48.215 169.065 48.505 169.110 ;
        RECT 49.580 169.050 49.900 169.110 ;
        RECT 57.400 169.050 57.720 169.310 ;
        RECT 63.010 169.250 63.150 169.790 ;
        RECT 65.310 169.790 76.030 169.930 ;
        RECT 65.310 169.635 65.450 169.790 ;
        RECT 76.720 169.730 77.040 169.990 ;
        RECT 88.770 169.930 88.910 170.130 ;
        RECT 79.110 169.790 88.910 169.930 ;
        RECT 65.235 169.405 65.525 169.635 ;
        RECT 67.060 169.590 67.380 169.650 ;
        RECT 73.040 169.590 73.360 169.650 ;
        RECT 79.110 169.590 79.250 169.790 ;
        RECT 89.140 169.730 89.460 169.990 ;
        RECT 89.690 169.930 89.830 170.130 ;
        RECT 90.995 170.130 94.980 170.270 ;
        RECT 90.995 170.085 91.285 170.130 ;
        RECT 94.660 170.070 94.980 170.130 ;
        RECT 95.580 170.270 95.900 170.330 ;
        RECT 97.970 170.315 98.110 170.470 ;
        RECT 97.895 170.270 98.185 170.315 ;
        RECT 95.580 170.130 98.185 170.270 ;
        RECT 95.580 170.070 95.900 170.130 ;
        RECT 97.895 170.085 98.185 170.130 ;
        RECT 98.340 170.070 98.660 170.330 ;
        RECT 98.815 170.270 99.105 170.315 ;
        RECT 99.260 170.270 99.580 170.330 ;
        RECT 98.815 170.130 99.580 170.270 ;
        RECT 98.815 170.085 99.105 170.130 ;
        RECT 99.260 170.070 99.580 170.130 ;
        RECT 99.720 170.070 100.040 170.330 ;
        RECT 102.020 170.070 102.340 170.330 ;
        RECT 102.480 170.070 102.800 170.330 ;
        RECT 102.955 170.085 103.245 170.315 ;
        RECT 103.400 170.270 103.720 170.330 ;
        RECT 103.875 170.270 104.165 170.315 ;
        RECT 104.870 170.270 105.010 170.470 ;
        RECT 108.090 170.315 108.230 170.470 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 103.400 170.130 105.010 170.270 ;
        RECT 91.440 169.930 91.760 169.990 ;
        RECT 91.915 169.930 92.205 169.975 ;
        RECT 100.180 169.930 100.500 169.990 ;
        RECT 89.690 169.790 91.210 169.930 ;
        RECT 67.060 169.450 79.250 169.590 ;
        RECT 80.860 169.590 81.180 169.650 ;
        RECT 82.025 169.590 82.315 169.635 ;
        RECT 80.860 169.450 82.315 169.590 ;
        RECT 67.060 169.390 67.380 169.450 ;
        RECT 73.040 169.390 73.360 169.450 ;
        RECT 80.860 169.390 81.180 169.450 ;
        RECT 82.025 169.405 82.315 169.450 ;
        RECT 85.890 169.590 86.180 169.635 ;
        RECT 88.670 169.590 88.960 169.635 ;
        RECT 90.530 169.590 90.820 169.635 ;
        RECT 85.890 169.450 90.820 169.590 ;
        RECT 91.070 169.590 91.210 169.790 ;
        RECT 91.440 169.790 92.205 169.930 ;
        RECT 91.440 169.730 91.760 169.790 ;
        RECT 91.915 169.745 92.205 169.790 ;
        RECT 92.450 169.790 100.500 169.930 ;
        RECT 92.450 169.590 92.590 169.790 ;
        RECT 100.180 169.730 100.500 169.790 ;
        RECT 101.560 169.930 101.880 169.990 ;
        RECT 103.030 169.930 103.170 170.085 ;
        RECT 103.400 170.070 103.720 170.130 ;
        RECT 103.875 170.085 104.165 170.130 ;
        RECT 108.015 170.085 108.305 170.315 ;
        RECT 108.460 170.270 108.780 170.330 ;
        RECT 108.935 170.270 109.225 170.315 ;
        RECT 108.460 170.130 109.225 170.270 ;
        RECT 108.460 170.070 108.780 170.130 ;
        RECT 108.935 170.085 109.225 170.130 ;
        RECT 109.380 170.070 109.700 170.330 ;
        RECT 109.855 170.085 110.145 170.315 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 107.095 169.930 107.385 169.975 ;
        RECT 101.560 169.790 103.170 169.930 ;
        RECT 101.560 169.730 101.880 169.790 ;
        RECT 91.070 169.450 92.590 169.590 ;
        RECT 103.030 169.590 103.170 169.790 ;
        RECT 105.790 169.790 107.385 169.930 ;
        RECT 105.790 169.590 105.930 169.790 ;
        RECT 107.095 169.745 107.385 169.790 ;
        RECT 103.030 169.450 105.930 169.590 ;
        RECT 106.620 169.590 106.940 169.650 ;
        RECT 109.380 169.590 109.700 169.650 ;
        RECT 106.620 169.450 109.700 169.590 ;
        RECT 85.890 169.405 86.180 169.450 ;
        RECT 88.670 169.405 88.960 169.450 ;
        RECT 90.530 169.405 90.820 169.450 ;
        RECT 106.620 169.390 106.940 169.450 ;
        RECT 109.380 169.390 109.700 169.450 ;
        RECT 65.680 169.250 66.000 169.310 ;
        RECT 63.010 169.110 66.000 169.250 ;
        RECT 65.680 169.050 66.000 169.110 ;
        RECT 67.520 169.250 67.840 169.310 ;
        RECT 72.595 169.250 72.885 169.295 ;
        RECT 74.880 169.250 75.200 169.310 ;
        RECT 67.520 169.110 75.200 169.250 ;
        RECT 67.520 169.050 67.840 169.110 ;
        RECT 72.595 169.065 72.885 169.110 ;
        RECT 74.880 169.050 75.200 169.110 ;
        RECT 79.955 169.250 80.245 169.295 ;
        RECT 86.840 169.250 87.160 169.310 ;
        RECT 79.955 169.110 87.160 169.250 ;
        RECT 79.955 169.065 80.245 169.110 ;
        RECT 86.840 169.050 87.160 169.110 ;
        RECT 96.515 169.250 96.805 169.295 ;
        RECT 98.340 169.250 98.660 169.310 ;
        RECT 96.515 169.110 98.660 169.250 ;
        RECT 96.515 169.065 96.805 169.110 ;
        RECT 98.340 169.050 98.660 169.110 ;
        RECT 99.260 169.250 99.580 169.310 ;
        RECT 100.655 169.250 100.945 169.295 ;
        RECT 99.260 169.110 100.945 169.250 ;
        RECT 99.260 169.050 99.580 169.110 ;
        RECT 100.655 169.065 100.945 169.110 ;
        RECT 102.020 169.250 102.340 169.310 ;
        RECT 109.930 169.250 110.070 170.085 ;
        RECT 102.020 169.110 110.070 169.250 ;
        RECT 111.235 169.250 111.525 169.295 ;
        RECT 111.680 169.250 112.000 169.310 ;
        RECT 111.235 169.110 112.000 169.250 ;
        RECT 102.020 169.050 102.340 169.110 ;
        RECT 111.235 169.065 111.525 169.110 ;
        RECT 111.680 169.050 112.000 169.110 ;
        RECT 26.970 168.430 113.450 168.910 ;
        RECT 27.500 168.230 27.820 168.290 ;
        RECT 31.655 168.230 31.945 168.275 ;
        RECT 27.500 168.090 31.945 168.230 ;
        RECT 27.500 168.030 27.820 168.090 ;
        RECT 31.655 168.045 31.945 168.090 ;
        RECT 37.635 168.230 37.925 168.275 ;
        RECT 40.840 168.230 41.160 168.290 ;
        RECT 37.635 168.090 41.160 168.230 ;
        RECT 37.635 168.045 37.925 168.090 ;
        RECT 40.840 168.030 41.160 168.090 ;
        RECT 44.150 168.090 51.190 168.230 ;
        RECT 44.150 167.950 44.290 168.090 ;
        RECT 44.060 167.890 44.380 167.950 ;
        RECT 39.550 167.750 44.380 167.890 ;
        RECT 29.355 167.550 29.645 167.595 ;
        RECT 31.640 167.550 31.960 167.610 ;
        RECT 29.355 167.410 31.960 167.550 ;
        RECT 29.355 167.365 29.645 167.410 ;
        RECT 31.640 167.350 31.960 167.410 ;
        RECT 32.560 167.550 32.880 167.610 ;
        RECT 34.875 167.550 35.165 167.595 ;
        RECT 36.240 167.550 36.560 167.610 ;
        RECT 32.560 167.410 36.560 167.550 ;
        RECT 32.560 167.350 32.880 167.410 ;
        RECT 34.875 167.365 35.165 167.410 ;
        RECT 36.240 167.350 36.560 167.410 ;
        RECT 30.260 167.010 30.580 167.270 ;
        RECT 36.700 167.010 37.020 167.270 ;
        RECT 38.080 167.010 38.400 167.270 ;
        RECT 39.550 167.255 39.690 167.750 ;
        RECT 44.060 167.690 44.380 167.750 ;
        RECT 45.870 167.890 46.160 167.935 ;
        RECT 48.650 167.890 48.940 167.935 ;
        RECT 50.510 167.890 50.800 167.935 ;
        RECT 45.870 167.750 50.800 167.890 ;
        RECT 51.050 167.890 51.190 168.090 ;
        RECT 51.420 168.030 51.740 168.290 ;
        RECT 57.415 168.230 57.705 168.275 ;
        RECT 64.760 168.230 65.080 168.290 ;
        RECT 57.415 168.090 65.080 168.230 ;
        RECT 57.415 168.045 57.705 168.090 ;
        RECT 64.760 168.030 65.080 168.090 ;
        RECT 65.680 168.230 66.000 168.290 ;
        RECT 67.060 168.230 67.380 168.290 ;
        RECT 65.680 168.090 67.380 168.230 ;
        RECT 65.680 168.030 66.000 168.090 ;
        RECT 67.060 168.030 67.380 168.090 ;
        RECT 67.520 168.230 67.840 168.290 ;
        RECT 81.780 168.230 82.100 168.290 ;
        RECT 67.520 168.090 68.210 168.230 ;
        RECT 67.520 168.030 67.840 168.090 ;
        RECT 53.260 167.890 53.580 167.950 ;
        RECT 59.700 167.890 60.020 167.950 ;
        RECT 60.620 167.890 60.940 167.950 ;
        RECT 51.050 167.750 60.020 167.890 ;
        RECT 45.870 167.705 46.160 167.750 ;
        RECT 48.650 167.705 48.940 167.750 ;
        RECT 50.510 167.705 50.800 167.750 ;
        RECT 53.260 167.690 53.580 167.750 ;
        RECT 59.700 167.690 60.020 167.750 ;
        RECT 60.250 167.750 60.940 167.890 ;
        RECT 41.300 167.350 41.620 167.610 ;
        RECT 42.680 167.550 43.000 167.610 ;
        RECT 49.135 167.550 49.425 167.595 ;
        RECT 49.580 167.550 49.900 167.610 ;
        RECT 42.680 167.410 48.890 167.550 ;
        RECT 42.680 167.350 43.000 167.410 ;
        RECT 39.015 167.025 39.305 167.255 ;
        RECT 39.475 167.025 39.765 167.255 ;
        RECT 39.935 167.210 40.225 167.255 ;
        RECT 44.520 167.210 44.840 167.270 ;
        RECT 39.935 167.070 44.840 167.210 ;
        RECT 39.935 167.025 40.225 167.070 ;
        RECT 31.195 166.870 31.485 166.915 ;
        RECT 32.100 166.870 32.420 166.930 ;
        RECT 31.195 166.730 32.420 166.870 ;
        RECT 31.195 166.685 31.485 166.730 ;
        RECT 32.100 166.670 32.420 166.730 ;
        RECT 33.955 166.870 34.245 166.915 ;
        RECT 34.860 166.870 35.180 166.930 ;
        RECT 39.090 166.870 39.230 167.025 ;
        RECT 44.520 167.010 44.840 167.070 ;
        RECT 45.870 167.210 46.160 167.255 ;
        RECT 48.750 167.210 48.890 167.410 ;
        RECT 49.135 167.410 49.900 167.550 ;
        RECT 49.135 167.365 49.425 167.410 ;
        RECT 49.580 167.350 49.900 167.410 ;
        RECT 54.640 167.350 54.960 167.610 ;
        RECT 50.975 167.210 51.265 167.255 ;
        RECT 45.870 167.070 48.405 167.210 ;
        RECT 48.750 167.070 51.265 167.210 ;
        RECT 45.870 167.025 46.160 167.070 ;
        RECT 48.190 166.915 48.405 167.070 ;
        RECT 50.975 167.025 51.265 167.070 ;
        RECT 52.800 167.210 53.120 167.270 ;
        RECT 55.560 167.210 55.880 167.270 ;
        RECT 52.800 167.070 55.880 167.210 ;
        RECT 52.800 167.010 53.120 167.070 ;
        RECT 55.560 167.010 55.880 167.070 ;
        RECT 56.495 167.210 56.785 167.255 ;
        RECT 57.400 167.210 57.720 167.270 ;
        RECT 59.240 167.255 59.560 167.270 ;
        RECT 59.790 167.255 59.930 167.690 ;
        RECT 60.250 167.255 60.390 167.750 ;
        RECT 60.620 167.690 60.940 167.750 ;
        RECT 61.080 167.890 61.400 167.950 ;
        RECT 62.015 167.890 62.305 167.935 ;
        RECT 61.080 167.750 62.305 167.890 ;
        RECT 61.080 167.690 61.400 167.750 ;
        RECT 62.015 167.705 62.305 167.750 ;
        RECT 61.540 167.550 61.860 167.610 ;
        RECT 61.540 167.410 64.990 167.550 ;
        RECT 61.540 167.350 61.860 167.410 ;
        RECT 62.920 167.255 63.240 167.270 ;
        RECT 56.495 167.070 57.720 167.210 ;
        RECT 56.495 167.025 56.785 167.070 ;
        RECT 57.400 167.010 57.720 167.070 ;
        RECT 59.155 167.025 59.560 167.255 ;
        RECT 59.715 167.025 60.005 167.255 ;
        RECT 60.175 167.025 60.465 167.255 ;
        RECT 61.065 167.195 61.355 167.255 ;
        RECT 61.630 167.195 62.690 167.210 ;
        RECT 61.065 167.070 62.690 167.195 ;
        RECT 61.065 167.055 61.770 167.070 ;
        RECT 61.065 167.025 61.355 167.055 ;
        RECT 59.240 167.010 59.560 167.025 ;
        RECT 44.010 166.870 44.300 166.915 ;
        RECT 47.270 166.870 47.560 166.915 ;
        RECT 33.955 166.730 39.230 166.870 ;
        RECT 41.390 166.730 47.560 166.870 ;
        RECT 33.955 166.685 34.245 166.730 ;
        RECT 34.860 166.670 35.180 166.730 ;
        RECT 29.800 166.530 30.120 166.590 ;
        RECT 32.560 166.530 32.880 166.590 ;
        RECT 29.800 166.390 32.880 166.530 ;
        RECT 29.800 166.330 30.120 166.390 ;
        RECT 32.560 166.330 32.880 166.390 ;
        RECT 33.495 166.530 33.785 166.575 ;
        RECT 35.780 166.530 36.100 166.590 ;
        RECT 33.495 166.390 36.100 166.530 ;
        RECT 33.495 166.345 33.785 166.390 ;
        RECT 35.780 166.330 36.100 166.390 ;
        RECT 39.000 166.530 39.320 166.590 ;
        RECT 41.390 166.530 41.530 166.730 ;
        RECT 44.010 166.685 44.300 166.730 ;
        RECT 47.270 166.685 47.560 166.730 ;
        RECT 48.190 166.870 48.480 166.915 ;
        RECT 50.050 166.870 50.340 166.915 ;
        RECT 48.190 166.730 50.340 166.870 ;
        RECT 48.190 166.685 48.480 166.730 ;
        RECT 50.050 166.685 50.340 166.730 ;
        RECT 50.500 166.870 50.820 166.930 ;
        RECT 53.275 166.870 53.565 166.915 ;
        RECT 50.500 166.730 53.565 166.870 ;
        RECT 50.500 166.670 50.820 166.730 ;
        RECT 53.275 166.685 53.565 166.730 ;
        RECT 54.640 166.870 54.960 166.930 ;
        RECT 57.875 166.870 58.165 166.915 ;
        RECT 54.640 166.730 58.165 166.870 ;
        RECT 54.640 166.670 54.960 166.730 ;
        RECT 57.875 166.685 58.165 166.730 ;
        RECT 42.220 166.575 42.540 166.590 ;
        RECT 39.000 166.390 41.530 166.530 ;
        RECT 39.000 166.330 39.320 166.390 ;
        RECT 42.005 166.345 42.540 166.575 ;
        RECT 42.220 166.330 42.540 166.345 ;
        RECT 44.520 166.530 44.840 166.590 ;
        RECT 51.420 166.530 51.740 166.590 ;
        RECT 44.520 166.390 51.740 166.530 ;
        RECT 44.520 166.330 44.840 166.390 ;
        RECT 51.420 166.330 51.740 166.390 ;
        RECT 52.340 166.530 52.660 166.590 ;
        RECT 53.735 166.530 54.025 166.575 ;
        RECT 52.340 166.390 54.025 166.530 ;
        RECT 52.340 166.330 52.660 166.390 ;
        RECT 53.735 166.345 54.025 166.390 ;
        RECT 55.560 166.530 55.880 166.590 ;
        RECT 62.550 166.530 62.690 167.070 ;
        RECT 62.920 167.025 63.455 167.255 ;
        RECT 62.920 167.010 63.240 167.025 ;
        RECT 63.840 167.010 64.160 167.270 ;
        RECT 64.420 167.195 64.710 167.240 ;
        RECT 64.850 167.195 64.990 167.410 ;
        RECT 67.520 167.350 67.840 167.610 ;
        RECT 64.420 167.055 64.990 167.195 ;
        RECT 64.420 167.010 64.710 167.055 ;
        RECT 65.235 167.025 65.525 167.255 ;
        RECT 65.680 167.210 66.000 167.270 ;
        RECT 66.155 167.210 66.445 167.255 ;
        RECT 68.070 167.210 68.210 168.090 ;
        RECT 69.910 168.090 82.100 168.230 ;
        RECT 69.910 167.255 70.050 168.090 ;
        RECT 81.780 168.030 82.100 168.090 ;
        RECT 82.240 168.230 82.560 168.290 ;
        RECT 85.935 168.230 86.225 168.275 ;
        RECT 82.240 168.090 86.225 168.230 ;
        RECT 82.240 168.030 82.560 168.090 ;
        RECT 85.935 168.045 86.225 168.090 ;
        RECT 91.915 168.230 92.205 168.275 ;
        RECT 93.280 168.230 93.600 168.290 ;
        RECT 91.915 168.090 93.600 168.230 ;
        RECT 91.915 168.045 92.205 168.090 ;
        RECT 93.280 168.030 93.600 168.090 ;
        RECT 94.660 168.230 94.980 168.290 ;
        RECT 95.595 168.230 95.885 168.275 ;
        RECT 94.660 168.090 95.885 168.230 ;
        RECT 94.660 168.030 94.980 168.090 ;
        RECT 95.595 168.045 95.885 168.090 ;
        RECT 97.420 168.230 97.740 168.290 ;
        RECT 102.480 168.230 102.800 168.290 ;
        RECT 106.620 168.230 106.940 168.290 ;
        RECT 97.420 168.090 106.940 168.230 ;
        RECT 97.420 168.030 97.740 168.090 ;
        RECT 102.480 168.030 102.800 168.090 ;
        RECT 106.620 168.030 106.940 168.090 ;
        RECT 70.280 167.890 70.600 167.950 ;
        RECT 75.800 167.890 76.120 167.950 ;
        RECT 70.280 167.750 76.120 167.890 ;
        RECT 70.280 167.690 70.600 167.750 ;
        RECT 72.135 167.550 72.425 167.595 ;
        RECT 73.040 167.550 73.360 167.610 ;
        RECT 72.135 167.410 73.360 167.550 ;
        RECT 72.135 167.365 72.425 167.410 ;
        RECT 73.040 167.350 73.360 167.410 ;
        RECT 68.915 167.210 69.205 167.255 ;
        RECT 65.680 167.070 66.445 167.210 ;
        RECT 65.310 166.870 65.450 167.025 ;
        RECT 65.680 167.010 66.000 167.070 ;
        RECT 66.155 167.025 66.445 167.070 ;
        RECT 66.690 167.070 69.205 167.210 ;
        RECT 66.690 166.870 66.830 167.070 ;
        RECT 68.915 167.025 69.205 167.070 ;
        RECT 69.835 167.025 70.125 167.255 ;
        RECT 70.280 167.010 70.600 167.270 ;
        RECT 70.755 167.210 71.045 167.255 ;
        RECT 71.660 167.210 71.980 167.270 ;
        RECT 73.960 167.210 74.280 167.270 ;
        RECT 74.510 167.255 74.650 167.750 ;
        RECT 75.800 167.690 76.120 167.750 ;
        RECT 80.370 167.890 80.660 167.935 ;
        RECT 83.150 167.890 83.440 167.935 ;
        RECT 85.010 167.890 85.300 167.935 ;
        RECT 80.370 167.750 85.300 167.890 ;
        RECT 80.370 167.705 80.660 167.750 ;
        RECT 83.150 167.705 83.440 167.750 ;
        RECT 85.010 167.705 85.300 167.750 ;
        RECT 89.140 167.890 89.460 167.950 ;
        RECT 97.880 167.890 98.200 167.950 ;
        RECT 89.140 167.750 98.200 167.890 ;
        RECT 89.140 167.690 89.460 167.750 ;
        RECT 97.880 167.690 98.200 167.750 ;
        RECT 98.800 167.690 99.120 167.950 ;
        RECT 99.720 167.890 100.040 167.950 ;
        RECT 99.350 167.750 100.040 167.890 ;
        RECT 79.940 167.550 80.260 167.610 ;
        RECT 74.970 167.410 80.260 167.550 ;
        RECT 74.970 167.255 75.110 167.410 ;
        RECT 79.940 167.350 80.260 167.410 ;
        RECT 88.695 167.550 88.985 167.595 ;
        RECT 91.440 167.550 91.760 167.610 ;
        RECT 88.695 167.410 91.760 167.550 ;
        RECT 88.695 167.365 88.985 167.410 ;
        RECT 70.755 167.070 74.280 167.210 ;
        RECT 70.755 167.025 71.045 167.070 ;
        RECT 65.310 166.730 66.830 166.870 ;
        RECT 67.060 166.870 67.380 166.930 ;
        RECT 70.830 166.870 70.970 167.025 ;
        RECT 71.660 167.010 71.980 167.070 ;
        RECT 73.960 167.010 74.280 167.070 ;
        RECT 74.435 167.025 74.725 167.255 ;
        RECT 74.895 167.025 75.185 167.255 ;
        RECT 75.815 167.025 76.105 167.255 ;
        RECT 80.370 167.210 80.660 167.255 ;
        RECT 83.160 167.210 83.480 167.270 ;
        RECT 83.635 167.210 83.925 167.255 ;
        RECT 80.370 167.070 82.905 167.210 ;
        RECT 80.370 167.025 80.660 167.070 ;
        RECT 67.060 166.730 70.970 166.870 ;
        RECT 65.310 166.530 65.450 166.730 ;
        RECT 67.060 166.670 67.380 166.730 ;
        RECT 72.580 166.670 72.900 166.930 ;
        RECT 55.560 166.390 65.450 166.530 ;
        RECT 73.960 166.530 74.280 166.590 ;
        RECT 74.510 166.530 74.650 167.025 ;
        RECT 75.890 166.870 76.030 167.025 ;
        RECT 74.970 166.730 76.030 166.870 ;
        RECT 77.180 166.870 77.500 166.930 ;
        RECT 82.690 166.915 82.905 167.070 ;
        RECT 83.160 167.070 83.925 167.210 ;
        RECT 83.160 167.010 83.480 167.070 ;
        RECT 83.635 167.025 83.925 167.070 ;
        RECT 85.000 167.210 85.320 167.270 ;
        RECT 85.475 167.210 85.765 167.255 ;
        RECT 85.000 167.070 85.765 167.210 ;
        RECT 85.000 167.010 85.320 167.070 ;
        RECT 85.475 167.025 85.765 167.070 ;
        RECT 86.840 167.010 87.160 167.270 ;
        RECT 78.510 166.870 78.800 166.915 ;
        RECT 81.770 166.870 82.060 166.915 ;
        RECT 77.180 166.730 82.060 166.870 ;
        RECT 74.970 166.590 75.110 166.730 ;
        RECT 77.180 166.670 77.500 166.730 ;
        RECT 78.510 166.685 78.800 166.730 ;
        RECT 81.770 166.685 82.060 166.730 ;
        RECT 82.690 166.870 82.980 166.915 ;
        RECT 84.550 166.870 84.840 166.915 ;
        RECT 88.770 166.870 88.910 167.365 ;
        RECT 91.440 167.350 91.760 167.410 ;
        RECT 95.135 167.550 95.425 167.595 ;
        RECT 98.890 167.550 99.030 167.690 ;
        RECT 95.135 167.410 99.030 167.550 ;
        RECT 95.135 167.365 95.425 167.410 ;
        RECT 89.140 167.010 89.460 167.270 ;
        RECT 89.615 167.210 89.905 167.255 ;
        RECT 91.900 167.210 92.220 167.270 ;
        RECT 89.615 167.070 92.220 167.210 ;
        RECT 89.615 167.025 89.905 167.070 ;
        RECT 91.900 167.010 92.220 167.070 ;
        RECT 96.975 167.025 97.265 167.255 ;
        RECT 82.690 166.730 84.840 166.870 ;
        RECT 82.690 166.685 82.980 166.730 ;
        RECT 84.550 166.685 84.840 166.730 ;
        RECT 85.090 166.730 88.910 166.870 ;
        RECT 90.980 166.870 91.300 166.930 ;
        RECT 95.580 166.870 95.900 166.930 ;
        RECT 97.050 166.870 97.190 167.025 ;
        RECT 97.420 167.010 97.740 167.270 ;
        RECT 97.970 167.255 98.110 167.410 ;
        RECT 97.895 167.025 98.185 167.255 ;
        RECT 98.800 167.210 99.120 167.270 ;
        RECT 99.350 167.210 99.490 167.750 ;
        RECT 99.720 167.690 100.040 167.750 ;
        RECT 105.355 167.890 105.645 167.935 ;
        RECT 108.475 167.890 108.765 167.935 ;
        RECT 110.365 167.890 110.655 167.935 ;
        RECT 105.355 167.750 110.655 167.890 ;
        RECT 105.355 167.705 105.645 167.750 ;
        RECT 108.475 167.705 108.765 167.750 ;
        RECT 110.365 167.705 110.655 167.750 ;
        RECT 111.220 167.350 111.540 167.610 ;
        RECT 98.800 167.070 99.490 167.210 ;
        RECT 99.735 167.210 100.025 167.255 ;
        RECT 100.180 167.210 100.500 167.270 ;
        RECT 99.735 167.070 100.500 167.210 ;
        RECT 98.800 167.010 99.120 167.070 ;
        RECT 99.735 167.025 100.025 167.070 ;
        RECT 100.180 167.010 100.500 167.070 ;
        RECT 101.115 167.210 101.405 167.255 ;
        RECT 102.940 167.210 103.260 167.270 ;
        RECT 101.115 167.070 103.260 167.210 ;
        RECT 101.115 167.025 101.405 167.070 ;
        RECT 102.940 167.010 103.260 167.070 ;
        RECT 90.980 166.730 97.190 166.870 ;
        RECT 101.560 166.870 101.880 166.930 ;
        RECT 104.275 166.915 104.565 167.230 ;
        RECT 105.355 167.210 105.645 167.255 ;
        RECT 108.935 167.210 109.225 167.255 ;
        RECT 110.770 167.210 111.060 167.255 ;
        RECT 105.355 167.070 111.060 167.210 ;
        RECT 105.355 167.025 105.645 167.070 ;
        RECT 108.935 167.025 109.225 167.070 ;
        RECT 110.770 167.025 111.060 167.070 ;
        RECT 103.975 166.870 104.565 166.915 ;
        RECT 107.215 166.870 107.865 166.915 ;
        RECT 101.560 166.730 107.865 166.870 ;
        RECT 73.960 166.390 74.650 166.530 ;
        RECT 55.560 166.330 55.880 166.390 ;
        RECT 73.960 166.330 74.280 166.390 ;
        RECT 74.880 166.330 75.200 166.590 ;
        RECT 76.720 166.575 77.040 166.590 ;
        RECT 76.505 166.345 77.040 166.575 ;
        RECT 76.720 166.330 77.040 166.345 ;
        RECT 79.020 166.530 79.340 166.590 ;
        RECT 85.090 166.530 85.230 166.730 ;
        RECT 90.980 166.670 91.300 166.730 ;
        RECT 95.580 166.670 95.900 166.730 ;
        RECT 101.560 166.670 101.880 166.730 ;
        RECT 103.975 166.685 104.265 166.730 ;
        RECT 107.215 166.685 107.865 166.730 ;
        RECT 109.855 166.870 110.145 166.915 ;
        RECT 111.680 166.870 112.000 166.930 ;
        RECT 109.855 166.730 112.000 166.870 ;
        RECT 109.855 166.685 110.145 166.730 ;
        RECT 111.680 166.670 112.000 166.730 ;
        RECT 79.020 166.390 85.230 166.530 ;
        RECT 91.455 166.530 91.745 166.575 ;
        RECT 100.180 166.530 100.500 166.590 ;
        RECT 91.455 166.390 100.500 166.530 ;
        RECT 79.020 166.330 79.340 166.390 ;
        RECT 91.455 166.345 91.745 166.390 ;
        RECT 100.180 166.330 100.500 166.390 ;
        RECT 102.020 166.530 102.340 166.590 ;
        RECT 102.495 166.530 102.785 166.575 ;
        RECT 102.020 166.390 102.785 166.530 ;
        RECT 102.020 166.330 102.340 166.390 ;
        RECT 102.495 166.345 102.785 166.390 ;
        RECT 26.970 165.710 113.450 166.190 ;
        RECT 29.800 165.510 30.120 165.570 ;
        RECT 32.560 165.510 32.880 165.570 ;
        RECT 39.000 165.510 39.320 165.570 ;
        RECT 40.395 165.510 40.685 165.555 ;
        RECT 29.800 165.370 37.390 165.510 ;
        RECT 29.800 165.310 30.120 165.370 ;
        RECT 32.560 165.310 32.880 165.370 ;
        RECT 27.960 165.170 28.280 165.230 ;
        RECT 30.670 165.170 30.960 165.215 ;
        RECT 33.930 165.170 34.220 165.215 ;
        RECT 27.960 165.030 34.220 165.170 ;
        RECT 27.960 164.970 28.280 165.030 ;
        RECT 30.670 164.985 30.960 165.030 ;
        RECT 33.930 164.985 34.220 165.030 ;
        RECT 34.850 165.170 35.140 165.215 ;
        RECT 36.710 165.170 37.000 165.215 ;
        RECT 34.850 165.030 37.000 165.170 ;
        RECT 37.250 165.170 37.390 165.370 ;
        RECT 39.000 165.370 40.685 165.510 ;
        RECT 39.000 165.310 39.320 165.370 ;
        RECT 40.395 165.325 40.685 165.370 ;
        RECT 42.220 165.510 42.540 165.570 ;
        RECT 48.215 165.510 48.505 165.555 ;
        RECT 50.500 165.510 50.820 165.570 ;
        RECT 56.940 165.510 57.260 165.570 ;
        RECT 69.820 165.510 70.140 165.570 ;
        RECT 42.220 165.370 47.970 165.510 ;
        RECT 42.220 165.310 42.540 165.370 ;
        RECT 41.300 165.170 41.620 165.230 ;
        RECT 44.980 165.170 45.300 165.230 ;
        RECT 37.250 165.030 41.070 165.170 ;
        RECT 34.850 164.985 35.140 165.030 ;
        RECT 36.710 164.985 37.000 165.030 ;
        RECT 32.530 164.830 32.820 164.875 ;
        RECT 34.850 164.830 35.065 164.985 ;
        RECT 32.530 164.690 35.065 164.830 ;
        RECT 35.795 164.830 36.085 164.875 ;
        RECT 38.080 164.830 38.400 164.890 ;
        RECT 35.795 164.690 38.400 164.830 ;
        RECT 32.530 164.645 32.820 164.690 ;
        RECT 35.795 164.645 36.085 164.690 ;
        RECT 38.080 164.630 38.400 164.690 ;
        RECT 39.000 164.630 39.320 164.890 ;
        RECT 36.240 164.490 36.560 164.550 ;
        RECT 37.635 164.490 37.925 164.535 ;
        RECT 40.380 164.490 40.700 164.550 ;
        RECT 36.240 164.350 40.700 164.490 ;
        RECT 40.930 164.490 41.070 165.030 ;
        RECT 41.300 165.030 45.300 165.170 ;
        RECT 47.830 165.170 47.970 165.370 ;
        RECT 48.215 165.370 50.820 165.510 ;
        RECT 48.215 165.325 48.505 165.370 ;
        RECT 50.500 165.310 50.820 165.370 ;
        RECT 52.890 165.370 56.710 165.510 ;
        RECT 52.340 165.170 52.660 165.230 ;
        RECT 47.830 165.030 52.660 165.170 ;
        RECT 41.300 164.970 41.620 165.030 ;
        RECT 44.980 164.970 45.300 165.030 ;
        RECT 52.340 164.970 52.660 165.030 ;
        RECT 42.695 164.830 42.985 164.875 ;
        RECT 44.060 164.830 44.380 164.890 ;
        RECT 42.695 164.690 44.380 164.830 ;
        RECT 42.695 164.645 42.985 164.690 ;
        RECT 44.060 164.630 44.380 164.690 ;
        RECT 50.055 164.645 50.345 164.875 ;
        RECT 51.420 164.830 51.740 164.890 ;
        RECT 52.890 164.875 53.030 165.370 ;
        RECT 54.180 165.170 54.500 165.230 ;
        RECT 56.570 165.170 56.710 165.370 ;
        RECT 56.940 165.370 82.930 165.510 ;
        RECT 56.940 165.310 57.260 165.370 ;
        RECT 69.820 165.310 70.140 165.370 ;
        RECT 59.240 165.170 59.560 165.230 ;
        RECT 61.540 165.215 61.860 165.230 ;
        RECT 54.180 165.030 56.250 165.170 ;
        RECT 56.570 165.030 59.560 165.170 ;
        RECT 54.180 164.970 54.500 165.030 ;
        RECT 52.815 164.830 53.105 164.875 ;
        RECT 51.420 164.690 53.105 164.830 ;
        RECT 43.155 164.490 43.445 164.535 ;
        RECT 40.930 164.350 43.445 164.490 ;
        RECT 36.240 164.290 36.560 164.350 ;
        RECT 37.635 164.305 37.925 164.350 ;
        RECT 40.380 164.290 40.700 164.350 ;
        RECT 43.155 164.305 43.445 164.350 ;
        RECT 45.455 164.490 45.745 164.535 ;
        RECT 45.455 164.350 48.890 164.490 ;
        RECT 45.455 164.305 45.745 164.350 ;
        RECT 32.530 164.150 32.820 164.195 ;
        RECT 35.310 164.150 35.600 164.195 ;
        RECT 37.170 164.150 37.460 164.195 ;
        RECT 32.530 164.010 37.460 164.150 ;
        RECT 32.530 163.965 32.820 164.010 ;
        RECT 35.310 163.965 35.600 164.010 ;
        RECT 37.170 163.965 37.460 164.010 ;
        RECT 38.080 163.950 38.400 164.210 ;
        RECT 44.980 164.150 45.300 164.210 ;
        RECT 48.200 164.150 48.520 164.210 ;
        RECT 44.980 164.010 48.520 164.150 ;
        RECT 44.980 163.950 45.300 164.010 ;
        RECT 48.200 163.950 48.520 164.010 ;
        RECT 28.665 163.810 28.955 163.855 ;
        RECT 33.020 163.810 33.340 163.870 ;
        RECT 35.780 163.810 36.100 163.870 ;
        RECT 46.820 163.810 47.140 163.870 ;
        RECT 28.665 163.670 47.140 163.810 ;
        RECT 48.750 163.810 48.890 164.350 ;
        RECT 49.120 164.290 49.440 164.550 ;
        RECT 50.130 164.490 50.270 164.645 ;
        RECT 51.420 164.630 51.740 164.690 ;
        RECT 52.815 164.645 53.105 164.690 ;
        RECT 53.260 164.630 53.580 164.890 ;
        RECT 53.720 164.630 54.040 164.890 ;
        RECT 54.655 164.830 54.945 164.875 ;
        RECT 55.115 164.830 55.405 164.875 ;
        RECT 55.560 164.830 55.880 164.890 ;
        RECT 56.110 164.875 56.250 165.030 ;
        RECT 57.030 164.875 57.170 165.030 ;
        RECT 59.240 164.970 59.560 165.030 ;
        RECT 61.490 165.170 61.860 165.215 ;
        RECT 64.750 165.170 65.040 165.215 ;
        RECT 61.490 165.030 65.040 165.170 ;
        RECT 61.490 164.985 61.860 165.030 ;
        RECT 64.750 164.985 65.040 165.030 ;
        RECT 65.670 165.170 65.960 165.215 ;
        RECT 67.530 165.170 67.820 165.215 ;
        RECT 65.670 165.030 67.820 165.170 ;
        RECT 65.670 164.985 65.960 165.030 ;
        RECT 67.530 164.985 67.820 165.030 ;
        RECT 61.540 164.970 61.860 164.985 ;
        RECT 54.655 164.690 55.880 164.830 ;
        RECT 54.655 164.645 54.945 164.690 ;
        RECT 55.115 164.645 55.405 164.690 ;
        RECT 55.560 164.630 55.880 164.690 ;
        RECT 56.035 164.645 56.325 164.875 ;
        RECT 56.495 164.645 56.785 164.875 ;
        RECT 56.955 164.645 57.245 164.875 ;
        RECT 63.350 164.830 63.640 164.875 ;
        RECT 65.670 164.830 65.885 164.985 ;
        RECT 70.740 164.970 71.060 165.230 ;
        RECT 73.500 165.170 73.820 165.230 ;
        RECT 72.670 165.030 73.820 165.170 ;
        RECT 63.350 164.690 65.885 164.830 ;
        RECT 63.350 164.645 63.640 164.690 ;
        RECT 51.880 164.490 52.200 164.550 ;
        RECT 50.130 164.350 52.200 164.490 ;
        RECT 51.880 164.290 52.200 164.350 ;
        RECT 53.810 164.150 53.950 164.630 ;
        RECT 54.180 164.490 54.500 164.550 ;
        RECT 56.570 164.490 56.710 164.645 ;
        RECT 68.440 164.630 68.760 164.890 ;
        RECT 70.295 164.830 70.585 164.875 ;
        RECT 71.200 164.830 71.520 164.890 ;
        RECT 70.295 164.690 71.520 164.830 ;
        RECT 70.295 164.645 70.585 164.690 ;
        RECT 71.200 164.630 71.520 164.690 ;
        RECT 71.660 164.830 71.980 164.890 ;
        RECT 72.670 164.875 72.810 165.030 ;
        RECT 73.500 164.970 73.820 165.030 ;
        RECT 76.720 165.170 77.040 165.230 ;
        RECT 79.480 165.170 79.800 165.230 ;
        RECT 76.720 165.030 79.800 165.170 ;
        RECT 82.790 165.170 82.930 165.370 ;
        RECT 83.160 165.310 83.480 165.570 ;
        RECT 85.015 165.510 85.305 165.555 ;
        RECT 85.460 165.510 85.780 165.570 ;
        RECT 85.015 165.370 85.780 165.510 ;
        RECT 85.015 165.325 85.305 165.370 ;
        RECT 85.460 165.310 85.780 165.370 ;
        RECT 92.820 165.510 93.140 165.570 ;
        RECT 95.120 165.510 95.440 165.570 ;
        RECT 92.820 165.370 95.440 165.510 ;
        RECT 92.820 165.310 93.140 165.370 ;
        RECT 95.120 165.310 95.440 165.370 ;
        RECT 97.880 165.510 98.200 165.570 ;
        RECT 100.655 165.510 100.945 165.555 ;
        RECT 110.300 165.510 110.620 165.570 ;
        RECT 97.880 165.370 100.945 165.510 ;
        RECT 97.880 165.310 98.200 165.370 ;
        RECT 100.655 165.325 100.945 165.370 ;
        RECT 108.550 165.370 110.620 165.510 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 97.420 165.170 97.740 165.230 ;
        RECT 82.790 165.030 97.740 165.170 ;
        RECT 76.720 164.970 77.040 165.030 ;
        RECT 79.480 164.970 79.800 165.030 ;
        RECT 72.135 164.830 72.425 164.875 ;
        RECT 71.660 164.690 72.425 164.830 ;
        RECT 71.660 164.630 71.980 164.690 ;
        RECT 72.135 164.645 72.425 164.690 ;
        RECT 72.595 164.645 72.885 164.875 ;
        RECT 73.055 164.645 73.345 164.875 ;
        RECT 73.975 164.830 74.265 164.875 ;
        RECT 74.880 164.830 75.200 164.890 ;
        RECT 73.975 164.690 75.200 164.830 ;
        RECT 73.975 164.645 74.265 164.690 ;
        RECT 54.180 164.350 56.710 164.490 ;
        RECT 64.760 164.490 65.080 164.550 ;
        RECT 66.615 164.490 66.905 164.535 ;
        RECT 64.760 164.350 66.905 164.490 ;
        RECT 54.180 164.290 54.500 164.350 ;
        RECT 64.760 164.290 65.080 164.350 ;
        RECT 66.615 164.305 66.905 164.350 ;
        RECT 67.060 164.490 67.380 164.550 ;
        RECT 73.130 164.490 73.270 164.645 ;
        RECT 74.880 164.630 75.200 164.690 ;
        RECT 75.340 164.830 75.660 164.890 ;
        RECT 76.275 164.830 76.565 164.875 ;
        RECT 75.340 164.690 76.565 164.830 ;
        RECT 75.340 164.630 75.660 164.690 ;
        RECT 76.275 164.645 76.565 164.690 ;
        RECT 76.810 164.490 76.950 164.970 ;
        RECT 77.180 164.630 77.500 164.890 ;
        RECT 77.640 164.630 77.960 164.890 ;
        RECT 79.940 164.830 80.260 164.890 ;
        RECT 80.860 164.830 81.180 164.890 ;
        RECT 79.940 164.690 81.180 164.830 ;
        RECT 83.620 164.830 83.940 164.890 ;
        RECT 84.555 164.830 84.845 164.875 ;
        RECT 85.460 164.830 85.780 164.890 ;
        RECT 79.940 164.630 80.260 164.690 ;
        RECT 80.860 164.630 81.180 164.690 ;
        RECT 82.255 164.565 82.545 164.795 ;
        RECT 83.620 164.690 85.780 164.830 ;
        RECT 83.620 164.630 83.940 164.690 ;
        RECT 84.555 164.645 84.845 164.690 ;
        RECT 85.460 164.630 85.780 164.690 ;
        RECT 85.920 164.630 86.240 164.890 ;
        RECT 88.220 164.630 88.540 164.890 ;
        RECT 89.600 164.630 89.920 164.890 ;
        RECT 91.440 164.630 91.760 164.890 ;
        RECT 91.990 164.875 92.130 165.030 ;
        RECT 91.915 164.645 92.205 164.875 ;
        RECT 92.360 164.630 92.680 164.890 ;
        RECT 93.295 164.645 93.585 164.875 ;
        RECT 94.200 164.830 94.520 164.890 ;
        RECT 95.670 164.875 95.810 165.030 ;
        RECT 97.420 164.970 97.740 165.030 ;
        RECT 104.730 165.170 105.020 165.215 ;
        RECT 107.990 165.170 108.280 165.215 ;
        RECT 108.550 165.170 108.690 165.370 ;
        RECT 110.300 165.310 110.620 165.370 ;
        RECT 104.730 165.030 108.690 165.170 ;
        RECT 108.910 165.170 109.200 165.215 ;
        RECT 110.770 165.170 111.060 165.215 ;
        RECT 108.910 165.030 111.060 165.170 ;
        RECT 104.730 164.985 105.020 165.030 ;
        RECT 107.990 164.985 108.280 165.030 ;
        RECT 108.910 164.985 109.200 165.030 ;
        RECT 110.770 164.985 111.060 165.030 ;
        RECT 95.135 164.830 95.425 164.875 ;
        RECT 94.200 164.690 95.425 164.830 ;
        RECT 67.060 164.350 71.890 164.490 ;
        RECT 73.130 164.350 76.950 164.490 ;
        RECT 67.060 164.290 67.380 164.350 ;
        RECT 50.130 164.010 53.950 164.150 ;
        RECT 63.350 164.150 63.640 164.195 ;
        RECT 66.130 164.150 66.420 164.195 ;
        RECT 67.990 164.150 68.280 164.195 ;
        RECT 63.350 164.010 68.280 164.150 ;
        RECT 50.130 163.810 50.270 164.010 ;
        RECT 63.350 163.965 63.640 164.010 ;
        RECT 66.130 163.965 66.420 164.010 ;
        RECT 67.990 163.965 68.280 164.010 ;
        RECT 69.375 164.150 69.665 164.195 ;
        RECT 71.200 164.150 71.520 164.210 ;
        RECT 69.375 164.010 71.520 164.150 ;
        RECT 71.750 164.150 71.890 164.350 ;
        RECT 78.560 164.290 78.880 164.550 ;
        RECT 81.795 164.150 82.085 164.195 ;
        RECT 82.330 164.150 82.470 164.565 ;
        RECT 89.155 164.490 89.445 164.535 ;
        RECT 92.820 164.490 93.140 164.550 ;
        RECT 71.750 164.010 72.350 164.150 ;
        RECT 69.375 163.965 69.665 164.010 ;
        RECT 71.200 163.950 71.520 164.010 ;
        RECT 48.750 163.670 50.270 163.810 ;
        RECT 50.500 163.810 50.820 163.870 ;
        RECT 50.975 163.810 51.265 163.855 ;
        RECT 50.500 163.670 51.265 163.810 ;
        RECT 28.665 163.625 28.955 163.670 ;
        RECT 33.020 163.610 33.340 163.670 ;
        RECT 35.780 163.610 36.100 163.670 ;
        RECT 46.820 163.610 47.140 163.670 ;
        RECT 50.500 163.610 50.820 163.670 ;
        RECT 50.975 163.625 51.265 163.670 ;
        RECT 51.420 163.610 51.740 163.870 ;
        RECT 58.320 163.610 58.640 163.870 ;
        RECT 59.700 163.855 60.020 163.870 ;
        RECT 59.485 163.625 60.020 163.855 ;
        RECT 72.210 163.810 72.350 164.010 ;
        RECT 81.795 164.010 82.470 164.150 ;
        RECT 86.470 164.350 88.910 164.490 ;
        RECT 81.795 163.965 82.085 164.010 ;
        RECT 75.355 163.810 75.645 163.855 ;
        RECT 86.470 163.810 86.610 164.350 ;
        RECT 87.300 163.950 87.620 164.210 ;
        RECT 88.770 164.150 88.910 164.350 ;
        RECT 89.155 164.350 93.140 164.490 ;
        RECT 89.155 164.305 89.445 164.350 ;
        RECT 92.820 164.290 93.140 164.350 ;
        RECT 93.370 164.490 93.510 164.645 ;
        RECT 94.200 164.630 94.520 164.690 ;
        RECT 95.135 164.645 95.425 164.690 ;
        RECT 95.595 164.645 95.885 164.875 ;
        RECT 96.040 164.630 96.360 164.890 ;
        RECT 96.975 164.645 97.265 164.875 ;
        RECT 97.050 164.490 97.190 164.645 ;
        RECT 98.340 164.630 98.660 164.890 ;
        RECT 99.720 164.630 100.040 164.890 ;
        RECT 100.180 164.830 100.500 164.890 ;
        RECT 101.575 164.830 101.865 164.875 ;
        RECT 100.180 164.690 101.865 164.830 ;
        RECT 100.180 164.630 100.500 164.690 ;
        RECT 101.575 164.645 101.865 164.690 ;
        RECT 106.590 164.830 106.880 164.875 ;
        RECT 108.910 164.830 109.125 164.985 ;
        RECT 106.590 164.690 109.125 164.830 ;
        RECT 111.220 164.830 111.540 164.890 ;
        RECT 111.695 164.830 111.985 164.875 ;
        RECT 111.220 164.690 111.985 164.830 ;
        RECT 106.590 164.645 106.880 164.690 ;
        RECT 111.220 164.630 111.540 164.690 ;
        RECT 111.695 164.645 111.985 164.690 ;
        RECT 98.800 164.490 99.120 164.550 ;
        RECT 93.370 164.350 99.120 164.490 ;
        RECT 93.370 164.150 93.510 164.350 ;
        RECT 98.800 164.290 99.120 164.350 ;
        RECT 99.275 164.490 99.565 164.535 ;
        RECT 106.160 164.490 106.480 164.550 ;
        RECT 99.275 164.350 106.480 164.490 ;
        RECT 99.275 164.305 99.565 164.350 ;
        RECT 106.160 164.290 106.480 164.350 ;
        RECT 109.855 164.490 110.145 164.535 ;
        RECT 110.300 164.490 110.620 164.550 ;
        RECT 109.855 164.350 110.620 164.490 ;
        RECT 109.855 164.305 110.145 164.350 ;
        RECT 110.300 164.290 110.620 164.350 ;
        RECT 88.770 164.010 93.510 164.150 ;
        RECT 106.590 164.150 106.880 164.195 ;
        RECT 109.370 164.150 109.660 164.195 ;
        RECT 111.230 164.150 111.520 164.195 ;
        RECT 106.590 164.010 111.520 164.150 ;
        RECT 106.590 163.965 106.880 164.010 ;
        RECT 109.370 163.965 109.660 164.010 ;
        RECT 111.230 163.965 111.520 164.010 ;
        RECT 72.210 163.670 86.610 163.810 ;
        RECT 86.855 163.810 87.145 163.855 ;
        RECT 88.680 163.810 89.000 163.870 ;
        RECT 86.855 163.670 89.000 163.810 ;
        RECT 75.355 163.625 75.645 163.670 ;
        RECT 86.855 163.625 87.145 163.670 ;
        RECT 59.700 163.610 60.020 163.625 ;
        RECT 88.680 163.610 89.000 163.670 ;
        RECT 89.140 163.610 89.460 163.870 ;
        RECT 90.075 163.810 90.365 163.855 ;
        RECT 90.980 163.810 91.300 163.870 ;
        RECT 90.075 163.670 91.300 163.810 ;
        RECT 90.075 163.625 90.365 163.670 ;
        RECT 90.980 163.610 91.300 163.670 ;
        RECT 93.755 163.810 94.045 163.855 ;
        RECT 94.660 163.810 94.980 163.870 ;
        RECT 93.755 163.670 94.980 163.810 ;
        RECT 93.755 163.625 94.045 163.670 ;
        RECT 94.660 163.610 94.980 163.670 ;
        RECT 97.420 163.610 97.740 163.870 ;
        RECT 98.340 163.610 98.660 163.870 ;
        RECT 98.800 163.810 99.120 163.870 ;
        RECT 102.020 163.810 102.340 163.870 ;
        RECT 98.800 163.670 102.340 163.810 ;
        RECT 98.800 163.610 99.120 163.670 ;
        RECT 102.020 163.610 102.340 163.670 ;
        RECT 102.725 163.810 103.015 163.855 ;
        RECT 104.780 163.810 105.100 163.870 ;
        RECT 102.725 163.670 105.100 163.810 ;
        RECT 102.725 163.625 103.015 163.670 ;
        RECT 104.780 163.610 105.100 163.670 ;
        RECT 26.970 162.990 113.450 163.470 ;
        RECT 35.335 162.790 35.625 162.835 ;
        RECT 39.000 162.790 39.320 162.850 ;
        RECT 35.335 162.650 39.320 162.790 ;
        RECT 35.335 162.605 35.625 162.650 ;
        RECT 39.000 162.590 39.320 162.650 ;
        RECT 39.460 162.790 39.780 162.850 ;
        RECT 41.760 162.790 42.080 162.850 ;
        RECT 39.460 162.650 47.510 162.790 ;
        RECT 39.460 162.590 39.780 162.650 ;
        RECT 41.760 162.590 42.080 162.650 ;
        RECT 36.720 162.450 37.010 162.495 ;
        RECT 38.580 162.450 38.870 162.495 ;
        RECT 41.360 162.450 41.650 162.495 ;
        RECT 36.720 162.310 41.650 162.450 ;
        RECT 36.720 162.265 37.010 162.310 ;
        RECT 38.580 162.265 38.870 162.310 ;
        RECT 41.360 162.265 41.650 162.310 ;
        RECT 26.120 162.110 26.440 162.170 ;
        RECT 31.180 162.110 31.500 162.170 ;
        RECT 26.120 161.970 31.500 162.110 ;
        RECT 26.120 161.910 26.440 161.970 ;
        RECT 31.180 161.910 31.500 161.970 ;
        RECT 32.560 161.910 32.880 162.170 ;
        RECT 33.020 161.910 33.340 162.170 ;
        RECT 36.240 161.910 36.560 162.170 ;
        RECT 37.620 162.110 37.940 162.170 ;
        RECT 38.095 162.110 38.385 162.155 ;
        RECT 37.620 161.970 38.385 162.110 ;
        RECT 37.620 161.910 37.940 161.970 ;
        RECT 38.095 161.925 38.385 161.970 ;
        RECT 39.000 162.110 39.320 162.170 ;
        RECT 45.915 162.110 46.205 162.155 ;
        RECT 39.000 161.970 46.205 162.110 ;
        RECT 39.000 161.910 39.320 161.970 ;
        RECT 45.915 161.925 46.205 161.970 ;
        RECT 47.370 162.110 47.510 162.650 ;
        RECT 64.300 162.590 64.620 162.850 ;
        RECT 69.360 162.790 69.680 162.850 ;
        RECT 72.595 162.790 72.885 162.835 ;
        RECT 69.360 162.650 72.885 162.790 ;
        RECT 69.360 162.590 69.680 162.650 ;
        RECT 72.595 162.605 72.885 162.650 ;
        RECT 79.495 162.790 79.785 162.835 ;
        RECT 84.540 162.790 84.860 162.850 ;
        RECT 79.495 162.650 84.860 162.790 ;
        RECT 79.495 162.605 79.785 162.650 ;
        RECT 84.540 162.590 84.860 162.650 ;
        RECT 85.920 162.790 86.240 162.850 ;
        RECT 86.855 162.790 87.145 162.835 ;
        RECT 98.800 162.790 99.120 162.850 ;
        RECT 85.920 162.650 87.145 162.790 ;
        RECT 85.920 162.590 86.240 162.650 ;
        RECT 86.855 162.605 87.145 162.650 ;
        RECT 90.610 162.650 99.120 162.790 ;
        RECT 56.495 162.450 56.785 162.495 ;
        RECT 61.540 162.450 61.860 162.510 ;
        RECT 56.495 162.310 61.860 162.450 ;
        RECT 56.495 162.265 56.785 162.310 ;
        RECT 61.540 162.250 61.860 162.310 ;
        RECT 70.280 162.450 70.600 162.510 ;
        RECT 74.420 162.450 74.740 162.510 ;
        RECT 70.280 162.310 74.740 162.450 ;
        RECT 70.280 162.250 70.600 162.310 ;
        RECT 67.980 162.110 68.300 162.170 ;
        RECT 70.740 162.110 71.060 162.170 ;
        RECT 47.370 161.970 68.300 162.110 ;
        RECT 29.800 161.570 30.120 161.830 ;
        RECT 30.260 161.570 30.580 161.830 ;
        RECT 41.360 161.770 41.650 161.815 ;
        RECT 39.115 161.630 41.650 161.770 ;
        RECT 28.420 161.430 28.740 161.490 ;
        RECT 30.350 161.430 30.490 161.570 ;
        RECT 39.115 161.475 39.330 161.630 ;
        RECT 41.360 161.585 41.650 161.630 ;
        RECT 45.440 161.570 45.760 161.830 ;
        RECT 47.370 161.815 47.510 161.970 ;
        RECT 47.295 161.585 47.585 161.815 ;
        RECT 47.755 161.585 48.045 161.815 ;
        RECT 28.420 161.290 30.490 161.430 ;
        RECT 37.180 161.430 37.470 161.475 ;
        RECT 39.040 161.430 39.330 161.475 ;
        RECT 37.180 161.290 39.330 161.430 ;
        RECT 28.420 161.230 28.740 161.290 ;
        RECT 37.180 161.245 37.470 161.290 ;
        RECT 39.040 161.245 39.330 161.290 ;
        RECT 39.960 161.430 40.250 161.475 ;
        RECT 42.220 161.430 42.540 161.490 ;
        RECT 43.220 161.430 43.510 161.475 ;
        RECT 39.960 161.290 43.510 161.430 ;
        RECT 45.530 161.430 45.670 161.570 ;
        RECT 47.830 161.430 47.970 161.585 ;
        RECT 48.200 161.570 48.520 161.830 ;
        RECT 49.135 161.770 49.425 161.815 ;
        RECT 49.580 161.770 49.900 161.830 ;
        RECT 51.510 161.815 51.650 161.970 ;
        RECT 67.980 161.910 68.300 161.970 ;
        RECT 70.600 161.910 71.060 162.110 ;
        RECT 71.660 162.110 71.980 162.170 ;
        RECT 73.590 162.155 73.730 162.310 ;
        RECT 74.420 162.250 74.740 162.310 ;
        RECT 71.660 161.970 72.810 162.110 ;
        RECT 71.660 161.910 71.980 161.970 ;
        RECT 49.135 161.630 49.900 161.770 ;
        RECT 49.135 161.585 49.425 161.630 ;
        RECT 49.580 161.570 49.900 161.630 ;
        RECT 51.435 161.585 51.725 161.815 ;
        RECT 51.895 161.585 52.185 161.815 ;
        RECT 51.970 161.430 52.110 161.585 ;
        RECT 52.340 161.570 52.660 161.830 ;
        RECT 52.800 161.770 53.120 161.830 ;
        RECT 53.275 161.770 53.565 161.815 ;
        RECT 52.800 161.630 53.565 161.770 ;
        RECT 52.800 161.570 53.120 161.630 ;
        RECT 53.275 161.585 53.565 161.630 ;
        RECT 53.720 161.770 54.040 161.830 ;
        RECT 56.035 161.770 56.325 161.815 ;
        RECT 53.720 161.630 56.325 161.770 ;
        RECT 53.720 161.570 54.040 161.630 ;
        RECT 56.035 161.585 56.325 161.630 ;
        RECT 56.110 161.430 56.250 161.585 ;
        RECT 58.780 161.570 59.100 161.830 ;
        RECT 59.240 161.570 59.560 161.830 ;
        RECT 59.700 161.570 60.020 161.830 ;
        RECT 60.635 161.770 60.925 161.815 ;
        RECT 61.080 161.770 61.400 161.830 ;
        RECT 67.060 161.770 67.380 161.830 ;
        RECT 70.600 161.770 70.740 161.910 ;
        RECT 60.635 161.630 67.380 161.770 ;
        RECT 60.635 161.585 60.925 161.630 ;
        RECT 61.080 161.570 61.400 161.630 ;
        RECT 67.060 161.570 67.380 161.630 ;
        RECT 67.610 161.630 70.740 161.770 ;
        RECT 67.610 161.430 67.750 161.630 ;
        RECT 72.120 161.570 72.440 161.830 ;
        RECT 72.670 161.770 72.810 161.970 ;
        RECT 73.515 161.925 73.805 162.155 ;
        RECT 73.975 162.110 74.265 162.155 ;
        RECT 75.340 162.110 75.660 162.170 ;
        RECT 73.975 161.970 75.660 162.110 ;
        RECT 73.975 161.925 74.265 161.970 ;
        RECT 75.340 161.910 75.660 161.970 ;
        RECT 75.800 162.110 76.120 162.170 ;
        RECT 79.940 162.110 80.260 162.170 ;
        RECT 83.160 162.110 83.480 162.170 ;
        RECT 75.800 161.970 76.950 162.110 ;
        RECT 75.800 161.910 76.120 161.970 ;
        RECT 76.810 161.815 76.950 161.970 ;
        RECT 77.270 161.970 80.260 162.110 ;
        RECT 77.270 161.815 77.410 161.970 ;
        RECT 79.940 161.910 80.260 161.970 ;
        RECT 80.950 161.970 83.480 162.110 ;
        RECT 76.275 161.770 76.565 161.815 ;
        RECT 72.670 161.630 76.565 161.770 ;
        RECT 76.275 161.585 76.565 161.630 ;
        RECT 76.735 161.585 77.025 161.815 ;
        RECT 77.195 161.585 77.485 161.815 ;
        RECT 78.115 161.585 78.405 161.815 ;
        RECT 79.035 161.770 79.325 161.815 ;
        RECT 80.950 161.770 81.090 161.970 ;
        RECT 83.160 161.910 83.480 161.970 ;
        RECT 84.080 161.910 84.400 162.170 ;
        RECT 90.610 162.155 90.750 162.650 ;
        RECT 98.800 162.590 99.120 162.650 ;
        RECT 99.720 162.790 100.040 162.850 ;
        RECT 101.115 162.790 101.405 162.835 ;
        RECT 99.720 162.650 101.405 162.790 ;
        RECT 99.720 162.590 100.040 162.650 ;
        RECT 101.115 162.605 101.405 162.650 ;
        RECT 105.700 162.790 106.020 162.850 ;
        RECT 109.840 162.790 110.160 162.850 ;
        RECT 105.700 162.650 110.160 162.790 ;
        RECT 105.700 162.590 106.020 162.650 ;
        RECT 109.840 162.590 110.160 162.650 ;
        RECT 90.535 161.925 90.825 162.155 ;
        RECT 93.280 161.910 93.600 162.170 ;
        RECT 100.180 162.110 100.500 162.170 ;
        RECT 95.670 161.970 100.500 162.110 ;
        RECT 79.035 161.630 81.090 161.770 ;
        RECT 81.335 161.770 81.625 161.815 ;
        RECT 81.795 161.770 82.085 161.815 ;
        RECT 84.540 161.770 84.860 161.830 ;
        RECT 81.335 161.630 84.860 161.770 ;
        RECT 79.035 161.585 79.325 161.630 ;
        RECT 81.335 161.585 81.625 161.630 ;
        RECT 81.795 161.585 82.085 161.630 ;
        RECT 67.980 161.430 68.300 161.490 ;
        RECT 45.530 161.290 55.330 161.430 ;
        RECT 56.110 161.290 68.300 161.430 ;
        RECT 39.960 161.245 40.250 161.290 ;
        RECT 42.220 161.230 42.540 161.290 ;
        RECT 43.220 161.245 43.510 161.290 ;
        RECT 31.180 160.890 31.500 161.150 ;
        RECT 33.495 161.090 33.785 161.135 ;
        RECT 44.060 161.090 44.380 161.150 ;
        RECT 45.225 161.090 45.515 161.135 ;
        RECT 33.495 160.950 45.515 161.090 ;
        RECT 33.495 160.905 33.785 160.950 ;
        RECT 44.060 160.890 44.380 160.950 ;
        RECT 45.225 160.905 45.515 160.950 ;
        RECT 49.580 161.090 49.900 161.150 ;
        RECT 50.055 161.090 50.345 161.135 ;
        RECT 49.580 160.950 50.345 161.090 ;
        RECT 49.580 160.890 49.900 160.950 ;
        RECT 50.055 160.905 50.345 160.950 ;
        RECT 54.195 161.090 54.485 161.135 ;
        RECT 54.640 161.090 54.960 161.150 ;
        RECT 54.195 160.950 54.960 161.090 ;
        RECT 55.190 161.090 55.330 161.290 ;
        RECT 67.980 161.230 68.300 161.290 ;
        RECT 70.740 161.230 71.060 161.490 ;
        RECT 75.340 161.430 75.660 161.490 ;
        RECT 78.190 161.430 78.330 161.585 ;
        RECT 84.540 161.570 84.860 161.630 ;
        RECT 85.460 161.770 85.780 161.830 ;
        RECT 87.775 161.770 88.065 161.815 ;
        RECT 85.460 161.630 88.065 161.770 ;
        RECT 85.460 161.570 85.780 161.630 ;
        RECT 87.775 161.585 88.065 161.630 ;
        RECT 95.120 161.570 95.440 161.830 ;
        RECT 95.670 161.815 95.810 161.970 ;
        RECT 95.595 161.585 95.885 161.815 ;
        RECT 96.040 161.570 96.360 161.830 ;
        RECT 96.975 161.770 97.265 161.815 ;
        RECT 97.895 161.770 98.185 161.815 ;
        RECT 96.975 161.630 98.185 161.770 ;
        RECT 96.975 161.585 97.265 161.630 ;
        RECT 97.895 161.585 98.185 161.630 ;
        RECT 75.340 161.290 78.330 161.430 ;
        RECT 78.560 161.430 78.880 161.490 ;
        RECT 85.015 161.430 85.305 161.475 ;
        RECT 78.560 161.290 85.305 161.430 ;
        RECT 75.340 161.230 75.660 161.290 ;
        RECT 78.560 161.230 78.880 161.290 ;
        RECT 85.015 161.245 85.305 161.290 ;
        RECT 96.500 161.430 96.820 161.490 ;
        RECT 97.970 161.430 98.110 161.585 ;
        RECT 98.800 161.570 99.120 161.830 ;
        RECT 99.350 161.815 99.490 161.970 ;
        RECT 100.180 161.910 100.500 161.970 ;
        RECT 102.020 162.110 102.340 162.170 ;
        RECT 106.175 162.110 106.465 162.155 ;
        RECT 102.020 161.970 106.465 162.110 ;
        RECT 102.020 161.910 102.340 161.970 ;
        RECT 106.175 161.925 106.465 161.970 ;
        RECT 99.275 161.585 99.565 161.815 ;
        RECT 99.735 161.585 100.025 161.815 ;
        RECT 104.780 161.770 105.100 161.830 ;
        RECT 107.095 161.770 107.385 161.815 ;
        RECT 104.780 161.630 107.385 161.770 ;
        RECT 96.500 161.290 98.110 161.430 ;
        RECT 96.500 161.230 96.820 161.290 ;
        RECT 56.940 161.090 57.260 161.150 ;
        RECT 55.190 160.950 57.260 161.090 ;
        RECT 54.195 160.905 54.485 160.950 ;
        RECT 54.640 160.890 54.960 160.950 ;
        RECT 56.940 160.890 57.260 160.950 ;
        RECT 57.400 160.890 57.720 161.150 ;
        RECT 72.120 161.090 72.440 161.150 ;
        RECT 73.975 161.090 74.265 161.135 ;
        RECT 72.120 160.950 74.265 161.090 ;
        RECT 72.120 160.890 72.440 160.950 ;
        RECT 73.975 160.905 74.265 160.950 ;
        RECT 74.880 160.890 75.200 161.150 ;
        RECT 80.860 160.890 81.180 161.150 ;
        RECT 82.240 160.890 82.560 161.150 ;
        RECT 83.620 161.090 83.940 161.150 ;
        RECT 84.555 161.090 84.845 161.135 ;
        RECT 83.620 160.950 84.845 161.090 ;
        RECT 83.620 160.890 83.940 160.950 ;
        RECT 84.555 160.905 84.845 160.950 ;
        RECT 88.235 161.090 88.525 161.135 ;
        RECT 91.440 161.090 91.760 161.150 ;
        RECT 88.235 160.950 91.760 161.090 ;
        RECT 88.235 160.905 88.525 160.950 ;
        RECT 91.440 160.890 91.760 160.950 ;
        RECT 91.900 161.090 92.220 161.150 ;
        RECT 93.755 161.090 94.045 161.135 ;
        RECT 91.900 160.950 94.045 161.090 ;
        RECT 91.900 160.890 92.220 160.950 ;
        RECT 93.755 160.905 94.045 160.950 ;
        RECT 97.880 161.090 98.200 161.150 ;
        RECT 99.810 161.090 99.950 161.585 ;
        RECT 104.780 161.570 105.100 161.630 ;
        RECT 107.095 161.585 107.385 161.630 ;
        RECT 109.840 161.570 110.160 161.830 ;
        RECT 102.480 161.430 102.800 161.490 ;
        RECT 102.955 161.430 103.245 161.475 ;
        RECT 107.555 161.430 107.845 161.475 ;
        RECT 102.480 161.290 107.845 161.430 ;
        RECT 102.480 161.230 102.800 161.290 ;
        RECT 102.955 161.245 103.245 161.290 ;
        RECT 107.555 161.245 107.845 161.290 ;
        RECT 97.880 160.950 99.950 161.090 ;
        RECT 97.880 160.890 98.200 160.950 ;
        RECT 103.400 160.890 103.720 161.150 ;
        RECT 105.255 161.090 105.545 161.135 ;
        RECT 107.080 161.090 107.400 161.150 ;
        RECT 105.255 160.950 107.400 161.090 ;
        RECT 105.255 160.905 105.545 160.950 ;
        RECT 107.080 160.890 107.400 160.950 ;
        RECT 109.380 160.890 109.700 161.150 ;
        RECT 110.760 160.890 111.080 161.150 ;
        RECT 26.970 160.270 113.450 160.750 ;
        RECT 39.000 160.070 39.320 160.130 ;
        RECT 45.900 160.070 46.220 160.130 ;
        RECT 48.200 160.070 48.520 160.130 ;
        RECT 29.430 159.930 39.320 160.070 ;
        RECT 29.430 159.435 29.570 159.930 ;
        RECT 39.000 159.870 39.320 159.930 ;
        RECT 39.780 159.930 43.370 160.070 ;
        RECT 33.480 159.530 33.800 159.790 ;
        RECT 37.635 159.730 37.925 159.775 ;
        RECT 39.780 159.730 39.920 159.930 ;
        RECT 42.220 159.730 42.540 159.790 ;
        RECT 34.950 159.590 37.925 159.730 ;
        RECT 29.355 159.205 29.645 159.435 ;
        RECT 30.735 159.390 31.025 159.435 ;
        RECT 29.890 159.250 31.025 159.390 ;
        RECT 29.890 158.710 30.030 159.250 ;
        RECT 30.735 159.205 31.025 159.250 ;
        RECT 32.115 159.390 32.405 159.435 ;
        RECT 34.950 159.390 35.090 159.590 ;
        RECT 37.635 159.545 37.925 159.590 ;
        RECT 39.550 159.590 39.920 159.730 ;
        RECT 40.930 159.590 42.540 159.730 ;
        RECT 32.115 159.250 35.090 159.390 ;
        RECT 37.175 159.390 37.465 159.435 ;
        RECT 38.540 159.390 38.860 159.450 ;
        RECT 37.175 159.250 38.860 159.390 ;
        RECT 32.115 159.205 32.405 159.250 ;
        RECT 37.175 159.205 37.465 159.250 ;
        RECT 38.540 159.190 38.860 159.250 ;
        RECT 39.000 159.190 39.320 159.450 ;
        RECT 39.550 159.435 39.690 159.590 ;
        RECT 39.475 159.205 39.765 159.435 ;
        RECT 39.920 159.190 40.240 159.450 ;
        RECT 40.930 159.435 41.070 159.590 ;
        RECT 42.220 159.530 42.540 159.590 ;
        RECT 43.230 159.730 43.370 159.930 ;
        RECT 45.900 159.930 48.520 160.070 ;
        RECT 45.900 159.870 46.220 159.930 ;
        RECT 48.200 159.870 48.520 159.930 ;
        RECT 59.700 160.070 60.020 160.130 ;
        RECT 60.175 160.070 60.465 160.115 ;
        RECT 59.700 159.930 60.465 160.070 ;
        RECT 59.700 159.870 60.020 159.930 ;
        RECT 60.175 159.885 60.465 159.930 ;
        RECT 64.760 159.870 65.080 160.130 ;
        RECT 77.195 160.070 77.485 160.115 ;
        RECT 88.220 160.070 88.540 160.130 ;
        RECT 77.195 159.930 88.540 160.070 ;
        RECT 77.195 159.885 77.485 159.930 ;
        RECT 88.220 159.870 88.540 159.930 ;
        RECT 106.635 160.070 106.925 160.115 ;
        RECT 109.840 160.070 110.160 160.130 ;
        RECT 106.635 159.930 110.160 160.070 ;
        RECT 106.635 159.885 106.925 159.930 ;
        RECT 109.840 159.870 110.160 159.930 ;
        RECT 45.440 159.730 45.760 159.790 ;
        RECT 50.060 159.730 50.350 159.775 ;
        RECT 51.920 159.730 52.210 159.775 ;
        RECT 43.230 159.590 45.760 159.730 ;
        RECT 40.855 159.205 41.145 159.435 ;
        RECT 41.760 159.390 42.080 159.450 ;
        RECT 43.230 159.435 43.370 159.590 ;
        RECT 45.440 159.530 45.760 159.590 ;
        RECT 47.370 159.590 49.810 159.730 ;
        RECT 42.695 159.390 42.985 159.435 ;
        RECT 41.760 159.250 42.985 159.390 ;
        RECT 41.760 159.190 42.080 159.250 ;
        RECT 42.695 159.205 42.985 159.250 ;
        RECT 43.155 159.205 43.445 159.435 ;
        RECT 43.615 159.390 43.905 159.435 ;
        RECT 44.060 159.390 44.380 159.450 ;
        RECT 43.615 159.250 44.380 159.390 ;
        RECT 43.615 159.205 43.905 159.250 ;
        RECT 44.060 159.190 44.380 159.250 ;
        RECT 44.520 159.190 44.840 159.450 ;
        RECT 45.900 159.390 46.220 159.450 ;
        RECT 46.375 159.390 46.665 159.435 ;
        RECT 45.900 159.250 46.665 159.390 ;
        RECT 45.900 159.190 46.220 159.250 ;
        RECT 46.375 159.205 46.665 159.250 ;
        RECT 46.820 159.190 47.140 159.450 ;
        RECT 47.370 159.435 47.510 159.590 ;
        RECT 47.295 159.205 47.585 159.435 ;
        RECT 48.200 159.190 48.520 159.450 ;
        RECT 49.670 159.390 49.810 159.590 ;
        RECT 50.060 159.590 52.210 159.730 ;
        RECT 50.060 159.545 50.350 159.590 ;
        RECT 51.920 159.545 52.210 159.590 ;
        RECT 52.840 159.730 53.130 159.775 ;
        RECT 54.640 159.730 54.960 159.790 ;
        RECT 56.100 159.730 56.390 159.775 ;
        RECT 52.840 159.590 56.390 159.730 ;
        RECT 52.840 159.545 53.130 159.590 ;
        RECT 51.995 159.390 52.210 159.545 ;
        RECT 54.640 159.530 54.960 159.590 ;
        RECT 56.100 159.545 56.390 159.590 ;
        RECT 59.240 159.730 59.560 159.790 ;
        RECT 68.915 159.730 69.205 159.775 ;
        RECT 72.120 159.730 72.440 159.790 ;
        RECT 59.240 159.590 65.910 159.730 ;
        RECT 59.240 159.530 59.560 159.590 ;
        RECT 54.240 159.390 54.530 159.435 ;
        RECT 60.635 159.390 60.925 159.435 ;
        RECT 63.855 159.390 64.145 159.435 ;
        RECT 49.670 159.250 51.650 159.390 ;
        RECT 51.995 159.250 54.530 159.390 ;
        RECT 30.275 159.050 30.565 159.095 ;
        RECT 32.560 159.050 32.880 159.110 ;
        RECT 30.275 158.910 32.880 159.050 ;
        RECT 30.275 158.865 30.565 158.910 ;
        RECT 32.560 158.850 32.880 158.910 ;
        RECT 33.035 159.050 33.325 159.095 ;
        RECT 33.480 159.050 33.800 159.110 ;
        RECT 33.035 158.910 33.800 159.050 ;
        RECT 33.035 158.865 33.325 158.910 ;
        RECT 33.480 158.850 33.800 158.910 ;
        RECT 33.955 159.050 34.245 159.095 ;
        RECT 36.240 159.050 36.560 159.110 ;
        RECT 33.955 158.910 36.560 159.050 ;
        RECT 33.955 158.865 34.245 158.910 ;
        RECT 36.240 158.850 36.560 158.910 ;
        RECT 37.620 159.050 37.940 159.110 ;
        RECT 49.135 159.050 49.425 159.095 ;
        RECT 37.620 158.910 49.425 159.050 ;
        RECT 37.620 158.850 37.940 158.910 ;
        RECT 49.135 158.865 49.425 158.910 ;
        RECT 50.960 158.850 51.280 159.110 ;
        RECT 51.510 159.050 51.650 159.250 ;
        RECT 54.240 159.205 54.530 159.250 ;
        RECT 58.180 159.250 60.925 159.390 ;
        RECT 55.560 159.050 55.880 159.110 ;
        RECT 58.180 159.095 58.320 159.250 ;
        RECT 60.635 159.205 60.925 159.250 ;
        RECT 62.550 159.250 64.145 159.390 ;
        RECT 58.105 159.050 58.395 159.095 ;
        RECT 51.510 158.910 58.395 159.050 ;
        RECT 55.560 158.850 55.880 158.910 ;
        RECT 58.105 158.865 58.395 158.910 ;
        RECT 59.715 159.050 60.005 159.095 ;
        RECT 59.715 158.910 62.230 159.050 ;
        RECT 59.715 158.865 60.005 158.910 ;
        RECT 44.995 158.710 45.285 158.755 ;
        RECT 29.890 158.570 45.285 158.710 ;
        RECT 44.995 158.525 45.285 158.570 ;
        RECT 49.600 158.710 49.890 158.755 ;
        RECT 51.460 158.710 51.750 158.755 ;
        RECT 54.240 158.710 54.530 158.755 ;
        RECT 49.600 158.570 54.530 158.710 ;
        RECT 49.600 158.525 49.890 158.570 ;
        RECT 51.460 158.525 51.750 158.570 ;
        RECT 54.240 158.525 54.530 158.570 ;
        RECT 27.960 158.370 28.280 158.430 ;
        RECT 28.435 158.370 28.725 158.415 ;
        RECT 27.960 158.230 28.725 158.370 ;
        RECT 27.960 158.170 28.280 158.230 ;
        RECT 28.435 158.185 28.725 158.230 ;
        RECT 30.260 158.170 30.580 158.430 ;
        RECT 30.720 158.370 31.040 158.430 ;
        RECT 31.195 158.370 31.485 158.415 ;
        RECT 30.720 158.230 31.485 158.370 ;
        RECT 30.720 158.170 31.040 158.230 ;
        RECT 31.195 158.185 31.485 158.230 ;
        RECT 32.100 158.170 32.420 158.430 ;
        RECT 37.160 158.370 37.480 158.430 ;
        RECT 41.315 158.370 41.605 158.415 ;
        RECT 37.160 158.230 41.605 158.370 ;
        RECT 37.160 158.170 37.480 158.230 ;
        RECT 41.315 158.185 41.605 158.230 ;
        RECT 43.600 158.370 43.920 158.430 ;
        RECT 52.800 158.370 53.120 158.430 ;
        RECT 43.600 158.230 53.120 158.370 ;
        RECT 62.090 158.370 62.230 158.910 ;
        RECT 62.550 158.755 62.690 159.250 ;
        RECT 63.855 159.205 64.145 159.250 ;
        RECT 65.770 158.755 65.910 159.590 ;
        RECT 68.915 159.590 72.440 159.730 ;
        RECT 68.915 159.545 69.205 159.590 ;
        RECT 72.120 159.530 72.440 159.590 ;
        RECT 73.975 159.730 74.265 159.775 ;
        RECT 77.885 159.730 78.175 159.775 ;
        RECT 78.560 159.730 78.880 159.790 ;
        RECT 73.975 159.590 77.410 159.730 ;
        RECT 73.975 159.545 74.265 159.590 ;
        RECT 66.615 159.390 66.905 159.435 ;
        RECT 69.360 159.390 69.680 159.450 ;
        RECT 66.615 159.250 69.680 159.390 ;
        RECT 66.615 159.205 66.905 159.250 ;
        RECT 69.360 159.190 69.680 159.250 ;
        RECT 69.835 159.390 70.125 159.435 ;
        RECT 71.660 159.390 71.980 159.450 ;
        RECT 69.835 159.250 71.980 159.390 ;
        RECT 69.835 159.205 70.125 159.250 ;
        RECT 71.660 159.190 71.980 159.250 ;
        RECT 75.815 159.205 76.105 159.435 ;
        RECT 76.275 159.205 76.565 159.435 ;
        RECT 77.270 159.390 77.410 159.590 ;
        RECT 77.885 159.590 78.880 159.730 ;
        RECT 77.885 159.545 78.175 159.590 ;
        RECT 78.560 159.530 78.880 159.590 ;
        RECT 79.890 159.730 80.180 159.775 ;
        RECT 80.860 159.730 81.180 159.790 ;
        RECT 83.150 159.730 83.440 159.775 ;
        RECT 79.890 159.590 83.440 159.730 ;
        RECT 79.890 159.545 80.180 159.590 ;
        RECT 80.860 159.530 81.180 159.590 ;
        RECT 83.150 159.545 83.440 159.590 ;
        RECT 84.070 159.730 84.360 159.775 ;
        RECT 85.930 159.730 86.220 159.775 ;
        RECT 84.070 159.590 86.220 159.730 ;
        RECT 84.070 159.545 84.360 159.590 ;
        RECT 85.930 159.545 86.220 159.590 ;
        RECT 81.750 159.390 82.040 159.435 ;
        RECT 84.070 159.390 84.285 159.545 ;
        RECT 88.680 159.530 89.000 159.790 ;
        RECT 91.440 159.775 91.760 159.790 ;
        RECT 90.975 159.730 91.760 159.775 ;
        RECT 94.575 159.730 94.865 159.775 ;
        RECT 90.975 159.590 94.865 159.730 ;
        RECT 90.975 159.545 91.760 159.590 ;
        RECT 91.440 159.530 91.760 159.545 ;
        RECT 94.275 159.545 94.865 159.590 ;
        RECT 96.500 159.730 96.820 159.790 ;
        RECT 102.480 159.730 102.800 159.790 ;
        RECT 111.220 159.730 111.540 159.790 ;
        RECT 96.500 159.590 99.950 159.730 ;
        RECT 77.270 159.250 80.630 159.390 ;
        RECT 66.140 159.050 66.460 159.110 ;
        RECT 75.890 159.050 76.030 159.205 ;
        RECT 66.140 158.910 76.030 159.050 ;
        RECT 76.350 159.050 76.490 159.205 ;
        RECT 80.490 159.050 80.630 159.250 ;
        RECT 81.750 159.250 84.285 159.390 ;
        RECT 87.780 159.390 88.070 159.435 ;
        RECT 89.615 159.390 89.905 159.435 ;
        RECT 93.195 159.390 93.485 159.435 ;
        RECT 87.780 159.250 93.485 159.390 ;
        RECT 81.750 159.205 82.040 159.250 ;
        RECT 87.780 159.205 88.070 159.250 ;
        RECT 89.615 159.205 89.905 159.250 ;
        RECT 93.195 159.205 93.485 159.250 ;
        RECT 94.275 159.230 94.565 159.545 ;
        RECT 96.500 159.530 96.820 159.590 ;
        RECT 97.880 159.190 98.200 159.450 ;
        RECT 99.810 159.435 99.950 159.590 ;
        RECT 101.190 159.590 111.910 159.730 ;
        RECT 98.355 159.205 98.645 159.435 ;
        RECT 98.815 159.205 99.105 159.435 ;
        RECT 99.735 159.390 100.025 159.435 ;
        RECT 100.180 159.390 100.500 159.450 ;
        RECT 101.190 159.435 101.330 159.590 ;
        RECT 102.480 159.530 102.800 159.590 ;
        RECT 111.220 159.530 111.540 159.590 ;
        RECT 99.735 159.250 100.500 159.390 ;
        RECT 99.735 159.205 100.025 159.250 ;
        RECT 84.080 159.050 84.400 159.110 ;
        RECT 76.350 158.910 80.170 159.050 ;
        RECT 80.490 158.910 84.400 159.050 ;
        RECT 66.140 158.850 66.460 158.910 ;
        RECT 62.475 158.525 62.765 158.755 ;
        RECT 65.695 158.710 65.985 158.755 ;
        RECT 67.060 158.710 67.380 158.770 ;
        RECT 65.695 158.570 67.380 158.710 ;
        RECT 65.695 158.525 65.985 158.570 ;
        RECT 67.060 158.510 67.380 158.570 ;
        RECT 70.755 158.710 71.045 158.755 ;
        RECT 76.260 158.710 76.580 158.770 ;
        RECT 70.755 158.570 76.580 158.710 ;
        RECT 70.755 158.525 71.045 158.570 ;
        RECT 76.260 158.510 76.580 158.570 ;
        RECT 63.840 158.370 64.160 158.430 ;
        RECT 67.535 158.370 67.825 158.415 ;
        RECT 62.090 158.230 67.825 158.370 ;
        RECT 43.600 158.170 43.920 158.230 ;
        RECT 52.800 158.170 53.120 158.230 ;
        RECT 63.840 158.170 64.160 158.230 ;
        RECT 67.535 158.185 67.825 158.230 ;
        RECT 69.360 158.370 69.680 158.430 ;
        RECT 74.895 158.370 75.185 158.415 ;
        RECT 69.360 158.230 75.185 158.370 ;
        RECT 80.030 158.370 80.170 158.910 ;
        RECT 84.080 158.850 84.400 158.910 ;
        RECT 85.015 159.050 85.305 159.095 ;
        RECT 85.460 159.050 85.780 159.110 ;
        RECT 85.015 158.910 85.780 159.050 ;
        RECT 85.015 158.865 85.305 158.910 ;
        RECT 85.460 158.850 85.780 158.910 ;
        RECT 86.855 159.050 87.145 159.095 ;
        RECT 87.300 159.050 87.620 159.110 ;
        RECT 86.855 158.910 87.620 159.050 ;
        RECT 86.855 158.865 87.145 158.910 ;
        RECT 87.300 158.850 87.620 158.910 ;
        RECT 92.360 159.050 92.680 159.110 ;
        RECT 96.040 159.050 96.360 159.110 ;
        RECT 92.360 158.910 96.360 159.050 ;
        RECT 92.360 158.850 92.680 158.910 ;
        RECT 96.040 158.850 96.360 158.910 ;
        RECT 96.500 159.050 96.820 159.110 ;
        RECT 98.430 159.050 98.570 159.205 ;
        RECT 96.500 158.910 98.570 159.050 ;
        RECT 96.500 158.850 96.820 158.910 ;
        RECT 81.750 158.710 82.040 158.755 ;
        RECT 84.530 158.710 84.820 158.755 ;
        RECT 86.390 158.710 86.680 158.755 ;
        RECT 81.750 158.570 86.680 158.710 ;
        RECT 81.750 158.525 82.040 158.570 ;
        RECT 84.530 158.525 84.820 158.570 ;
        RECT 86.390 158.525 86.680 158.570 ;
        RECT 88.185 158.710 88.475 158.755 ;
        RECT 90.075 158.710 90.365 158.755 ;
        RECT 93.195 158.710 93.485 158.755 ;
        RECT 88.185 158.570 93.485 158.710 ;
        RECT 98.890 158.710 99.030 159.205 ;
        RECT 100.180 159.190 100.500 159.250 ;
        RECT 101.115 159.205 101.405 159.435 ;
        RECT 101.560 159.190 101.880 159.450 ;
        RECT 104.780 159.190 105.100 159.450 ;
        RECT 107.080 159.190 107.400 159.450 ;
        RECT 111.770 159.435 111.910 159.590 ;
        RECT 111.695 159.205 111.985 159.435 ;
        RECT 102.020 159.050 102.340 159.110 ;
        RECT 103.415 159.050 103.705 159.095 ;
        RECT 102.020 158.910 103.705 159.050 ;
        RECT 102.020 158.850 102.340 158.910 ;
        RECT 103.415 158.865 103.705 158.910 ;
        RECT 104.320 158.850 104.640 159.110 ;
        RECT 104.870 158.710 105.010 159.190 ;
        RECT 110.315 159.050 110.605 159.095 ;
        RECT 111.220 159.050 111.540 159.110 ;
        RECT 110.315 158.910 111.540 159.050 ;
        RECT 110.315 158.865 110.605 158.910 ;
        RECT 111.220 158.850 111.540 158.910 ;
        RECT 98.890 158.570 105.010 158.710 ;
        RECT 88.185 158.525 88.475 158.570 ;
        RECT 90.075 158.525 90.365 158.570 ;
        RECT 93.195 158.525 93.485 158.570 ;
        RECT 87.760 158.370 88.080 158.430 ;
        RECT 80.030 158.230 88.080 158.370 ;
        RECT 69.360 158.170 69.680 158.230 ;
        RECT 74.895 158.185 75.185 158.230 ;
        RECT 87.760 158.170 88.080 158.230 ;
        RECT 89.600 158.370 89.920 158.430 ;
        RECT 96.515 158.370 96.805 158.415 ;
        RECT 89.600 158.230 96.805 158.370 ;
        RECT 89.600 158.170 89.920 158.230 ;
        RECT 96.515 158.185 96.805 158.230 ;
        RECT 97.420 158.370 97.740 158.430 ;
        RECT 101.100 158.370 101.420 158.430 ;
        RECT 97.420 158.230 101.420 158.370 ;
        RECT 97.420 158.170 97.740 158.230 ;
        RECT 101.100 158.170 101.420 158.230 ;
        RECT 107.080 158.370 107.400 158.430 ;
        RECT 111.235 158.370 111.525 158.415 ;
        RECT 107.080 158.230 111.525 158.370 ;
        RECT 107.080 158.170 107.400 158.230 ;
        RECT 111.235 158.185 111.525 158.230 ;
        RECT 26.970 157.550 113.450 158.030 ;
        RECT 30.260 157.150 30.580 157.410 ;
        RECT 33.480 157.350 33.800 157.410 ;
        RECT 30.810 157.210 33.800 157.350 ;
        RECT 26.580 157.010 26.900 157.070 ;
        RECT 30.810 157.010 30.950 157.210 ;
        RECT 33.480 157.150 33.800 157.210 ;
        RECT 36.700 157.350 37.020 157.410 ;
        RECT 37.175 157.350 37.465 157.395 ;
        RECT 39.935 157.350 40.225 157.395 ;
        RECT 36.700 157.210 37.465 157.350 ;
        RECT 36.700 157.150 37.020 157.210 ;
        RECT 37.175 157.165 37.465 157.210 ;
        RECT 38.630 157.210 40.225 157.350 ;
        RECT 26.580 156.870 30.950 157.010 ;
        RECT 31.180 157.010 31.500 157.070 ;
        RECT 38.630 157.010 38.770 157.210 ;
        RECT 39.935 157.165 40.225 157.210 ;
        RECT 41.760 157.150 42.080 157.410 ;
        RECT 44.060 157.150 44.380 157.410 ;
        RECT 44.520 157.350 44.840 157.410 ;
        RECT 48.215 157.350 48.505 157.395 ;
        RECT 44.520 157.210 48.505 157.350 ;
        RECT 44.520 157.150 44.840 157.210 ;
        RECT 48.215 157.165 48.505 157.210 ;
        RECT 50.960 157.350 51.280 157.410 ;
        RECT 51.895 157.350 52.185 157.395 ;
        RECT 50.960 157.210 52.185 157.350 ;
        RECT 50.960 157.150 51.280 157.210 ;
        RECT 51.895 157.165 52.185 157.210 ;
        RECT 52.430 157.210 55.330 157.350 ;
        RECT 52.430 157.010 52.570 157.210 ;
        RECT 31.180 156.870 38.770 157.010 ;
        RECT 46.910 156.870 52.570 157.010 ;
        RECT 26.580 156.810 26.900 156.870 ;
        RECT 31.180 156.810 31.500 156.870 ;
        RECT 28.420 156.670 28.740 156.730 ;
        RECT 33.955 156.670 34.245 156.715 ;
        RECT 35.780 156.670 36.100 156.730 ;
        RECT 28.420 156.530 33.250 156.670 ;
        RECT 28.420 156.470 28.740 156.530 ;
        RECT 29.430 156.375 29.570 156.530 ;
        RECT 28.895 156.145 29.185 156.375 ;
        RECT 29.355 156.145 29.645 156.375 ;
        RECT 29.800 156.330 30.120 156.390 ;
        RECT 32.575 156.330 32.865 156.375 ;
        RECT 29.800 156.190 32.865 156.330 ;
        RECT 33.110 156.330 33.250 156.530 ;
        RECT 33.955 156.530 36.100 156.670 ;
        RECT 33.955 156.485 34.245 156.530 ;
        RECT 35.780 156.470 36.100 156.530 ;
        RECT 38.080 156.470 38.400 156.730 ;
        RECT 40.840 156.470 41.160 156.730 ;
        RECT 43.600 156.470 43.920 156.730 ;
        RECT 44.520 156.670 44.840 156.730 ;
        RECT 46.910 156.670 47.050 156.870 ;
        RECT 53.275 156.825 53.565 157.055 ;
        RECT 50.960 156.670 51.280 156.730 ;
        RECT 44.520 156.530 47.050 156.670 ;
        RECT 44.520 156.470 44.840 156.530 ;
        RECT 34.860 156.330 35.180 156.390 ;
        RECT 33.110 156.190 35.180 156.330 ;
        RECT 28.970 155.990 29.110 156.145 ;
        RECT 29.800 156.130 30.120 156.190 ;
        RECT 32.575 156.145 32.865 156.190 ;
        RECT 34.860 156.130 35.180 156.190 ;
        RECT 35.320 156.330 35.640 156.390 ;
        RECT 36.240 156.330 36.560 156.390 ;
        RECT 35.320 156.190 36.560 156.330 ;
        RECT 35.320 156.130 35.640 156.190 ;
        RECT 36.240 156.130 36.560 156.190 ;
        RECT 37.160 156.130 37.480 156.390 ;
        RECT 39.920 156.130 40.240 156.390 ;
        RECT 41.300 156.130 41.620 156.390 ;
        RECT 42.680 156.130 43.000 156.390 ;
        RECT 44.075 156.330 44.365 156.375 ;
        RECT 44.075 156.190 45.670 156.330 ;
        RECT 44.075 156.145 44.365 156.190 ;
        RECT 32.100 155.990 32.420 156.050 ;
        RECT 33.035 155.990 33.325 156.035 ;
        RECT 28.970 155.850 33.325 155.990 ;
        RECT 32.100 155.790 32.420 155.850 ;
        RECT 33.035 155.805 33.325 155.850 ;
        RECT 38.555 155.990 38.845 156.035 ;
        RECT 44.535 155.990 44.825 156.035 ;
        RECT 38.555 155.850 44.825 155.990 ;
        RECT 38.555 155.805 38.845 155.850 ;
        RECT 44.535 155.805 44.825 155.850 ;
        RECT 28.420 155.650 28.740 155.710 ;
        RECT 30.735 155.650 31.025 155.695 ;
        RECT 28.420 155.510 31.025 155.650 ;
        RECT 28.420 155.450 28.740 155.510 ;
        RECT 30.735 155.465 31.025 155.510 ;
        RECT 36.255 155.650 36.545 155.695 ;
        RECT 38.080 155.650 38.400 155.710 ;
        RECT 36.255 155.510 38.400 155.650 ;
        RECT 36.255 155.465 36.545 155.510 ;
        RECT 38.080 155.450 38.400 155.510 ;
        RECT 39.015 155.650 39.305 155.695 ;
        RECT 43.600 155.650 43.920 155.710 ;
        RECT 39.015 155.510 43.920 155.650 ;
        RECT 45.530 155.650 45.670 156.190 ;
        RECT 45.900 156.130 46.220 156.390 ;
        RECT 46.360 156.130 46.680 156.390 ;
        RECT 46.910 156.375 47.050 156.530 ;
        RECT 50.590 156.530 51.280 156.670 ;
        RECT 46.835 156.145 47.125 156.375 ;
        RECT 47.740 156.130 48.060 156.390 ;
        RECT 49.495 156.330 49.785 156.375 ;
        RECT 49.210 156.190 49.785 156.330 ;
        RECT 45.990 155.990 46.130 156.130 ;
        RECT 49.210 155.990 49.350 156.190 ;
        RECT 49.495 156.145 49.785 156.190 ;
        RECT 50.040 156.130 50.360 156.390 ;
        RECT 50.590 156.375 50.730 156.530 ;
        RECT 50.960 156.470 51.280 156.530 ;
        RECT 50.515 156.145 50.805 156.375 ;
        RECT 51.435 156.330 51.725 156.375 ;
        RECT 52.340 156.330 52.660 156.390 ;
        RECT 51.435 156.190 52.660 156.330 ;
        RECT 51.435 156.145 51.725 156.190 ;
        RECT 52.340 156.130 52.660 156.190 ;
        RECT 52.815 156.330 53.105 156.375 ;
        RECT 53.350 156.330 53.490 156.825 ;
        RECT 55.190 156.375 55.330 157.210 ;
        RECT 66.140 157.150 66.460 157.410 ;
        RECT 67.060 157.350 67.380 157.410 ;
        RECT 74.420 157.350 74.740 157.410 ;
        RECT 67.060 157.210 74.740 157.350 ;
        RECT 67.060 157.150 67.380 157.210 ;
        RECT 74.420 157.150 74.740 157.210 ;
        RECT 75.355 157.350 75.645 157.395 ;
        RECT 80.860 157.350 81.180 157.410 ;
        RECT 75.355 157.210 81.180 157.350 ;
        RECT 75.355 157.165 75.645 157.210 ;
        RECT 80.860 157.150 81.180 157.210 ;
        RECT 83.620 157.150 83.940 157.410 ;
        RECT 89.600 157.150 89.920 157.410 ;
        RECT 91.900 157.150 92.220 157.410 ;
        RECT 99.720 157.350 100.040 157.410 ;
        RECT 102.725 157.350 103.015 157.395 ;
        RECT 104.320 157.350 104.640 157.410 ;
        RECT 99.720 157.210 104.640 157.350 ;
        RECT 99.720 157.150 100.040 157.210 ;
        RECT 102.725 157.165 103.015 157.210 ;
        RECT 104.320 157.150 104.640 157.210 ;
        RECT 58.780 157.010 59.100 157.070 ;
        RECT 69.835 157.010 70.125 157.055 ;
        RECT 56.110 156.870 70.125 157.010 ;
        RECT 55.560 156.470 55.880 156.730 ;
        RECT 52.815 156.190 53.490 156.330 ;
        RECT 52.815 156.145 53.105 156.190 ;
        RECT 55.115 156.145 55.405 156.375 ;
        RECT 56.110 155.990 56.250 156.870 ;
        RECT 58.780 156.810 59.100 156.870 ;
        RECT 69.835 156.825 70.125 156.870 ;
        RECT 71.675 157.010 71.965 157.055 ;
        RECT 82.700 157.010 83.020 157.070 ;
        RECT 95.120 157.010 95.440 157.070 ;
        RECT 97.880 157.010 98.200 157.070 ;
        RECT 71.675 156.870 77.870 157.010 ;
        RECT 71.675 156.825 71.965 156.870 ;
        RECT 56.495 156.670 56.785 156.715 ;
        RECT 63.395 156.670 63.685 156.715 ;
        RECT 63.840 156.670 64.160 156.730 ;
        RECT 56.495 156.530 64.160 156.670 ;
        RECT 69.910 156.670 70.050 156.825 ;
        RECT 75.800 156.670 76.120 156.730 ;
        RECT 69.910 156.530 76.120 156.670 ;
        RECT 56.495 156.485 56.785 156.530 ;
        RECT 59.330 156.375 59.470 156.530 ;
        RECT 63.395 156.485 63.685 156.530 ;
        RECT 63.840 156.470 64.160 156.530 ;
        RECT 75.800 156.470 76.120 156.530 ;
        RECT 76.260 156.670 76.580 156.730 ;
        RECT 76.260 156.530 77.410 156.670 ;
        RECT 76.260 156.470 76.580 156.530 ;
        RECT 58.335 156.330 58.625 156.375 ;
        RECT 45.990 155.850 56.250 155.990 ;
        RECT 56.800 156.190 58.625 156.330 ;
        RECT 53.260 155.650 53.580 155.710 ;
        RECT 45.530 155.510 53.580 155.650 ;
        RECT 39.015 155.465 39.305 155.510 ;
        RECT 43.600 155.450 43.920 155.510 ;
        RECT 53.260 155.450 53.580 155.510 ;
        RECT 56.020 155.650 56.340 155.710 ;
        RECT 56.800 155.650 56.940 156.190 ;
        RECT 58.335 156.145 58.625 156.190 ;
        RECT 59.255 156.145 59.545 156.375 ;
        RECT 60.160 156.130 60.480 156.390 ;
        RECT 61.630 156.190 67.290 156.330 ;
        RECT 59.715 155.990 60.005 156.035 ;
        RECT 61.630 155.990 61.770 156.190 ;
        RECT 59.715 155.850 61.770 155.990 ;
        RECT 62.000 155.990 62.320 156.050 ;
        RECT 64.315 155.990 64.605 156.035 ;
        RECT 62.000 155.850 64.605 155.990 ;
        RECT 67.150 155.990 67.290 156.190 ;
        RECT 67.520 156.130 67.840 156.390 ;
        RECT 68.915 156.145 69.205 156.375 ;
        RECT 69.820 156.330 70.140 156.390 ;
        RECT 70.755 156.330 71.045 156.375 ;
        RECT 69.820 156.190 71.045 156.330 ;
        RECT 68.990 155.990 69.130 156.145 ;
        RECT 69.820 156.130 70.140 156.190 ;
        RECT 70.755 156.145 71.045 156.190 ;
        RECT 73.040 156.330 73.360 156.390 ;
        RECT 77.270 156.375 77.410 156.530 ;
        RECT 77.730 156.390 77.870 156.870 ;
        RECT 82.700 156.870 92.130 157.010 ;
        RECT 82.700 156.810 83.020 156.870 ;
        RECT 80.415 156.670 80.705 156.715 ;
        RECT 84.080 156.670 84.400 156.730 ;
        RECT 91.990 156.715 92.130 156.870 ;
        RECT 95.120 156.870 98.200 157.010 ;
        RECT 95.120 156.810 95.440 156.870 ;
        RECT 97.880 156.810 98.200 156.870 ;
        RECT 78.190 156.530 79.710 156.670 ;
        RECT 73.975 156.330 74.265 156.375 ;
        RECT 73.040 156.190 74.265 156.330 ;
        RECT 73.040 156.130 73.360 156.190 ;
        RECT 73.975 156.145 74.265 156.190 ;
        RECT 74.435 156.330 74.725 156.375 ;
        RECT 74.435 156.190 76.950 156.330 ;
        RECT 74.435 156.145 74.725 156.190 ;
        RECT 71.660 155.990 71.980 156.050 ;
        RECT 67.150 155.850 68.670 155.990 ;
        RECT 68.990 155.850 71.980 155.990 ;
        RECT 59.715 155.805 60.005 155.850 ;
        RECT 62.000 155.790 62.320 155.850 ;
        RECT 64.315 155.805 64.605 155.850 ;
        RECT 56.020 155.510 56.940 155.650 ;
        RECT 56.020 155.450 56.340 155.510 ;
        RECT 61.080 155.450 61.400 155.710 ;
        RECT 63.855 155.650 64.145 155.695 ;
        RECT 65.680 155.650 66.000 155.710 ;
        RECT 63.855 155.510 66.000 155.650 ;
        RECT 63.855 155.465 64.145 155.510 ;
        RECT 65.680 155.450 66.000 155.510 ;
        RECT 67.060 155.450 67.380 155.710 ;
        RECT 68.530 155.650 68.670 155.850 ;
        RECT 71.660 155.790 71.980 155.850 ;
        RECT 75.355 155.990 75.645 156.035 ;
        RECT 75.815 155.990 76.105 156.035 ;
        RECT 75.355 155.850 76.105 155.990 ;
        RECT 76.810 155.990 76.950 156.190 ;
        RECT 77.195 156.145 77.485 156.375 ;
        RECT 77.640 156.130 77.960 156.390 ;
        RECT 78.190 156.375 78.330 156.530 ;
        RECT 79.570 156.390 79.710 156.530 ;
        RECT 80.415 156.530 84.400 156.670 ;
        RECT 80.415 156.485 80.705 156.530 ;
        RECT 84.080 156.470 84.400 156.530 ;
        RECT 91.915 156.485 92.205 156.715 ;
        RECT 93.740 156.670 94.060 156.730 ;
        RECT 99.810 156.670 99.950 157.150 ;
        RECT 106.590 157.010 106.880 157.055 ;
        RECT 109.370 157.010 109.660 157.055 ;
        RECT 111.230 157.010 111.520 157.055 ;
        RECT 106.590 156.870 111.520 157.010 ;
        RECT 106.590 156.825 106.880 156.870 ;
        RECT 109.370 156.825 109.660 156.870 ;
        RECT 111.230 156.825 111.520 156.870 ;
        RECT 93.740 156.530 95.810 156.670 ;
        RECT 93.740 156.470 94.060 156.530 ;
        RECT 78.115 156.145 78.405 156.375 ;
        RECT 78.560 156.330 78.880 156.390 ;
        RECT 79.035 156.330 79.325 156.375 ;
        RECT 78.560 156.190 79.325 156.330 ;
        RECT 78.560 156.130 78.880 156.190 ;
        RECT 79.035 156.145 79.325 156.190 ;
        RECT 79.480 156.330 79.800 156.390 ;
        RECT 80.875 156.330 81.165 156.375 ;
        RECT 79.480 156.190 81.165 156.330 ;
        RECT 79.480 156.130 79.800 156.190 ;
        RECT 80.875 156.145 81.165 156.190 ;
        RECT 86.855 156.145 87.145 156.375 ;
        RECT 88.680 156.330 89.000 156.390 ;
        RECT 89.155 156.330 89.445 156.375 ;
        RECT 88.680 156.190 89.445 156.330 ;
        RECT 80.400 155.990 80.720 156.050 ;
        RECT 76.810 155.850 80.720 155.990 ;
        RECT 86.930 155.990 87.070 156.145 ;
        RECT 88.680 156.130 89.000 156.190 ;
        RECT 89.155 156.145 89.445 156.190 ;
        RECT 89.615 156.330 89.905 156.375 ;
        RECT 90.060 156.330 90.380 156.390 ;
        RECT 89.615 156.190 90.380 156.330 ;
        RECT 89.615 156.145 89.905 156.190 ;
        RECT 90.060 156.130 90.380 156.190 ;
        RECT 90.590 156.330 90.880 156.375 ;
        RECT 91.440 156.330 91.760 156.390 ;
        RECT 90.590 156.190 91.760 156.330 ;
        RECT 90.590 156.145 90.880 156.190 ;
        RECT 91.440 156.130 91.760 156.190 ;
        RECT 92.375 156.330 92.665 156.375 ;
        RECT 94.200 156.330 94.520 156.390 ;
        RECT 92.375 156.190 94.520 156.330 ;
        RECT 92.375 156.145 92.665 156.190 ;
        RECT 94.200 156.130 94.520 156.190 ;
        RECT 95.120 156.130 95.440 156.390 ;
        RECT 95.670 156.375 95.810 156.530 ;
        RECT 96.590 156.530 99.950 156.670 ;
        RECT 109.855 156.670 110.145 156.715 ;
        RECT 110.760 156.670 111.080 156.730 ;
        RECT 109.855 156.530 111.080 156.670 ;
        RECT 95.595 156.145 95.885 156.375 ;
        RECT 96.055 156.315 96.345 156.375 ;
        RECT 96.590 156.315 96.730 156.530 ;
        RECT 109.855 156.485 110.145 156.530 ;
        RECT 110.760 156.470 111.080 156.530 ;
        RECT 96.055 156.175 96.730 156.315 ;
        RECT 96.975 156.330 97.265 156.375 ;
        RECT 97.420 156.330 97.740 156.390 ;
        RECT 96.975 156.190 97.740 156.330 ;
        RECT 96.055 156.145 96.345 156.175 ;
        RECT 96.975 156.145 97.265 156.190 ;
        RECT 90.995 155.990 91.285 156.035 ;
        RECT 93.755 155.990 94.045 156.035 ;
        RECT 86.930 155.850 90.805 155.990 ;
        RECT 75.355 155.805 75.645 155.850 ;
        RECT 75.815 155.805 76.105 155.850 ;
        RECT 80.400 155.790 80.720 155.850 ;
        RECT 69.820 155.650 70.140 155.710 ;
        RECT 68.530 155.510 70.140 155.650 ;
        RECT 69.820 155.450 70.140 155.510 ;
        RECT 73.055 155.650 73.345 155.695 ;
        RECT 79.480 155.650 79.800 155.710 ;
        RECT 73.055 155.510 79.800 155.650 ;
        RECT 73.055 155.465 73.345 155.510 ;
        RECT 79.480 155.450 79.800 155.510 ;
        RECT 81.335 155.650 81.625 155.695 ;
        RECT 81.780 155.650 82.100 155.710 ;
        RECT 81.335 155.510 82.100 155.650 ;
        RECT 81.335 155.465 81.625 155.510 ;
        RECT 81.780 155.450 82.100 155.510 ;
        RECT 83.175 155.650 83.465 155.695 ;
        RECT 86.380 155.650 86.700 155.710 ;
        RECT 83.175 155.510 86.700 155.650 ;
        RECT 83.175 155.465 83.465 155.510 ;
        RECT 86.380 155.450 86.700 155.510 ;
        RECT 87.760 155.650 88.080 155.710 ;
        RECT 88.235 155.650 88.525 155.695 ;
        RECT 87.760 155.510 88.525 155.650 ;
        RECT 90.665 155.650 90.805 155.850 ;
        RECT 90.995 155.850 94.045 155.990 ;
        RECT 90.995 155.805 91.285 155.850 ;
        RECT 93.755 155.805 94.045 155.850 ;
        RECT 92.360 155.650 92.680 155.710 ;
        RECT 90.665 155.510 92.680 155.650 ;
        RECT 87.760 155.450 88.080 155.510 ;
        RECT 88.235 155.465 88.525 155.510 ;
        RECT 92.360 155.450 92.680 155.510 ;
        RECT 93.295 155.650 93.585 155.695 ;
        RECT 95.120 155.650 95.440 155.710 ;
        RECT 93.295 155.510 95.440 155.650 ;
        RECT 95.670 155.650 95.810 156.145 ;
        RECT 97.420 156.130 97.740 156.190 ;
        RECT 97.880 156.330 98.200 156.390 ;
        RECT 98.815 156.330 99.105 156.375 ;
        RECT 97.880 156.190 99.105 156.330 ;
        RECT 97.880 156.130 98.200 156.190 ;
        RECT 98.815 156.145 99.105 156.190 ;
        RECT 99.260 156.130 99.580 156.390 ;
        RECT 99.735 156.145 100.025 156.375 ;
        RECT 100.180 156.330 100.500 156.390 ;
        RECT 100.655 156.330 100.945 156.375 ;
        RECT 100.180 156.190 100.945 156.330 ;
        RECT 99.810 155.990 99.950 156.145 ;
        RECT 100.180 156.130 100.500 156.190 ;
        RECT 100.655 156.145 100.945 156.190 ;
        RECT 101.115 156.330 101.405 156.375 ;
        RECT 102.480 156.330 102.800 156.390 ;
        RECT 101.115 156.190 102.800 156.330 ;
        RECT 101.115 156.145 101.405 156.190 ;
        RECT 102.480 156.130 102.800 156.190 ;
        RECT 106.590 156.330 106.880 156.375 ;
        RECT 111.695 156.330 111.985 156.375 ;
        RECT 106.590 156.190 109.125 156.330 ;
        RECT 106.590 156.145 106.880 156.190 ;
        RECT 98.890 155.850 99.950 155.990 ;
        RECT 104.730 155.990 105.020 156.035 ;
        RECT 107.080 155.990 107.400 156.050 ;
        RECT 108.910 156.035 109.125 156.190 ;
        RECT 111.310 156.190 111.985 156.330 ;
        RECT 107.990 155.990 108.280 156.035 ;
        RECT 104.730 155.850 108.280 155.990 ;
        RECT 98.890 155.710 99.030 155.850 ;
        RECT 104.730 155.805 105.020 155.850 ;
        RECT 107.080 155.790 107.400 155.850 ;
        RECT 107.990 155.805 108.280 155.850 ;
        RECT 108.910 155.990 109.200 156.035 ;
        RECT 110.770 155.990 111.060 156.035 ;
        RECT 108.910 155.850 111.060 155.990 ;
        RECT 108.910 155.805 109.200 155.850 ;
        RECT 110.770 155.805 111.060 155.850 ;
        RECT 96.040 155.650 96.360 155.710 ;
        RECT 95.670 155.510 96.360 155.650 ;
        RECT 93.295 155.465 93.585 155.510 ;
        RECT 95.120 155.450 95.440 155.510 ;
        RECT 96.040 155.450 96.360 155.510 ;
        RECT 97.435 155.650 97.725 155.695 ;
        RECT 97.880 155.650 98.200 155.710 ;
        RECT 97.435 155.510 98.200 155.650 ;
        RECT 97.435 155.465 97.725 155.510 ;
        RECT 97.880 155.450 98.200 155.510 ;
        RECT 98.800 155.450 99.120 155.710 ;
        RECT 101.560 155.450 101.880 155.710 ;
        RECT 110.300 155.650 110.620 155.710 ;
        RECT 111.310 155.650 111.450 156.190 ;
        RECT 111.695 156.145 111.985 156.190 ;
        RECT 110.300 155.510 111.450 155.650 ;
        RECT 110.300 155.450 110.620 155.510 ;
        RECT 26.970 154.830 113.450 155.310 ;
        RECT 31.640 154.630 31.960 154.690 ;
        RECT 33.020 154.630 33.340 154.690 ;
        RECT 31.640 154.490 33.340 154.630 ;
        RECT 31.640 154.430 31.960 154.490 ;
        RECT 33.020 154.430 33.340 154.490 ;
        RECT 35.780 154.630 36.100 154.690 ;
        RECT 39.460 154.630 39.780 154.690 ;
        RECT 42.695 154.630 42.985 154.675 ;
        RECT 43.140 154.630 43.460 154.690 ;
        RECT 35.780 154.490 37.390 154.630 ;
        RECT 35.780 154.430 36.100 154.490 ;
        RECT 37.250 154.350 37.390 154.490 ;
        RECT 39.460 154.490 43.460 154.630 ;
        RECT 39.460 154.430 39.780 154.490 ;
        RECT 42.695 154.445 42.985 154.490 ;
        RECT 43.140 154.430 43.460 154.490 ;
        RECT 44.060 154.630 44.380 154.690 ;
        RECT 49.135 154.630 49.425 154.675 ;
        RECT 44.060 154.490 49.425 154.630 ;
        RECT 44.060 154.430 44.380 154.490 ;
        RECT 49.135 154.445 49.425 154.490 ;
        RECT 50.960 154.630 51.280 154.690 ;
        RECT 51.665 154.630 51.955 154.675 ;
        RECT 54.640 154.630 54.960 154.690 ;
        RECT 62.000 154.630 62.320 154.690 ;
        RECT 50.960 154.490 62.320 154.630 ;
        RECT 50.960 154.430 51.280 154.490 ;
        RECT 51.665 154.445 51.955 154.490 ;
        RECT 54.640 154.430 54.960 154.490 ;
        RECT 62.000 154.430 62.320 154.490 ;
        RECT 85.460 154.630 85.780 154.690 ;
        RECT 88.235 154.630 88.525 154.675 ;
        RECT 85.460 154.490 88.525 154.630 ;
        RECT 85.460 154.430 85.780 154.490 ;
        RECT 88.235 154.445 88.525 154.490 ;
        RECT 94.660 154.430 94.980 154.690 ;
        RECT 97.420 154.430 97.740 154.690 ;
        RECT 97.895 154.630 98.185 154.675 ;
        RECT 99.260 154.630 99.580 154.690 ;
        RECT 97.895 154.490 99.580 154.630 ;
        RECT 97.895 154.445 98.185 154.490 ;
        RECT 99.260 154.430 99.580 154.490 ;
        RECT 99.735 154.445 100.025 154.675 ;
        RECT 29.340 154.290 29.660 154.350 ;
        RECT 30.670 154.290 30.960 154.335 ;
        RECT 33.930 154.290 34.220 154.335 ;
        RECT 29.340 154.150 34.220 154.290 ;
        RECT 29.340 154.090 29.660 154.150 ;
        RECT 30.670 154.105 30.960 154.150 ;
        RECT 33.930 154.105 34.220 154.150 ;
        RECT 34.850 154.290 35.140 154.335 ;
        RECT 36.710 154.290 37.000 154.335 ;
        RECT 34.850 154.150 37.000 154.290 ;
        RECT 34.850 154.105 35.140 154.150 ;
        RECT 36.710 154.105 37.000 154.150 ;
        RECT 37.160 154.290 37.480 154.350 ;
        RECT 38.095 154.290 38.385 154.335 ;
        RECT 44.980 154.290 45.300 154.350 ;
        RECT 37.160 154.150 43.830 154.290 ;
        RECT 32.530 153.950 32.820 153.995 ;
        RECT 34.850 153.950 35.065 154.105 ;
        RECT 37.160 154.090 37.480 154.150 ;
        RECT 38.095 154.105 38.385 154.150 ;
        RECT 32.530 153.810 35.065 153.950 ;
        RECT 32.530 153.765 32.820 153.810 ;
        RECT 35.780 153.750 36.100 154.010 ;
        RECT 37.620 153.750 37.940 154.010 ;
        RECT 39.935 153.950 40.225 153.995 ;
        RECT 42.220 153.950 42.540 154.010 ;
        RECT 39.935 153.810 42.540 153.950 ;
        RECT 39.935 153.765 40.225 153.810 ;
        RECT 42.220 153.750 42.540 153.810 ;
        RECT 39.000 153.610 39.320 153.670 ;
        RECT 43.690 153.655 43.830 154.150 ;
        RECT 44.150 154.150 45.300 154.290 ;
        RECT 44.150 154.010 44.290 154.150 ;
        RECT 44.980 154.090 45.300 154.150 ;
        RECT 46.360 154.290 46.680 154.350 ;
        RECT 67.060 154.335 67.380 154.350 ;
        RECT 53.670 154.290 53.960 154.335 ;
        RECT 56.930 154.290 57.220 154.335 ;
        RECT 46.360 154.150 57.220 154.290 ;
        RECT 46.360 154.090 46.680 154.150 ;
        RECT 53.670 154.105 53.960 154.150 ;
        RECT 56.930 154.105 57.220 154.150 ;
        RECT 57.850 154.290 58.140 154.335 ;
        RECT 59.710 154.290 60.000 154.335 ;
        RECT 57.850 154.150 60.000 154.290 ;
        RECT 57.850 154.105 58.140 154.150 ;
        RECT 59.710 154.105 60.000 154.150 ;
        RECT 63.495 154.290 63.785 154.335 ;
        RECT 66.735 154.290 67.385 154.335 ;
        RECT 63.495 154.150 67.385 154.290 ;
        RECT 63.495 154.105 64.085 154.150 ;
        RECT 66.735 154.105 67.385 154.150 ;
        RECT 44.060 153.750 44.380 154.010 ;
        RECT 45.440 153.950 45.760 154.010 ;
        RECT 45.915 153.950 46.205 153.995 ;
        RECT 45.440 153.810 46.205 153.950 ;
        RECT 45.440 153.750 45.760 153.810 ;
        RECT 45.915 153.765 46.205 153.810 ;
        RECT 46.820 153.750 47.140 154.010 ;
        RECT 47.295 153.950 47.585 153.995 ;
        RECT 49.580 153.950 49.900 154.010 ;
        RECT 47.295 153.810 49.900 153.950 ;
        RECT 47.295 153.765 47.585 153.810 ;
        RECT 49.580 153.750 49.900 153.810 ;
        RECT 50.040 153.950 50.360 154.010 ;
        RECT 51.880 153.950 52.200 154.010 ;
        RECT 55.530 153.950 55.820 153.995 ;
        RECT 57.850 153.950 58.065 154.105 ;
        RECT 50.040 153.810 54.870 153.950 ;
        RECT 50.040 153.750 50.360 153.810 ;
        RECT 51.880 153.750 52.200 153.810 ;
        RECT 43.155 153.610 43.445 153.655 ;
        RECT 39.000 153.470 43.445 153.610 ;
        RECT 39.000 153.410 39.320 153.470 ;
        RECT 43.155 153.425 43.445 153.470 ;
        RECT 43.615 153.425 43.905 153.655 ;
        RECT 44.980 153.610 45.300 153.670 ;
        RECT 50.975 153.610 51.265 153.655 ;
        RECT 54.180 153.610 54.500 153.670 ;
        RECT 44.980 153.470 51.265 153.610 ;
        RECT 44.980 153.410 45.300 153.470 ;
        RECT 50.975 153.425 51.265 153.470 ;
        RECT 51.510 153.470 54.500 153.610 ;
        RECT 32.530 153.270 32.820 153.315 ;
        RECT 35.310 153.270 35.600 153.315 ;
        RECT 37.170 153.270 37.460 153.315 ;
        RECT 32.530 153.130 37.460 153.270 ;
        RECT 32.530 153.085 32.820 153.130 ;
        RECT 35.310 153.085 35.600 153.130 ;
        RECT 37.170 153.085 37.460 153.130 ;
        RECT 42.680 153.270 43.000 153.330 ;
        RECT 51.510 153.270 51.650 153.470 ;
        RECT 54.180 153.410 54.500 153.470 ;
        RECT 42.680 153.130 51.650 153.270 ;
        RECT 42.680 153.070 43.000 153.130 ;
        RECT 28.665 152.930 28.955 152.975 ;
        RECT 32.100 152.930 32.420 152.990 ;
        RECT 28.665 152.790 32.420 152.930 ;
        RECT 28.665 152.745 28.955 152.790 ;
        RECT 32.100 152.730 32.420 152.790 ;
        RECT 36.240 152.930 36.560 152.990 ;
        RECT 39.460 152.930 39.780 152.990 ;
        RECT 36.240 152.790 39.780 152.930 ;
        RECT 36.240 152.730 36.560 152.790 ;
        RECT 39.460 152.730 39.780 152.790 ;
        RECT 40.840 152.730 41.160 152.990 ;
        RECT 45.900 152.730 46.220 152.990 ;
        RECT 46.820 152.930 47.140 152.990 ;
        RECT 48.215 152.930 48.505 152.975 ;
        RECT 46.820 152.790 48.505 152.930 ;
        RECT 54.730 152.930 54.870 153.810 ;
        RECT 55.530 153.810 58.065 153.950 ;
        RECT 58.795 153.950 59.085 153.995 ;
        RECT 61.080 153.950 61.400 154.010 ;
        RECT 58.795 153.810 61.400 153.950 ;
        RECT 55.530 153.765 55.820 153.810 ;
        RECT 58.795 153.765 59.085 153.810 ;
        RECT 61.080 153.750 61.400 153.810 ;
        RECT 63.795 153.790 64.085 154.105 ;
        RECT 67.060 154.090 67.380 154.105 ;
        RECT 69.360 154.090 69.680 154.350 ;
        RECT 73.975 154.290 74.265 154.335 ;
        RECT 74.895 154.290 75.185 154.335 ;
        RECT 73.975 154.150 75.185 154.290 ;
        RECT 73.975 154.105 74.265 154.150 ;
        RECT 74.895 154.105 75.185 154.150 ;
        RECT 80.810 154.290 81.100 154.335 ;
        RECT 82.240 154.290 82.560 154.350 ;
        RECT 84.070 154.290 84.360 154.335 ;
        RECT 80.810 154.150 84.360 154.290 ;
        RECT 80.810 154.105 81.100 154.150 ;
        RECT 82.240 154.090 82.560 154.150 ;
        RECT 84.070 154.105 84.360 154.150 ;
        RECT 84.990 154.290 85.280 154.335 ;
        RECT 86.850 154.290 87.140 154.335 ;
        RECT 84.990 154.150 87.140 154.290 ;
        RECT 84.990 154.105 85.280 154.150 ;
        RECT 86.850 154.105 87.140 154.150 ;
        RECT 89.615 154.290 89.905 154.335 ;
        RECT 92.375 154.290 92.665 154.335 ;
        RECT 94.750 154.290 94.890 154.430 ;
        RECT 97.510 154.290 97.650 154.430 ;
        RECT 89.615 154.150 92.665 154.290 ;
        RECT 89.615 154.105 89.905 154.150 ;
        RECT 92.375 154.105 92.665 154.150 ;
        RECT 93.830 154.150 94.890 154.290 ;
        RECT 95.670 154.150 97.650 154.290 ;
        RECT 64.875 153.950 65.165 153.995 ;
        RECT 68.455 153.950 68.745 153.995 ;
        RECT 70.290 153.950 70.580 153.995 ;
        RECT 64.875 153.810 70.580 153.950 ;
        RECT 64.875 153.765 65.165 153.810 ;
        RECT 68.455 153.765 68.745 153.810 ;
        RECT 70.290 153.765 70.580 153.810 ;
        RECT 72.580 153.750 72.900 154.010 ;
        RECT 76.260 153.750 76.580 154.010 ;
        RECT 76.720 153.750 77.040 154.010 ;
        RECT 77.195 153.765 77.485 153.995 ;
        RECT 78.115 153.950 78.405 153.995 ;
        RECT 78.560 153.950 78.880 154.010 ;
        RECT 79.940 153.950 80.260 154.010 ;
        RECT 78.115 153.810 80.260 153.950 ;
        RECT 78.115 153.765 78.405 153.810 ;
        RECT 56.480 153.610 56.800 153.670 ;
        RECT 60.635 153.610 60.925 153.655 ;
        RECT 56.480 153.470 60.925 153.610 ;
        RECT 56.480 153.410 56.800 153.470 ;
        RECT 60.635 153.425 60.925 153.470 ;
        RECT 70.740 153.410 71.060 153.670 ;
        RECT 73.515 153.610 73.805 153.655 ;
        RECT 75.340 153.610 75.660 153.670 ;
        RECT 73.515 153.470 75.660 153.610 ;
        RECT 73.515 153.425 73.805 153.470 ;
        RECT 75.340 153.410 75.660 153.470 ;
        RECT 55.530 153.270 55.820 153.315 ;
        RECT 58.310 153.270 58.600 153.315 ;
        RECT 60.170 153.270 60.460 153.315 ;
        RECT 55.530 153.130 60.460 153.270 ;
        RECT 55.530 153.085 55.820 153.130 ;
        RECT 58.310 153.085 58.600 153.130 ;
        RECT 60.170 153.085 60.460 153.130 ;
        RECT 64.875 153.270 65.165 153.315 ;
        RECT 67.995 153.270 68.285 153.315 ;
        RECT 69.885 153.270 70.175 153.315 ;
        RECT 64.875 153.130 70.175 153.270 ;
        RECT 64.875 153.085 65.165 153.130 ;
        RECT 67.995 153.085 68.285 153.130 ;
        RECT 69.885 153.085 70.175 153.130 ;
        RECT 56.940 152.930 57.260 152.990 ;
        RECT 54.730 152.790 57.260 152.930 ;
        RECT 46.820 152.730 47.140 152.790 ;
        RECT 48.215 152.745 48.505 152.790 ;
        RECT 56.940 152.730 57.260 152.790 ;
        RECT 62.000 152.730 62.320 152.990 ;
        RECT 71.660 152.730 71.980 152.990 ;
        RECT 73.960 152.730 74.280 152.990 ;
        RECT 77.270 152.930 77.410 153.765 ;
        RECT 78.560 153.750 78.880 153.810 ;
        RECT 79.940 153.750 80.260 153.810 ;
        RECT 82.670 153.950 82.960 153.995 ;
        RECT 84.990 153.950 85.205 154.105 ;
        RECT 82.670 153.810 85.205 153.950 ;
        RECT 86.380 153.950 86.700 154.010 ;
        RECT 89.155 153.950 89.445 153.995 ;
        RECT 86.380 153.810 89.445 153.950 ;
        RECT 82.670 153.765 82.960 153.810 ;
        RECT 86.380 153.750 86.700 153.810 ;
        RECT 89.155 153.765 89.445 153.810 ;
        RECT 90.520 153.750 90.840 154.010 ;
        RECT 90.980 153.750 91.300 154.010 ;
        RECT 93.830 153.995 93.970 154.150 ;
        RECT 93.755 153.765 94.045 153.995 ;
        RECT 94.215 153.765 94.505 153.995 ;
        RECT 85.920 153.410 86.240 153.670 ;
        RECT 86.840 153.610 87.160 153.670 ;
        RECT 87.775 153.610 88.065 153.655 ;
        RECT 86.840 153.470 88.065 153.610 ;
        RECT 94.290 153.610 94.430 153.765 ;
        RECT 94.660 153.750 94.980 154.010 ;
        RECT 95.670 153.995 95.810 154.150 ;
        RECT 95.595 153.765 95.885 153.995 ;
        RECT 97.435 153.950 97.725 153.995 ;
        RECT 98.800 153.950 99.120 154.010 ;
        RECT 97.435 153.810 99.120 153.950 ;
        RECT 99.810 153.950 99.950 154.445 ;
        RECT 101.560 154.290 101.880 154.350 ;
        RECT 104.730 154.290 105.020 154.335 ;
        RECT 107.990 154.290 108.280 154.335 ;
        RECT 101.560 154.150 108.280 154.290 ;
        RECT 101.560 154.090 101.880 154.150 ;
        RECT 104.730 154.105 105.020 154.150 ;
        RECT 107.990 154.105 108.280 154.150 ;
        RECT 108.910 154.290 109.200 154.335 ;
        RECT 110.770 154.290 111.060 154.335 ;
        RECT 108.910 154.150 111.060 154.290 ;
        RECT 108.910 154.105 109.200 154.150 ;
        RECT 110.770 154.105 111.060 154.150 ;
        RECT 101.115 153.950 101.405 153.995 ;
        RECT 99.810 153.810 101.405 153.950 ;
        RECT 97.435 153.765 97.725 153.810 ;
        RECT 98.800 153.750 99.120 153.810 ;
        RECT 101.115 153.765 101.405 153.810 ;
        RECT 106.590 153.950 106.880 153.995 ;
        RECT 108.910 153.950 109.125 154.105 ;
        RECT 106.590 153.810 109.125 153.950 ;
        RECT 106.590 153.765 106.880 153.810 ;
        RECT 96.040 153.610 96.360 153.670 ;
        RECT 94.290 153.470 96.360 153.610 ;
        RECT 86.840 153.410 87.160 153.470 ;
        RECT 87.775 153.425 88.065 153.470 ;
        RECT 96.040 153.410 96.360 153.470 ;
        RECT 96.500 153.610 96.820 153.670 ;
        RECT 99.260 153.610 99.580 153.670 ;
        RECT 109.855 153.610 110.145 153.655 ;
        RECT 96.500 153.470 99.580 153.610 ;
        RECT 96.500 153.410 96.820 153.470 ;
        RECT 99.260 153.410 99.580 153.470 ;
        RECT 105.100 153.470 110.145 153.610 ;
        RECT 82.670 153.270 82.960 153.315 ;
        RECT 85.450 153.270 85.740 153.315 ;
        RECT 87.310 153.270 87.600 153.315 ;
        RECT 82.670 153.130 87.600 153.270 ;
        RECT 82.670 153.085 82.960 153.130 ;
        RECT 85.450 153.085 85.740 153.130 ;
        RECT 87.310 153.085 87.600 153.130 ;
        RECT 102.035 153.270 102.325 153.315 ;
        RECT 105.100 153.270 105.240 153.470 ;
        RECT 109.855 153.425 110.145 153.470 ;
        RECT 110.300 153.610 110.620 153.670 ;
        RECT 111.695 153.610 111.985 153.655 ;
        RECT 110.300 153.470 111.985 153.610 ;
        RECT 110.300 153.410 110.620 153.470 ;
        RECT 111.695 153.425 111.985 153.470 ;
        RECT 102.035 153.130 105.240 153.270 ;
        RECT 106.590 153.270 106.880 153.315 ;
        RECT 109.370 153.270 109.660 153.315 ;
        RECT 111.230 153.270 111.520 153.315 ;
        RECT 106.590 153.130 111.520 153.270 ;
        RECT 102.035 153.085 102.325 153.130 ;
        RECT 106.590 153.085 106.880 153.130 ;
        RECT 109.370 153.085 109.660 153.130 ;
        RECT 111.230 153.085 111.520 153.130 ;
        RECT 78.805 152.930 79.095 152.975 ;
        RECT 81.780 152.930 82.100 152.990 ;
        RECT 77.270 152.790 82.100 152.930 ;
        RECT 78.805 152.745 79.095 152.790 ;
        RECT 81.780 152.730 82.100 152.790 ;
        RECT 90.520 152.730 90.840 152.990 ;
        RECT 91.900 152.730 92.220 152.990 ;
        RECT 92.360 152.930 92.680 152.990 ;
        RECT 94.660 152.930 94.980 152.990 ;
        RECT 92.360 152.790 94.980 152.930 ;
        RECT 92.360 152.730 92.680 152.790 ;
        RECT 94.660 152.730 94.980 152.790 ;
        RECT 98.800 152.930 99.120 152.990 ;
        RECT 102.725 152.930 103.015 152.975 ;
        RECT 103.400 152.930 103.720 152.990 ;
        RECT 98.800 152.790 103.720 152.930 ;
        RECT 98.800 152.730 99.120 152.790 ;
        RECT 102.725 152.745 103.015 152.790 ;
        RECT 103.400 152.730 103.720 152.790 ;
        RECT 26.970 152.110 113.450 152.590 ;
        RECT 28.880 151.910 29.200 151.970 ;
        RECT 31.655 151.910 31.945 151.955 ;
        RECT 28.880 151.770 31.945 151.910 ;
        RECT 28.880 151.710 29.200 151.770 ;
        RECT 31.655 151.725 31.945 151.770 ;
        RECT 36.330 151.770 44.750 151.910 ;
        RECT 31.195 151.570 31.485 151.615 ;
        RECT 36.330 151.570 36.470 151.770 ;
        RECT 31.195 151.430 36.470 151.570 ;
        RECT 36.720 151.570 37.010 151.615 ;
        RECT 38.580 151.570 38.870 151.615 ;
        RECT 41.360 151.570 41.650 151.615 ;
        RECT 36.720 151.430 41.650 151.570 ;
        RECT 44.610 151.570 44.750 151.770 ;
        RECT 46.360 151.710 46.680 151.970 ;
        RECT 47.755 151.725 48.045 151.955 ;
        RECT 50.960 151.910 51.280 151.970 ;
        RECT 48.750 151.770 51.280 151.910 ;
        RECT 47.830 151.570 47.970 151.725 ;
        RECT 44.610 151.430 47.970 151.570 ;
        RECT 31.195 151.385 31.485 151.430 ;
        RECT 36.720 151.385 37.010 151.430 ;
        RECT 38.580 151.385 38.870 151.430 ;
        RECT 41.360 151.385 41.650 151.430 ;
        RECT 28.880 151.230 29.200 151.290 ;
        RECT 34.875 151.230 35.165 151.275 ;
        RECT 37.160 151.230 37.480 151.290 ;
        RECT 28.880 151.090 30.490 151.230 ;
        RECT 28.880 151.030 29.200 151.090 ;
        RECT 30.350 150.950 30.490 151.090 ;
        RECT 34.875 151.090 37.480 151.230 ;
        RECT 34.875 151.045 35.165 151.090 ;
        RECT 37.160 151.030 37.480 151.090 ;
        RECT 42.680 151.230 43.000 151.290 ;
        RECT 48.750 151.275 48.890 151.770 ;
        RECT 50.960 151.710 51.280 151.770 ;
        RECT 67.520 151.910 67.840 151.970 ;
        RECT 72.580 151.910 72.900 151.970 ;
        RECT 67.520 151.770 72.900 151.910 ;
        RECT 67.520 151.710 67.840 151.770 ;
        RECT 72.580 151.710 72.900 151.770 ;
        RECT 79.035 151.910 79.325 151.955 ;
        RECT 85.920 151.910 86.240 151.970 ;
        RECT 79.035 151.770 86.240 151.910 ;
        RECT 79.035 151.725 79.325 151.770 ;
        RECT 85.920 151.710 86.240 151.770 ;
        RECT 90.520 151.710 90.840 151.970 ;
        RECT 97.420 151.710 97.740 151.970 ;
        RECT 100.640 151.710 100.960 151.970 ;
        RECT 110.760 151.710 111.080 151.970 ;
        RECT 53.735 151.570 54.025 151.615 ;
        RECT 56.020 151.570 56.340 151.630 ;
        RECT 53.735 151.430 56.340 151.570 ;
        RECT 53.735 151.385 54.025 151.430 ;
        RECT 56.020 151.370 56.340 151.430 ;
        RECT 67.030 151.570 67.320 151.615 ;
        RECT 69.810 151.570 70.100 151.615 ;
        RECT 71.670 151.570 71.960 151.615 ;
        RECT 67.030 151.430 71.960 151.570 ;
        RECT 67.030 151.385 67.320 151.430 ;
        RECT 69.810 151.385 70.100 151.430 ;
        RECT 71.670 151.385 71.960 151.430 ;
        RECT 73.975 151.385 74.265 151.615 ;
        RECT 79.495 151.385 79.785 151.615 ;
        RECT 84.540 151.570 84.860 151.630 ;
        RECT 90.980 151.570 91.300 151.630 ;
        RECT 84.540 151.430 91.300 151.570 ;
        RECT 45.225 151.230 45.515 151.275 ;
        RECT 42.680 151.090 45.515 151.230 ;
        RECT 42.680 151.030 43.000 151.090 ;
        RECT 45.225 151.045 45.515 151.090 ;
        RECT 48.675 151.045 48.965 151.275 ;
        RECT 50.975 151.230 51.265 151.275 ;
        RECT 54.640 151.230 54.960 151.290 ;
        RECT 58.335 151.230 58.625 151.275 ;
        RECT 62.000 151.230 62.320 151.290 ;
        RECT 50.975 151.090 54.960 151.230 ;
        RECT 50.975 151.045 51.265 151.090 ;
        RECT 54.640 151.030 54.960 151.090 ;
        RECT 56.570 151.090 62.320 151.230 ;
        RECT 29.815 150.705 30.105 150.935 ;
        RECT 29.890 150.210 30.030 150.705 ;
        RECT 30.260 150.690 30.580 150.950 ;
        RECT 32.100 150.890 32.420 150.950 ;
        RECT 33.495 150.890 33.785 150.935 ;
        RECT 32.100 150.750 33.785 150.890 ;
        RECT 32.100 150.690 32.420 150.750 ;
        RECT 33.495 150.705 33.785 150.750 ;
        RECT 33.955 150.890 34.245 150.935 ;
        RECT 35.780 150.890 36.100 150.950 ;
        RECT 33.955 150.750 36.100 150.890 ;
        RECT 33.955 150.705 34.245 150.750 ;
        RECT 35.780 150.690 36.100 150.750 ;
        RECT 36.240 150.690 36.560 150.950 ;
        RECT 38.080 150.690 38.400 150.950 ;
        RECT 41.360 150.890 41.650 150.935 ;
        RECT 39.115 150.750 41.650 150.890 ;
        RECT 39.115 150.595 39.330 150.750 ;
        RECT 41.360 150.705 41.650 150.750 ;
        RECT 45.915 150.890 46.205 150.935 ;
        RECT 46.360 150.890 46.680 150.950 ;
        RECT 45.915 150.750 46.680 150.890 ;
        RECT 45.915 150.705 46.205 150.750 ;
        RECT 46.360 150.690 46.680 150.750 ;
        RECT 49.135 150.890 49.425 150.935 ;
        RECT 49.580 150.890 49.900 150.950 ;
        RECT 49.135 150.750 49.900 150.890 ;
        RECT 49.135 150.705 49.425 150.750 ;
        RECT 49.580 150.690 49.900 150.750 ;
        RECT 53.720 150.890 54.040 150.950 ;
        RECT 56.570 150.935 56.710 151.090 ;
        RECT 58.335 151.045 58.625 151.090 ;
        RECT 62.000 151.030 62.320 151.090 ;
        RECT 70.295 151.230 70.585 151.275 ;
        RECT 74.050 151.230 74.190 151.385 ;
        RECT 70.295 151.090 74.190 151.230 ;
        RECT 70.295 151.045 70.585 151.090 ;
        RECT 55.575 150.890 55.865 150.935 ;
        RECT 53.720 150.750 55.865 150.890 ;
        RECT 53.720 150.690 54.040 150.750 ;
        RECT 55.575 150.705 55.865 150.750 ;
        RECT 56.035 150.705 56.325 150.935 ;
        RECT 56.495 150.705 56.785 150.935 ;
        RECT 57.415 150.890 57.705 150.935 ;
        RECT 59.240 150.890 59.560 150.950 ;
        RECT 57.415 150.750 59.560 150.890 ;
        RECT 57.415 150.705 57.705 150.750 ;
        RECT 37.180 150.550 37.470 150.595 ;
        RECT 39.040 150.550 39.330 150.595 ;
        RECT 37.180 150.410 39.330 150.550 ;
        RECT 37.180 150.365 37.470 150.410 ;
        RECT 39.040 150.365 39.330 150.410 ;
        RECT 39.920 150.595 40.240 150.610 ;
        RECT 39.920 150.550 40.250 150.595 ;
        RECT 43.220 150.550 43.510 150.595 ;
        RECT 39.920 150.410 43.510 150.550 ;
        RECT 39.920 150.365 40.250 150.410 ;
        RECT 43.220 150.365 43.510 150.410 ;
        RECT 47.755 150.550 48.045 150.595 ;
        RECT 54.195 150.550 54.485 150.595 ;
        RECT 47.755 150.410 54.485 150.550 ;
        RECT 56.110 150.550 56.250 150.705 ;
        RECT 57.860 150.550 58.180 150.610 ;
        RECT 56.110 150.410 58.180 150.550 ;
        RECT 47.755 150.365 48.045 150.410 ;
        RECT 54.195 150.365 54.485 150.410 ;
        RECT 39.920 150.350 40.240 150.365 ;
        RECT 57.860 150.350 58.180 150.410 ;
        RECT 30.260 150.210 30.580 150.270 ;
        RECT 29.890 150.070 30.580 150.210 ;
        RECT 30.260 150.010 30.580 150.070 ;
        RECT 31.180 150.210 31.500 150.270 ;
        RECT 45.900 150.210 46.220 150.270 ;
        RECT 31.180 150.070 46.220 150.210 ;
        RECT 31.180 150.010 31.500 150.070 ;
        RECT 45.900 150.010 46.220 150.070 ;
        RECT 50.055 150.210 50.345 150.255 ;
        RECT 52.340 150.210 52.660 150.270 ;
        RECT 50.055 150.070 52.660 150.210 ;
        RECT 50.055 150.025 50.345 150.070 ;
        RECT 52.340 150.010 52.660 150.070 ;
        RECT 55.560 150.210 55.880 150.270 ;
        RECT 58.410 150.210 58.550 150.750 ;
        RECT 59.240 150.690 59.560 150.750 ;
        RECT 63.165 150.890 63.455 150.935 ;
        RECT 66.140 150.890 66.460 150.950 ;
        RECT 63.165 150.750 66.460 150.890 ;
        RECT 63.165 150.705 63.455 150.750 ;
        RECT 66.140 150.690 66.460 150.750 ;
        RECT 67.030 150.890 67.320 150.935 ;
        RECT 70.740 150.890 71.060 150.950 ;
        RECT 72.120 150.890 72.440 150.950 ;
        RECT 67.030 150.750 69.565 150.890 ;
        RECT 67.030 150.705 67.320 150.750 ;
        RECT 69.350 150.595 69.565 150.750 ;
        RECT 70.740 150.750 72.440 150.890 ;
        RECT 70.740 150.690 71.060 150.750 ;
        RECT 72.120 150.690 72.440 150.750 ;
        RECT 72.580 150.690 72.900 150.950 ;
        RECT 74.420 150.890 74.740 150.950 ;
        RECT 74.895 150.890 75.185 150.935 ;
        RECT 74.420 150.750 75.185 150.890 ;
        RECT 74.420 150.690 74.740 150.750 ;
        RECT 74.895 150.705 75.185 150.750 ;
        RECT 78.115 150.890 78.405 150.935 ;
        RECT 79.570 150.890 79.710 151.385 ;
        RECT 84.540 151.370 84.860 151.430 ;
        RECT 90.980 151.370 91.300 151.430 ;
        RECT 94.660 151.570 94.980 151.630 ;
        RECT 97.895 151.570 98.185 151.615 ;
        RECT 94.660 151.430 98.185 151.570 ;
        RECT 94.660 151.370 94.980 151.430 ;
        RECT 97.895 151.385 98.185 151.430 ;
        RECT 99.260 151.570 99.580 151.630 ;
        RECT 99.260 151.430 102.250 151.570 ;
        RECT 99.260 151.370 99.580 151.430 ;
        RECT 102.110 151.290 102.250 151.430 ;
        RECT 105.255 151.385 105.545 151.615 ;
        RECT 109.395 151.570 109.685 151.615 ;
        RECT 111.680 151.570 112.000 151.630 ;
        RECT 109.395 151.430 112.000 151.570 ;
        RECT 109.395 151.385 109.685 151.430 ;
        RECT 81.780 151.030 82.100 151.290 ;
        RECT 82.715 151.230 83.005 151.275 ;
        RECT 84.080 151.230 84.400 151.290 ;
        RECT 91.915 151.230 92.205 151.275 ;
        RECT 96.500 151.230 96.820 151.290 ;
        RECT 82.715 151.090 96.820 151.230 ;
        RECT 82.715 151.045 83.005 151.090 ;
        RECT 84.080 151.030 84.400 151.090 ;
        RECT 91.915 151.045 92.205 151.090 ;
        RECT 96.500 151.030 96.820 151.090 ;
        RECT 96.960 151.030 97.280 151.290 ;
        RECT 102.020 151.030 102.340 151.290 ;
        RECT 78.115 150.750 79.710 150.890 ;
        RECT 78.115 150.705 78.405 150.750 ;
        RECT 84.540 150.690 84.860 150.950 ;
        RECT 85.000 150.690 85.320 150.950 ;
        RECT 88.680 150.690 89.000 150.950 ;
        RECT 89.615 150.705 89.905 150.935 ;
        RECT 95.580 150.890 95.900 150.950 ;
        RECT 96.055 150.890 96.345 150.935 ;
        RECT 95.580 150.750 96.345 150.890 ;
        RECT 65.170 150.550 65.460 150.595 ;
        RECT 68.430 150.550 68.720 150.595 ;
        RECT 69.350 150.550 69.640 150.595 ;
        RECT 71.210 150.550 71.500 150.595 ;
        RECT 65.170 150.410 69.130 150.550 ;
        RECT 65.170 150.365 65.460 150.410 ;
        RECT 68.430 150.365 68.720 150.410 ;
        RECT 55.560 150.070 58.550 150.210 ;
        RECT 61.095 150.210 61.385 150.255 ;
        RECT 65.680 150.210 66.000 150.270 ;
        RECT 61.095 150.070 66.000 150.210 ;
        RECT 68.990 150.210 69.130 150.410 ;
        RECT 69.350 150.410 71.500 150.550 ;
        RECT 69.350 150.365 69.640 150.410 ;
        RECT 71.210 150.365 71.500 150.410 ;
        RECT 73.500 150.550 73.820 150.610 ;
        RECT 89.690 150.550 89.830 150.705 ;
        RECT 95.580 150.690 95.900 150.750 ;
        RECT 96.055 150.705 96.345 150.750 ;
        RECT 97.435 150.890 97.725 150.935 ;
        RECT 97.880 150.890 98.200 150.950 ;
        RECT 97.435 150.750 98.200 150.890 ;
        RECT 97.435 150.705 97.725 150.750 ;
        RECT 97.880 150.690 98.200 150.750 ;
        RECT 98.815 150.890 99.105 150.935 ;
        RECT 99.260 150.890 99.580 150.950 ;
        RECT 98.815 150.750 99.580 150.890 ;
        RECT 98.815 150.705 99.105 150.750 ;
        RECT 99.260 150.690 99.580 150.750 ;
        RECT 99.720 150.690 100.040 150.950 ;
        RECT 100.180 150.690 100.500 150.950 ;
        RECT 103.400 150.690 103.720 150.950 ;
        RECT 105.330 150.890 105.470 151.385 ;
        RECT 111.680 151.370 112.000 151.430 ;
        RECT 111.220 151.230 111.540 151.290 ;
        RECT 108.550 151.090 111.540 151.230 ;
        RECT 108.550 150.935 108.690 151.090 ;
        RECT 111.220 151.030 111.540 151.090 ;
        RECT 106.635 150.890 106.925 150.935 ;
        RECT 105.330 150.750 106.925 150.890 ;
        RECT 106.635 150.705 106.925 150.750 ;
        RECT 108.475 150.705 108.765 150.935 ;
        RECT 109.840 150.690 110.160 150.950 ;
        RECT 91.440 150.550 91.760 150.610 ;
        RECT 73.500 150.410 91.760 150.550 ;
        RECT 73.500 150.350 73.820 150.410 ;
        RECT 91.440 150.350 91.760 150.410 ;
        RECT 92.835 150.550 93.125 150.595 ;
        RECT 94.200 150.550 94.520 150.610 ;
        RECT 100.270 150.550 100.410 150.690 ;
        RECT 110.760 150.550 111.080 150.610 ;
        RECT 92.835 150.410 98.110 150.550 ;
        RECT 100.270 150.410 111.080 150.550 ;
        RECT 92.835 150.365 93.125 150.410 ;
        RECT 94.200 150.350 94.520 150.410 ;
        RECT 73.055 150.210 73.345 150.255 ;
        RECT 68.990 150.070 73.345 150.210 ;
        RECT 55.560 150.010 55.880 150.070 ;
        RECT 61.095 150.025 61.385 150.070 ;
        RECT 65.680 150.010 66.000 150.070 ;
        RECT 73.055 150.025 73.345 150.070 ;
        RECT 81.335 150.210 81.625 150.255 ;
        RECT 82.240 150.210 82.560 150.270 ;
        RECT 81.335 150.070 82.560 150.210 ;
        RECT 81.335 150.025 81.625 150.070 ;
        RECT 82.240 150.010 82.560 150.070 ;
        RECT 83.620 150.210 83.940 150.270 ;
        RECT 84.095 150.210 84.385 150.255 ;
        RECT 83.620 150.070 84.385 150.210 ;
        RECT 83.620 150.010 83.940 150.070 ;
        RECT 84.095 150.025 84.385 150.070 ;
        RECT 85.920 150.010 86.240 150.270 ;
        RECT 86.380 150.210 86.700 150.270 ;
        RECT 92.375 150.210 92.665 150.255 ;
        RECT 86.380 150.070 92.665 150.210 ;
        RECT 86.380 150.010 86.700 150.070 ;
        RECT 92.375 150.025 92.665 150.070 ;
        RECT 94.660 150.010 94.980 150.270 ;
        RECT 95.135 150.210 95.425 150.255 ;
        RECT 96.500 150.210 96.820 150.270 ;
        RECT 95.135 150.070 96.820 150.210 ;
        RECT 97.970 150.210 98.110 150.410 ;
        RECT 110.760 150.350 111.080 150.410 ;
        RECT 102.480 150.210 102.800 150.270 ;
        RECT 102.955 150.210 103.245 150.255 ;
        RECT 97.970 150.070 103.245 150.210 ;
        RECT 95.135 150.025 95.425 150.070 ;
        RECT 96.500 150.010 96.820 150.070 ;
        RECT 102.480 150.010 102.800 150.070 ;
        RECT 102.955 150.025 103.245 150.070 ;
        RECT 107.555 150.210 107.845 150.255 ;
        RECT 108.460 150.210 108.780 150.270 ;
        RECT 107.555 150.070 108.780 150.210 ;
        RECT 107.555 150.025 107.845 150.070 ;
        RECT 108.460 150.010 108.780 150.070 ;
        RECT 26.970 149.390 113.450 149.870 ;
        RECT 27.040 149.190 27.360 149.250 ;
        RECT 40.840 149.190 41.160 149.250 ;
        RECT 27.040 149.050 41.160 149.190 ;
        RECT 27.040 148.990 27.360 149.050 ;
        RECT 40.840 148.990 41.160 149.050 ;
        RECT 41.760 149.190 42.080 149.250 ;
        RECT 52.800 149.190 53.120 149.250 ;
        RECT 41.760 149.050 53.120 149.190 ;
        RECT 41.760 148.990 42.080 149.050 ;
        RECT 52.800 148.990 53.120 149.050 ;
        RECT 53.260 149.190 53.580 149.250 ;
        RECT 60.175 149.190 60.465 149.235 ;
        RECT 53.260 149.050 60.465 149.190 ;
        RECT 53.260 148.990 53.580 149.050 ;
        RECT 60.175 149.005 60.465 149.050 ;
        RECT 61.540 149.190 61.860 149.250 ;
        RECT 61.540 149.050 62.230 149.190 ;
        RECT 61.540 148.990 61.860 149.050 ;
        RECT 30.670 148.850 30.960 148.895 ;
        RECT 31.640 148.850 31.960 148.910 ;
        RECT 33.930 148.850 34.220 148.895 ;
        RECT 30.670 148.710 34.220 148.850 ;
        RECT 30.670 148.665 30.960 148.710 ;
        RECT 31.640 148.650 31.960 148.710 ;
        RECT 33.930 148.665 34.220 148.710 ;
        RECT 34.850 148.850 35.140 148.895 ;
        RECT 36.710 148.850 37.000 148.895 ;
        RECT 34.850 148.710 37.000 148.850 ;
        RECT 34.850 148.665 35.140 148.710 ;
        RECT 36.710 148.665 37.000 148.710 ;
        RECT 39.920 148.850 40.240 148.910 ;
        RECT 49.595 148.850 49.885 148.895 ;
        RECT 52.355 148.850 52.645 148.895 ;
        RECT 61.080 148.850 61.400 148.910 ;
        RECT 39.920 148.710 47.510 148.850 ;
        RECT 32.530 148.510 32.820 148.555 ;
        RECT 34.850 148.510 35.065 148.665 ;
        RECT 39.920 148.650 40.240 148.710 ;
        RECT 47.370 148.555 47.510 148.710 ;
        RECT 49.595 148.710 52.645 148.850 ;
        RECT 49.595 148.665 49.885 148.710 ;
        RECT 52.355 148.665 52.645 148.710 ;
        RECT 54.730 148.710 61.400 148.850 ;
        RECT 32.530 148.370 35.065 148.510 ;
        RECT 32.530 148.325 32.820 148.370 ;
        RECT 46.835 148.325 47.125 148.555 ;
        RECT 47.295 148.325 47.585 148.555 ;
        RECT 50.975 148.510 51.265 148.555 ;
        RECT 51.420 148.510 51.740 148.570 ;
        RECT 50.975 148.370 51.740 148.510 ;
        RECT 50.975 148.325 51.265 148.370 ;
        RECT 29.340 148.170 29.660 148.230 ;
        RECT 35.795 148.170 36.085 148.215 ;
        RECT 29.340 148.030 36.085 148.170 ;
        RECT 29.340 147.970 29.660 148.030 ;
        RECT 35.795 147.985 36.085 148.030 ;
        RECT 36.240 148.170 36.560 148.230 ;
        RECT 37.620 148.170 37.940 148.230 ;
        RECT 46.910 148.170 47.050 148.325 ;
        RECT 51.420 148.310 51.740 148.370 ;
        RECT 53.720 148.310 54.040 148.570 ;
        RECT 54.730 148.555 54.870 148.710 ;
        RECT 61.080 148.650 61.400 148.710 ;
        RECT 62.090 148.850 62.230 149.050 ;
        RECT 65.680 148.990 66.000 149.250 ;
        RECT 77.180 149.190 77.500 149.250 ;
        RECT 81.780 149.190 82.100 149.250 ;
        RECT 66.230 149.050 77.500 149.190 ;
        RECT 66.230 148.850 66.370 149.050 ;
        RECT 77.180 148.990 77.500 149.050 ;
        RECT 80.950 149.050 82.100 149.190 ;
        RECT 62.090 148.710 66.370 148.850 ;
        RECT 66.600 148.850 66.920 148.910 ;
        RECT 68.915 148.850 69.205 148.895 ;
        RECT 69.820 148.850 70.140 148.910 ;
        RECT 70.295 148.850 70.585 148.895 ;
        RECT 66.600 148.710 70.585 148.850 ;
        RECT 54.195 148.325 54.485 148.555 ;
        RECT 54.655 148.325 54.945 148.555 ;
        RECT 49.580 148.170 49.900 148.230 ;
        RECT 36.240 148.030 40.610 148.170 ;
        RECT 46.910 148.030 49.900 148.170 ;
        RECT 36.240 147.970 36.560 148.030 ;
        RECT 37.620 147.970 37.940 148.030 ;
        RECT 32.530 147.830 32.820 147.875 ;
        RECT 35.310 147.830 35.600 147.875 ;
        RECT 37.170 147.830 37.460 147.875 ;
        RECT 32.530 147.690 37.460 147.830 ;
        RECT 32.530 147.645 32.820 147.690 ;
        RECT 35.310 147.645 35.600 147.690 ;
        RECT 37.170 147.645 37.460 147.690 ;
        RECT 40.470 147.550 40.610 148.030 ;
        RECT 49.580 147.970 49.900 148.030 ;
        RECT 50.515 148.170 50.805 148.215 ;
        RECT 51.880 148.170 52.200 148.230 ;
        RECT 50.515 148.030 52.200 148.170 ;
        RECT 50.515 147.985 50.805 148.030 ;
        RECT 51.880 147.970 52.200 148.030 ;
        RECT 53.260 148.170 53.580 148.230 ;
        RECT 54.270 148.170 54.410 148.325 ;
        RECT 55.560 148.310 55.880 148.570 ;
        RECT 57.400 148.310 57.720 148.570 ;
        RECT 57.860 148.310 58.180 148.570 ;
        RECT 58.335 148.325 58.625 148.555 ;
        RECT 59.240 148.510 59.560 148.570 ;
        RECT 59.240 148.370 60.390 148.510 ;
        RECT 53.260 148.030 54.410 148.170 ;
        RECT 53.260 147.970 53.580 148.030 ;
        RECT 45.440 147.830 45.760 147.890 ;
        RECT 58.410 147.830 58.550 148.325 ;
        RECT 59.240 148.310 59.560 148.370 ;
        RECT 59.240 147.830 59.560 147.890 ;
        RECT 45.440 147.690 55.330 147.830 ;
        RECT 58.410 147.690 59.560 147.830 ;
        RECT 60.250 147.830 60.390 148.370 ;
        RECT 61.540 148.310 61.860 148.570 ;
        RECT 62.090 148.555 62.230 148.710 ;
        RECT 66.600 148.650 66.920 148.710 ;
        RECT 68.915 148.665 69.205 148.710 ;
        RECT 69.820 148.650 70.140 148.710 ;
        RECT 70.295 148.665 70.585 148.710 ;
        RECT 70.740 148.850 71.060 148.910 ;
        RECT 73.500 148.850 73.820 148.910 ;
        RECT 70.740 148.710 73.820 148.850 ;
        RECT 70.740 148.650 71.060 148.710 ;
        RECT 73.500 148.650 73.820 148.710 ;
        RECT 73.975 148.850 74.265 148.895 ;
        RECT 75.355 148.850 75.645 148.895 ;
        RECT 80.950 148.850 81.090 149.050 ;
        RECT 81.780 148.990 82.100 149.050 ;
        RECT 87.760 149.190 88.080 149.250 ;
        RECT 101.345 149.190 101.635 149.235 ;
        RECT 102.480 149.190 102.800 149.250 ;
        RECT 87.760 149.050 99.030 149.190 ;
        RECT 87.760 148.990 88.080 149.050 ;
        RECT 73.975 148.710 75.645 148.850 ;
        RECT 73.975 148.665 74.265 148.710 ;
        RECT 75.355 148.665 75.645 148.710 ;
        RECT 76.350 148.710 81.090 148.850 ;
        RECT 81.270 148.850 81.560 148.895 ;
        RECT 83.620 148.850 83.940 148.910 ;
        RECT 84.530 148.850 84.820 148.895 ;
        RECT 81.270 148.710 84.820 148.850 ;
        RECT 62.015 148.325 62.305 148.555 ;
        RECT 62.460 148.310 62.780 148.570 ;
        RECT 63.380 148.310 63.700 148.570 ;
        RECT 71.200 148.510 71.520 148.570 ;
        RECT 72.595 148.510 72.885 148.555 ;
        RECT 63.930 148.370 70.740 148.510 ;
        RECT 61.630 148.170 61.770 148.310 ;
        RECT 63.930 148.170 64.070 148.370 ;
        RECT 61.630 148.030 64.070 148.170 ;
        RECT 64.760 147.970 65.080 148.230 ;
        RECT 65.235 148.170 65.525 148.215 ;
        RECT 66.140 148.170 66.460 148.230 ;
        RECT 65.235 148.030 66.460 148.170 ;
        RECT 70.600 148.170 70.740 148.370 ;
        RECT 71.200 148.370 72.885 148.510 ;
        RECT 71.200 148.310 71.520 148.370 ;
        RECT 72.595 148.325 72.885 148.370 ;
        RECT 73.055 148.510 73.345 148.555 ;
        RECT 76.350 148.510 76.490 148.710 ;
        RECT 81.270 148.665 81.560 148.710 ;
        RECT 83.620 148.650 83.940 148.710 ;
        RECT 84.530 148.665 84.820 148.710 ;
        RECT 85.450 148.850 85.740 148.895 ;
        RECT 87.310 148.850 87.600 148.895 ;
        RECT 85.450 148.710 87.600 148.850 ;
        RECT 85.450 148.665 85.740 148.710 ;
        RECT 87.310 148.665 87.600 148.710 ;
        RECT 90.930 148.850 91.220 148.895 ;
        RECT 92.360 148.850 92.680 148.910 ;
        RECT 94.190 148.850 94.480 148.895 ;
        RECT 90.930 148.710 94.480 148.850 ;
        RECT 90.930 148.665 91.220 148.710 ;
        RECT 73.055 148.370 76.490 148.510 ;
        RECT 73.055 148.325 73.345 148.370 ;
        RECT 76.720 148.310 77.040 148.570 ;
        RECT 77.180 148.310 77.500 148.570 ;
        RECT 77.640 148.310 77.960 148.570 ;
        RECT 78.575 148.510 78.865 148.555 ;
        RECT 79.940 148.510 80.260 148.570 ;
        RECT 78.575 148.370 80.260 148.510 ;
        RECT 78.575 148.325 78.865 148.370 ;
        RECT 79.940 148.310 80.260 148.370 ;
        RECT 83.130 148.510 83.420 148.555 ;
        RECT 85.450 148.510 85.665 148.665 ;
        RECT 92.360 148.650 92.680 148.710 ;
        RECT 94.190 148.665 94.480 148.710 ;
        RECT 95.110 148.850 95.400 148.895 ;
        RECT 96.970 148.850 97.260 148.895 ;
        RECT 95.110 148.710 97.260 148.850 ;
        RECT 95.110 148.665 95.400 148.710 ;
        RECT 96.970 148.665 97.260 148.710 ;
        RECT 83.130 148.370 85.665 148.510 ;
        RECT 85.920 148.510 86.240 148.570 ;
        RECT 86.395 148.510 86.685 148.555 ;
        RECT 85.920 148.370 86.685 148.510 ;
        RECT 83.130 148.325 83.420 148.370 ;
        RECT 85.920 148.310 86.240 148.370 ;
        RECT 86.395 148.325 86.685 148.370 ;
        RECT 92.790 148.510 93.080 148.555 ;
        RECT 95.110 148.510 95.325 148.665 ;
        RECT 92.790 148.370 95.325 148.510 ;
        RECT 92.790 148.325 93.080 148.370 ;
        RECT 96.040 148.310 96.360 148.570 ;
        RECT 98.355 148.325 98.645 148.555 ;
        RECT 76.810 148.170 76.950 148.310 ;
        RECT 70.600 148.030 76.950 148.170 ;
        RECT 77.270 148.170 77.410 148.310 ;
        RECT 80.400 148.170 80.720 148.230 ;
        RECT 77.270 148.030 80.720 148.170 ;
        RECT 65.235 147.985 65.525 148.030 ;
        RECT 66.140 147.970 66.460 148.030 ;
        RECT 80.400 147.970 80.720 148.030 ;
        RECT 87.300 148.170 87.620 148.230 ;
        RECT 88.235 148.170 88.525 148.215 ;
        RECT 96.960 148.170 97.280 148.230 ;
        RECT 97.895 148.170 98.185 148.215 ;
        RECT 87.300 148.030 98.185 148.170 ;
        RECT 87.300 147.970 87.620 148.030 ;
        RECT 88.235 147.985 88.525 148.030 ;
        RECT 96.960 147.970 97.280 148.030 ;
        RECT 97.895 147.985 98.185 148.030 ;
        RECT 63.380 147.830 63.700 147.890 ;
        RECT 60.250 147.690 63.700 147.830 ;
        RECT 45.440 147.630 45.760 147.690 ;
        RECT 28.665 147.490 28.955 147.535 ;
        RECT 29.800 147.490 30.120 147.550 ;
        RECT 33.940 147.490 34.260 147.550 ;
        RECT 28.665 147.350 34.260 147.490 ;
        RECT 28.665 147.305 28.955 147.350 ;
        RECT 29.800 147.290 30.120 147.350 ;
        RECT 33.940 147.290 34.260 147.350 ;
        RECT 40.380 147.290 40.700 147.550 ;
        RECT 46.820 147.490 47.140 147.550 ;
        RECT 48.215 147.490 48.505 147.535 ;
        RECT 46.820 147.350 48.505 147.490 ;
        RECT 46.820 147.290 47.140 147.350 ;
        RECT 48.215 147.305 48.505 147.350 ;
        RECT 50.500 147.290 50.820 147.550 ;
        RECT 51.880 147.290 52.200 147.550 ;
        RECT 55.190 147.490 55.330 147.690 ;
        RECT 59.240 147.630 59.560 147.690 ;
        RECT 63.380 147.630 63.700 147.690 ;
        RECT 67.535 147.830 67.825 147.875 ;
        RECT 74.420 147.830 74.740 147.890 ;
        RECT 67.535 147.690 74.740 147.830 ;
        RECT 67.535 147.645 67.825 147.690 ;
        RECT 74.420 147.630 74.740 147.690 ;
        RECT 83.130 147.830 83.420 147.875 ;
        RECT 85.910 147.830 86.200 147.875 ;
        RECT 87.770 147.830 88.060 147.875 ;
        RECT 83.130 147.690 88.060 147.830 ;
        RECT 83.130 147.645 83.420 147.690 ;
        RECT 85.910 147.645 86.200 147.690 ;
        RECT 87.770 147.645 88.060 147.690 ;
        RECT 92.790 147.830 93.080 147.875 ;
        RECT 95.570 147.830 95.860 147.875 ;
        RECT 97.430 147.830 97.720 147.875 ;
        RECT 92.790 147.690 97.720 147.830 ;
        RECT 92.790 147.645 93.080 147.690 ;
        RECT 95.570 147.645 95.860 147.690 ;
        RECT 97.430 147.645 97.720 147.690 ;
        RECT 98.430 147.830 98.570 148.325 ;
        RECT 98.890 148.170 99.030 149.050 ;
        RECT 101.345 149.050 102.800 149.190 ;
        RECT 101.345 149.005 101.635 149.050 ;
        RECT 102.480 148.990 102.800 149.050 ;
        RECT 106.160 149.190 106.480 149.250 ;
        RECT 111.235 149.190 111.525 149.235 ;
        RECT 106.160 149.050 111.525 149.190 ;
        RECT 106.160 148.990 106.480 149.050 ;
        RECT 111.235 149.005 111.525 149.050 ;
        RECT 103.350 148.850 103.640 148.895 ;
        RECT 104.780 148.850 105.100 148.910 ;
        RECT 106.610 148.850 106.900 148.895 ;
        RECT 103.350 148.710 106.900 148.850 ;
        RECT 103.350 148.665 103.640 148.710 ;
        RECT 104.780 148.650 105.100 148.710 ;
        RECT 106.610 148.665 106.900 148.710 ;
        RECT 107.530 148.850 107.820 148.895 ;
        RECT 109.390 148.850 109.680 148.895 ;
        RECT 107.530 148.710 109.680 148.850 ;
        RECT 107.530 148.665 107.820 148.710 ;
        RECT 109.390 148.665 109.680 148.710 ;
        RECT 105.210 148.510 105.500 148.555 ;
        RECT 107.530 148.510 107.745 148.665 ;
        RECT 105.210 148.370 107.745 148.510 ;
        RECT 105.210 148.325 105.500 148.370 ;
        RECT 108.460 148.310 108.780 148.570 ;
        RECT 110.760 148.310 111.080 148.570 ;
        RECT 109.380 148.170 109.700 148.230 ;
        RECT 98.890 148.030 109.700 148.170 ;
        RECT 109.380 147.970 109.700 148.030 ;
        RECT 110.300 147.970 110.620 148.230 ;
        RECT 102.940 147.830 103.260 147.890 ;
        RECT 98.430 147.690 103.260 147.830 ;
        RECT 56.035 147.490 56.325 147.535 ;
        RECT 55.190 147.350 56.325 147.490 ;
        RECT 56.035 147.305 56.325 147.350 ;
        RECT 56.940 147.490 57.260 147.550 ;
        RECT 68.455 147.490 68.745 147.535 ;
        RECT 70.280 147.490 70.600 147.550 ;
        RECT 56.940 147.350 70.600 147.490 ;
        RECT 56.940 147.290 57.260 147.350 ;
        RECT 68.455 147.305 68.745 147.350 ;
        RECT 70.280 147.290 70.600 147.350 ;
        RECT 70.740 147.290 71.060 147.550 ;
        RECT 71.675 147.490 71.965 147.535 ;
        RECT 73.040 147.490 73.360 147.550 ;
        RECT 71.675 147.350 73.360 147.490 ;
        RECT 71.675 147.305 71.965 147.350 ;
        RECT 73.040 147.290 73.360 147.350 ;
        RECT 73.975 147.490 74.265 147.535 ;
        RECT 75.800 147.490 76.120 147.550 ;
        RECT 73.975 147.350 76.120 147.490 ;
        RECT 73.975 147.305 74.265 147.350 ;
        RECT 75.800 147.290 76.120 147.350 ;
        RECT 77.640 147.490 77.960 147.550 ;
        RECT 79.265 147.490 79.555 147.535 ;
        RECT 82.240 147.490 82.560 147.550 ;
        RECT 77.640 147.350 82.560 147.490 ;
        RECT 77.640 147.290 77.960 147.350 ;
        RECT 79.265 147.305 79.555 147.350 ;
        RECT 82.240 147.290 82.560 147.350 ;
        RECT 86.380 147.490 86.700 147.550 ;
        RECT 88.925 147.490 89.215 147.535 ;
        RECT 86.380 147.350 89.215 147.490 ;
        RECT 86.380 147.290 86.700 147.350 ;
        RECT 88.925 147.305 89.215 147.350 ;
        RECT 90.980 147.490 91.300 147.550 ;
        RECT 98.430 147.490 98.570 147.690 ;
        RECT 102.940 147.630 103.260 147.690 ;
        RECT 105.210 147.830 105.500 147.875 ;
        RECT 107.990 147.830 108.280 147.875 ;
        RECT 109.850 147.830 110.140 147.875 ;
        RECT 105.210 147.690 110.140 147.830 ;
        RECT 105.210 147.645 105.500 147.690 ;
        RECT 107.990 147.645 108.280 147.690 ;
        RECT 109.850 147.645 110.140 147.690 ;
        RECT 90.980 147.350 98.570 147.490 ;
        RECT 90.980 147.290 91.300 147.350 ;
        RECT 98.800 147.290 99.120 147.550 ;
        RECT 26.970 146.670 113.450 147.150 ;
        RECT 31.180 146.270 31.500 146.530 ;
        RECT 34.860 146.270 35.180 146.530 ;
        RECT 39.920 146.270 40.240 146.530 ;
        RECT 70.740 146.470 71.060 146.530 ;
        RECT 40.470 146.330 71.060 146.470 ;
        RECT 34.950 146.130 35.090 146.270 ;
        RECT 40.470 146.130 40.610 146.330 ;
        RECT 70.740 146.270 71.060 146.330 ;
        RECT 74.420 146.470 74.740 146.530 ;
        RECT 74.895 146.470 75.185 146.515 ;
        RECT 74.420 146.330 75.185 146.470 ;
        RECT 74.420 146.270 74.740 146.330 ;
        RECT 74.895 146.285 75.185 146.330 ;
        RECT 84.555 146.470 84.845 146.515 ;
        RECT 85.000 146.470 85.320 146.530 ;
        RECT 84.555 146.330 85.320 146.470 ;
        RECT 84.555 146.285 84.845 146.330 ;
        RECT 85.000 146.270 85.320 146.330 ;
        RECT 92.360 146.270 92.680 146.530 ;
        RECT 97.420 146.270 97.740 146.530 ;
        RECT 104.780 146.270 105.100 146.530 ;
        RECT 108.475 146.470 108.765 146.515 ;
        RECT 105.790 146.330 108.765 146.470 ;
        RECT 34.950 145.990 40.610 146.130 ;
        RECT 44.490 146.130 44.780 146.175 ;
        RECT 47.270 146.130 47.560 146.175 ;
        RECT 49.130 146.130 49.420 146.175 ;
        RECT 44.490 145.990 49.420 146.130 ;
        RECT 44.490 145.945 44.780 145.990 ;
        RECT 47.270 145.945 47.560 145.990 ;
        RECT 49.130 145.945 49.420 145.990 ;
        RECT 63.380 146.130 63.700 146.190 ;
        RECT 79.940 146.130 80.260 146.190 ;
        RECT 84.080 146.130 84.400 146.190 ;
        RECT 63.380 145.990 80.260 146.130 ;
        RECT 63.380 145.930 63.700 145.990 ;
        RECT 79.940 145.930 80.260 145.990 ;
        RECT 81.870 145.990 84.400 146.130 ;
        RECT 28.880 145.790 29.200 145.850 ;
        RECT 28.880 145.650 30.490 145.790 ;
        RECT 28.880 145.590 29.200 145.650 ;
        RECT 30.350 145.495 30.490 145.650 ;
        RECT 33.940 145.590 34.260 145.850 ;
        RECT 34.860 145.790 35.180 145.850 ;
        RECT 36.715 145.790 37.005 145.835 ;
        RECT 37.160 145.790 37.480 145.850 ;
        RECT 34.860 145.650 37.480 145.790 ;
        RECT 34.860 145.590 35.180 145.650 ;
        RECT 36.715 145.605 37.005 145.650 ;
        RECT 37.160 145.590 37.480 145.650 ;
        RECT 46.820 145.790 47.140 145.850 ;
        RECT 47.755 145.790 48.045 145.835 ;
        RECT 46.820 145.650 48.045 145.790 ;
        RECT 46.820 145.590 47.140 145.650 ;
        RECT 47.755 145.605 48.045 145.650 ;
        RECT 50.500 145.590 50.820 145.850 ;
        RECT 53.260 145.790 53.580 145.850 ;
        RECT 57.860 145.790 58.180 145.850 ;
        RECT 63.470 145.790 63.610 145.930 ;
        RECT 53.260 145.650 59.930 145.790 ;
        RECT 53.260 145.590 53.580 145.650 ;
        RECT 29.815 145.265 30.105 145.495 ;
        RECT 30.275 145.450 30.565 145.495 ;
        RECT 31.640 145.450 31.960 145.510 ;
        RECT 30.275 145.310 31.960 145.450 ;
        RECT 30.275 145.265 30.565 145.310 ;
        RECT 29.890 145.110 30.030 145.265 ;
        RECT 31.640 145.250 31.960 145.310 ;
        RECT 32.100 145.450 32.420 145.510 ;
        RECT 33.495 145.450 33.785 145.495 ;
        RECT 32.100 145.310 33.785 145.450 ;
        RECT 32.100 145.250 32.420 145.310 ;
        RECT 33.495 145.265 33.785 145.310 ;
        RECT 44.490 145.450 44.780 145.495 ;
        RECT 44.490 145.310 47.025 145.450 ;
        RECT 44.490 145.265 44.780 145.310 ;
        RECT 38.095 145.110 38.385 145.155 ;
        RECT 39.000 145.110 39.320 145.170 ;
        RECT 42.680 145.155 43.000 145.170 ;
        RECT 46.810 145.155 47.025 145.310 ;
        RECT 49.595 145.265 49.885 145.495 ;
        RECT 54.195 145.450 54.485 145.495 ;
        RECT 54.640 145.450 54.960 145.510 ;
        RECT 55.650 145.495 55.790 145.650 ;
        RECT 57.860 145.590 58.180 145.650 ;
        RECT 54.195 145.310 54.960 145.450 ;
        RECT 54.195 145.265 54.485 145.310 ;
        RECT 40.625 145.110 40.915 145.155 ;
        RECT 29.890 144.970 40.915 145.110 ;
        RECT 38.095 144.925 38.385 144.970 ;
        RECT 39.000 144.910 39.320 144.970 ;
        RECT 40.625 144.925 40.915 144.970 ;
        RECT 42.630 145.110 43.000 145.155 ;
        RECT 45.890 145.110 46.180 145.155 ;
        RECT 42.630 144.970 46.180 145.110 ;
        RECT 42.630 144.925 43.000 144.970 ;
        RECT 45.890 144.925 46.180 144.970 ;
        RECT 46.810 145.110 47.100 145.155 ;
        RECT 48.670 145.110 48.960 145.155 ;
        RECT 46.810 144.970 48.960 145.110 ;
        RECT 49.670 145.110 49.810 145.265 ;
        RECT 54.640 145.250 54.960 145.310 ;
        RECT 55.115 145.265 55.405 145.495 ;
        RECT 55.575 145.265 55.865 145.495 ;
        RECT 56.035 145.450 56.325 145.495 ;
        RECT 57.400 145.450 57.720 145.510 ;
        RECT 59.790 145.495 59.930 145.650 ;
        RECT 61.170 145.650 63.610 145.790 ;
        RECT 65.220 145.790 65.540 145.850 ;
        RECT 65.220 145.650 67.290 145.790 ;
        RECT 61.170 145.495 61.310 145.650 ;
        RECT 65.220 145.590 65.540 145.650 ;
        RECT 59.255 145.450 59.545 145.495 ;
        RECT 56.035 145.310 59.545 145.450 ;
        RECT 56.035 145.265 56.325 145.310 ;
        RECT 50.040 145.110 50.360 145.170 ;
        RECT 49.670 144.970 50.360 145.110 ;
        RECT 46.810 144.925 47.100 144.970 ;
        RECT 48.670 144.925 48.960 144.970 ;
        RECT 42.680 144.910 43.000 144.925 ;
        RECT 50.040 144.910 50.360 144.970 ;
        RECT 51.435 145.110 51.725 145.155 ;
        RECT 53.260 145.110 53.580 145.170 ;
        RECT 51.435 144.970 53.580 145.110 ;
        RECT 51.435 144.925 51.725 144.970 ;
        RECT 53.260 144.910 53.580 144.970 ;
        RECT 28.880 144.770 29.200 144.830 ;
        RECT 31.655 144.770 31.945 144.815 ;
        RECT 28.880 144.630 31.945 144.770 ;
        RECT 28.880 144.570 29.200 144.630 ;
        RECT 31.655 144.585 31.945 144.630 ;
        RECT 37.620 144.770 37.940 144.830 ;
        RECT 44.060 144.770 44.380 144.830 ;
        RECT 51.895 144.770 52.185 144.815 ;
        RECT 37.620 144.630 52.185 144.770 ;
        RECT 37.620 144.570 37.940 144.630 ;
        RECT 44.060 144.570 44.380 144.630 ;
        RECT 51.895 144.585 52.185 144.630 ;
        RECT 53.720 144.570 54.040 144.830 ;
        RECT 55.190 144.770 55.330 145.265 ;
        RECT 57.400 145.250 57.720 145.310 ;
        RECT 59.255 145.265 59.545 145.310 ;
        RECT 59.715 145.265 60.005 145.495 ;
        RECT 60.175 145.265 60.465 145.495 ;
        RECT 61.095 145.265 61.385 145.495 ;
        RECT 62.935 145.450 63.225 145.495 ;
        RECT 66.600 145.450 66.920 145.510 ;
        RECT 62.935 145.310 66.920 145.450 ;
        RECT 62.935 145.265 63.225 145.310 ;
        RECT 60.250 145.110 60.390 145.265 ;
        RECT 66.600 145.250 66.920 145.310 ;
        RECT 66.140 145.110 66.460 145.170 ;
        RECT 60.250 144.970 66.460 145.110 ;
        RECT 66.140 144.910 66.460 144.970 ;
        RECT 67.150 144.830 67.290 145.650 ;
        RECT 75.340 145.590 75.660 145.850 ;
        RECT 76.720 145.790 77.040 145.850 ;
        RECT 80.400 145.790 80.720 145.850 ;
        RECT 81.870 145.835 82.010 145.990 ;
        RECT 84.080 145.930 84.400 145.990 ;
        RECT 85.460 146.130 85.780 146.190 ;
        RECT 91.440 146.130 91.760 146.190 ;
        RECT 99.260 146.130 99.580 146.190 ;
        RECT 103.860 146.130 104.180 146.190 ;
        RECT 105.790 146.130 105.930 146.330 ;
        RECT 108.475 146.285 108.765 146.330 ;
        RECT 85.460 145.990 88.450 146.130 ;
        RECT 85.460 145.930 85.780 145.990 ;
        RECT 76.720 145.650 78.330 145.790 ;
        RECT 76.720 145.590 77.040 145.650 ;
        RECT 69.360 145.250 69.680 145.510 ;
        RECT 69.820 145.250 70.140 145.510 ;
        RECT 73.515 145.265 73.805 145.495 ;
        RECT 70.740 145.110 71.060 145.170 ;
        RECT 71.675 145.110 71.965 145.155 ;
        RECT 70.740 144.970 71.965 145.110 ;
        RECT 73.590 145.110 73.730 145.265 ;
        RECT 74.880 145.250 75.200 145.510 ;
        RECT 77.640 145.450 77.960 145.510 ;
        RECT 78.190 145.495 78.330 145.650 ;
        RECT 78.650 145.650 80.720 145.790 ;
        RECT 78.650 145.495 78.790 145.650 ;
        RECT 80.400 145.590 80.720 145.650 ;
        RECT 81.795 145.605 82.085 145.835 ;
        RECT 82.240 145.590 82.560 145.850 ;
        RECT 86.380 145.790 86.700 145.850 ;
        RECT 88.310 145.835 88.450 145.990 ;
        RECT 91.440 145.990 94.430 146.130 ;
        RECT 91.440 145.930 91.760 145.990 ;
        RECT 82.790 145.650 86.700 145.790 ;
        RECT 75.890 145.310 77.960 145.450 ;
        RECT 75.340 145.110 75.660 145.170 ;
        RECT 75.890 145.110 76.030 145.310 ;
        RECT 77.640 145.250 77.960 145.310 ;
        RECT 78.115 145.265 78.405 145.495 ;
        RECT 78.575 145.265 78.865 145.495 ;
        RECT 79.035 145.265 79.325 145.495 ;
        RECT 73.590 144.970 76.030 145.110 ;
        RECT 76.275 145.110 76.565 145.155 ;
        RECT 76.735 145.110 77.025 145.155 ;
        RECT 76.275 144.970 77.025 145.110 ;
        RECT 79.110 145.110 79.250 145.265 ;
        RECT 79.940 145.250 80.260 145.510 ;
        RECT 82.790 145.495 82.930 145.650 ;
        RECT 86.380 145.590 86.700 145.650 ;
        RECT 88.235 145.605 88.525 145.835 ;
        RECT 89.600 145.790 89.920 145.850 ;
        RECT 93.295 145.790 93.585 145.835 ;
        RECT 89.600 145.650 93.585 145.790 ;
        RECT 89.600 145.590 89.920 145.650 ;
        RECT 93.295 145.605 93.585 145.650 ;
        RECT 94.290 145.790 94.430 145.990 ;
        RECT 96.590 145.990 101.790 146.130 ;
        RECT 96.590 145.790 96.730 145.990 ;
        RECT 99.260 145.930 99.580 145.990 ;
        RECT 94.290 145.650 96.730 145.790 ;
        RECT 82.715 145.450 83.005 145.495 ;
        RECT 80.490 145.310 83.005 145.450 ;
        RECT 80.490 145.110 80.630 145.310 ;
        RECT 82.715 145.265 83.005 145.310 ;
        RECT 85.015 145.265 85.305 145.495 ;
        RECT 91.440 145.435 91.760 145.510 ;
        RECT 94.290 145.495 94.430 145.650 ;
        RECT 91.915 145.435 92.205 145.495 ;
        RECT 91.440 145.295 92.205 145.435 ;
        RECT 79.110 144.970 80.630 145.110 ;
        RECT 81.780 145.110 82.100 145.170 ;
        RECT 85.090 145.110 85.230 145.265 ;
        RECT 91.440 145.250 91.760 145.295 ;
        RECT 91.915 145.265 92.205 145.295 ;
        RECT 94.215 145.265 94.505 145.495 ;
        RECT 95.135 145.265 95.425 145.495 ;
        RECT 89.155 145.110 89.445 145.155 ;
        RECT 95.210 145.110 95.350 145.265 ;
        RECT 95.580 145.250 95.900 145.510 ;
        RECT 96.590 145.495 96.730 145.650 ;
        RECT 98.340 145.590 98.660 145.850 ;
        RECT 100.195 145.790 100.485 145.835 ;
        RECT 100.640 145.790 100.960 145.850 ;
        RECT 100.195 145.650 100.960 145.790 ;
        RECT 100.195 145.605 100.485 145.650 ;
        RECT 100.640 145.590 100.960 145.650 ;
        RECT 96.515 145.265 96.805 145.495 ;
        RECT 99.260 145.250 99.580 145.510 ;
        RECT 101.650 145.495 101.790 145.990 ;
        RECT 103.860 145.990 105.930 146.130 ;
        RECT 103.860 145.930 104.180 145.990 ;
        RECT 106.620 145.930 106.940 146.190 ;
        RECT 108.920 146.130 109.240 146.190 ;
        RECT 110.760 146.130 111.080 146.190 ;
        RECT 108.920 145.990 111.080 146.130 ;
        RECT 108.920 145.930 109.240 145.990 ;
        RECT 110.760 145.930 111.080 145.990 ;
        RECT 106.710 145.790 106.850 145.930 ;
        RECT 106.710 145.650 109.610 145.790 ;
        RECT 101.575 145.265 101.865 145.495 ;
        RECT 102.020 145.250 102.340 145.510 ;
        RECT 102.940 145.450 103.260 145.510 ;
        RECT 104.320 145.450 104.640 145.510 ;
        RECT 102.940 145.310 104.640 145.450 ;
        RECT 102.940 145.250 103.260 145.310 ;
        RECT 104.320 145.250 104.640 145.310 ;
        RECT 106.635 145.265 106.925 145.495 ;
        RECT 81.780 144.970 85.230 145.110 ;
        RECT 85.550 144.970 89.445 145.110 ;
        RECT 70.740 144.910 71.060 144.970 ;
        RECT 71.675 144.925 71.965 144.970 ;
        RECT 75.340 144.910 75.660 144.970 ;
        RECT 76.275 144.925 76.565 144.970 ;
        RECT 76.735 144.925 77.025 144.970 ;
        RECT 81.780 144.910 82.100 144.970 ;
        RECT 56.940 144.770 57.260 144.830 ;
        RECT 55.190 144.630 57.260 144.770 ;
        RECT 56.940 144.570 57.260 144.630 ;
        RECT 57.400 144.570 57.720 144.830 ;
        RECT 57.860 144.570 58.180 144.830 ;
        RECT 63.395 144.770 63.685 144.815 ;
        RECT 65.220 144.770 65.540 144.830 ;
        RECT 63.395 144.630 65.540 144.770 ;
        RECT 63.395 144.585 63.685 144.630 ;
        RECT 65.220 144.570 65.540 144.630 ;
        RECT 65.680 144.570 66.000 144.830 ;
        RECT 67.060 144.570 67.380 144.830 ;
        RECT 67.995 144.770 68.285 144.815 ;
        RECT 73.500 144.770 73.820 144.830 ;
        RECT 67.995 144.630 73.820 144.770 ;
        RECT 67.995 144.585 68.285 144.630 ;
        RECT 73.500 144.570 73.820 144.630 ;
        RECT 73.975 144.770 74.265 144.815 ;
        RECT 77.640 144.770 77.960 144.830 ;
        RECT 73.975 144.630 77.960 144.770 ;
        RECT 73.975 144.585 74.265 144.630 ;
        RECT 77.640 144.570 77.960 144.630 ;
        RECT 79.940 144.770 80.260 144.830 ;
        RECT 85.550 144.770 85.690 144.970 ;
        RECT 89.155 144.925 89.445 144.970 ;
        RECT 89.690 144.970 95.350 145.110 ;
        RECT 99.720 145.110 100.040 145.170 ;
        RECT 106.710 145.110 106.850 145.265 ;
        RECT 108.920 145.250 109.240 145.510 ;
        RECT 109.470 145.495 109.610 145.650 ;
        RECT 109.395 145.265 109.685 145.495 ;
        RECT 111.680 145.250 112.000 145.510 ;
        RECT 99.720 144.970 106.850 145.110 ;
        RECT 107.170 144.970 110.530 145.110 ;
        RECT 89.690 144.830 89.830 144.970 ;
        RECT 99.720 144.910 100.040 144.970 ;
        RECT 79.940 144.630 85.690 144.770 ;
        RECT 79.940 144.570 80.260 144.630 ;
        RECT 85.920 144.570 86.240 144.830 ;
        RECT 89.600 144.570 89.920 144.830 ;
        RECT 91.455 144.770 91.745 144.815 ;
        RECT 97.420 144.770 97.740 144.830 ;
        RECT 91.455 144.630 97.740 144.770 ;
        RECT 91.455 144.585 91.745 144.630 ;
        RECT 97.420 144.570 97.740 144.630 ;
        RECT 100.655 144.770 100.945 144.815 ;
        RECT 101.560 144.770 101.880 144.830 ;
        RECT 100.655 144.630 101.880 144.770 ;
        RECT 100.655 144.585 100.945 144.630 ;
        RECT 101.560 144.570 101.880 144.630 ;
        RECT 103.400 144.570 103.720 144.830 ;
        RECT 105.700 144.770 106.020 144.830 ;
        RECT 107.170 144.770 107.310 144.970 ;
        RECT 105.700 144.630 107.310 144.770 ;
        RECT 107.555 144.770 107.845 144.815 ;
        RECT 109.380 144.770 109.700 144.830 ;
        RECT 110.390 144.815 110.530 144.970 ;
        RECT 107.555 144.630 109.700 144.770 ;
        RECT 105.700 144.570 106.020 144.630 ;
        RECT 107.555 144.585 107.845 144.630 ;
        RECT 109.380 144.570 109.700 144.630 ;
        RECT 110.315 144.585 110.605 144.815 ;
        RECT 110.760 144.570 111.080 144.830 ;
        RECT 26.970 143.950 113.450 144.430 ;
        RECT 29.585 143.750 29.875 143.795 ;
        RECT 32.100 143.750 32.420 143.810 ;
        RECT 29.585 143.610 32.420 143.750 ;
        RECT 29.585 143.565 29.875 143.610 ;
        RECT 32.100 143.550 32.420 143.610 ;
        RECT 36.240 143.750 36.560 143.810 ;
        RECT 51.420 143.750 51.740 143.810 ;
        RECT 58.795 143.750 59.085 143.795 ;
        RECT 59.240 143.750 59.560 143.810 ;
        RECT 36.240 143.610 47.970 143.750 ;
        RECT 36.240 143.550 36.560 143.610 ;
        RECT 31.590 143.410 31.880 143.455 ;
        RECT 34.850 143.410 35.140 143.455 ;
        RECT 31.590 143.270 35.140 143.410 ;
        RECT 31.590 143.225 31.880 143.270 ;
        RECT 34.850 143.225 35.140 143.270 ;
        RECT 35.770 143.410 36.060 143.455 ;
        RECT 37.630 143.410 37.920 143.455 ;
        RECT 35.770 143.270 37.920 143.410 ;
        RECT 35.770 143.225 36.060 143.270 ;
        RECT 37.630 143.225 37.920 143.270 ;
        RECT 41.250 143.410 41.540 143.455 ;
        RECT 44.510 143.410 44.800 143.455 ;
        RECT 41.250 143.270 44.800 143.410 ;
        RECT 41.250 143.225 41.540 143.270 ;
        RECT 44.510 143.225 44.800 143.270 ;
        RECT 45.430 143.410 45.720 143.455 ;
        RECT 47.290 143.410 47.580 143.455 ;
        RECT 45.430 143.270 47.580 143.410 ;
        RECT 45.430 143.225 45.720 143.270 ;
        RECT 47.290 143.225 47.580 143.270 ;
        RECT 29.800 143.070 30.120 143.130 ;
        RECT 31.730 143.070 31.870 143.225 ;
        RECT 29.800 142.930 31.870 143.070 ;
        RECT 33.450 143.070 33.740 143.115 ;
        RECT 35.770 143.070 35.985 143.225 ;
        RECT 41.390 143.070 41.530 143.225 ;
        RECT 33.450 142.930 35.985 143.070 ;
        RECT 36.330 142.930 41.530 143.070 ;
        RECT 43.110 143.070 43.400 143.115 ;
        RECT 45.430 143.070 45.645 143.225 ;
        RECT 43.110 142.930 45.645 143.070 ;
        RECT 46.375 143.070 46.665 143.115 ;
        RECT 47.830 143.070 47.970 143.610 ;
        RECT 51.420 143.610 59.560 143.750 ;
        RECT 51.420 143.550 51.740 143.610 ;
        RECT 58.795 143.565 59.085 143.610 ;
        RECT 59.240 143.550 59.560 143.610 ;
        RECT 62.000 143.750 62.320 143.810 ;
        RECT 63.165 143.750 63.455 143.795 ;
        RECT 65.680 143.750 66.000 143.810 ;
        RECT 62.000 143.610 66.000 143.750 ;
        RECT 62.000 143.550 62.320 143.610 ;
        RECT 63.165 143.565 63.455 143.610 ;
        RECT 65.680 143.550 66.000 143.610 ;
        RECT 72.595 143.565 72.885 143.795 ;
        RECT 53.720 143.410 54.040 143.470 ;
        RECT 56.940 143.410 57.260 143.470 ;
        RECT 63.840 143.410 64.160 143.470 ;
        RECT 65.220 143.455 65.540 143.470 ;
        RECT 53.720 143.270 56.710 143.410 ;
        RECT 53.720 143.210 54.040 143.270 ;
        RECT 46.375 142.930 47.970 143.070 ;
        RECT 50.040 143.070 50.360 143.130 ;
        RECT 54.655 143.070 54.945 143.115 ;
        RECT 56.020 143.070 56.340 143.130 ;
        RECT 56.570 143.115 56.710 143.270 ;
        RECT 56.940 143.270 64.160 143.410 ;
        RECT 56.940 143.210 57.260 143.270 ;
        RECT 63.840 143.210 64.160 143.270 ;
        RECT 65.170 143.410 65.540 143.455 ;
        RECT 68.430 143.410 68.720 143.455 ;
        RECT 65.170 143.270 68.720 143.410 ;
        RECT 65.170 143.225 65.540 143.270 ;
        RECT 68.430 143.225 68.720 143.270 ;
        RECT 69.350 143.410 69.640 143.455 ;
        RECT 71.210 143.410 71.500 143.455 ;
        RECT 69.350 143.270 71.500 143.410 ;
        RECT 69.350 143.225 69.640 143.270 ;
        RECT 71.210 143.225 71.500 143.270 ;
        RECT 65.220 143.210 65.540 143.225 ;
        RECT 50.040 142.930 56.340 143.070 ;
        RECT 29.800 142.870 30.120 142.930 ;
        RECT 33.450 142.885 33.740 142.930 ;
        RECT 27.500 142.730 27.820 142.790 ;
        RECT 36.330 142.730 36.470 142.930 ;
        RECT 43.110 142.885 43.400 142.930 ;
        RECT 46.375 142.885 46.665 142.930 ;
        RECT 50.040 142.870 50.360 142.930 ;
        RECT 54.655 142.885 54.945 142.930 ;
        RECT 56.020 142.870 56.340 142.930 ;
        RECT 56.495 142.885 56.785 143.115 ;
        RECT 59.255 143.070 59.545 143.115 ;
        RECT 61.080 143.070 61.400 143.130 ;
        RECT 59.255 142.930 61.400 143.070 ;
        RECT 59.255 142.885 59.545 142.930 ;
        RECT 61.080 142.870 61.400 142.930 ;
        RECT 67.030 143.070 67.320 143.115 ;
        RECT 69.350 143.070 69.565 143.225 ;
        RECT 67.030 142.930 69.565 143.070 ;
        RECT 70.295 143.070 70.585 143.115 ;
        RECT 72.670 143.070 72.810 143.565 ;
        RECT 79.940 143.550 80.260 143.810 ;
        RECT 81.780 143.550 82.100 143.810 ;
        RECT 86.855 143.750 87.145 143.795 ;
        RECT 87.300 143.750 87.620 143.810 ;
        RECT 86.855 143.610 87.620 143.750 ;
        RECT 86.855 143.565 87.145 143.610 ;
        RECT 87.300 143.550 87.620 143.610 ;
        RECT 94.675 143.750 94.965 143.795 ;
        RECT 96.040 143.750 96.360 143.810 ;
        RECT 94.675 143.610 96.360 143.750 ;
        RECT 94.675 143.565 94.965 143.610 ;
        RECT 96.040 143.550 96.360 143.610 ;
        RECT 99.720 143.550 100.040 143.810 ;
        RECT 75.340 143.410 75.660 143.470 ;
        RECT 79.495 143.410 79.785 143.455 ;
        RECT 89.600 143.410 89.920 143.470 ;
        RECT 97.435 143.410 97.725 143.455 ;
        RECT 100.640 143.410 100.960 143.470 ;
        RECT 102.265 143.410 102.555 143.455 ;
        RECT 75.340 143.270 83.850 143.410 ;
        RECT 75.340 143.210 75.660 143.270 ;
        RECT 79.495 143.225 79.785 143.270 ;
        RECT 70.295 142.930 72.810 143.070 ;
        RECT 67.030 142.885 67.320 142.930 ;
        RECT 70.295 142.885 70.585 142.930 ;
        RECT 73.500 142.870 73.820 143.130 ;
        RECT 76.720 143.070 77.040 143.130 ;
        RECT 77.195 143.070 77.485 143.115 ;
        RECT 82.240 143.070 82.560 143.130 ;
        RECT 83.710 143.115 83.850 143.270 ;
        RECT 89.600 143.270 97.725 143.410 ;
        RECT 89.600 143.210 89.920 143.270 ;
        RECT 97.435 143.225 97.725 143.270 ;
        RECT 99.350 143.270 102.555 143.410 ;
        RECT 99.350 143.130 99.490 143.270 ;
        RECT 100.640 143.210 100.960 143.270 ;
        RECT 102.265 143.225 102.555 143.270 ;
        RECT 103.400 143.410 103.720 143.470 ;
        RECT 104.270 143.410 104.560 143.455 ;
        RECT 107.530 143.410 107.820 143.455 ;
        RECT 103.400 143.270 107.820 143.410 ;
        RECT 103.400 143.210 103.720 143.270 ;
        RECT 104.270 143.225 104.560 143.270 ;
        RECT 107.530 143.225 107.820 143.270 ;
        RECT 108.450 143.410 108.740 143.455 ;
        RECT 110.310 143.410 110.600 143.455 ;
        RECT 108.450 143.270 110.600 143.410 ;
        RECT 108.450 143.225 108.740 143.270 ;
        RECT 110.310 143.225 110.600 143.270 ;
        RECT 83.175 143.070 83.465 143.115 ;
        RECT 76.720 142.930 79.250 143.070 ;
        RECT 76.720 142.870 77.040 142.930 ;
        RECT 77.195 142.885 77.485 142.930 ;
        RECT 27.500 142.590 36.470 142.730 ;
        RECT 27.500 142.530 27.820 142.590 ;
        RECT 36.700 142.530 37.020 142.790 ;
        RECT 38.555 142.730 38.845 142.775 ;
        RECT 40.380 142.730 40.700 142.790 ;
        RECT 48.215 142.730 48.505 142.775 ;
        RECT 38.555 142.590 48.505 142.730 ;
        RECT 38.555 142.545 38.845 142.590 ;
        RECT 40.380 142.530 40.700 142.590 ;
        RECT 48.215 142.545 48.505 142.590 ;
        RECT 58.335 142.730 58.625 142.775 ;
        RECT 64.300 142.730 64.620 142.790 ;
        RECT 58.335 142.590 64.620 142.730 ;
        RECT 58.335 142.545 58.625 142.590 ;
        RECT 64.300 142.530 64.620 142.590 ;
        RECT 72.120 142.730 72.440 142.790 ;
        RECT 76.810 142.730 76.950 142.870 ;
        RECT 72.120 142.590 76.950 142.730 ;
        RECT 78.100 142.730 78.420 142.790 ;
        RECT 78.575 142.730 78.865 142.775 ;
        RECT 78.100 142.590 78.865 142.730 ;
        RECT 79.110 142.730 79.250 142.930 ;
        RECT 82.240 142.930 83.465 143.070 ;
        RECT 82.240 142.870 82.560 142.930 ;
        RECT 83.175 142.885 83.465 142.930 ;
        RECT 83.635 142.885 83.925 143.115 ;
        RECT 93.280 142.870 93.600 143.130 ;
        RECT 93.755 143.070 94.045 143.115 ;
        RECT 94.660 143.070 94.980 143.130 ;
        RECT 93.755 142.930 94.980 143.070 ;
        RECT 93.755 142.885 94.045 142.930 ;
        RECT 94.660 142.870 94.980 142.930 ;
        RECT 97.895 143.070 98.185 143.115 ;
        RECT 99.260 143.070 99.580 143.130 ;
        RECT 97.895 142.930 99.580 143.070 ;
        RECT 97.895 142.885 98.185 142.930 ;
        RECT 99.260 142.870 99.580 142.930 ;
        RECT 101.575 142.885 101.865 143.115 ;
        RECT 106.130 143.070 106.420 143.115 ;
        RECT 108.450 143.070 108.665 143.225 ;
        RECT 106.130 142.930 108.665 143.070 ;
        RECT 106.130 142.885 106.420 142.930 ;
        RECT 86.840 142.730 87.160 142.790 ;
        RECT 79.110 142.590 87.160 142.730 ;
        RECT 72.120 142.530 72.440 142.590 ;
        RECT 78.100 142.530 78.420 142.590 ;
        RECT 78.575 142.545 78.865 142.590 ;
        RECT 86.840 142.530 87.160 142.590 ;
        RECT 96.040 142.730 96.360 142.790 ;
        RECT 96.515 142.730 96.805 142.775 ;
        RECT 96.040 142.590 96.805 142.730 ;
        RECT 96.040 142.530 96.360 142.590 ;
        RECT 96.515 142.545 96.805 142.590 ;
        RECT 97.420 142.730 97.740 142.790 ;
        RECT 101.650 142.730 101.790 142.885 ;
        RECT 109.380 142.870 109.700 143.130 ;
        RECT 97.420 142.590 101.790 142.730 ;
        RECT 110.300 142.730 110.620 142.790 ;
        RECT 111.235 142.730 111.525 142.775 ;
        RECT 110.300 142.590 111.525 142.730 ;
        RECT 97.420 142.530 97.740 142.590 ;
        RECT 110.300 142.530 110.620 142.590 ;
        RECT 111.235 142.545 111.525 142.590 ;
        RECT 33.450 142.390 33.740 142.435 ;
        RECT 36.230 142.390 36.520 142.435 ;
        RECT 38.090 142.390 38.380 142.435 ;
        RECT 33.450 142.250 38.380 142.390 ;
        RECT 33.450 142.205 33.740 142.250 ;
        RECT 36.230 142.205 36.520 142.250 ;
        RECT 38.090 142.205 38.380 142.250 ;
        RECT 43.110 142.390 43.400 142.435 ;
        RECT 45.890 142.390 46.180 142.435 ;
        RECT 47.750 142.390 48.040 142.435 ;
        RECT 43.110 142.250 48.040 142.390 ;
        RECT 43.110 142.205 43.400 142.250 ;
        RECT 45.890 142.205 46.180 142.250 ;
        RECT 47.750 142.205 48.040 142.250 ;
        RECT 67.030 142.390 67.320 142.435 ;
        RECT 69.810 142.390 70.100 142.435 ;
        RECT 71.670 142.390 71.960 142.435 ;
        RECT 67.030 142.250 71.960 142.390 ;
        RECT 67.030 142.205 67.320 142.250 ;
        RECT 69.810 142.205 70.100 142.250 ;
        RECT 71.670 142.205 71.960 142.250 ;
        RECT 73.960 142.390 74.280 142.450 ;
        RECT 82.255 142.390 82.545 142.435 ;
        RECT 73.960 142.250 82.545 142.390 ;
        RECT 73.960 142.190 74.280 142.250 ;
        RECT 82.255 142.205 82.545 142.250 ;
        RECT 89.140 142.390 89.460 142.450 ;
        RECT 101.560 142.390 101.880 142.450 ;
        RECT 89.140 142.250 101.880 142.390 ;
        RECT 89.140 142.190 89.460 142.250 ;
        RECT 101.560 142.190 101.880 142.250 ;
        RECT 106.130 142.390 106.420 142.435 ;
        RECT 108.910 142.390 109.200 142.435 ;
        RECT 110.770 142.390 111.060 142.435 ;
        RECT 106.130 142.250 111.060 142.390 ;
        RECT 106.130 142.205 106.420 142.250 ;
        RECT 108.910 142.205 109.200 142.250 ;
        RECT 110.770 142.205 111.060 142.250 ;
        RECT 30.260 142.050 30.580 142.110 ;
        RECT 31.180 142.050 31.500 142.110 ;
        RECT 33.020 142.050 33.340 142.110 ;
        RECT 39.245 142.050 39.535 142.095 ;
        RECT 30.260 141.910 39.535 142.050 ;
        RECT 30.260 141.850 30.580 141.910 ;
        RECT 31.180 141.850 31.500 141.910 ;
        RECT 33.020 141.850 33.340 141.910 ;
        RECT 39.245 141.865 39.535 141.910 ;
        RECT 43.600 142.050 43.920 142.110 ;
        RECT 44.520 142.050 44.840 142.110 ;
        RECT 43.600 141.910 44.840 142.050 ;
        RECT 43.600 141.850 43.920 141.910 ;
        RECT 44.520 141.850 44.840 141.910 ;
        RECT 46.820 142.050 47.140 142.110 ;
        RECT 55.575 142.050 55.865 142.095 ;
        RECT 46.820 141.910 55.865 142.050 ;
        RECT 46.820 141.850 47.140 141.910 ;
        RECT 55.575 141.865 55.865 141.910 ;
        RECT 59.240 142.050 59.560 142.110 ;
        RECT 61.095 142.050 61.385 142.095 ;
        RECT 59.240 141.910 61.385 142.050 ;
        RECT 59.240 141.850 59.560 141.910 ;
        RECT 61.095 141.865 61.385 141.910 ;
        RECT 77.640 142.050 77.960 142.110 ;
        RECT 83.620 142.050 83.940 142.110 ;
        RECT 77.640 141.910 83.940 142.050 ;
        RECT 77.640 141.850 77.960 141.910 ;
        RECT 83.620 141.850 83.940 141.910 ;
        RECT 95.120 142.050 95.440 142.110 ;
        RECT 100.655 142.050 100.945 142.095 ;
        RECT 95.120 141.910 100.945 142.050 ;
        RECT 95.120 141.850 95.440 141.910 ;
        RECT 100.655 141.865 100.945 141.910 ;
        RECT 26.970 141.230 113.450 141.710 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 37.620 141.030 37.940 141.090 ;
        RECT 39.705 141.030 39.995 141.075 ;
        RECT 29.430 140.890 35.550 141.030 ;
        RECT 29.430 140.395 29.570 140.890 ;
        RECT 32.560 140.690 32.880 140.750 ;
        RECT 34.860 140.690 35.180 140.750 ;
        RECT 32.560 140.550 35.180 140.690 ;
        RECT 32.560 140.490 32.880 140.550 ;
        RECT 29.355 140.165 29.645 140.395 ;
        RECT 32.100 140.350 32.420 140.410 ;
        RECT 34.490 140.395 34.630 140.550 ;
        RECT 34.860 140.490 35.180 140.550 ;
        RECT 33.955 140.350 34.245 140.395 ;
        RECT 32.100 140.210 34.245 140.350 ;
        RECT 32.100 140.150 32.420 140.210 ;
        RECT 33.955 140.165 34.245 140.210 ;
        RECT 34.415 140.165 34.705 140.395 ;
        RECT 35.410 140.350 35.550 140.890 ;
        RECT 37.620 140.890 39.995 141.030 ;
        RECT 37.620 140.830 37.940 140.890 ;
        RECT 39.705 140.845 39.995 140.890 ;
        RECT 42.220 141.030 42.540 141.090 ;
        RECT 42.220 140.890 49.810 141.030 ;
        RECT 42.220 140.830 42.540 140.890 ;
        RECT 37.160 140.690 37.480 140.750 ;
        RECT 38.540 140.690 38.860 140.750 ;
        RECT 37.160 140.550 38.860 140.690 ;
        RECT 37.160 140.490 37.480 140.550 ;
        RECT 38.540 140.490 38.860 140.550 ;
        RECT 43.570 140.690 43.860 140.735 ;
        RECT 46.350 140.690 46.640 140.735 ;
        RECT 48.210 140.690 48.500 140.735 ;
        RECT 43.570 140.550 48.500 140.690 ;
        RECT 49.670 140.690 49.810 140.890 ;
        RECT 56.480 140.830 56.800 141.090 ;
        RECT 59.700 140.830 60.020 141.090 ;
        RECT 70.740 141.030 71.060 141.090 ;
        RECT 60.250 140.890 71.060 141.030 ;
        RECT 60.250 140.690 60.390 140.890 ;
        RECT 70.740 140.830 71.060 140.890 ;
        RECT 74.880 141.030 75.200 141.090 ;
        RECT 84.080 141.030 84.400 141.090 ;
        RECT 74.880 140.890 84.400 141.030 ;
        RECT 74.880 140.830 75.200 140.890 ;
        RECT 84.080 140.830 84.400 140.890 ;
        RECT 88.005 141.030 88.295 141.075 ;
        RECT 89.600 141.030 89.920 141.090 ;
        RECT 88.005 140.890 89.920 141.030 ;
        RECT 88.005 140.845 88.295 140.890 ;
        RECT 89.600 140.830 89.920 140.890 ;
        RECT 49.670 140.550 60.390 140.690 ;
        RECT 60.635 140.690 60.925 140.735 ;
        RECT 66.600 140.690 66.920 140.750 ;
        RECT 60.635 140.550 66.920 140.690 ;
        RECT 43.570 140.505 43.860 140.550 ;
        RECT 46.350 140.505 46.640 140.550 ;
        RECT 48.210 140.505 48.500 140.550 ;
        RECT 60.635 140.505 60.925 140.550 ;
        RECT 66.600 140.490 66.920 140.550 ;
        RECT 81.750 140.690 82.040 140.735 ;
        RECT 84.530 140.690 84.820 140.735 ;
        RECT 86.390 140.690 86.680 140.735 ;
        RECT 81.750 140.550 86.680 140.690 ;
        RECT 81.750 140.505 82.040 140.550 ;
        RECT 84.530 140.505 84.820 140.550 ;
        RECT 86.390 140.505 86.680 140.550 ;
        RECT 91.870 140.690 92.160 140.735 ;
        RECT 94.650 140.690 94.940 140.735 ;
        RECT 96.510 140.690 96.800 140.735 ;
        RECT 91.870 140.550 96.800 140.690 ;
        RECT 91.870 140.505 92.160 140.550 ;
        RECT 94.650 140.505 94.940 140.550 ;
        RECT 96.510 140.505 96.800 140.550 ;
        RECT 106.130 140.690 106.420 140.735 ;
        RECT 108.910 140.690 109.200 140.735 ;
        RECT 110.770 140.690 111.060 140.735 ;
        RECT 106.130 140.550 111.060 140.690 ;
        RECT 106.130 140.505 106.420 140.550 ;
        RECT 108.910 140.505 109.200 140.550 ;
        RECT 110.770 140.505 111.060 140.550 ;
        RECT 42.220 140.350 42.540 140.410 ;
        RECT 35.410 140.210 42.540 140.350 ;
        RECT 42.220 140.150 42.540 140.210 ;
        RECT 46.820 140.150 47.140 140.410 ;
        RECT 48.675 140.350 48.965 140.395 ;
        RECT 50.040 140.350 50.360 140.410 ;
        RECT 48.675 140.210 50.360 140.350 ;
        RECT 48.675 140.165 48.965 140.210 ;
        RECT 50.040 140.150 50.360 140.210 ;
        RECT 54.180 140.350 54.500 140.410 ;
        RECT 58.795 140.350 59.085 140.395 ;
        RECT 54.180 140.210 59.085 140.350 ;
        RECT 54.180 140.150 54.500 140.210 ;
        RECT 58.795 140.165 59.085 140.210 ;
        RECT 64.300 140.350 64.620 140.410 ;
        RECT 67.060 140.350 67.380 140.410 ;
        RECT 64.300 140.210 67.380 140.350 ;
        RECT 64.300 140.150 64.620 140.210 ;
        RECT 67.060 140.150 67.380 140.210 ;
        RECT 76.720 140.150 77.040 140.410 ;
        RECT 77.885 140.350 78.175 140.395 ;
        RECT 79.940 140.350 80.260 140.410 ;
        RECT 82.700 140.350 83.020 140.410 ;
        RECT 77.885 140.210 83.020 140.350 ;
        RECT 77.885 140.165 78.175 140.210 ;
        RECT 79.940 140.150 80.260 140.210 ;
        RECT 82.700 140.150 83.020 140.210 ;
        RECT 85.015 140.350 85.305 140.395 ;
        RECT 85.920 140.350 86.240 140.410 ;
        RECT 85.015 140.210 86.240 140.350 ;
        RECT 85.015 140.165 85.305 140.210 ;
        RECT 85.920 140.150 86.240 140.210 ;
        RECT 86.840 140.150 87.160 140.410 ;
        RECT 95.120 140.150 95.440 140.410 ;
        RECT 96.040 140.150 96.360 140.410 ;
        RECT 96.960 140.150 97.280 140.410 ;
        RECT 98.355 140.165 98.645 140.395 ;
        RECT 30.275 140.010 30.565 140.055 ;
        RECT 31.640 140.010 31.960 140.070 ;
        RECT 30.275 139.870 31.960 140.010 ;
        RECT 30.275 139.825 30.565 139.870 ;
        RECT 31.640 139.810 31.960 139.870 ;
        RECT 33.020 140.010 33.340 140.070 ;
        RECT 33.495 140.010 33.785 140.055 ;
        RECT 33.020 139.870 33.785 140.010 ;
        RECT 33.020 139.810 33.340 139.870 ;
        RECT 33.495 139.825 33.785 139.870 ;
        RECT 39.015 140.010 39.305 140.055 ;
        RECT 40.380 140.010 40.700 140.070 ;
        RECT 39.015 139.870 40.700 140.010 ;
        RECT 39.015 139.825 39.305 139.870 ;
        RECT 40.380 139.810 40.700 139.870 ;
        RECT 43.570 140.010 43.860 140.055 ;
        RECT 43.570 139.870 46.105 140.010 ;
        RECT 43.570 139.825 43.860 139.870 ;
        RECT 31.195 139.670 31.485 139.715 ;
        RECT 41.710 139.670 42.000 139.715 ;
        RECT 43.140 139.670 43.460 139.730 ;
        RECT 45.890 139.715 46.105 139.870 ;
        RECT 49.120 139.810 49.440 140.070 ;
        RECT 57.860 140.010 58.180 140.070 ;
        RECT 58.335 140.010 58.625 140.055 ;
        RECT 57.860 139.870 58.625 140.010 ;
        RECT 57.860 139.810 58.180 139.870 ;
        RECT 58.335 139.825 58.625 139.870 ;
        RECT 59.715 140.010 60.005 140.055 ;
        RECT 60.620 140.010 60.940 140.070 ;
        RECT 59.715 139.870 60.940 140.010 ;
        RECT 59.715 139.825 60.005 139.870 ;
        RECT 60.620 139.810 60.940 139.870 ;
        RECT 62.015 139.825 62.305 140.055 ;
        RECT 65.235 140.010 65.525 140.055 ;
        RECT 65.680 140.010 66.000 140.070 ;
        RECT 65.235 139.870 66.000 140.010 ;
        RECT 65.235 139.825 65.525 139.870 ;
        RECT 44.970 139.670 45.260 139.715 ;
        RECT 31.195 139.530 41.530 139.670 ;
        RECT 31.195 139.485 31.485 139.530 ;
        RECT 30.260 139.330 30.580 139.390 ;
        RECT 31.655 139.330 31.945 139.375 ;
        RECT 30.260 139.190 31.945 139.330 ;
        RECT 41.390 139.330 41.530 139.530 ;
        RECT 41.710 139.530 45.260 139.670 ;
        RECT 41.710 139.485 42.000 139.530 ;
        RECT 43.140 139.470 43.460 139.530 ;
        RECT 44.970 139.485 45.260 139.530 ;
        RECT 45.890 139.670 46.180 139.715 ;
        RECT 47.750 139.670 48.040 139.715 ;
        RECT 45.890 139.530 48.040 139.670 ;
        RECT 62.090 139.670 62.230 139.825 ;
        RECT 65.680 139.810 66.000 139.870 ;
        RECT 68.440 139.810 68.760 140.070 ;
        RECT 81.750 140.010 82.040 140.055 ;
        RECT 91.870 140.010 92.160 140.055 ;
        RECT 96.130 140.010 96.270 140.150 ;
        RECT 98.430 140.010 98.570 140.165 ;
        RECT 99.260 140.150 99.580 140.410 ;
        RECT 110.300 140.350 110.620 140.410 ;
        RECT 111.235 140.350 111.525 140.395 ;
        RECT 110.300 140.210 111.525 140.350 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 110.300 140.150 110.620 140.210 ;
        RECT 111.235 140.165 111.525 140.210 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 81.750 139.870 84.285 140.010 ;
        RECT 81.750 139.825 82.040 139.870 ;
        RECT 83.160 139.715 83.480 139.730 ;
        RECT 79.890 139.670 80.180 139.715 ;
        RECT 83.150 139.670 83.480 139.715 ;
        RECT 62.090 139.530 65.910 139.670 ;
        RECT 45.890 139.485 46.180 139.530 ;
        RECT 47.750 139.485 48.040 139.530 ;
        RECT 65.770 139.390 65.910 139.530 ;
        RECT 79.890 139.530 83.480 139.670 ;
        RECT 79.890 139.485 80.180 139.530 ;
        RECT 83.150 139.485 83.480 139.530 ;
        RECT 84.070 139.715 84.285 139.870 ;
        RECT 91.870 139.870 94.405 140.010 ;
        RECT 96.130 139.870 98.570 140.010 ;
        RECT 106.130 140.010 106.420 140.055 ;
        RECT 106.130 139.870 108.665 140.010 ;
        RECT 91.870 139.825 92.160 139.870 ;
        RECT 84.070 139.670 84.360 139.715 ;
        RECT 85.930 139.670 86.220 139.715 ;
        RECT 84.070 139.530 86.220 139.670 ;
        RECT 84.070 139.485 84.360 139.530 ;
        RECT 85.930 139.485 86.220 139.530 ;
        RECT 90.010 139.670 90.300 139.715 ;
        RECT 90.980 139.670 91.300 139.730 ;
        RECT 94.190 139.715 94.405 139.870 ;
        RECT 106.130 139.825 106.420 139.870 ;
        RECT 102.020 139.715 102.340 139.730 ;
        RECT 93.270 139.670 93.560 139.715 ;
        RECT 90.010 139.530 93.560 139.670 ;
        RECT 90.010 139.485 90.300 139.530 ;
        RECT 83.160 139.470 83.480 139.485 ;
        RECT 90.980 139.470 91.300 139.530 ;
        RECT 93.270 139.485 93.560 139.530 ;
        RECT 94.190 139.670 94.480 139.715 ;
        RECT 96.050 139.670 96.340 139.715 ;
        RECT 102.020 139.670 102.555 139.715 ;
        RECT 94.190 139.530 96.340 139.670 ;
        RECT 94.190 139.485 94.480 139.530 ;
        RECT 96.050 139.485 96.340 139.530 ;
        RECT 99.810 139.530 102.555 139.670 ;
        RECT 49.580 139.330 49.900 139.390 ;
        RECT 41.390 139.190 49.900 139.330 ;
        RECT 30.260 139.130 30.580 139.190 ;
        RECT 31.655 139.145 31.945 139.190 ;
        RECT 49.580 139.130 49.900 139.190 ;
        RECT 62.000 139.330 62.320 139.390 ;
        RECT 62.475 139.330 62.765 139.375 ;
        RECT 62.000 139.190 62.765 139.330 ;
        RECT 62.000 139.130 62.320 139.190 ;
        RECT 62.475 139.145 62.765 139.190 ;
        RECT 63.840 139.330 64.160 139.390 ;
        RECT 64.760 139.330 65.080 139.390 ;
        RECT 63.840 139.190 65.080 139.330 ;
        RECT 63.840 139.130 64.160 139.190 ;
        RECT 64.760 139.130 65.080 139.190 ;
        RECT 65.680 139.130 66.000 139.390 ;
        RECT 67.075 139.330 67.365 139.375 ;
        RECT 73.960 139.330 74.280 139.390 ;
        RECT 67.075 139.190 74.280 139.330 ;
        RECT 67.075 139.145 67.365 139.190 ;
        RECT 73.960 139.130 74.280 139.190 ;
        RECT 99.260 139.330 99.580 139.390 ;
        RECT 99.810 139.375 99.950 139.530 ;
        RECT 102.020 139.485 102.555 139.530 ;
        RECT 104.270 139.670 104.560 139.715 ;
        RECT 105.700 139.670 106.020 139.730 ;
        RECT 108.450 139.715 108.665 139.870 ;
        RECT 109.380 139.810 109.700 140.070 ;
        RECT 107.530 139.670 107.820 139.715 ;
        RECT 104.270 139.530 107.820 139.670 ;
        RECT 104.270 139.485 104.560 139.530 ;
        RECT 102.020 139.470 102.340 139.485 ;
        RECT 105.700 139.470 106.020 139.530 ;
        RECT 107.530 139.485 107.820 139.530 ;
        RECT 108.450 139.670 108.740 139.715 ;
        RECT 110.310 139.670 110.600 139.715 ;
        RECT 108.450 139.530 110.600 139.670 ;
        RECT 108.450 139.485 108.740 139.530 ;
        RECT 110.310 139.485 110.600 139.530 ;
        RECT 99.735 139.330 100.025 139.375 ;
        RECT 99.260 139.190 100.025 139.330 ;
        RECT 99.260 139.130 99.580 139.190 ;
        RECT 99.735 139.145 100.025 139.190 ;
        RECT 101.560 139.130 101.880 139.390 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 26.970 138.510 113.450 138.990 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 37.620 138.310 37.940 138.370 ;
        RECT 43.600 138.310 43.920 138.370 ;
        RECT 61.080 138.355 61.400 138.370 ;
        RECT 37.620 138.170 42.450 138.310 ;
        RECT 37.620 138.110 37.940 138.170 ;
        RECT 31.295 137.970 31.585 138.015 ;
        RECT 34.535 137.970 35.185 138.015 ;
        RECT 31.295 137.830 35.185 137.970 ;
        RECT 31.295 137.785 31.885 137.830 ;
        RECT 34.535 137.785 35.185 137.830 ;
        RECT 35.780 137.970 36.100 138.030 ;
        RECT 37.175 137.970 37.465 138.015 ;
        RECT 35.780 137.830 37.465 137.970 ;
        RECT 31.595 137.690 31.885 137.785 ;
        RECT 35.780 137.770 36.100 137.830 ;
        RECT 37.175 137.785 37.465 137.830 ;
        RECT 39.940 137.970 40.230 138.015 ;
        RECT 41.800 137.970 42.090 138.015 ;
        RECT 39.940 137.830 42.090 137.970 ;
        RECT 42.310 137.970 42.450 138.170 ;
        RECT 43.600 138.170 46.590 138.310 ;
        RECT 43.600 138.110 43.920 138.170 ;
        RECT 42.720 137.970 43.010 138.015 ;
        RECT 45.980 137.970 46.270 138.015 ;
        RECT 42.310 137.830 46.270 137.970 ;
        RECT 46.450 137.970 46.590 138.170 ;
        RECT 49.670 138.170 52.570 138.310 ;
        RECT 49.670 137.970 49.810 138.170 ;
        RECT 46.450 137.830 49.810 137.970 ;
        RECT 50.060 137.970 50.350 138.015 ;
        RECT 51.920 137.970 52.210 138.015 ;
        RECT 50.060 137.830 52.210 137.970 ;
        RECT 52.430 137.970 52.570 138.170 ;
        RECT 60.865 138.125 61.400 138.355 ;
        RECT 72.595 138.310 72.885 138.355 ;
        RECT 74.420 138.310 74.740 138.370 ;
        RECT 72.595 138.170 74.740 138.310 ;
        RECT 72.595 138.125 72.885 138.170 ;
        RECT 61.080 138.110 61.400 138.125 ;
        RECT 74.420 138.110 74.740 138.170 ;
        RECT 75.430 138.170 81.090 138.310 ;
        RECT 52.840 137.970 53.130 138.015 ;
        RECT 56.100 137.970 56.390 138.015 ;
        RECT 52.430 137.830 56.390 137.970 ;
        RECT 39.940 137.785 40.230 137.830 ;
        RECT 41.800 137.785 42.090 137.830 ;
        RECT 42.720 137.785 43.010 137.830 ;
        RECT 45.980 137.785 46.270 137.830 ;
        RECT 50.060 137.785 50.350 137.830 ;
        RECT 51.920 137.785 52.210 137.830 ;
        RECT 52.840 137.785 53.130 137.830 ;
        RECT 56.100 137.785 56.390 137.830 ;
        RECT 62.870 137.970 63.160 138.015 ;
        RECT 65.220 137.970 65.540 138.030 ;
        RECT 66.130 137.970 66.420 138.015 ;
        RECT 62.870 137.830 66.420 137.970 ;
        RECT 62.870 137.785 63.160 137.830 ;
        RECT 31.595 137.470 31.960 137.690 ;
        RECT 31.640 137.430 31.960 137.470 ;
        RECT 32.675 137.630 32.965 137.675 ;
        RECT 36.255 137.630 36.545 137.675 ;
        RECT 38.090 137.630 38.380 137.675 ;
        RECT 32.675 137.490 38.380 137.630 ;
        RECT 41.875 137.630 42.090 137.785 ;
        RECT 44.120 137.630 44.410 137.675 ;
        RECT 41.875 137.490 44.410 137.630 ;
        RECT 51.995 137.630 52.210 137.785 ;
        RECT 65.220 137.770 65.540 137.830 ;
        RECT 66.130 137.785 66.420 137.830 ;
        RECT 67.050 137.970 67.340 138.015 ;
        RECT 68.910 137.970 69.200 138.015 ;
        RECT 75.430 137.970 75.570 138.170 ;
        RECT 67.050 137.830 69.200 137.970 ;
        RECT 67.050 137.785 67.340 137.830 ;
        RECT 68.910 137.785 69.200 137.830 ;
        RECT 71.290 137.830 75.570 137.970 ;
        RECT 75.800 137.970 76.120 138.030 ;
        RECT 79.035 137.970 79.325 138.015 ;
        RECT 75.800 137.830 79.325 137.970 ;
        RECT 80.950 137.970 81.090 138.170 ;
        RECT 81.320 138.110 81.640 138.370 ;
        RECT 83.160 138.110 83.480 138.370 ;
        RECT 85.935 138.310 86.225 138.355 ;
        RECT 88.680 138.310 89.000 138.370 ;
        RECT 93.755 138.310 94.045 138.355 ;
        RECT 85.935 138.170 94.045 138.310 ;
        RECT 85.935 138.125 86.225 138.170 ;
        RECT 88.680 138.110 89.000 138.170 ;
        RECT 93.755 138.125 94.045 138.170 ;
        RECT 97.435 138.310 97.725 138.355 ;
        RECT 98.340 138.310 98.660 138.370 ;
        RECT 100.180 138.310 100.500 138.370 ;
        RECT 100.885 138.310 101.175 138.355 ;
        RECT 97.435 138.170 101.175 138.310 ;
        RECT 97.435 138.125 97.725 138.170 ;
        RECT 98.340 138.110 98.660 138.170 ;
        RECT 100.180 138.110 100.500 138.170 ;
        RECT 100.885 138.125 101.175 138.170 ;
        RECT 109.380 138.310 109.700 138.370 ;
        RECT 110.315 138.310 110.605 138.355 ;
        RECT 109.380 138.170 110.605 138.310 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 109.380 138.110 109.700 138.170 ;
        RECT 110.315 138.125 110.605 138.170 ;
        RECT 83.250 137.970 83.390 138.110 ;
        RECT 89.155 137.970 89.445 138.015 ;
        RECT 80.950 137.830 82.930 137.970 ;
        RECT 83.250 137.830 89.445 137.970 ;
        RECT 54.240 137.630 54.530 137.675 ;
        RECT 51.995 137.490 54.530 137.630 ;
        RECT 32.675 137.445 32.965 137.490 ;
        RECT 36.255 137.445 36.545 137.490 ;
        RECT 38.090 137.445 38.380 137.490 ;
        RECT 44.120 137.445 44.410 137.490 ;
        RECT 54.240 137.445 54.530 137.490 ;
        RECT 59.240 137.430 59.560 137.690 ;
        RECT 64.730 137.630 65.020 137.675 ;
        RECT 67.050 137.630 67.265 137.785 ;
        RECT 71.290 137.675 71.430 137.830 ;
        RECT 75.800 137.770 76.120 137.830 ;
        RECT 79.035 137.785 79.325 137.830 ;
        RECT 64.730 137.490 67.265 137.630 ;
        RECT 64.730 137.445 65.020 137.490 ;
        RECT 71.215 137.445 71.505 137.675 ;
        RECT 71.675 137.630 71.965 137.675 ;
        RECT 71.675 137.490 72.810 137.630 ;
        RECT 71.675 137.445 71.965 137.490 ;
        RECT 26.580 137.290 26.900 137.350 ;
        RECT 28.435 137.290 28.725 137.335 ;
        RECT 26.580 137.150 28.725 137.290 ;
        RECT 26.580 137.090 26.900 137.150 ;
        RECT 28.435 137.105 28.725 137.150 ;
        RECT 38.555 137.290 38.845 137.335 ;
        RECT 39.015 137.290 39.305 137.335 ;
        RECT 40.380 137.290 40.700 137.350 ;
        RECT 38.555 137.150 40.700 137.290 ;
        RECT 38.555 137.105 38.845 137.150 ;
        RECT 39.015 137.105 39.305 137.150 ;
        RECT 40.380 137.090 40.700 137.150 ;
        RECT 40.840 137.090 41.160 137.350 ;
        RECT 49.135 137.290 49.425 137.335 ;
        RECT 50.040 137.290 50.360 137.350 ;
        RECT 49.135 137.150 50.360 137.290 ;
        RECT 49.135 137.105 49.425 137.150 ;
        RECT 50.040 137.090 50.360 137.150 ;
        RECT 50.960 137.090 51.280 137.350 ;
        RECT 67.980 137.090 68.300 137.350 ;
        RECT 69.835 137.290 70.125 137.335 ;
        RECT 72.120 137.290 72.440 137.350 ;
        RECT 69.835 137.150 72.440 137.290 ;
        RECT 69.835 137.105 70.125 137.150 ;
        RECT 72.120 137.090 72.440 137.150 ;
        RECT 32.675 136.950 32.965 136.995 ;
        RECT 35.795 136.950 36.085 136.995 ;
        RECT 37.685 136.950 37.975 136.995 ;
        RECT 32.675 136.810 37.975 136.950 ;
        RECT 32.675 136.765 32.965 136.810 ;
        RECT 35.795 136.765 36.085 136.810 ;
        RECT 37.685 136.765 37.975 136.810 ;
        RECT 39.480 136.950 39.770 136.995 ;
        RECT 41.340 136.950 41.630 136.995 ;
        RECT 44.120 136.950 44.410 136.995 ;
        RECT 39.480 136.810 44.410 136.950 ;
        RECT 39.480 136.765 39.770 136.810 ;
        RECT 41.340 136.765 41.630 136.810 ;
        RECT 44.120 136.765 44.410 136.810 ;
        RECT 49.600 136.950 49.890 136.995 ;
        RECT 51.460 136.950 51.750 136.995 ;
        RECT 54.240 136.950 54.530 136.995 ;
        RECT 49.600 136.810 54.530 136.950 ;
        RECT 49.600 136.765 49.890 136.810 ;
        RECT 51.460 136.765 51.750 136.810 ;
        RECT 54.240 136.765 54.530 136.810 ;
        RECT 64.730 136.950 65.020 136.995 ;
        RECT 67.510 136.950 67.800 136.995 ;
        RECT 69.370 136.950 69.660 136.995 ;
        RECT 72.670 136.950 72.810 137.490 ;
        RECT 73.960 137.430 74.280 137.690 ;
        RECT 75.340 137.630 75.660 137.690 ;
        RECT 76.735 137.630 77.025 137.675 ;
        RECT 75.340 137.490 77.025 137.630 ;
        RECT 75.340 137.430 75.660 137.490 ;
        RECT 76.735 137.445 77.025 137.490 ;
        RECT 78.100 137.630 78.420 137.690 ;
        RECT 79.955 137.630 80.245 137.675 ;
        RECT 82.240 137.630 82.560 137.690 ;
        RECT 78.100 137.620 81.090 137.630 ;
        RECT 81.870 137.620 82.560 137.630 ;
        RECT 78.100 137.490 82.560 137.620 ;
        RECT 78.100 137.430 78.420 137.490 ;
        RECT 79.955 137.445 80.245 137.490 ;
        RECT 80.950 137.480 82.010 137.490 ;
        RECT 82.240 137.430 82.560 137.490 ;
        RECT 74.880 137.290 75.200 137.350 ;
        RECT 75.815 137.290 76.105 137.335 ;
        RECT 74.880 137.150 76.105 137.290 ;
        RECT 74.880 137.090 75.200 137.150 ;
        RECT 75.815 137.105 76.105 137.150 ;
        RECT 76.275 137.290 76.565 137.335 ;
        RECT 76.275 137.150 79.710 137.290 ;
        RECT 76.275 137.105 76.565 137.150 ;
        RECT 78.100 136.950 78.420 137.010 ;
        RECT 64.730 136.810 69.660 136.950 ;
        RECT 64.730 136.765 65.020 136.810 ;
        RECT 67.510 136.765 67.800 136.810 ;
        RECT 69.370 136.765 69.660 136.810 ;
        RECT 69.910 136.810 78.420 136.950 ;
        RECT 79.570 136.950 79.710 137.150 ;
        RECT 80.875 137.105 81.165 137.335 ;
        RECT 82.790 137.290 82.930 137.830 ;
        RECT 89.155 137.785 89.445 137.830 ;
        RECT 102.890 137.970 103.180 138.015 ;
        RECT 103.400 137.970 103.720 138.030 ;
        RECT 106.150 137.970 106.440 138.015 ;
        RECT 102.890 137.830 106.440 137.970 ;
        RECT 102.890 137.785 103.180 137.830 ;
        RECT 103.400 137.770 103.720 137.830 ;
        RECT 106.150 137.785 106.440 137.830 ;
        RECT 107.070 137.970 107.360 138.015 ;
        RECT 108.930 137.970 109.220 138.015 ;
        RECT 107.070 137.830 109.220 137.970 ;
        RECT 107.070 137.785 107.360 137.830 ;
        RECT 108.930 137.785 109.220 137.830 ;
        RECT 83.160 137.430 83.480 137.690 ;
        RECT 86.395 137.630 86.685 137.675 ;
        RECT 85.090 137.490 86.685 137.630 ;
        RECT 84.540 137.290 84.860 137.350 ;
        RECT 85.090 137.290 85.230 137.490 ;
        RECT 86.395 137.445 86.685 137.490 ;
        RECT 87.760 137.630 88.080 137.690 ;
        RECT 89.615 137.630 89.905 137.675 ;
        RECT 90.075 137.630 90.365 137.675 ;
        RECT 87.760 137.490 90.365 137.630 ;
        RECT 87.760 137.430 88.080 137.490 ;
        RECT 89.615 137.445 89.905 137.490 ;
        RECT 90.075 137.445 90.365 137.490 ;
        RECT 93.295 137.630 93.585 137.675 ;
        RECT 95.580 137.630 95.900 137.690 ;
        RECT 97.880 137.630 98.200 137.690 ;
        RECT 93.295 137.490 98.200 137.630 ;
        RECT 93.295 137.445 93.585 137.490 ;
        RECT 95.580 137.430 95.900 137.490 ;
        RECT 97.880 137.430 98.200 137.490 ;
        RECT 104.750 137.630 105.040 137.675 ;
        RECT 107.070 137.630 107.285 137.785 ;
        RECT 104.750 137.490 107.285 137.630 ;
        RECT 107.540 137.630 107.860 137.690 ;
        RECT 108.015 137.630 108.305 137.675 ;
        RECT 107.540 137.490 108.305 137.630 ;
        RECT 104.750 137.445 105.040 137.490 ;
        RECT 107.540 137.430 107.860 137.490 ;
        RECT 108.015 137.445 108.305 137.490 ;
        RECT 111.235 137.445 111.525 137.675 ;
        RECT 82.790 137.150 85.230 137.290 ;
        RECT 85.475 137.290 85.765 137.335 ;
        RECT 92.375 137.290 92.665 137.335 ;
        RECT 96.040 137.290 96.360 137.350 ;
        RECT 96.515 137.290 96.805 137.335 ;
        RECT 85.475 137.150 96.805 137.290 ;
        RECT 80.950 136.950 81.090 137.105 ;
        RECT 84.540 137.090 84.860 137.150 ;
        RECT 85.475 137.105 85.765 137.150 ;
        RECT 92.375 137.105 92.665 137.150 ;
        RECT 83.160 136.950 83.480 137.010 ;
        RECT 79.570 136.810 83.480 136.950 ;
        RECT 69.910 136.670 70.050 136.810 ;
        RECT 78.100 136.750 78.420 136.810 ;
        RECT 83.160 136.750 83.480 136.810 ;
        RECT 84.080 136.950 84.400 137.010 ;
        RECT 85.550 136.950 85.690 137.105 ;
        RECT 96.040 137.090 96.360 137.150 ;
        RECT 96.515 137.105 96.805 137.150 ;
        RECT 106.620 137.290 106.940 137.350 ;
        RECT 109.855 137.290 110.145 137.335 ;
        RECT 110.300 137.290 110.620 137.350 ;
        RECT 106.620 137.150 110.620 137.290 ;
        RECT 106.620 137.090 106.940 137.150 ;
        RECT 109.855 137.105 110.145 137.150 ;
        RECT 110.300 137.090 110.620 137.150 ;
        RECT 84.080 136.810 85.690 136.950 ;
        RECT 104.750 136.950 105.040 136.995 ;
        RECT 107.530 136.950 107.820 136.995 ;
        RECT 109.390 136.950 109.680 136.995 ;
        RECT 104.750 136.810 109.680 136.950 ;
        RECT 84.080 136.750 84.400 136.810 ;
        RECT 104.750 136.765 105.040 136.810 ;
        RECT 107.530 136.765 107.820 136.810 ;
        RECT 109.390 136.765 109.680 136.810 ;
        RECT 34.400 136.610 34.720 136.670 ;
        RECT 38.080 136.610 38.400 136.670 ;
        RECT 34.400 136.470 38.400 136.610 ;
        RECT 34.400 136.410 34.720 136.470 ;
        RECT 38.080 136.410 38.400 136.470 ;
        RECT 42.220 136.610 42.540 136.670 ;
        RECT 47.985 136.610 48.275 136.655 ;
        RECT 53.260 136.610 53.580 136.670 ;
        RECT 42.220 136.470 53.580 136.610 ;
        RECT 42.220 136.410 42.540 136.470 ;
        RECT 47.985 136.425 48.275 136.470 ;
        RECT 53.260 136.410 53.580 136.470 ;
        RECT 57.860 136.655 58.180 136.670 ;
        RECT 57.860 136.425 58.395 136.655 ;
        RECT 60.175 136.610 60.465 136.655 ;
        RECT 60.620 136.610 60.940 136.670 ;
        RECT 60.175 136.470 60.940 136.610 ;
        RECT 60.175 136.425 60.465 136.470 ;
        RECT 57.860 136.410 58.180 136.425 ;
        RECT 60.620 136.410 60.940 136.470 ;
        RECT 69.820 136.410 70.140 136.670 ;
        RECT 70.280 136.610 70.600 136.670 ;
        RECT 73.055 136.610 73.345 136.655 ;
        RECT 70.280 136.470 73.345 136.610 ;
        RECT 70.280 136.410 70.600 136.470 ;
        RECT 73.055 136.425 73.345 136.470 ;
        RECT 78.575 136.610 78.865 136.655 ;
        RECT 86.380 136.610 86.700 136.670 ;
        RECT 78.575 136.470 86.700 136.610 ;
        RECT 78.575 136.425 78.865 136.470 ;
        RECT 86.380 136.410 86.700 136.470 ;
        RECT 88.235 136.610 88.525 136.655 ;
        RECT 88.680 136.610 89.000 136.670 ;
        RECT 88.235 136.470 89.000 136.610 ;
        RECT 88.235 136.425 88.525 136.470 ;
        RECT 88.680 136.410 89.000 136.470 ;
        RECT 90.520 136.410 90.840 136.670 ;
        RECT 95.580 136.410 95.900 136.670 ;
        RECT 99.720 136.410 100.040 136.670 ;
        RECT 101.560 136.610 101.880 136.670 ;
        RECT 111.310 136.610 111.450 137.445 ;
        RECT 101.560 136.470 111.450 136.610 ;
        RECT 101.560 136.410 101.880 136.470 ;
        RECT 26.970 135.790 113.450 136.270 ;
        RECT 30.275 135.590 30.565 135.635 ;
        RECT 42.680 135.590 43.000 135.650 ;
        RECT 30.275 135.450 43.000 135.590 ;
        RECT 30.275 135.405 30.565 135.450 ;
        RECT 42.680 135.390 43.000 135.450 ;
        RECT 45.440 135.590 45.760 135.650 ;
        RECT 47.985 135.590 48.275 135.635 ;
        RECT 45.440 135.450 48.275 135.590 ;
        RECT 45.440 135.390 45.760 135.450 ;
        RECT 47.985 135.405 48.275 135.450 ;
        RECT 49.580 135.590 49.900 135.650 ;
        RECT 49.580 135.450 58.090 135.590 ;
        RECT 49.580 135.390 49.900 135.450 ;
        RECT 29.355 135.250 29.645 135.295 ;
        RECT 34.400 135.250 34.720 135.310 ;
        RECT 29.355 135.110 34.720 135.250 ;
        RECT 29.355 135.065 29.645 135.110 ;
        RECT 34.400 135.050 34.720 135.110 ;
        RECT 34.875 135.065 35.165 135.295 ;
        RECT 39.480 135.250 39.770 135.295 ;
        RECT 41.340 135.250 41.630 135.295 ;
        RECT 44.120 135.250 44.410 135.295 ;
        RECT 39.480 135.110 44.410 135.250 ;
        RECT 39.480 135.065 39.770 135.110 ;
        RECT 41.340 135.065 41.630 135.110 ;
        RECT 44.120 135.065 44.410 135.110 ;
        RECT 52.770 135.250 53.060 135.295 ;
        RECT 55.550 135.250 55.840 135.295 ;
        RECT 57.410 135.250 57.700 135.295 ;
        RECT 52.770 135.110 57.700 135.250 ;
        RECT 57.950 135.250 58.090 135.450 ;
        RECT 59.255 135.405 59.545 135.635 ;
        RECT 62.245 135.590 62.535 135.635 ;
        RECT 64.760 135.590 65.080 135.650 ;
        RECT 62.245 135.450 65.080 135.590 ;
        RECT 62.245 135.405 62.535 135.450 ;
        RECT 59.330 135.250 59.470 135.405 ;
        RECT 64.760 135.390 65.080 135.450 ;
        RECT 71.905 135.590 72.195 135.635 ;
        RECT 75.340 135.590 75.660 135.650 ;
        RECT 88.220 135.635 88.540 135.650 ;
        RECT 97.880 135.635 98.200 135.650 ;
        RECT 71.905 135.450 75.660 135.590 ;
        RECT 71.905 135.405 72.195 135.450 ;
        RECT 75.340 135.390 75.660 135.450 ;
        RECT 88.005 135.405 88.540 135.635 ;
        RECT 97.665 135.405 98.200 135.635 ;
        RECT 88.220 135.390 88.540 135.405 ;
        RECT 97.880 135.390 98.200 135.405 ;
        RECT 105.700 135.590 106.020 135.650 ;
        RECT 107.555 135.590 107.845 135.635 ;
        RECT 105.700 135.450 107.845 135.590 ;
        RECT 105.700 135.390 106.020 135.450 ;
        RECT 107.555 135.405 107.845 135.450 ;
        RECT 57.950 135.110 59.470 135.250 ;
        RECT 66.110 135.250 66.400 135.295 ;
        RECT 68.890 135.250 69.180 135.295 ;
        RECT 70.750 135.250 71.040 135.295 ;
        RECT 66.110 135.110 71.040 135.250 ;
        RECT 52.770 135.065 53.060 135.110 ;
        RECT 55.550 135.065 55.840 135.110 ;
        RECT 57.410 135.065 57.700 135.110 ;
        RECT 66.110 135.065 66.400 135.110 ;
        RECT 68.890 135.065 69.180 135.110 ;
        RECT 70.750 135.065 71.040 135.110 ;
        RECT 75.770 135.250 76.060 135.295 ;
        RECT 78.550 135.250 78.840 135.295 ;
        RECT 80.410 135.250 80.700 135.295 ;
        RECT 85.475 135.250 85.765 135.295 ;
        RECT 75.770 135.110 80.700 135.250 ;
        RECT 75.770 135.065 76.060 135.110 ;
        RECT 78.550 135.065 78.840 135.110 ;
        RECT 80.410 135.065 80.700 135.110 ;
        RECT 82.330 135.110 85.765 135.250 ;
        RECT 26.120 134.910 26.440 134.970 ;
        RECT 26.120 134.770 30.030 134.910 ;
        RECT 26.120 134.710 26.440 134.770 ;
        RECT 27.040 134.570 27.360 134.630 ;
        RECT 29.890 134.615 30.030 134.770 ;
        RECT 32.100 134.710 32.420 134.970 ;
        RECT 28.435 134.570 28.725 134.615 ;
        RECT 27.040 134.430 28.725 134.570 ;
        RECT 27.040 134.370 27.360 134.430 ;
        RECT 28.435 134.385 28.725 134.430 ;
        RECT 29.815 134.385 30.105 134.615 ;
        RECT 31.180 134.570 31.500 134.630 ;
        RECT 32.575 134.570 32.865 134.615 ;
        RECT 31.180 134.430 32.865 134.570 ;
        RECT 34.950 134.570 35.090 135.065 ;
        RECT 35.320 134.910 35.640 134.970 ;
        RECT 37.175 134.910 37.465 134.955 ;
        RECT 35.320 134.770 37.465 134.910 ;
        RECT 35.320 134.710 35.640 134.770 ;
        RECT 37.175 134.725 37.465 134.770 ;
        RECT 44.520 134.910 44.840 134.970 ;
        RECT 48.905 134.910 49.195 134.955 ;
        RECT 50.040 134.910 50.360 134.970 ;
        RECT 44.520 134.770 50.360 134.910 ;
        RECT 44.520 134.710 44.840 134.770 ;
        RECT 48.905 134.725 49.195 134.770 ;
        RECT 50.040 134.710 50.360 134.770 ;
        RECT 56.480 134.910 56.800 134.970 ;
        RECT 57.875 134.910 58.165 134.955 ;
        RECT 56.480 134.770 58.165 134.910 ;
        RECT 56.480 134.710 56.800 134.770 ;
        RECT 57.875 134.725 58.165 134.770 ;
        RECT 60.160 134.710 60.480 134.970 ;
        RECT 69.375 134.910 69.665 134.955 ;
        RECT 70.280 134.910 70.600 134.970 ;
        RECT 69.375 134.770 70.600 134.910 ;
        RECT 69.375 134.725 69.665 134.770 ;
        RECT 70.280 134.710 70.600 134.770 ;
        RECT 71.215 134.910 71.505 134.955 ;
        RECT 72.120 134.910 72.440 134.970 ;
        RECT 71.215 134.770 72.440 134.910 ;
        RECT 71.215 134.725 71.505 134.770 ;
        RECT 72.120 134.710 72.440 134.770 ;
        RECT 76.720 134.910 77.040 134.970 ;
        RECT 79.035 134.910 79.325 134.955 ;
        RECT 82.330 134.910 82.470 135.110 ;
        RECT 85.475 135.065 85.765 135.110 ;
        RECT 91.870 135.250 92.160 135.295 ;
        RECT 94.650 135.250 94.940 135.295 ;
        RECT 96.510 135.250 96.800 135.295 ;
        RECT 91.870 135.110 96.800 135.250 ;
        RECT 91.870 135.065 92.160 135.110 ;
        RECT 94.650 135.065 94.940 135.110 ;
        RECT 96.510 135.065 96.800 135.110 ;
        RECT 101.530 135.250 101.820 135.295 ;
        RECT 104.310 135.250 104.600 135.295 ;
        RECT 106.170 135.250 106.460 135.295 ;
        RECT 101.530 135.110 106.460 135.250 ;
        RECT 101.530 135.065 101.820 135.110 ;
        RECT 104.310 135.065 104.600 135.110 ;
        RECT 106.170 135.065 106.460 135.110 ;
        RECT 76.720 134.770 78.790 134.910 ;
        RECT 76.720 134.710 77.040 134.770 ;
        RECT 38.080 134.570 38.400 134.630 ;
        RECT 34.950 134.430 38.400 134.570 ;
        RECT 31.180 134.370 31.500 134.430 ;
        RECT 32.575 134.385 32.865 134.430 ;
        RECT 38.080 134.370 38.400 134.430 ;
        RECT 38.540 134.370 38.860 134.630 ;
        RECT 39.015 134.570 39.305 134.615 ;
        RECT 40.380 134.570 40.700 134.630 ;
        RECT 39.015 134.430 40.700 134.570 ;
        RECT 39.015 134.385 39.305 134.430 ;
        RECT 40.380 134.370 40.700 134.430 ;
        RECT 40.855 134.570 41.145 134.615 ;
        RECT 41.300 134.570 41.620 134.630 ;
        RECT 44.120 134.570 44.410 134.615 ;
        RECT 40.855 134.430 41.620 134.570 ;
        RECT 40.855 134.385 41.145 134.430 ;
        RECT 41.300 134.370 41.620 134.430 ;
        RECT 41.875 134.430 44.410 134.570 ;
        RECT 41.875 134.275 42.090 134.430 ;
        RECT 44.120 134.385 44.410 134.430 ;
        RECT 52.770 134.570 53.060 134.615 ;
        RECT 52.770 134.430 55.305 134.570 ;
        RECT 52.770 134.385 53.060 134.430 ;
        RECT 33.035 134.230 33.325 134.275 ;
        RECT 39.940 134.230 40.230 134.275 ;
        RECT 41.800 134.230 42.090 134.275 ;
        RECT 33.035 134.090 39.690 134.230 ;
        RECT 33.035 134.045 33.325 134.090 ;
        RECT 39.550 133.890 39.690 134.090 ;
        RECT 39.940 134.090 42.090 134.230 ;
        RECT 39.940 134.045 40.230 134.090 ;
        RECT 41.800 134.045 42.090 134.090 ;
        RECT 42.680 134.275 43.000 134.290 ;
        RECT 54.180 134.275 54.500 134.290 ;
        RECT 42.680 134.230 43.010 134.275 ;
        RECT 45.980 134.230 46.270 134.275 ;
        RECT 42.680 134.090 46.270 134.230 ;
        RECT 42.680 134.045 43.010 134.090 ;
        RECT 45.980 134.045 46.270 134.090 ;
        RECT 50.910 134.230 51.200 134.275 ;
        RECT 54.170 134.230 54.500 134.275 ;
        RECT 50.910 134.090 54.500 134.230 ;
        RECT 50.910 134.045 51.200 134.090 ;
        RECT 54.170 134.045 54.500 134.090 ;
        RECT 55.090 134.275 55.305 134.430 ;
        RECT 56.020 134.370 56.340 134.630 ;
        RECT 58.320 134.570 58.640 134.630 ;
        RECT 59.255 134.570 59.545 134.615 ;
        RECT 58.320 134.430 59.545 134.570 ;
        RECT 58.320 134.370 58.640 134.430 ;
        RECT 59.255 134.385 59.545 134.430 ;
        RECT 66.110 134.570 66.400 134.615 ;
        RECT 75.770 134.570 76.060 134.615 ;
        RECT 78.650 134.570 78.790 134.770 ;
        RECT 79.035 134.770 82.470 134.910 ;
        RECT 79.035 134.725 79.325 134.770 ;
        RECT 84.080 134.710 84.400 134.970 ;
        RECT 96.960 134.910 97.280 134.970 ;
        RECT 96.960 134.770 104.550 134.910 ;
        RECT 96.960 134.710 97.280 134.770 ;
        RECT 80.875 134.570 81.165 134.615 ;
        RECT 66.110 134.430 68.645 134.570 ;
        RECT 66.110 134.385 66.400 134.430 ;
        RECT 55.090 134.230 55.380 134.275 ;
        RECT 56.950 134.230 57.240 134.275 ;
        RECT 55.090 134.090 57.240 134.230 ;
        RECT 55.090 134.045 55.380 134.090 ;
        RECT 56.950 134.045 57.240 134.090 ;
        RECT 57.400 134.230 57.720 134.290 ;
        RECT 60.635 134.230 60.925 134.275 ;
        RECT 57.400 134.090 60.925 134.230 ;
        RECT 42.680 134.030 43.000 134.045 ;
        RECT 54.180 134.030 54.500 134.045 ;
        RECT 57.400 134.030 57.720 134.090 ;
        RECT 60.635 134.045 60.925 134.090 ;
        RECT 62.000 134.230 62.320 134.290 ;
        RECT 68.430 134.275 68.645 134.430 ;
        RECT 75.770 134.430 78.305 134.570 ;
        RECT 78.650 134.430 81.165 134.570 ;
        RECT 75.770 134.385 76.060 134.430 ;
        RECT 73.960 134.275 74.280 134.290 ;
        RECT 78.090 134.275 78.305 134.430 ;
        RECT 80.875 134.385 81.165 134.430 ;
        RECT 86.380 134.370 86.700 134.630 ;
        RECT 91.870 134.570 92.160 134.615 ;
        RECT 91.870 134.430 94.405 134.570 ;
        RECT 91.870 134.385 92.160 134.430 ;
        RECT 64.250 134.230 64.540 134.275 ;
        RECT 67.510 134.230 67.800 134.275 ;
        RECT 62.000 134.090 67.800 134.230 ;
        RECT 62.000 134.030 62.320 134.090 ;
        RECT 64.250 134.045 64.540 134.090 ;
        RECT 67.510 134.045 67.800 134.090 ;
        RECT 68.430 134.230 68.720 134.275 ;
        RECT 70.290 134.230 70.580 134.275 ;
        RECT 68.430 134.090 70.580 134.230 ;
        RECT 68.430 134.045 68.720 134.090 ;
        RECT 70.290 134.045 70.580 134.090 ;
        RECT 73.910 134.230 74.280 134.275 ;
        RECT 77.170 134.230 77.460 134.275 ;
        RECT 73.910 134.090 77.460 134.230 ;
        RECT 73.910 134.045 74.280 134.090 ;
        RECT 77.170 134.045 77.460 134.090 ;
        RECT 78.090 134.230 78.380 134.275 ;
        RECT 79.950 134.230 80.240 134.275 ;
        RECT 78.090 134.090 80.240 134.230 ;
        RECT 78.090 134.045 78.380 134.090 ;
        RECT 79.950 134.045 80.240 134.090 ;
        RECT 83.635 134.230 83.925 134.275 ;
        RECT 84.540 134.230 84.860 134.290 ;
        RECT 83.635 134.090 84.860 134.230 ;
        RECT 83.635 134.045 83.925 134.090 ;
        RECT 73.960 134.030 74.280 134.045 ;
        RECT 84.540 134.030 84.860 134.090 ;
        RECT 90.010 134.230 90.300 134.275 ;
        RECT 90.520 134.230 90.840 134.290 ;
        RECT 94.190 134.275 94.405 134.430 ;
        RECT 95.120 134.370 95.440 134.630 ;
        RECT 101.530 134.570 101.820 134.615 ;
        RECT 104.410 134.570 104.550 134.770 ;
        RECT 104.780 134.710 105.100 134.970 ;
        RECT 106.620 134.570 106.940 134.630 ;
        RECT 101.530 134.430 104.065 134.570 ;
        RECT 104.410 134.430 106.940 134.570 ;
        RECT 101.530 134.385 101.820 134.430 ;
        RECT 93.270 134.230 93.560 134.275 ;
        RECT 90.010 134.090 93.560 134.230 ;
        RECT 90.010 134.045 90.300 134.090 ;
        RECT 90.520 134.030 90.840 134.090 ;
        RECT 93.270 134.045 93.560 134.090 ;
        RECT 94.190 134.230 94.480 134.275 ;
        RECT 96.050 134.230 96.340 134.275 ;
        RECT 94.190 134.090 96.340 134.230 ;
        RECT 94.190 134.045 94.480 134.090 ;
        RECT 96.050 134.045 96.340 134.090 ;
        RECT 98.800 134.230 99.120 134.290 ;
        RECT 103.850 134.275 104.065 134.430 ;
        RECT 106.620 134.370 106.940 134.430 ;
        RECT 107.095 134.385 107.385 134.615 ;
        RECT 111.220 134.570 111.540 134.630 ;
        RECT 111.695 134.570 111.985 134.615 ;
        RECT 111.220 134.430 111.985 134.570 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 99.670 134.230 99.960 134.275 ;
        RECT 102.930 134.230 103.220 134.275 ;
        RECT 98.800 134.090 103.220 134.230 ;
        RECT 98.800 134.030 99.120 134.090 ;
        RECT 99.670 134.045 99.960 134.090 ;
        RECT 102.930 134.045 103.220 134.090 ;
        RECT 103.850 134.230 104.140 134.275 ;
        RECT 105.710 134.230 106.000 134.275 ;
        RECT 103.850 134.090 106.000 134.230 ;
        RECT 103.850 134.045 104.140 134.090 ;
        RECT 105.710 134.045 106.000 134.090 ;
        RECT 46.820 133.890 47.140 133.950 ;
        RECT 39.550 133.750 47.140 133.890 ;
        RECT 46.820 133.690 47.140 133.750 ;
        RECT 55.560 133.890 55.880 133.950 ;
        RECT 58.335 133.890 58.625 133.935 ;
        RECT 55.560 133.750 58.625 133.890 ;
        RECT 55.560 133.690 55.880 133.750 ;
        RECT 58.335 133.705 58.625 133.750 ;
        RECT 79.480 133.890 79.800 133.950 ;
        RECT 81.335 133.890 81.625 133.935 ;
        RECT 79.480 133.750 81.625 133.890 ;
        RECT 79.480 133.690 79.800 133.750 ;
        RECT 81.335 133.705 81.625 133.750 ;
        RECT 83.160 133.690 83.480 133.950 ;
        RECT 104.320 133.890 104.640 133.950 ;
        RECT 107.170 133.890 107.310 134.385 ;
        RECT 111.220 134.370 111.540 134.430 ;
        RECT 111.695 134.385 111.985 134.430 ;
        RECT 104.320 133.750 107.310 133.890 ;
        RECT 104.320 133.690 104.640 133.750 ;
        RECT 110.760 133.690 111.080 133.950 ;
        RECT 26.970 133.070 113.450 133.550 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 29.340 132.670 29.660 132.930 ;
        RECT 33.940 132.870 34.260 132.930 ;
        RECT 38.080 132.870 38.400 132.930 ;
        RECT 33.940 132.730 38.400 132.870 ;
        RECT 33.940 132.670 34.260 132.730 ;
        RECT 38.080 132.670 38.400 132.730 ;
        RECT 42.220 132.670 42.540 132.930 ;
        RECT 42.695 132.870 42.985 132.915 ;
        RECT 45.440 132.870 45.760 132.930 ;
        RECT 46.375 132.870 46.665 132.915 ;
        RECT 42.695 132.730 46.665 132.870 ;
        RECT 42.695 132.685 42.985 132.730 ;
        RECT 45.440 132.670 45.760 132.730 ;
        RECT 46.375 132.685 46.665 132.730 ;
        RECT 46.820 132.670 47.140 132.930 ;
        RECT 50.040 132.870 50.360 132.930 ;
        RECT 50.515 132.870 50.805 132.915 ;
        RECT 50.040 132.730 50.805 132.870 ;
        RECT 50.040 132.670 50.360 132.730 ;
        RECT 50.515 132.685 50.805 132.730 ;
        RECT 50.975 132.870 51.265 132.915 ;
        RECT 51.420 132.870 51.740 132.930 ;
        RECT 53.505 132.870 53.795 132.915 ;
        RECT 58.320 132.870 58.640 132.930 ;
        RECT 50.975 132.730 53.795 132.870 ;
        RECT 50.975 132.685 51.265 132.730 ;
        RECT 51.420 132.670 51.740 132.730 ;
        RECT 53.505 132.685 53.795 132.730 ;
        RECT 54.270 132.730 58.640 132.870 ;
        RECT 32.100 132.530 32.420 132.590 ;
        RECT 32.675 132.530 32.965 132.575 ;
        RECT 35.915 132.530 36.565 132.575 ;
        RECT 32.100 132.390 36.565 132.530 ;
        RECT 46.910 132.530 47.050 132.670 ;
        RECT 54.270 132.530 54.410 132.730 ;
        RECT 58.320 132.670 58.640 132.730 ;
        RECT 61.080 132.870 61.400 132.930 ;
        RECT 64.315 132.870 64.605 132.915 ;
        RECT 61.080 132.730 64.605 132.870 ;
        RECT 61.080 132.670 61.400 132.730 ;
        RECT 64.315 132.685 64.605 132.730 ;
        RECT 64.760 132.670 65.080 132.930 ;
        RECT 66.615 132.685 66.905 132.915 ;
        RECT 46.910 132.390 54.410 132.530 ;
        RECT 54.640 132.530 54.960 132.590 ;
        RECT 55.510 132.530 55.800 132.575 ;
        RECT 58.770 132.530 59.060 132.575 ;
        RECT 54.640 132.390 59.060 132.530 ;
        RECT 32.100 132.330 32.420 132.390 ;
        RECT 32.675 132.345 33.265 132.390 ;
        RECT 35.915 132.345 36.565 132.390 ;
        RECT 28.420 131.990 28.740 132.250 ;
        RECT 29.815 132.190 30.105 132.235 ;
        RECT 31.180 132.190 31.500 132.250 ;
        RECT 29.815 132.050 31.500 132.190 ;
        RECT 29.815 132.005 30.105 132.050 ;
        RECT 31.180 131.990 31.500 132.050 ;
        RECT 32.975 132.030 33.265 132.345 ;
        RECT 54.640 132.330 54.960 132.390 ;
        RECT 55.510 132.345 55.800 132.390 ;
        RECT 58.770 132.345 59.060 132.390 ;
        RECT 59.690 132.530 59.980 132.575 ;
        RECT 61.550 132.530 61.840 132.575 ;
        RECT 59.690 132.390 61.840 132.530 ;
        RECT 59.690 132.345 59.980 132.390 ;
        RECT 61.550 132.345 61.840 132.390 ;
        RECT 34.055 132.190 34.345 132.235 ;
        RECT 37.635 132.190 37.925 132.235 ;
        RECT 39.470 132.190 39.760 132.235 ;
        RECT 50.500 132.190 50.820 132.250 ;
        RECT 34.055 132.050 39.760 132.190 ;
        RECT 34.055 132.005 34.345 132.050 ;
        RECT 37.635 132.005 37.925 132.050 ;
        RECT 39.470 132.005 39.760 132.050 ;
        RECT 47.370 132.050 50.820 132.190 ;
        RECT 38.540 131.650 38.860 131.910 ;
        RECT 39.935 131.850 40.225 131.895 ;
        RECT 40.380 131.850 40.700 131.910 ;
        RECT 39.935 131.710 40.700 131.850 ;
        RECT 39.935 131.665 40.225 131.710 ;
        RECT 40.380 131.650 40.700 131.710 ;
        RECT 41.760 131.850 42.080 131.910 ;
        RECT 47.370 131.895 47.510 132.050 ;
        RECT 50.500 131.990 50.820 132.050 ;
        RECT 57.370 132.190 57.660 132.235 ;
        RECT 59.690 132.190 59.905 132.345 ;
        RECT 57.370 132.050 59.905 132.190 ;
        RECT 57.370 132.005 57.660 132.050 ;
        RECT 60.620 131.990 60.940 132.250 ;
        RECT 66.690 132.190 66.830 132.685 ;
        RECT 67.980 132.670 68.300 132.930 ;
        RECT 73.515 132.870 73.805 132.915 ;
        RECT 73.960 132.870 74.280 132.930 ;
        RECT 83.160 132.870 83.480 132.930 ;
        RECT 84.540 132.915 84.860 132.930 ;
        RECT 83.865 132.870 84.155 132.915 ;
        RECT 73.515 132.730 74.280 132.870 ;
        RECT 73.515 132.685 73.805 132.730 ;
        RECT 73.960 132.670 74.280 132.730 ;
        RECT 75.430 132.730 78.330 132.870 ;
        RECT 72.135 132.530 72.425 132.575 ;
        RECT 75.430 132.530 75.570 132.730 ;
        RECT 72.135 132.390 75.570 132.530 ;
        RECT 75.820 132.530 76.110 132.575 ;
        RECT 77.680 132.530 77.970 132.575 ;
        RECT 75.820 132.390 77.970 132.530 ;
        RECT 78.190 132.530 78.330 132.730 ;
        RECT 83.160 132.730 84.155 132.870 ;
        RECT 83.160 132.670 83.480 132.730 ;
        RECT 83.865 132.685 84.155 132.730 ;
        RECT 84.540 132.685 85.075 132.915 ;
        RECT 84.540 132.670 84.860 132.685 ;
        RECT 95.120 132.670 95.440 132.930 ;
        RECT 97.895 132.870 98.185 132.915 ;
        RECT 98.340 132.870 98.660 132.930 ;
        RECT 97.895 132.730 98.660 132.870 ;
        RECT 97.895 132.685 98.185 132.730 ;
        RECT 98.340 132.670 98.660 132.730 ;
        RECT 99.735 132.870 100.025 132.915 ;
        RECT 99.735 132.730 101.330 132.870 ;
        RECT 99.735 132.685 100.025 132.730 ;
        RECT 78.600 132.530 78.890 132.575 ;
        RECT 81.860 132.530 82.150 132.575 ;
        RECT 78.190 132.390 82.150 132.530 ;
        RECT 72.135 132.345 72.425 132.390 ;
        RECT 75.820 132.345 76.110 132.390 ;
        RECT 77.680 132.345 77.970 132.390 ;
        RECT 78.600 132.345 78.890 132.390 ;
        RECT 81.860 132.345 82.150 132.390 ;
        RECT 85.920 132.530 86.240 132.590 ;
        RECT 86.790 132.530 87.080 132.575 ;
        RECT 90.050 132.530 90.340 132.575 ;
        RECT 85.920 132.390 90.340 132.530 ;
        RECT 67.075 132.190 67.365 132.235 ;
        RECT 66.690 132.050 67.365 132.190 ;
        RECT 67.075 132.005 67.365 132.050 ;
        RECT 71.675 132.005 71.965 132.235 ;
        RECT 73.055 132.005 73.345 132.235 ;
        RECT 74.895 132.190 75.185 132.235 ;
        RECT 76.260 132.190 76.580 132.250 ;
        RECT 74.895 132.050 76.580 132.190 ;
        RECT 77.755 132.190 77.970 132.345 ;
        RECT 85.920 132.330 86.240 132.390 ;
        RECT 86.790 132.345 87.080 132.390 ;
        RECT 90.050 132.345 90.340 132.390 ;
        RECT 90.970 132.530 91.260 132.575 ;
        RECT 92.830 132.530 93.120 132.575 ;
        RECT 96.960 132.530 97.280 132.590 ;
        RECT 90.970 132.390 93.120 132.530 ;
        RECT 90.970 132.345 91.260 132.390 ;
        RECT 92.830 132.345 93.120 132.390 ;
        RECT 93.830 132.390 97.280 132.530 ;
        RECT 80.000 132.190 80.290 132.235 ;
        RECT 77.755 132.050 80.290 132.190 ;
        RECT 74.895 132.005 75.185 132.050 ;
        RECT 43.615 131.850 43.905 131.895 ;
        RECT 47.295 131.850 47.585 131.895 ;
        RECT 41.760 131.710 47.585 131.850 ;
        RECT 41.760 131.650 42.080 131.710 ;
        RECT 43.615 131.665 43.905 131.710 ;
        RECT 47.295 131.665 47.585 131.710 ;
        RECT 50.055 131.665 50.345 131.895 ;
        RECT 56.480 131.850 56.800 131.910 ;
        RECT 62.475 131.850 62.765 131.895 ;
        RECT 56.480 131.710 62.765 131.850 ;
        RECT 34.055 131.510 34.345 131.555 ;
        RECT 37.175 131.510 37.465 131.555 ;
        RECT 39.065 131.510 39.355 131.555 ;
        RECT 34.055 131.370 39.355 131.510 ;
        RECT 50.130 131.510 50.270 131.665 ;
        RECT 56.480 131.650 56.800 131.710 ;
        RECT 62.475 131.665 62.765 131.710 ;
        RECT 63.855 131.665 64.145 131.895 ;
        RECT 68.900 131.850 69.220 131.910 ;
        RECT 71.750 131.850 71.890 132.005 ;
        RECT 73.130 131.850 73.270 132.005 ;
        RECT 76.260 131.990 76.580 132.050 ;
        RECT 80.000 132.005 80.290 132.050 ;
        RECT 88.650 132.190 88.940 132.235 ;
        RECT 90.970 132.190 91.185 132.345 ;
        RECT 93.830 132.235 93.970 132.390 ;
        RECT 96.960 132.330 97.280 132.390 ;
        RECT 88.650 132.050 91.185 132.190 ;
        RECT 88.650 132.005 88.940 132.050 ;
        RECT 93.755 132.005 94.045 132.235 ;
        RECT 94.215 132.190 94.505 132.235 ;
        RECT 95.580 132.190 95.900 132.250 ;
        RECT 94.215 132.050 95.900 132.190 ;
        RECT 94.215 132.005 94.505 132.050 ;
        RECT 95.580 131.990 95.900 132.050 ;
        RECT 99.720 132.190 100.040 132.250 ;
        RECT 100.655 132.190 100.945 132.235 ;
        RECT 99.720 132.050 100.945 132.190 ;
        RECT 101.190 132.190 101.330 132.730 ;
        RECT 101.575 132.685 101.865 132.915 ;
        RECT 101.650 132.530 101.790 132.685 ;
        RECT 103.400 132.670 103.720 132.930 ;
        RECT 104.320 132.870 104.640 132.930 ;
        RECT 106.175 132.870 106.465 132.915 ;
        RECT 107.080 132.870 107.400 132.930 ;
        RECT 108.935 132.870 109.225 132.915 ;
        RECT 104.320 132.730 105.930 132.870 ;
        RECT 104.320 132.670 104.640 132.730 ;
        RECT 104.780 132.530 105.100 132.590 ;
        RECT 101.650 132.390 105.100 132.530 ;
        RECT 105.790 132.530 105.930 132.730 ;
        RECT 106.175 132.730 107.400 132.870 ;
        RECT 106.175 132.685 106.465 132.730 ;
        RECT 107.080 132.670 107.400 132.730 ;
        RECT 107.630 132.730 109.225 132.870 ;
        RECT 107.630 132.530 107.770 132.730 ;
        RECT 108.935 132.685 109.225 132.730 ;
        RECT 110.775 132.530 111.065 132.575 ;
        RECT 105.790 132.390 107.770 132.530 ;
        RECT 109.470 132.390 111.065 132.530 ;
        RECT 104.780 132.330 105.100 132.390 ;
        RECT 101.190 132.050 102.710 132.190 ;
        RECT 99.720 131.990 100.040 132.050 ;
        RECT 100.655 132.005 100.945 132.050 ;
        RECT 68.900 131.710 73.270 131.850 ;
        RECT 75.800 131.850 76.120 131.910 ;
        RECT 76.735 131.850 77.025 131.895 ;
        RECT 75.800 131.710 77.025 131.850 ;
        RECT 57.370 131.510 57.660 131.555 ;
        RECT 60.150 131.510 60.440 131.555 ;
        RECT 62.010 131.510 62.300 131.555 ;
        RECT 50.130 131.370 56.940 131.510 ;
        RECT 34.055 131.325 34.345 131.370 ;
        RECT 37.175 131.325 37.465 131.370 ;
        RECT 39.065 131.325 39.355 131.370 ;
        RECT 38.080 131.170 38.400 131.230 ;
        RECT 40.395 131.170 40.685 131.215 ;
        RECT 38.080 131.030 40.685 131.170 ;
        RECT 38.080 130.970 38.400 131.030 ;
        RECT 40.395 130.985 40.685 131.030 ;
        RECT 44.520 130.970 44.840 131.230 ;
        RECT 52.815 131.170 53.105 131.215 ;
        RECT 55.560 131.170 55.880 131.230 ;
        RECT 52.815 131.030 55.880 131.170 ;
        RECT 56.800 131.170 56.940 131.370 ;
        RECT 57.370 131.370 62.300 131.510 ;
        RECT 57.370 131.325 57.660 131.370 ;
        RECT 60.150 131.325 60.440 131.370 ;
        RECT 62.010 131.325 62.300 131.370 ;
        RECT 63.930 131.510 64.070 131.665 ;
        RECT 68.900 131.650 69.220 131.710 ;
        RECT 75.800 131.650 76.120 131.710 ;
        RECT 76.735 131.665 77.025 131.710 ;
        RECT 89.600 131.850 89.920 131.910 ;
        RECT 91.915 131.850 92.205 131.895 ;
        RECT 89.600 131.710 92.205 131.850 ;
        RECT 89.600 131.650 89.920 131.710 ;
        RECT 91.915 131.665 92.205 131.710 ;
        RECT 96.040 131.850 96.360 131.910 ;
        RECT 96.515 131.850 96.805 131.895 ;
        RECT 96.040 131.710 96.805 131.850 ;
        RECT 96.040 131.650 96.360 131.710 ;
        RECT 96.515 131.665 96.805 131.710 ;
        RECT 97.435 131.850 97.725 131.895 ;
        RECT 99.260 131.850 99.580 131.910 ;
        RECT 97.435 131.710 99.580 131.850 ;
        RECT 102.570 131.850 102.710 132.050 ;
        RECT 102.940 131.990 103.260 132.250 ;
        RECT 105.255 132.190 105.545 132.235 ;
        RECT 103.490 132.050 105.545 132.190 ;
        RECT 106.635 132.180 106.925 132.235 ;
        RECT 103.490 131.850 103.630 132.050 ;
        RECT 105.255 132.005 105.545 132.050 ;
        RECT 106.525 132.040 106.925 132.180 ;
        RECT 106.635 132.005 106.925 132.040 ;
        RECT 107.080 132.190 107.400 132.250 ;
        RECT 109.470 132.190 109.610 132.390 ;
        RECT 110.775 132.345 111.065 132.390 ;
        RECT 107.080 132.050 109.610 132.190 ;
        RECT 102.570 131.710 103.630 131.850 ;
        RECT 106.710 131.850 106.850 132.005 ;
        RECT 107.080 131.990 107.400 132.050 ;
        RECT 109.840 131.990 110.160 132.250 ;
        RECT 110.315 132.190 110.605 132.235 ;
        RECT 110.315 132.050 110.990 132.190 ;
        RECT 110.315 132.005 110.605 132.050 ;
        RECT 110.850 131.850 110.990 132.050 ;
        RECT 106.710 131.710 110.990 131.850 ;
        RECT 97.435 131.665 97.725 131.710 ;
        RECT 99.260 131.650 99.580 131.710 ;
        RECT 110.390 131.570 110.530 131.710 ;
        RECT 67.060 131.510 67.380 131.570 ;
        RECT 63.930 131.370 67.380 131.510 ;
        RECT 63.930 131.170 64.070 131.370 ;
        RECT 67.060 131.310 67.380 131.370 ;
        RECT 75.360 131.510 75.650 131.555 ;
        RECT 77.220 131.510 77.510 131.555 ;
        RECT 80.000 131.510 80.290 131.555 ;
        RECT 75.360 131.370 80.290 131.510 ;
        RECT 75.360 131.325 75.650 131.370 ;
        RECT 77.220 131.325 77.510 131.370 ;
        RECT 80.000 131.325 80.290 131.370 ;
        RECT 88.650 131.510 88.940 131.555 ;
        RECT 91.430 131.510 91.720 131.555 ;
        RECT 93.290 131.510 93.580 131.555 ;
        RECT 88.650 131.370 93.580 131.510 ;
        RECT 88.650 131.325 88.940 131.370 ;
        RECT 91.430 131.325 91.720 131.370 ;
        RECT 93.290 131.325 93.580 131.370 ;
        RECT 110.300 131.310 110.620 131.570 ;
        RECT 56.800 131.030 64.070 131.170 ;
        RECT 74.880 131.170 75.200 131.230 ;
        RECT 106.160 131.170 106.480 131.230 ;
        RECT 74.880 131.030 106.480 131.170 ;
        RECT 52.815 130.985 53.105 131.030 ;
        RECT 55.560 130.970 55.880 131.030 ;
        RECT 74.880 130.970 75.200 131.030 ;
        RECT 106.160 130.970 106.480 131.030 ;
        RECT 106.620 131.170 106.940 131.230 ;
        RECT 107.095 131.170 107.385 131.215 ;
        RECT 106.620 131.030 107.385 131.170 ;
        RECT 106.620 130.970 106.940 131.030 ;
        RECT 107.095 130.985 107.385 131.030 ;
        RECT 26.970 130.350 113.450 130.830 ;
        RECT 34.875 130.150 35.165 130.195 ;
        RECT 34.875 130.010 37.390 130.150 ;
        RECT 34.875 129.965 35.165 130.010 ;
        RECT 29.355 129.810 29.645 129.855 ;
        RECT 36.700 129.810 37.020 129.870 ;
        RECT 29.355 129.670 37.020 129.810 ;
        RECT 37.250 129.810 37.390 130.010 ;
        RECT 37.620 129.950 37.940 130.210 ;
        RECT 50.960 130.150 51.280 130.210 ;
        RECT 39.090 130.010 51.280 130.150 ;
        RECT 39.090 129.810 39.230 130.010 ;
        RECT 50.960 129.950 51.280 130.010 ;
        RECT 54.640 129.950 54.960 130.210 ;
        RECT 56.020 130.150 56.340 130.210 ;
        RECT 56.495 130.150 56.785 130.195 ;
        RECT 56.020 130.010 56.785 130.150 ;
        RECT 56.020 129.950 56.340 130.010 ;
        RECT 56.495 129.965 56.785 130.010 ;
        RECT 59.700 130.150 60.020 130.210 ;
        RECT 60.175 130.150 60.465 130.195 ;
        RECT 59.700 130.010 60.465 130.150 ;
        RECT 59.700 129.950 60.020 130.010 ;
        RECT 60.175 129.965 60.465 130.010 ;
        RECT 64.775 130.150 65.065 130.195 ;
        RECT 65.220 130.150 65.540 130.210 ;
        RECT 64.775 130.010 65.540 130.150 ;
        RECT 64.775 129.965 65.065 130.010 ;
        RECT 65.220 129.950 65.540 130.010 ;
        RECT 68.900 130.150 69.220 130.210 ;
        RECT 68.900 130.010 85.690 130.150 ;
        RECT 68.900 129.950 69.220 130.010 ;
        RECT 37.250 129.670 39.230 129.810 ;
        RECT 39.475 129.810 39.765 129.855 ;
        RECT 40.840 129.810 41.160 129.870 ;
        RECT 39.475 129.670 41.160 129.810 ;
        RECT 29.355 129.625 29.645 129.670 ;
        RECT 36.700 129.610 37.020 129.670 ;
        RECT 39.475 129.625 39.765 129.670 ;
        RECT 40.840 129.610 41.160 129.670 ;
        RECT 41.300 129.610 41.620 129.870 ;
        RECT 42.680 129.810 43.000 129.870 ;
        RECT 41.850 129.670 43.000 129.810 ;
        RECT 26.120 129.470 26.440 129.530 ;
        RECT 35.320 129.470 35.640 129.530 ;
        RECT 40.395 129.470 40.685 129.515 ;
        RECT 41.850 129.470 41.990 129.670 ;
        RECT 42.680 129.610 43.000 129.670 ;
        RECT 46.935 129.810 47.225 129.855 ;
        RECT 50.055 129.810 50.345 129.855 ;
        RECT 51.945 129.810 52.235 129.855 ;
        RECT 46.935 129.670 52.235 129.810 ;
        RECT 46.935 129.625 47.225 129.670 ;
        RECT 50.055 129.625 50.345 129.670 ;
        RECT 51.945 129.625 52.235 129.670 ;
        RECT 75.800 129.810 76.120 129.870 ;
        RECT 77.655 129.810 77.945 129.855 ;
        RECT 80.400 129.810 80.720 129.870 ;
        RECT 75.800 129.670 77.945 129.810 ;
        RECT 75.800 129.610 76.120 129.670 ;
        RECT 77.655 129.625 77.945 129.670 ;
        RECT 78.190 129.670 80.720 129.810 ;
        RECT 44.520 129.470 44.840 129.530 ;
        RECT 26.120 129.330 30.030 129.470 ;
        RECT 26.120 129.270 26.440 129.330 ;
        RECT 28.435 129.130 28.725 129.175 ;
        RECT 28.880 129.130 29.200 129.190 ;
        RECT 28.435 128.990 29.200 129.130 ;
        RECT 28.435 128.945 28.725 128.990 ;
        RECT 28.880 128.930 29.200 128.990 ;
        RECT 29.340 129.130 29.660 129.190 ;
        RECT 29.890 129.175 30.030 129.330 ;
        RECT 31.730 129.330 40.150 129.470 ;
        RECT 31.730 129.175 31.870 129.330 ;
        RECT 35.320 129.270 35.640 129.330 ;
        RECT 29.815 129.130 30.105 129.175 ;
        RECT 31.655 129.130 31.945 129.175 ;
        RECT 29.340 128.990 31.945 129.130 ;
        RECT 29.340 128.930 29.660 128.990 ;
        RECT 29.815 128.945 30.105 128.990 ;
        RECT 31.655 128.945 31.945 128.990 ;
        RECT 33.940 128.930 34.260 129.190 ;
        RECT 37.250 129.175 37.390 129.330 ;
        RECT 37.175 128.945 37.465 129.175 ;
        RECT 38.080 129.130 38.400 129.190 ;
        RECT 40.010 129.175 40.150 129.330 ;
        RECT 40.395 129.330 41.990 129.470 ;
        RECT 42.310 129.330 44.840 129.470 ;
        RECT 40.395 129.285 40.685 129.330 ;
        RECT 42.310 129.175 42.450 129.330 ;
        RECT 44.520 129.270 44.840 129.330 ;
        RECT 52.815 129.470 53.105 129.515 ;
        RECT 57.400 129.470 57.720 129.530 ;
        RECT 52.815 129.330 57.720 129.470 ;
        RECT 52.815 129.285 53.105 129.330 ;
        RECT 57.400 129.270 57.720 129.330 ;
        RECT 58.320 129.270 58.640 129.530 ;
        RECT 69.820 129.470 70.140 129.530 ;
        RECT 78.190 129.470 78.330 129.670 ;
        RECT 80.400 129.610 80.720 129.670 ;
        RECT 85.550 129.810 85.690 130.010 ;
        RECT 85.920 129.950 86.240 130.210 ;
        RECT 89.600 129.950 89.920 130.210 ;
        RECT 90.535 130.150 90.825 130.195 ;
        RECT 90.980 130.150 91.300 130.210 ;
        RECT 102.940 130.150 103.260 130.210 ;
        RECT 90.535 130.010 91.300 130.150 ;
        RECT 90.535 129.965 90.825 130.010 ;
        RECT 90.980 129.950 91.300 130.010 ;
        RECT 91.530 130.010 103.260 130.150 ;
        RECT 87.760 129.810 88.080 129.870 ;
        RECT 85.550 129.670 88.080 129.810 ;
        RECT 79.480 129.470 79.800 129.530 ;
        RECT 59.330 129.330 70.140 129.470 ;
        RECT 38.555 129.130 38.845 129.175 ;
        RECT 38.080 128.990 38.845 129.130 ;
        RECT 38.080 128.930 38.400 128.990 ;
        RECT 38.555 128.945 38.845 128.990 ;
        RECT 39.935 128.945 40.225 129.175 ;
        RECT 42.235 128.945 42.525 129.175 ;
        RECT 42.695 129.130 42.985 129.175 ;
        RECT 44.980 129.130 45.300 129.190 ;
        RECT 42.695 128.990 45.300 129.130 ;
        RECT 42.695 128.945 42.985 128.990 ;
        RECT 44.980 128.930 45.300 128.990 ;
        RECT 32.115 128.790 32.405 128.835 ;
        RECT 39.000 128.790 39.320 128.850 ;
        RECT 32.115 128.650 39.320 128.790 ;
        RECT 32.115 128.605 32.405 128.650 ;
        RECT 39.000 128.590 39.320 128.650 ;
        RECT 39.460 128.790 39.780 128.850 ;
        RECT 45.855 128.835 46.145 129.150 ;
        RECT 46.935 129.130 47.225 129.175 ;
        RECT 50.515 129.130 50.805 129.175 ;
        RECT 52.350 129.130 52.640 129.175 ;
        RECT 46.935 128.990 52.640 129.130 ;
        RECT 46.935 128.945 47.225 128.990 ;
        RECT 50.515 128.945 50.805 128.990 ;
        RECT 52.350 128.945 52.640 128.990 ;
        RECT 53.720 129.130 54.040 129.190 ;
        RECT 54.195 129.130 54.485 129.175 ;
        RECT 53.720 128.990 54.485 129.130 ;
        RECT 53.720 128.930 54.040 128.990 ;
        RECT 54.195 128.945 54.485 128.990 ;
        RECT 55.560 128.930 55.880 129.190 ;
        RECT 59.330 129.175 59.470 129.330 ;
        RECT 69.820 129.270 70.140 129.330 ;
        RECT 76.350 129.330 78.330 129.470 ;
        RECT 78.650 129.330 79.800 129.470 ;
        RECT 56.955 128.945 57.245 129.175 ;
        RECT 59.255 128.945 59.545 129.175 ;
        RECT 65.235 129.130 65.525 129.175 ;
        RECT 65.680 129.130 66.000 129.190 ;
        RECT 65.235 128.990 66.000 129.130 ;
        RECT 65.235 128.945 65.525 128.990 ;
        RECT 45.555 128.790 46.145 128.835 ;
        RECT 48.795 128.790 49.445 128.835 ;
        RECT 39.460 128.650 49.445 128.790 ;
        RECT 39.460 128.590 39.780 128.650 ;
        RECT 45.555 128.605 45.845 128.650 ;
        RECT 48.795 128.605 49.445 128.650 ;
        RECT 50.960 128.790 51.280 128.850 ;
        RECT 51.435 128.790 51.725 128.835 ;
        RECT 50.960 128.650 51.725 128.790 ;
        RECT 50.960 128.590 51.280 128.650 ;
        RECT 51.435 128.605 51.725 128.650 ;
        RECT 52.800 128.790 53.120 128.850 ;
        RECT 57.030 128.790 57.170 128.945 ;
        RECT 65.680 128.930 66.000 128.990 ;
        RECT 71.660 129.130 71.980 129.190 ;
        RECT 76.350 129.175 76.490 129.330 ;
        RECT 78.650 129.175 78.790 129.330 ;
        RECT 79.480 129.270 79.800 129.330 ;
        RECT 74.895 129.130 75.185 129.175 ;
        RECT 71.660 128.990 75.185 129.130 ;
        RECT 71.660 128.930 71.980 128.990 ;
        RECT 74.895 128.945 75.185 128.990 ;
        RECT 76.275 128.945 76.565 129.175 ;
        RECT 78.575 128.945 78.865 129.175 ;
        RECT 79.035 129.130 79.325 129.175 ;
        RECT 79.940 129.130 80.260 129.190 ;
        RECT 85.550 129.175 85.690 129.670 ;
        RECT 87.760 129.610 88.080 129.670 ;
        RECT 79.035 128.990 80.260 129.130 ;
        RECT 79.035 128.945 79.325 128.990 ;
        RECT 79.940 128.930 80.260 128.990 ;
        RECT 85.475 128.945 85.765 129.175 ;
        RECT 88.680 128.930 89.000 129.190 ;
        RECT 90.075 129.130 90.365 129.175 ;
        RECT 91.530 129.130 91.670 130.010 ;
        RECT 102.940 129.950 103.260 130.010 ;
        RECT 106.160 130.150 106.480 130.210 ;
        RECT 110.760 130.150 111.080 130.210 ;
        RECT 106.160 130.010 111.080 130.150 ;
        RECT 106.160 129.950 106.480 130.010 ;
        RECT 110.760 129.950 111.080 130.010 ;
        RECT 96.960 129.810 97.280 129.870 ;
        RECT 102.445 129.810 102.735 129.855 ;
        RECT 104.335 129.810 104.625 129.855 ;
        RECT 107.455 129.810 107.745 129.855 ;
        RECT 96.960 129.670 101.790 129.810 ;
        RECT 96.960 129.610 97.280 129.670 ;
        RECT 91.900 129.470 92.220 129.530 ;
        RECT 91.900 129.330 93.510 129.470 ;
        RECT 91.900 129.270 92.220 129.330 ;
        RECT 93.370 129.175 93.510 129.330 ;
        RECT 97.050 129.330 100.410 129.470 ;
        RECT 90.075 128.990 91.670 129.130 ;
        RECT 90.075 128.945 90.365 128.990 ;
        RECT 92.835 128.945 93.125 129.175 ;
        RECT 93.295 128.945 93.585 129.175 ;
        RECT 52.800 128.650 57.170 128.790 ;
        RECT 75.340 128.790 75.660 128.850 ;
        RECT 80.415 128.790 80.705 128.835 ;
        RECT 86.840 128.790 87.160 128.850 ;
        RECT 92.910 128.790 93.050 128.945 ;
        RECT 94.660 128.930 94.980 129.190 ;
        RECT 97.050 129.175 97.190 129.330 ;
        RECT 96.975 129.130 97.265 129.175 ;
        RECT 95.210 128.990 97.265 129.130 ;
        RECT 95.210 128.790 95.350 128.990 ;
        RECT 96.975 128.945 97.265 128.990 ;
        RECT 98.340 128.930 98.660 129.190 ;
        RECT 100.270 129.175 100.410 129.330 ;
        RECT 101.650 129.175 101.790 129.670 ;
        RECT 102.445 129.670 107.745 129.810 ;
        RECT 102.445 129.625 102.735 129.670 ;
        RECT 104.335 129.625 104.625 129.670 ;
        RECT 107.455 129.625 107.745 129.670 ;
        RECT 100.195 129.130 100.485 129.175 ;
        RECT 100.195 128.990 101.330 129.130 ;
        RECT 100.195 128.945 100.485 128.990 ;
        RECT 98.800 128.790 99.120 128.850 ;
        RECT 75.340 128.650 77.410 128.790 ;
        RECT 52.800 128.590 53.120 128.650 ;
        RECT 75.340 128.590 75.660 128.650 ;
        RECT 30.275 128.450 30.565 128.495 ;
        RECT 43.140 128.450 43.460 128.510 ;
        RECT 30.275 128.310 43.460 128.450 ;
        RECT 30.275 128.265 30.565 128.310 ;
        RECT 43.140 128.250 43.460 128.310 ;
        RECT 57.860 128.250 58.180 128.510 ;
        RECT 75.800 128.250 76.120 128.510 ;
        RECT 77.270 128.495 77.410 128.650 ;
        RECT 80.415 128.650 95.350 128.790 ;
        RECT 95.670 128.650 99.120 128.790 ;
        RECT 80.415 128.605 80.705 128.650 ;
        RECT 86.840 128.590 87.160 128.650 ;
        RECT 77.195 128.265 77.485 128.495 ;
        RECT 91.440 128.450 91.760 128.510 ;
        RECT 92.375 128.450 92.665 128.495 ;
        RECT 91.440 128.310 92.665 128.450 ;
        RECT 91.440 128.250 91.760 128.310 ;
        RECT 92.375 128.265 92.665 128.310 ;
        RECT 94.215 128.450 94.505 128.495 ;
        RECT 95.120 128.450 95.440 128.510 ;
        RECT 95.670 128.495 95.810 128.650 ;
        RECT 98.800 128.590 99.120 128.650 ;
        RECT 94.215 128.310 95.440 128.450 ;
        RECT 94.215 128.265 94.505 128.310 ;
        RECT 95.120 128.250 95.440 128.310 ;
        RECT 95.595 128.265 95.885 128.495 ;
        RECT 96.040 128.450 96.360 128.510 ;
        RECT 96.515 128.450 96.805 128.495 ;
        RECT 96.040 128.310 96.805 128.450 ;
        RECT 96.040 128.250 96.360 128.310 ;
        RECT 96.515 128.265 96.805 128.310 ;
        RECT 99.260 128.250 99.580 128.510 ;
        RECT 100.640 128.250 100.960 128.510 ;
        RECT 101.190 128.450 101.330 128.990 ;
        RECT 101.575 128.945 101.865 129.175 ;
        RECT 102.040 129.130 102.330 129.175 ;
        RECT 103.875 129.130 104.165 129.175 ;
        RECT 107.455 129.130 107.745 129.175 ;
        RECT 102.040 128.990 107.745 129.130 ;
        RECT 102.040 128.945 102.330 128.990 ;
        RECT 103.875 128.945 104.165 128.990 ;
        RECT 107.455 128.945 107.745 128.990 ;
        RECT 102.955 128.790 103.245 128.835 ;
        RECT 104.320 128.790 104.640 128.850 ;
        RECT 102.955 128.650 104.640 128.790 ;
        RECT 102.955 128.605 103.245 128.650 ;
        RECT 104.320 128.590 104.640 128.650 ;
        RECT 105.235 128.790 105.885 128.835 ;
        RECT 106.620 128.790 106.940 128.850 ;
        RECT 108.535 128.835 108.825 129.150 ;
        RECT 108.535 128.790 109.125 128.835 ;
        RECT 105.235 128.650 109.125 128.790 ;
        RECT 105.235 128.605 105.885 128.650 ;
        RECT 106.620 128.590 106.940 128.650 ;
        RECT 108.835 128.605 109.125 128.650 ;
        RECT 111.695 128.790 111.985 128.835 ;
        RECT 113.980 128.790 114.300 128.850 ;
        RECT 111.695 128.650 114.300 128.790 ;
        RECT 111.695 128.605 111.985 128.650 ;
        RECT 113.980 128.590 114.300 128.650 ;
        RECT 110.300 128.450 110.620 128.510 ;
        RECT 101.190 128.310 110.620 128.450 ;
        RECT 110.300 128.250 110.620 128.310 ;
        RECT 26.970 127.630 113.450 128.110 ;
        RECT 29.355 127.430 29.645 127.475 ;
        RECT 29.800 127.430 30.120 127.490 ;
        RECT 29.355 127.290 30.120 127.430 ;
        RECT 29.355 127.245 29.645 127.290 ;
        RECT 29.800 127.230 30.120 127.290 ;
        RECT 31.195 127.430 31.485 127.475 ;
        RECT 36.240 127.430 36.560 127.490 ;
        RECT 31.195 127.290 36.560 127.430 ;
        RECT 31.195 127.245 31.485 127.290 ;
        RECT 36.240 127.230 36.560 127.290 ;
        RECT 36.715 127.430 37.005 127.475 ;
        RECT 39.000 127.430 39.320 127.490 ;
        RECT 43.600 127.430 43.920 127.490 ;
        RECT 36.715 127.290 38.770 127.430 ;
        RECT 36.715 127.245 37.005 127.290 ;
        RECT 27.960 127.090 28.280 127.150 ;
        RECT 37.160 127.090 37.480 127.150 ;
        RECT 38.630 127.135 38.770 127.290 ;
        RECT 39.000 127.290 43.920 127.430 ;
        RECT 39.000 127.230 39.320 127.290 ;
        RECT 43.600 127.230 43.920 127.290 ;
        RECT 53.735 127.430 54.025 127.475 ;
        RECT 54.180 127.430 54.500 127.490 ;
        RECT 53.735 127.290 54.500 127.430 ;
        RECT 53.735 127.245 54.025 127.290 ;
        RECT 54.180 127.230 54.500 127.290 ;
        RECT 58.780 127.430 59.100 127.490 ;
        RECT 99.260 127.430 99.580 127.490 ;
        RECT 104.320 127.430 104.640 127.490 ;
        RECT 58.780 127.290 66.370 127.430 ;
        RECT 58.780 127.230 59.100 127.290 ;
        RECT 40.840 127.135 41.160 127.150 ;
        RECT 27.960 126.950 34.630 127.090 ;
        RECT 27.960 126.890 28.280 126.950 ;
        RECT 29.340 126.750 29.660 126.810 ;
        RECT 29.815 126.750 30.105 126.795 ;
        RECT 29.340 126.610 30.105 126.750 ;
        RECT 29.340 126.550 29.660 126.610 ;
        RECT 29.815 126.565 30.105 126.610 ;
        RECT 30.260 126.550 30.580 126.810 ;
        RECT 30.720 126.750 31.040 126.810 ;
        RECT 34.490 126.795 34.630 126.950 ;
        RECT 35.870 126.950 37.480 127.090 ;
        RECT 35.870 126.795 36.010 126.950 ;
        RECT 37.160 126.890 37.480 126.950 ;
        RECT 38.555 126.905 38.845 127.135 ;
        RECT 40.835 127.090 41.485 127.135 ;
        RECT 44.435 127.090 44.725 127.135 ;
        RECT 40.835 126.950 44.725 127.090 ;
        RECT 40.835 126.905 41.485 126.950 ;
        RECT 44.135 126.905 44.725 126.950 ;
        RECT 57.415 127.090 57.705 127.135 ;
        RECT 57.860 127.090 58.180 127.150 ;
        RECT 57.415 126.950 58.180 127.090 ;
        RECT 57.415 126.905 57.705 126.950 ;
        RECT 40.840 126.890 41.160 126.905 ;
        RECT 33.035 126.750 33.325 126.795 ;
        RECT 30.720 126.610 33.325 126.750 ;
        RECT 30.720 126.550 31.040 126.610 ;
        RECT 33.035 126.565 33.325 126.610 ;
        RECT 34.415 126.565 34.705 126.795 ;
        RECT 35.795 126.565 36.085 126.795 ;
        RECT 37.640 126.750 37.930 126.795 ;
        RECT 39.475 126.750 39.765 126.795 ;
        RECT 43.055 126.750 43.345 126.795 ;
        RECT 37.640 126.610 43.345 126.750 ;
        RECT 37.640 126.565 37.930 126.610 ;
        RECT 39.475 126.565 39.765 126.610 ;
        RECT 43.055 126.565 43.345 126.610 ;
        RECT 44.135 126.590 44.425 126.905 ;
        RECT 57.860 126.890 58.180 126.950 ;
        RECT 59.695 127.090 60.345 127.135 ;
        RECT 60.620 127.090 60.940 127.150 ;
        RECT 66.230 127.135 66.370 127.290 ;
        RECT 99.260 127.290 103.170 127.430 ;
        RECT 99.260 127.230 99.580 127.290 ;
        RECT 63.295 127.090 63.585 127.135 ;
        RECT 59.695 126.950 63.585 127.090 ;
        RECT 59.695 126.905 60.345 126.950 ;
        RECT 60.620 126.890 60.940 126.950 ;
        RECT 62.995 126.905 63.585 126.950 ;
        RECT 66.155 126.905 66.445 127.135 ;
        RECT 75.800 127.090 76.120 127.150 ;
        RECT 76.275 127.090 76.565 127.135 ;
        RECT 75.800 126.950 76.565 127.090 ;
        RECT 51.895 126.750 52.185 126.795 ;
        RECT 53.720 126.750 54.040 126.810 ;
        RECT 54.195 126.750 54.485 126.795 ;
        RECT 51.895 126.610 54.485 126.750 ;
        RECT 51.895 126.565 52.185 126.610 ;
        RECT 53.720 126.550 54.040 126.610 ;
        RECT 54.195 126.565 54.485 126.610 ;
        RECT 54.655 126.750 54.945 126.795 ;
        RECT 55.100 126.750 55.420 126.810 ;
        RECT 54.655 126.610 55.420 126.750 ;
        RECT 54.655 126.565 54.945 126.610 ;
        RECT 55.100 126.550 55.420 126.610 ;
        RECT 56.500 126.750 56.790 126.795 ;
        RECT 58.335 126.750 58.625 126.795 ;
        RECT 61.915 126.750 62.205 126.795 ;
        RECT 56.500 126.610 62.205 126.750 ;
        RECT 56.500 126.565 56.790 126.610 ;
        RECT 58.335 126.565 58.625 126.610 ;
        RECT 61.915 126.565 62.205 126.610 ;
        RECT 62.995 126.590 63.285 126.905 ;
        RECT 75.800 126.890 76.120 126.950 ;
        RECT 76.275 126.905 76.565 126.950 ;
        RECT 78.555 127.090 79.205 127.135 ;
        RECT 82.155 127.090 82.445 127.135 ;
        RECT 84.080 127.090 84.400 127.150 ;
        RECT 78.555 126.950 84.400 127.090 ;
        RECT 78.555 126.905 79.205 126.950 ;
        RECT 81.855 126.905 82.445 126.950 ;
        RECT 66.600 126.550 66.920 126.810 ;
        RECT 67.995 126.565 68.285 126.795 ;
        RECT 69.375 126.565 69.665 126.795 ;
        RECT 37.175 126.410 37.465 126.455 ;
        RECT 40.380 126.410 40.700 126.470 ;
        RECT 41.300 126.410 41.620 126.470 ;
        RECT 37.175 126.270 41.620 126.410 ;
        RECT 37.175 126.225 37.465 126.270 ;
        RECT 40.380 126.210 40.700 126.270 ;
        RECT 41.300 126.210 41.620 126.270 ;
        RECT 47.295 126.225 47.585 126.455 ;
        RECT 33.955 126.070 34.245 126.115 ;
        RECT 35.780 126.070 36.100 126.130 ;
        RECT 33.955 125.930 36.100 126.070 ;
        RECT 33.955 125.885 34.245 125.930 ;
        RECT 35.780 125.870 36.100 125.930 ;
        RECT 38.045 126.070 38.335 126.115 ;
        RECT 39.935 126.070 40.225 126.115 ;
        RECT 43.055 126.070 43.345 126.115 ;
        RECT 38.045 125.930 43.345 126.070 ;
        RECT 38.045 125.885 38.335 125.930 ;
        RECT 39.935 125.885 40.225 125.930 ;
        RECT 43.055 125.885 43.345 125.930 ;
        RECT 35.320 125.530 35.640 125.790 ;
        RECT 40.380 125.730 40.700 125.790 ;
        RECT 47.370 125.730 47.510 126.225 ;
        RECT 50.500 126.210 50.820 126.470 ;
        RECT 56.035 126.410 56.325 126.455 ;
        RECT 57.400 126.410 57.720 126.470 ;
        RECT 61.080 126.410 61.400 126.470 ;
        RECT 56.035 126.270 61.400 126.410 ;
        RECT 56.035 126.225 56.325 126.270 ;
        RECT 57.400 126.210 57.720 126.270 ;
        RECT 61.080 126.210 61.400 126.270 ;
        RECT 64.760 126.410 65.080 126.470 ;
        RECT 68.070 126.410 68.210 126.565 ;
        RECT 64.760 126.270 68.210 126.410 ;
        RECT 64.760 126.210 65.080 126.270 ;
        RECT 52.340 126.070 52.660 126.130 ;
        RECT 56.905 126.070 57.195 126.115 ;
        RECT 58.795 126.070 59.085 126.115 ;
        RECT 61.915 126.070 62.205 126.115 ;
        RECT 69.450 126.070 69.590 126.565 ;
        RECT 73.040 126.550 73.360 126.810 ;
        RECT 75.360 126.750 75.650 126.795 ;
        RECT 77.195 126.750 77.485 126.795 ;
        RECT 80.775 126.750 81.065 126.795 ;
        RECT 75.360 126.610 81.065 126.750 ;
        RECT 75.360 126.565 75.650 126.610 ;
        RECT 77.195 126.565 77.485 126.610 ;
        RECT 80.775 126.565 81.065 126.610 ;
        RECT 81.855 126.590 82.145 126.905 ;
        RECT 84.080 126.890 84.400 126.950 ;
        RECT 90.635 127.090 90.925 127.135 ;
        RECT 91.440 127.090 91.760 127.150 ;
        RECT 93.875 127.090 94.525 127.135 ;
        RECT 90.635 126.950 94.525 127.090 ;
        RECT 90.635 126.905 91.225 126.950 ;
        RECT 83.620 126.750 83.940 126.810 ;
        RECT 86.395 126.750 86.685 126.795 ;
        RECT 83.620 126.610 86.685 126.750 ;
        RECT 83.620 126.550 83.940 126.610 ;
        RECT 86.395 126.565 86.685 126.610 ;
        RECT 90.935 126.590 91.225 126.905 ;
        RECT 91.440 126.890 91.760 126.950 ;
        RECT 93.875 126.905 94.525 126.950 ;
        RECT 95.120 127.090 95.440 127.150 ;
        RECT 96.515 127.090 96.805 127.135 ;
        RECT 95.120 126.950 96.805 127.090 ;
        RECT 95.120 126.890 95.440 126.950 ;
        RECT 96.515 126.905 96.805 126.950 ;
        RECT 96.960 127.090 97.280 127.150 ;
        RECT 103.030 127.135 103.170 127.290 ;
        RECT 104.320 127.290 111.910 127.430 ;
        RECT 104.320 127.230 104.640 127.290 ;
        RECT 96.960 126.950 101.330 127.090 ;
        RECT 96.960 126.890 97.280 126.950 ;
        RECT 97.970 126.810 98.110 126.950 ;
        RECT 92.015 126.750 92.305 126.795 ;
        RECT 95.595 126.750 95.885 126.795 ;
        RECT 97.430 126.750 97.720 126.795 ;
        RECT 92.015 126.610 97.720 126.750 ;
        RECT 92.015 126.565 92.305 126.610 ;
        RECT 95.595 126.565 95.885 126.610 ;
        RECT 97.430 126.565 97.720 126.610 ;
        RECT 97.880 126.550 98.200 126.810 ;
        RECT 99.275 126.565 99.565 126.795 ;
        RECT 74.895 126.410 75.185 126.455 ;
        RECT 76.260 126.410 76.580 126.470 ;
        RECT 74.895 126.270 76.580 126.410 ;
        RECT 74.895 126.225 75.185 126.270 ;
        RECT 76.260 126.210 76.580 126.270 ;
        RECT 76.720 126.410 77.040 126.470 ;
        RECT 85.015 126.410 85.305 126.455 ;
        RECT 76.720 126.270 85.305 126.410 ;
        RECT 76.720 126.210 77.040 126.270 ;
        RECT 85.015 126.225 85.305 126.270 ;
        RECT 87.775 126.225 88.065 126.455 ;
        RECT 96.500 126.410 96.820 126.470 ;
        RECT 99.350 126.410 99.490 126.565 ;
        RECT 96.500 126.270 99.490 126.410 ;
        RECT 101.190 126.410 101.330 126.950 ;
        RECT 102.955 126.905 103.245 127.135 ;
        RECT 105.235 127.090 105.885 127.135 ;
        RECT 108.835 127.090 109.125 127.135 ;
        RECT 109.840 127.090 110.160 127.150 ;
        RECT 111.770 127.135 111.910 127.290 ;
        RECT 105.235 126.950 110.160 127.090 ;
        RECT 105.235 126.905 105.885 126.950 ;
        RECT 108.535 126.905 109.125 126.950 ;
        RECT 102.040 126.750 102.330 126.795 ;
        RECT 103.875 126.750 104.165 126.795 ;
        RECT 107.455 126.750 107.745 126.795 ;
        RECT 102.040 126.610 107.745 126.750 ;
        RECT 102.040 126.565 102.330 126.610 ;
        RECT 103.875 126.565 104.165 126.610 ;
        RECT 107.455 126.565 107.745 126.610 ;
        RECT 108.535 126.590 108.825 126.905 ;
        RECT 109.840 126.890 110.160 126.950 ;
        RECT 111.695 126.905 111.985 127.135 ;
        RECT 101.575 126.410 101.865 126.455 ;
        RECT 101.190 126.270 101.865 126.410 ;
        RECT 52.340 125.930 56.710 126.070 ;
        RECT 52.340 125.870 52.660 125.930 ;
        RECT 40.380 125.590 47.510 125.730 ;
        RECT 55.575 125.730 55.865 125.775 ;
        RECT 56.020 125.730 56.340 125.790 ;
        RECT 55.575 125.590 56.340 125.730 ;
        RECT 56.570 125.730 56.710 125.930 ;
        RECT 56.905 125.930 62.205 126.070 ;
        RECT 56.905 125.885 57.195 125.930 ;
        RECT 58.795 125.885 59.085 125.930 ;
        RECT 61.915 125.885 62.205 125.930 ;
        RECT 63.010 125.930 69.590 126.070 ;
        RECT 75.765 126.070 76.055 126.115 ;
        RECT 77.655 126.070 77.945 126.115 ;
        RECT 80.775 126.070 81.065 126.115 ;
        RECT 75.765 125.930 81.065 126.070 ;
        RECT 87.850 126.070 87.990 126.225 ;
        RECT 96.500 126.210 96.820 126.270 ;
        RECT 101.575 126.225 101.865 126.270 ;
        RECT 90.980 126.070 91.300 126.130 ;
        RECT 87.850 125.930 91.300 126.070 ;
        RECT 63.010 125.730 63.150 125.930 ;
        RECT 75.765 125.885 76.055 125.930 ;
        RECT 77.655 125.885 77.945 125.930 ;
        RECT 80.775 125.885 81.065 125.930 ;
        RECT 90.980 125.870 91.300 125.930 ;
        RECT 92.015 126.070 92.305 126.115 ;
        RECT 95.135 126.070 95.425 126.115 ;
        RECT 97.025 126.070 97.315 126.115 ;
        RECT 92.015 125.930 97.315 126.070 ;
        RECT 92.015 125.885 92.305 125.930 ;
        RECT 95.135 125.885 95.425 125.930 ;
        RECT 97.025 125.885 97.315 125.930 ;
        RECT 102.445 126.070 102.735 126.115 ;
        RECT 104.335 126.070 104.625 126.115 ;
        RECT 107.455 126.070 107.745 126.115 ;
        RECT 102.445 125.930 107.745 126.070 ;
        RECT 102.445 125.885 102.735 125.930 ;
        RECT 104.335 125.885 104.625 125.930 ;
        RECT 107.455 125.885 107.745 125.930 ;
        RECT 56.570 125.590 63.150 125.730 ;
        RECT 40.380 125.530 40.700 125.590 ;
        RECT 55.575 125.545 55.865 125.590 ;
        RECT 56.020 125.530 56.340 125.590 ;
        RECT 67.520 125.530 67.840 125.790 ;
        RECT 68.455 125.730 68.745 125.775 ;
        RECT 68.900 125.730 69.220 125.790 ;
        RECT 68.455 125.590 69.220 125.730 ;
        RECT 68.455 125.545 68.745 125.590 ;
        RECT 68.900 125.530 69.220 125.590 ;
        RECT 70.280 125.530 70.600 125.790 ;
        RECT 73.960 125.530 74.280 125.790 ;
        RECT 87.300 125.530 87.620 125.790 ;
        RECT 98.340 125.530 98.660 125.790 ;
        RECT 26.970 124.910 113.450 125.390 ;
        RECT 27.500 124.710 27.820 124.770 ;
        RECT 28.895 124.710 29.185 124.755 ;
        RECT 27.500 124.570 29.185 124.710 ;
        RECT 27.500 124.510 27.820 124.570 ;
        RECT 28.895 124.525 29.185 124.570 ;
        RECT 31.640 124.710 31.960 124.770 ;
        RECT 32.115 124.710 32.405 124.755 ;
        RECT 31.640 124.570 32.405 124.710 ;
        RECT 31.640 124.510 31.960 124.570 ;
        RECT 32.115 124.525 32.405 124.570 ;
        RECT 38.540 124.510 38.860 124.770 ;
        RECT 39.460 124.510 39.780 124.770 ;
        RECT 44.060 124.710 44.380 124.770 ;
        RECT 40.930 124.570 44.380 124.710 ;
        RECT 40.930 124.370 41.070 124.570 ;
        RECT 44.060 124.510 44.380 124.570 ;
        RECT 76.260 124.710 76.580 124.770 ;
        RECT 84.080 124.710 84.400 124.770 ;
        RECT 85.015 124.710 85.305 124.755 ;
        RECT 76.260 124.570 82.470 124.710 ;
        RECT 76.260 124.510 76.580 124.570 ;
        RECT 38.630 124.230 41.070 124.370 ;
        RECT 41.265 124.370 41.555 124.415 ;
        RECT 43.155 124.370 43.445 124.415 ;
        RECT 46.275 124.370 46.565 124.415 ;
        RECT 41.265 124.230 46.565 124.370 ;
        RECT 32.100 124.030 32.420 124.090 ;
        RECT 33.495 124.030 33.785 124.075 ;
        RECT 32.100 123.890 33.785 124.030 ;
        RECT 32.100 123.830 32.420 123.890 ;
        RECT 33.495 123.845 33.785 123.890 ;
        RECT 29.340 123.490 29.660 123.750 ;
        RECT 32.575 123.690 32.865 123.735 ;
        RECT 33.035 123.690 33.325 123.735 ;
        RECT 34.415 123.690 34.705 123.735 ;
        RECT 36.255 123.690 36.545 123.735 ;
        RECT 32.575 123.550 36.545 123.690 ;
        RECT 32.575 123.505 32.865 123.550 ;
        RECT 33.035 123.505 33.325 123.550 ;
        RECT 34.415 123.505 34.705 123.550 ;
        RECT 36.255 123.505 36.545 123.550 ;
        RECT 37.635 123.690 37.925 123.735 ;
        RECT 38.630 123.690 38.770 124.230 ;
        RECT 41.265 124.185 41.555 124.230 ;
        RECT 43.155 124.185 43.445 124.230 ;
        RECT 46.275 124.185 46.565 124.230 ;
        RECT 55.215 124.370 55.505 124.415 ;
        RECT 58.335 124.370 58.625 124.415 ;
        RECT 60.225 124.370 60.515 124.415 ;
        RECT 55.215 124.230 60.515 124.370 ;
        RECT 55.215 124.185 55.505 124.230 ;
        RECT 58.335 124.185 58.625 124.230 ;
        RECT 60.225 124.185 60.515 124.230 ;
        RECT 66.255 124.370 66.545 124.415 ;
        RECT 69.375 124.370 69.665 124.415 ;
        RECT 71.265 124.370 71.555 124.415 ;
        RECT 76.350 124.370 76.490 124.510 ;
        RECT 66.255 124.230 71.555 124.370 ;
        RECT 66.255 124.185 66.545 124.230 ;
        RECT 69.375 124.185 69.665 124.230 ;
        RECT 71.265 124.185 71.555 124.230 ;
        RECT 72.210 124.230 76.490 124.370 ;
        RECT 76.835 124.370 77.125 124.415 ;
        RECT 79.955 124.370 80.245 124.415 ;
        RECT 81.845 124.370 82.135 124.415 ;
        RECT 76.835 124.230 82.135 124.370 ;
        RECT 50.500 124.030 50.820 124.090 ;
        RECT 40.010 123.890 50.820 124.030 ;
        RECT 37.635 123.550 38.770 123.690 ;
        RECT 39.015 123.690 39.305 123.735 ;
        RECT 40.010 123.690 40.150 123.890 ;
        RECT 50.500 123.830 50.820 123.890 ;
        RECT 50.975 124.030 51.265 124.075 ;
        RECT 53.720 124.030 54.040 124.090 ;
        RECT 50.975 123.890 54.040 124.030 ;
        RECT 50.975 123.845 51.265 123.890 ;
        RECT 53.720 123.830 54.040 123.890 ;
        RECT 56.020 124.030 56.340 124.090 ;
        RECT 59.715 124.030 60.005 124.075 ;
        RECT 56.020 123.890 60.005 124.030 ;
        RECT 56.020 123.830 56.340 123.890 ;
        RECT 59.715 123.845 60.005 123.890 ;
        RECT 61.080 123.830 61.400 124.090 ;
        RECT 67.520 124.030 67.840 124.090 ;
        RECT 72.210 124.075 72.350 124.230 ;
        RECT 76.835 124.185 77.125 124.230 ;
        RECT 79.955 124.185 80.245 124.230 ;
        RECT 81.845 124.185 82.135 124.230 ;
        RECT 70.755 124.030 71.045 124.075 ;
        RECT 67.520 123.890 71.045 124.030 ;
        RECT 67.520 123.830 67.840 123.890 ;
        RECT 70.755 123.845 71.045 123.890 ;
        RECT 72.135 123.845 72.425 124.075 ;
        RECT 75.340 124.030 75.660 124.090 ;
        RECT 81.335 124.030 81.625 124.075 ;
        RECT 75.340 123.890 81.625 124.030 ;
        RECT 82.330 124.030 82.470 124.570 ;
        RECT 84.080 124.570 85.305 124.710 ;
        RECT 84.080 124.510 84.400 124.570 ;
        RECT 85.015 124.525 85.305 124.570 ;
        RECT 101.100 124.710 101.420 124.770 ;
        RECT 109.395 124.710 109.685 124.755 ;
        RECT 109.840 124.710 110.160 124.770 ;
        RECT 101.100 124.570 108.230 124.710 ;
        RECT 101.100 124.510 101.420 124.570 ;
        RECT 92.015 124.370 92.305 124.415 ;
        RECT 95.135 124.370 95.425 124.415 ;
        RECT 97.025 124.370 97.315 124.415 ;
        RECT 92.015 124.230 97.315 124.370 ;
        RECT 92.015 124.185 92.305 124.230 ;
        RECT 95.135 124.185 95.425 124.230 ;
        RECT 97.025 124.185 97.315 124.230 ;
        RECT 102.595 124.370 102.885 124.415 ;
        RECT 105.715 124.370 106.005 124.415 ;
        RECT 107.605 124.370 107.895 124.415 ;
        RECT 102.595 124.230 107.895 124.370 ;
        RECT 102.595 124.185 102.885 124.230 ;
        RECT 105.715 124.185 106.005 124.230 ;
        RECT 107.605 124.185 107.895 124.230 ;
        RECT 82.715 124.030 83.005 124.075 ;
        RECT 82.330 123.890 83.005 124.030 ;
        RECT 75.340 123.830 75.660 123.890 ;
        RECT 81.335 123.845 81.625 123.890 ;
        RECT 82.715 123.845 83.005 123.890 ;
        RECT 87.300 124.030 87.620 124.090 ;
        RECT 96.515 124.030 96.805 124.075 ;
        RECT 87.300 123.890 96.805 124.030 ;
        RECT 87.300 123.830 87.620 123.890 ;
        RECT 96.515 123.845 96.805 123.890 ;
        RECT 97.880 123.830 98.200 124.090 ;
        RECT 98.800 124.030 99.120 124.090 ;
        RECT 107.095 124.030 107.385 124.075 ;
        RECT 98.800 123.890 107.385 124.030 ;
        RECT 108.090 124.030 108.230 124.570 ;
        RECT 109.395 124.570 110.160 124.710 ;
        RECT 109.395 124.525 109.685 124.570 ;
        RECT 109.840 124.510 110.160 124.570 ;
        RECT 108.090 123.890 111.450 124.030 ;
        RECT 98.800 123.830 99.120 123.890 ;
        RECT 107.095 123.845 107.385 123.890 ;
        RECT 39.015 123.550 40.150 123.690 ;
        RECT 37.635 123.505 37.925 123.550 ;
        RECT 39.015 123.505 39.305 123.550 ;
        RECT 40.395 123.505 40.685 123.735 ;
        RECT 40.860 123.690 41.150 123.735 ;
        RECT 42.695 123.690 42.985 123.735 ;
        RECT 46.275 123.690 46.565 123.735 ;
        RECT 40.860 123.550 46.565 123.690 ;
        RECT 40.860 123.505 41.150 123.550 ;
        RECT 42.695 123.505 42.985 123.550 ;
        RECT 46.275 123.505 46.565 123.550 ;
        RECT 47.280 123.710 47.600 123.750 ;
        RECT 36.330 123.350 36.470 123.505 ;
        RECT 39.090 123.350 39.230 123.505 ;
        RECT 36.330 123.210 39.230 123.350 ;
        RECT 40.470 123.350 40.610 123.505 ;
        RECT 47.280 123.490 47.645 123.710 ;
        RECT 41.300 123.350 41.620 123.410 ;
        RECT 47.355 123.395 47.645 123.490 ;
        RECT 40.470 123.210 41.620 123.350 ;
        RECT 41.300 123.150 41.620 123.210 ;
        RECT 41.775 123.165 42.065 123.395 ;
        RECT 44.055 123.350 44.705 123.395 ;
        RECT 47.355 123.350 47.945 123.395 ;
        RECT 44.055 123.210 47.945 123.350 ;
        RECT 44.055 123.165 44.705 123.210 ;
        RECT 47.655 123.165 47.945 123.210 ;
        RECT 49.580 123.350 49.900 123.410 ;
        RECT 54.135 123.395 54.425 123.710 ;
        RECT 55.215 123.690 55.505 123.735 ;
        RECT 58.795 123.690 59.085 123.735 ;
        RECT 60.630 123.690 60.920 123.735 ;
        RECT 55.215 123.550 60.920 123.690 ;
        RECT 55.215 123.505 55.505 123.550 ;
        RECT 58.795 123.505 59.085 123.550 ;
        RECT 60.630 123.505 60.920 123.550 ;
        RECT 50.515 123.350 50.805 123.395 ;
        RECT 49.580 123.210 50.805 123.350 ;
        RECT 34.860 122.810 35.180 123.070 ;
        RECT 36.715 123.010 37.005 123.055 ;
        RECT 40.840 123.010 41.160 123.070 ;
        RECT 36.715 122.870 41.160 123.010 ;
        RECT 41.850 123.010 41.990 123.165 ;
        RECT 49.580 123.150 49.900 123.210 ;
        RECT 50.515 123.165 50.805 123.210 ;
        RECT 53.835 123.350 54.425 123.395 ;
        RECT 56.020 123.350 56.340 123.410 ;
        RECT 57.075 123.350 57.725 123.395 ;
        RECT 53.835 123.210 57.725 123.350 ;
        RECT 53.835 123.165 54.125 123.210 ;
        RECT 56.020 123.150 56.340 123.210 ;
        RECT 57.075 123.165 57.725 123.210 ;
        RECT 62.000 123.150 62.320 123.410 ;
        RECT 65.175 123.395 65.465 123.710 ;
        RECT 66.255 123.690 66.545 123.735 ;
        RECT 69.835 123.690 70.125 123.735 ;
        RECT 71.670 123.690 71.960 123.735 ;
        RECT 66.255 123.550 71.960 123.690 ;
        RECT 66.255 123.505 66.545 123.550 ;
        RECT 69.835 123.505 70.125 123.550 ;
        RECT 71.670 123.505 71.960 123.550 ;
        RECT 64.875 123.350 65.465 123.395 ;
        RECT 65.680 123.350 66.000 123.410 ;
        RECT 68.115 123.350 68.765 123.395 ;
        RECT 64.875 123.210 68.765 123.350 ;
        RECT 64.875 123.165 65.165 123.210 ;
        RECT 65.680 123.150 66.000 123.210 ;
        RECT 68.115 123.165 68.765 123.210 ;
        RECT 72.580 123.150 72.900 123.410 ;
        RECT 75.755 123.395 76.045 123.710 ;
        RECT 76.835 123.690 77.125 123.735 ;
        RECT 80.415 123.690 80.705 123.735 ;
        RECT 82.250 123.690 82.540 123.735 ;
        RECT 76.835 123.550 82.540 123.690 ;
        RECT 76.835 123.505 77.125 123.550 ;
        RECT 80.415 123.505 80.705 123.550 ;
        RECT 82.250 123.505 82.540 123.550 ;
        RECT 84.095 123.690 84.385 123.735 ;
        RECT 85.475 123.690 85.765 123.735 ;
        RECT 86.840 123.690 87.160 123.750 ;
        RECT 84.095 123.550 87.160 123.690 ;
        RECT 84.095 123.505 84.385 123.550 ;
        RECT 85.475 123.505 85.765 123.550 ;
        RECT 86.840 123.490 87.160 123.550 ;
        RECT 75.455 123.350 76.045 123.395 ;
        RECT 78.695 123.350 79.345 123.395 ;
        RECT 83.635 123.350 83.925 123.395 ;
        RECT 75.455 123.210 83.925 123.350 ;
        RECT 75.455 123.165 75.745 123.210 ;
        RECT 78.695 123.165 79.345 123.210 ;
        RECT 83.635 123.165 83.925 123.210 ;
        RECT 87.775 123.165 88.065 123.395 ;
        RECT 88.220 123.350 88.540 123.410 ;
        RECT 90.935 123.395 91.225 123.710 ;
        RECT 92.015 123.690 92.305 123.735 ;
        RECT 95.595 123.690 95.885 123.735 ;
        RECT 97.430 123.690 97.720 123.735 ;
        RECT 92.015 123.550 97.720 123.690 ;
        RECT 92.015 123.505 92.305 123.550 ;
        RECT 95.595 123.505 95.885 123.550 ;
        RECT 97.430 123.505 97.720 123.550 ;
        RECT 90.635 123.350 91.225 123.395 ;
        RECT 93.875 123.350 94.525 123.395 ;
        RECT 88.220 123.210 94.525 123.350 ;
        RECT 53.260 123.010 53.580 123.070 ;
        RECT 41.850 122.870 53.580 123.010 ;
        RECT 36.715 122.825 37.005 122.870 ;
        RECT 40.840 122.810 41.160 122.870 ;
        RECT 53.260 122.810 53.580 122.870 ;
        RECT 86.380 122.810 86.700 123.070 ;
        RECT 86.840 123.010 87.160 123.070 ;
        RECT 87.850 123.010 87.990 123.165 ;
        RECT 88.220 123.150 88.540 123.210 ;
        RECT 90.635 123.165 90.925 123.210 ;
        RECT 93.875 123.165 94.525 123.210 ;
        RECT 98.355 123.350 98.645 123.395 ;
        RECT 100.180 123.350 100.500 123.410 ;
        RECT 98.355 123.210 100.500 123.350 ;
        RECT 98.355 123.165 98.645 123.210 ;
        RECT 100.180 123.150 100.500 123.210 ;
        RECT 100.640 123.350 100.960 123.410 ;
        RECT 101.515 123.395 101.805 123.710 ;
        RECT 102.595 123.690 102.885 123.735 ;
        RECT 106.175 123.690 106.465 123.735 ;
        RECT 108.010 123.690 108.300 123.735 ;
        RECT 102.595 123.550 108.300 123.690 ;
        RECT 102.595 123.505 102.885 123.550 ;
        RECT 106.175 123.505 106.465 123.550 ;
        RECT 108.010 123.505 108.300 123.550 ;
        RECT 108.475 123.505 108.765 123.735 ;
        RECT 109.855 123.690 110.145 123.735 ;
        RECT 110.300 123.690 110.620 123.750 ;
        RECT 111.310 123.735 111.450 123.890 ;
        RECT 109.855 123.550 110.620 123.690 ;
        RECT 109.855 123.505 110.145 123.550 ;
        RECT 101.215 123.350 101.805 123.395 ;
        RECT 104.455 123.350 105.105 123.395 ;
        RECT 108.550 123.350 108.690 123.505 ;
        RECT 110.300 123.490 110.620 123.550 ;
        RECT 111.235 123.505 111.525 123.735 ;
        RECT 111.680 123.350 112.000 123.410 ;
        RECT 100.640 123.210 105.105 123.350 ;
        RECT 100.640 123.150 100.960 123.210 ;
        RECT 101.215 123.165 101.505 123.210 ;
        RECT 104.455 123.165 105.105 123.210 ;
        RECT 108.090 123.210 112.000 123.350 ;
        RECT 86.840 122.870 87.990 123.010 ;
        RECT 97.880 123.010 98.200 123.070 ;
        RECT 108.090 123.010 108.230 123.210 ;
        RECT 111.680 123.150 112.000 123.210 ;
        RECT 97.880 122.870 108.230 123.010 ;
        RECT 86.840 122.810 87.160 122.870 ;
        RECT 97.880 122.810 98.200 122.870 ;
        RECT 110.300 122.810 110.620 123.070 ;
        RECT 26.970 122.190 113.450 122.670 ;
        RECT 35.320 121.990 35.640 122.050 ;
        RECT 47.280 121.990 47.600 122.050 ;
        RECT 47.755 121.990 48.045 122.035 ;
        RECT 35.320 121.850 45.210 121.990 ;
        RECT 35.320 121.790 35.640 121.850 ;
        RECT 34.860 121.650 35.180 121.710 ;
        RECT 45.070 121.695 45.210 121.850 ;
        RECT 47.280 121.850 48.045 121.990 ;
        RECT 47.280 121.790 47.600 121.850 ;
        RECT 47.755 121.805 48.045 121.850 ;
        RECT 50.960 121.790 51.280 122.050 ;
        RECT 53.260 121.790 53.580 122.050 ;
        RECT 56.020 121.790 56.340 122.050 ;
        RECT 60.620 121.790 60.940 122.050 ;
        RECT 62.935 121.990 63.225 122.035 ;
        RECT 65.680 121.990 66.000 122.050 ;
        RECT 62.935 121.850 66.000 121.990 ;
        RECT 62.935 121.805 63.225 121.850 ;
        RECT 65.680 121.790 66.000 121.850 ;
        RECT 69.360 121.990 69.680 122.050 ;
        RECT 75.815 121.990 76.105 122.035 ;
        RECT 69.360 121.850 76.105 121.990 ;
        RECT 69.360 121.790 69.680 121.850 ;
        RECT 75.815 121.805 76.105 121.850 ;
        RECT 88.220 121.790 88.540 122.050 ;
        RECT 109.840 121.990 110.160 122.050 ;
        RECT 101.650 121.850 110.160 121.990 ;
        RECT 39.115 121.650 39.405 121.695 ;
        RECT 42.355 121.650 43.005 121.695 ;
        RECT 34.860 121.510 43.005 121.650 ;
        RECT 34.860 121.450 35.180 121.510 ;
        RECT 39.115 121.465 39.705 121.510 ;
        RECT 42.355 121.465 43.005 121.510 ;
        RECT 44.995 121.465 45.285 121.695 ;
        RECT 46.360 121.650 46.680 121.710 ;
        RECT 66.715 121.650 67.005 121.695 ;
        RECT 68.900 121.650 69.220 121.710 ;
        RECT 69.955 121.650 70.605 121.695 ;
        RECT 46.360 121.510 50.270 121.650 ;
        RECT 39.415 121.150 39.705 121.465 ;
        RECT 46.360 121.450 46.680 121.510 ;
        RECT 50.130 121.355 50.270 121.510 ;
        RECT 66.715 121.510 70.605 121.650 ;
        RECT 66.715 121.465 67.305 121.510 ;
        RECT 40.495 121.310 40.785 121.355 ;
        RECT 44.075 121.310 44.365 121.355 ;
        RECT 45.910 121.310 46.200 121.355 ;
        RECT 40.495 121.170 46.200 121.310 ;
        RECT 40.495 121.125 40.785 121.170 ;
        RECT 44.075 121.125 44.365 121.170 ;
        RECT 45.910 121.125 46.200 121.170 ;
        RECT 48.215 121.125 48.505 121.355 ;
        RECT 50.055 121.125 50.345 121.355 ;
        RECT 51.880 121.310 52.200 121.370 ;
        RECT 54.195 121.310 54.485 121.355 ;
        RECT 51.880 121.170 54.485 121.310 ;
        RECT 35.780 120.970 36.100 121.030 ;
        RECT 36.255 120.970 36.545 121.015 ;
        RECT 35.780 120.830 36.545 120.970 ;
        RECT 35.780 120.770 36.100 120.830 ;
        RECT 36.255 120.785 36.545 120.830 ;
        RECT 41.300 120.970 41.620 121.030 ;
        RECT 46.375 120.970 46.665 121.015 ;
        RECT 41.300 120.830 46.665 120.970 ;
        RECT 48.290 120.970 48.430 121.125 ;
        RECT 51.880 121.110 52.200 121.170 ;
        RECT 54.195 121.125 54.485 121.170 ;
        RECT 56.495 121.310 56.785 121.355 ;
        RECT 60.175 121.310 60.465 121.355 ;
        RECT 62.475 121.310 62.765 121.355 ;
        RECT 64.760 121.310 65.080 121.370 ;
        RECT 56.495 121.170 65.080 121.310 ;
        RECT 56.495 121.125 56.785 121.170 ;
        RECT 60.175 121.125 60.465 121.170 ;
        RECT 62.475 121.125 62.765 121.170 ;
        RECT 50.500 120.970 50.820 121.030 ;
        RECT 56.570 120.970 56.710 121.125 ;
        RECT 64.760 121.110 65.080 121.170 ;
        RECT 67.015 121.150 67.305 121.465 ;
        RECT 68.900 121.450 69.220 121.510 ;
        RECT 69.955 121.465 70.605 121.510 ;
        RECT 73.960 121.650 74.280 121.710 ;
        RECT 78.115 121.650 78.405 121.695 ;
        RECT 73.960 121.510 78.405 121.650 ;
        RECT 73.960 121.450 74.280 121.510 ;
        RECT 78.115 121.465 78.405 121.510 ;
        RECT 80.395 121.650 81.045 121.695 ;
        RECT 83.995 121.650 84.285 121.695 ;
        RECT 86.380 121.650 86.700 121.710 ;
        RECT 96.040 121.695 96.360 121.710 ;
        RECT 80.395 121.510 86.700 121.650 ;
        RECT 80.395 121.465 81.045 121.510 ;
        RECT 83.695 121.465 84.285 121.510 ;
        RECT 68.095 121.310 68.385 121.355 ;
        RECT 71.675 121.310 71.965 121.355 ;
        RECT 73.510 121.310 73.800 121.355 ;
        RECT 68.095 121.170 73.800 121.310 ;
        RECT 68.095 121.125 68.385 121.170 ;
        RECT 71.675 121.125 71.965 121.170 ;
        RECT 73.510 121.125 73.800 121.170 ;
        RECT 74.880 121.310 75.200 121.370 ;
        RECT 76.275 121.310 76.565 121.355 ;
        RECT 74.880 121.170 76.565 121.310 ;
        RECT 74.880 121.110 75.200 121.170 ;
        RECT 76.275 121.125 76.565 121.170 ;
        RECT 76.720 121.110 77.040 121.370 ;
        RECT 77.200 121.310 77.490 121.355 ;
        RECT 79.035 121.310 79.325 121.355 ;
        RECT 82.615 121.310 82.905 121.355 ;
        RECT 77.200 121.170 82.905 121.310 ;
        RECT 77.200 121.125 77.490 121.170 ;
        RECT 79.035 121.125 79.325 121.170 ;
        RECT 82.615 121.125 82.905 121.170 ;
        RECT 83.695 121.150 83.985 121.465 ;
        RECT 86.380 121.450 86.700 121.510 ;
        RECT 92.475 121.650 92.765 121.695 ;
        RECT 95.715 121.650 96.365 121.695 ;
        RECT 92.475 121.510 96.365 121.650 ;
        RECT 92.475 121.465 93.065 121.510 ;
        RECT 95.715 121.465 96.365 121.510 ;
        RECT 87.300 121.310 87.620 121.370 ;
        RECT 87.775 121.310 88.065 121.355 ;
        RECT 87.300 121.170 88.065 121.310 ;
        RECT 87.300 121.110 87.620 121.170 ;
        RECT 87.775 121.125 88.065 121.170 ;
        RECT 92.775 121.150 93.065 121.465 ;
        RECT 96.040 121.450 96.360 121.465 ;
        RECT 98.340 121.450 98.660 121.710 ;
        RECT 101.650 121.695 101.790 121.850 ;
        RECT 109.840 121.790 110.160 121.850 ;
        RECT 101.575 121.465 101.865 121.695 ;
        RECT 104.435 121.650 104.725 121.695 ;
        RECT 107.675 121.650 108.325 121.695 ;
        RECT 104.435 121.510 108.325 121.650 ;
        RECT 104.435 121.465 105.025 121.510 ;
        RECT 107.675 121.465 108.325 121.510 ;
        RECT 104.735 121.370 105.025 121.465 ;
        RECT 110.300 121.450 110.620 121.710 ;
        RECT 93.855 121.310 94.145 121.355 ;
        RECT 97.435 121.310 97.725 121.355 ;
        RECT 99.270 121.310 99.560 121.355 ;
        RECT 93.855 121.170 99.560 121.310 ;
        RECT 93.855 121.125 94.145 121.170 ;
        RECT 97.435 121.125 97.725 121.170 ;
        RECT 99.270 121.125 99.560 121.170 ;
        RECT 104.735 121.150 105.100 121.370 ;
        RECT 104.780 121.110 105.100 121.150 ;
        RECT 105.815 121.310 106.105 121.355 ;
        RECT 109.395 121.310 109.685 121.355 ;
        RECT 111.230 121.310 111.520 121.355 ;
        RECT 105.815 121.170 111.520 121.310 ;
        RECT 105.815 121.125 106.105 121.170 ;
        RECT 109.395 121.125 109.685 121.170 ;
        RECT 111.230 121.125 111.520 121.170 ;
        RECT 111.680 121.110 112.000 121.370 ;
        RECT 48.290 120.830 56.710 120.970 ;
        RECT 63.855 120.970 64.145 121.015 ;
        RECT 67.520 120.970 67.840 121.030 ;
        RECT 63.855 120.830 67.840 120.970 ;
        RECT 41.300 120.770 41.620 120.830 ;
        RECT 46.375 120.785 46.665 120.830 ;
        RECT 50.500 120.770 50.820 120.830 ;
        RECT 63.855 120.785 64.145 120.830 ;
        RECT 67.520 120.770 67.840 120.830 ;
        RECT 70.280 120.970 70.600 121.030 ;
        RECT 72.595 120.970 72.885 121.015 ;
        RECT 70.280 120.830 72.885 120.970 ;
        RECT 70.280 120.770 70.600 120.830 ;
        RECT 72.595 120.785 72.885 120.830 ;
        RECT 73.975 120.970 74.265 121.015 ;
        RECT 76.810 120.970 76.950 121.110 ;
        RECT 73.975 120.830 76.950 120.970 ;
        RECT 81.780 120.970 82.100 121.030 ;
        RECT 86.855 120.970 87.145 121.015 ;
        RECT 81.780 120.830 87.145 120.970 ;
        RECT 73.975 120.785 74.265 120.830 ;
        RECT 81.780 120.770 82.100 120.830 ;
        RECT 86.855 120.785 87.145 120.830 ;
        RECT 89.615 120.970 89.905 121.015 ;
        RECT 95.580 120.970 95.900 121.030 ;
        RECT 89.615 120.830 95.900 120.970 ;
        RECT 89.615 120.785 89.905 120.830 ;
        RECT 95.580 120.770 95.900 120.830 ;
        RECT 97.880 120.970 98.200 121.030 ;
        RECT 99.735 120.970 100.025 121.015 ;
        RECT 97.880 120.830 100.025 120.970 ;
        RECT 97.880 120.770 98.200 120.830 ;
        RECT 99.735 120.785 100.025 120.830 ;
        RECT 40.495 120.630 40.785 120.675 ;
        RECT 43.615 120.630 43.905 120.675 ;
        RECT 45.505 120.630 45.795 120.675 ;
        RECT 40.495 120.490 45.795 120.630 ;
        RECT 40.495 120.445 40.785 120.490 ;
        RECT 43.615 120.445 43.905 120.490 ;
        RECT 45.505 120.445 45.795 120.490 ;
        RECT 68.095 120.630 68.385 120.675 ;
        RECT 71.215 120.630 71.505 120.675 ;
        RECT 73.105 120.630 73.395 120.675 ;
        RECT 68.095 120.490 73.395 120.630 ;
        RECT 68.095 120.445 68.385 120.490 ;
        RECT 71.215 120.445 71.505 120.490 ;
        RECT 73.105 120.445 73.395 120.490 ;
        RECT 77.605 120.630 77.895 120.675 ;
        RECT 79.495 120.630 79.785 120.675 ;
        RECT 82.615 120.630 82.905 120.675 ;
        RECT 77.605 120.490 82.905 120.630 ;
        RECT 77.605 120.445 77.895 120.490 ;
        RECT 79.495 120.445 79.785 120.490 ;
        RECT 82.615 120.445 82.905 120.490 ;
        RECT 93.855 120.630 94.145 120.675 ;
        RECT 96.975 120.630 97.265 120.675 ;
        RECT 98.865 120.630 99.155 120.675 ;
        RECT 93.855 120.490 99.155 120.630 ;
        RECT 93.855 120.445 94.145 120.490 ;
        RECT 96.975 120.445 97.265 120.490 ;
        RECT 98.865 120.445 99.155 120.490 ;
        RECT 105.815 120.630 106.105 120.675 ;
        RECT 108.935 120.630 109.225 120.675 ;
        RECT 110.825 120.630 111.115 120.675 ;
        RECT 105.815 120.490 111.115 120.630 ;
        RECT 105.815 120.445 106.105 120.490 ;
        RECT 108.935 120.445 109.225 120.490 ;
        RECT 110.825 120.445 111.115 120.490 ;
        RECT 26.970 119.470 113.450 119.950 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 46.850 206.760 47.110 207.080 ;
        RECT 99.750 206.760 100.010 207.080 ;
        RECT 40.400 206.225 40.680 206.595 ;
        RECT 39.030 204.380 39.290 204.700 ;
        RECT 32.510 203.845 34.390 204.215 ;
        RECT 39.090 203.000 39.230 204.380 ;
        RECT 39.950 203.360 40.210 203.680 ;
        RECT 40.010 203.195 40.150 203.360 ;
        RECT 32.590 202.680 32.850 203.000 ;
        RECT 39.030 202.680 39.290 203.000 ;
        RECT 39.940 202.825 40.220 203.195 ;
        RECT 27.530 201.660 27.790 201.980 ;
        RECT 32.130 201.660 32.390 201.980 ;
        RECT 27.590 201.180 27.730 201.660 ;
        RECT 32.190 201.180 32.330 201.660 ;
        RECT 27.130 201.040 27.730 201.180 ;
        RECT 30.810 201.040 32.330 201.180 ;
        RECT 26.610 200.300 26.870 200.620 ;
        RECT 25.230 199.960 25.490 200.280 ;
        RECT 25.290 171.040 25.430 199.960 ;
        RECT 26.150 196.900 26.410 197.220 ;
        RECT 26.210 185.660 26.350 196.900 ;
        RECT 26.150 185.340 26.410 185.660 ;
        RECT 26.150 183.300 26.410 183.620 ;
        RECT 26.210 177.840 26.350 183.300 ;
        RECT 26.150 177.520 26.410 177.840 ;
        RECT 25.230 170.720 25.490 171.040 ;
        RECT 26.150 161.880 26.410 162.200 ;
        RECT 26.210 135.000 26.350 161.880 ;
        RECT 26.670 157.100 26.810 200.300 ;
        RECT 27.130 181.580 27.270 201.040 ;
        RECT 28.450 199.620 28.710 199.940 ;
        RECT 29.370 199.620 29.630 199.940 ;
        RECT 27.990 196.560 28.250 196.880 ;
        RECT 27.530 191.800 27.790 192.120 ;
        RECT 27.070 181.260 27.330 181.580 ;
        RECT 27.070 177.520 27.330 177.840 ;
        RECT 27.130 174.780 27.270 177.520 ;
        RECT 27.070 174.460 27.330 174.780 ;
        RECT 27.590 168.320 27.730 191.800 ;
        RECT 27.530 168.000 27.790 168.320 ;
        RECT 28.050 165.260 28.190 196.560 ;
        RECT 28.510 178.860 28.650 199.620 ;
        RECT 29.430 197.560 29.570 199.620 ;
        RECT 29.830 198.940 30.090 199.260 ;
        RECT 30.290 198.940 30.550 199.260 ;
        RECT 29.370 197.240 29.630 197.560 ;
        RECT 28.910 194.180 29.170 194.500 ;
        RECT 28.970 184.300 29.110 194.180 ;
        RECT 29.430 189.400 29.570 197.240 ;
        RECT 29.370 189.080 29.630 189.400 ;
        RECT 28.910 183.980 29.170 184.300 ;
        RECT 29.430 183.530 29.570 189.080 ;
        RECT 28.970 183.390 29.570 183.530 ;
        RECT 28.970 181.435 29.110 183.390 ;
        RECT 29.370 182.620 29.630 182.940 ;
        RECT 28.900 181.065 29.180 181.435 ;
        RECT 28.910 180.920 29.170 181.065 ;
        RECT 28.450 178.540 28.710 178.860 ;
        RECT 28.910 177.860 29.170 178.180 ;
        RECT 28.450 175.140 28.710 175.460 ;
        RECT 28.510 170.360 28.650 175.140 ;
        RECT 28.450 170.040 28.710 170.360 ;
        RECT 27.990 164.940 28.250 165.260 ;
        RECT 28.450 161.200 28.710 161.520 ;
        RECT 27.990 158.140 28.250 158.460 ;
        RECT 26.610 156.780 26.870 157.100 ;
        RECT 27.070 148.960 27.330 149.280 ;
        RECT 26.610 137.060 26.870 137.380 ;
        RECT 26.150 134.680 26.410 135.000 ;
        RECT 26.210 129.560 26.350 134.680 ;
        RECT 26.150 129.240 26.410 129.560 ;
        RECT 26.670 108.580 26.810 137.060 ;
        RECT 27.130 134.660 27.270 148.960 ;
        RECT 27.530 142.500 27.790 142.820 ;
        RECT 27.070 134.340 27.330 134.660 ;
        RECT 27.590 124.800 27.730 142.500 ;
        RECT 28.050 127.180 28.190 158.140 ;
        RECT 28.510 156.760 28.650 161.200 ;
        RECT 28.450 156.440 28.710 156.760 ;
        RECT 28.450 155.420 28.710 155.740 ;
        RECT 28.510 132.280 28.650 155.420 ;
        RECT 28.970 152.000 29.110 177.860 ;
        RECT 29.430 154.380 29.570 182.620 ;
        RECT 29.890 175.800 30.030 198.940 ;
        RECT 30.350 191.690 30.490 198.940 ;
        RECT 30.810 192.460 30.950 201.040 ;
        RECT 32.650 199.940 32.790 202.680 ;
        RECT 32.590 199.850 32.850 199.940 ;
        RECT 32.190 199.710 32.850 199.850 ;
        RECT 31.210 198.940 31.470 199.260 ;
        RECT 30.750 192.140 31.010 192.460 ;
        RECT 30.350 191.550 30.950 191.690 ;
        RECT 30.290 190.780 30.550 191.100 ;
        RECT 29.830 175.480 30.090 175.800 ;
        RECT 29.830 172.420 30.090 172.740 ;
        RECT 29.890 167.210 30.030 172.420 ;
        RECT 30.350 170.360 30.490 190.780 ;
        RECT 30.810 176.480 30.950 191.550 ;
        RECT 31.270 187.020 31.410 198.940 ;
        RECT 32.190 197.900 32.330 199.710 ;
        RECT 32.590 199.620 32.850 199.710 ;
        RECT 34.890 199.620 35.150 199.940 ;
        RECT 36.270 199.620 36.530 199.940 ;
        RECT 38.110 199.620 38.370 199.940 ;
        RECT 32.510 198.405 34.390 198.775 ;
        RECT 32.130 197.580 32.390 197.900 ;
        RECT 33.510 197.240 33.770 197.560 ;
        RECT 31.670 196.900 31.930 197.220 ;
        RECT 31.730 195.520 31.870 196.900 ;
        RECT 32.130 196.220 32.390 196.540 ;
        RECT 31.670 195.200 31.930 195.520 ;
        RECT 32.190 189.060 32.330 196.220 ;
        RECT 33.040 194.665 33.320 195.035 ;
        RECT 33.570 194.840 33.710 197.240 ;
        RECT 33.970 196.395 34.230 196.540 ;
        RECT 33.960 196.025 34.240 196.395 ;
        RECT 33.050 194.520 33.310 194.665 ;
        RECT 33.510 194.520 33.770 194.840 ;
        RECT 32.510 192.965 34.390 193.335 ;
        RECT 33.050 190.780 33.310 191.100 ;
        RECT 33.110 189.400 33.250 190.780 ;
        RECT 32.590 189.080 32.850 189.400 ;
        RECT 33.050 189.080 33.310 189.400 ;
        RECT 31.670 188.740 31.930 189.060 ;
        RECT 32.130 188.740 32.390 189.060 ;
        RECT 31.210 186.700 31.470 187.020 ;
        RECT 31.210 183.640 31.470 183.960 ;
        RECT 30.750 176.160 31.010 176.480 ;
        RECT 31.270 175.880 31.410 183.640 ;
        RECT 30.810 175.740 31.410 175.880 ;
        RECT 30.290 170.040 30.550 170.360 ;
        RECT 30.290 167.210 30.550 167.300 ;
        RECT 29.890 167.070 30.550 167.210 ;
        RECT 30.290 166.980 30.550 167.070 ;
        RECT 29.830 166.300 30.090 166.620 ;
        RECT 29.890 165.600 30.030 166.300 ;
        RECT 29.830 165.280 30.090 165.600 ;
        RECT 30.350 161.860 30.490 166.980 ;
        RECT 29.830 161.540 30.090 161.860 ;
        RECT 30.290 161.540 30.550 161.860 ;
        RECT 29.890 156.420 30.030 161.540 ;
        RECT 30.810 158.995 30.950 175.740 ;
        RECT 31.210 174.460 31.470 174.780 ;
        RECT 31.270 162.200 31.410 174.460 ;
        RECT 31.730 173.420 31.870 188.740 ;
        RECT 32.650 188.290 32.790 189.080 ;
        RECT 32.190 188.150 32.790 188.290 ;
        RECT 32.190 183.960 32.330 188.150 ;
        RECT 32.510 187.525 34.390 187.895 ;
        RECT 33.970 185.340 34.230 185.660 ;
        RECT 32.130 183.640 32.390 183.960 ;
        RECT 34.030 182.940 34.170 185.340 ;
        RECT 34.950 184.640 35.090 199.620 ;
        RECT 35.350 198.940 35.610 199.260 ;
        RECT 34.890 184.320 35.150 184.640 ;
        RECT 33.970 182.620 34.230 182.940 ;
        RECT 32.510 182.085 34.390 182.455 ;
        RECT 33.050 181.600 33.310 181.920 ;
        RECT 33.110 180.755 33.250 181.600 ;
        RECT 33.040 180.385 33.320 180.755 ;
        RECT 35.410 180.220 35.550 198.940 ;
        RECT 35.810 194.180 36.070 194.500 ;
        RECT 35.870 183.620 36.010 194.180 ;
        RECT 36.330 190.080 36.470 199.620 ;
        RECT 38.170 199.115 38.310 199.620 ;
        RECT 39.950 199.280 40.210 199.600 ;
        RECT 38.100 198.745 38.380 199.115 ;
        RECT 38.570 198.940 38.830 199.260 ;
        RECT 39.030 198.940 39.290 199.260 ;
        RECT 37.650 196.220 37.910 196.540 ;
        RECT 36.730 194.180 36.990 194.500 ;
        RECT 36.790 190.080 36.930 194.180 ;
        RECT 37.190 193.500 37.450 193.820 ;
        RECT 36.270 189.760 36.530 190.080 ;
        RECT 36.730 189.760 36.990 190.080 ;
        RECT 36.720 189.225 37.000 189.595 ;
        RECT 36.790 189.060 36.930 189.225 ;
        RECT 36.730 188.740 36.990 189.060 ;
        RECT 37.250 188.915 37.390 193.500 ;
        RECT 37.180 188.545 37.460 188.915 ;
        RECT 36.270 188.060 36.530 188.380 ;
        RECT 36.730 188.060 36.990 188.380 ;
        RECT 37.190 188.060 37.450 188.380 ;
        RECT 35.810 183.300 36.070 183.620 ;
        RECT 35.350 179.900 35.610 180.220 ;
        RECT 32.130 178.200 32.390 178.520 ;
        RECT 31.670 173.100 31.930 173.420 ;
        RECT 32.190 172.740 32.330 178.200 ;
        RECT 35.350 177.860 35.610 178.180 ;
        RECT 34.890 177.180 35.150 177.500 ;
        RECT 32.510 176.645 34.390 177.015 ;
        RECT 34.430 172.760 34.690 173.080 ;
        RECT 32.130 172.420 32.390 172.740 ;
        RECT 34.490 172.595 34.630 172.760 ;
        RECT 34.420 172.225 34.700 172.595 ;
        RECT 32.510 171.205 34.390 171.575 ;
        RECT 34.950 171.040 35.090 177.180 ;
        RECT 34.890 170.720 35.150 171.040 ;
        RECT 31.670 167.320 31.930 167.640 ;
        RECT 32.590 167.320 32.850 167.640 ;
        RECT 31.210 161.880 31.470 162.200 ;
        RECT 31.210 160.860 31.470 161.180 ;
        RECT 30.740 158.625 31.020 158.995 ;
        RECT 30.290 158.140 30.550 158.460 ;
        RECT 30.750 158.140 31.010 158.460 ;
        RECT 30.350 157.440 30.490 158.140 ;
        RECT 30.290 157.120 30.550 157.440 ;
        RECT 29.830 156.100 30.090 156.420 ;
        RECT 29.370 154.060 29.630 154.380 ;
        RECT 28.910 151.680 29.170 152.000 ;
        RECT 28.910 151.000 29.170 151.320 ;
        RECT 28.970 145.880 29.110 151.000 ;
        RECT 29.370 147.940 29.630 148.260 ;
        RECT 28.910 145.560 29.170 145.880 ;
        RECT 28.910 144.540 29.170 144.860 ;
        RECT 28.450 131.960 28.710 132.280 ;
        RECT 28.970 129.220 29.110 144.540 ;
        RECT 29.430 132.960 29.570 147.940 ;
        RECT 29.890 147.580 30.030 156.100 ;
        RECT 30.280 153.865 30.560 154.235 ;
        RECT 30.350 150.980 30.490 153.865 ;
        RECT 30.290 150.660 30.550 150.980 ;
        RECT 30.290 149.980 30.550 150.300 ;
        RECT 29.830 147.260 30.090 147.580 ;
        RECT 29.830 142.840 30.090 143.160 ;
        RECT 29.370 132.640 29.630 132.960 ;
        RECT 28.910 128.900 29.170 129.220 ;
        RECT 29.370 128.900 29.630 129.220 ;
        RECT 27.990 126.860 28.250 127.180 ;
        RECT 29.430 126.840 29.570 128.900 ;
        RECT 29.890 127.520 30.030 142.840 ;
        RECT 30.350 142.140 30.490 149.980 ;
        RECT 30.290 141.820 30.550 142.140 ;
        RECT 30.290 139.100 30.550 139.420 ;
        RECT 29.830 127.200 30.090 127.520 ;
        RECT 30.350 126.840 30.490 139.100 ;
        RECT 30.810 126.840 30.950 158.140 ;
        RECT 31.270 157.100 31.410 160.860 ;
        RECT 31.210 156.780 31.470 157.100 ;
        RECT 31.200 155.905 31.480 156.275 ;
        RECT 31.270 152.880 31.410 155.905 ;
        RECT 31.730 154.720 31.870 167.320 ;
        RECT 32.130 166.640 32.390 166.960 ;
        RECT 32.190 158.460 32.330 166.640 ;
        RECT 32.650 166.620 32.790 167.320 ;
        RECT 34.950 166.960 35.090 170.720 ;
        RECT 34.890 166.640 35.150 166.960 ;
        RECT 32.590 166.300 32.850 166.620 ;
        RECT 32.510 165.765 34.390 166.135 ;
        RECT 32.590 165.280 32.850 165.600 ;
        RECT 32.650 162.200 32.790 165.280 ;
        RECT 33.050 163.580 33.310 163.900 ;
        RECT 33.110 162.200 33.250 163.580 ;
        RECT 32.590 161.880 32.850 162.200 ;
        RECT 33.050 161.880 33.310 162.200 ;
        RECT 32.510 160.325 34.390 160.695 ;
        RECT 33.510 159.730 33.770 159.820 ;
        RECT 33.510 159.590 34.170 159.730 ;
        RECT 33.510 159.500 33.770 159.590 ;
        RECT 32.590 158.995 32.850 159.140 ;
        RECT 32.580 158.625 32.860 158.995 ;
        RECT 33.510 158.820 33.770 159.140 ;
        RECT 32.130 158.140 32.390 158.460 ;
        RECT 33.570 157.440 33.710 158.820 ;
        RECT 34.030 158.315 34.170 159.590 ;
        RECT 33.960 157.945 34.240 158.315 ;
        RECT 33.510 157.120 33.770 157.440 ;
        RECT 35.410 156.420 35.550 177.860 ;
        RECT 35.810 177.520 36.070 177.840 ;
        RECT 35.870 175.200 36.010 177.520 ;
        RECT 36.330 176.140 36.470 188.060 ;
        RECT 36.790 182.795 36.930 188.060 ;
        RECT 36.720 182.425 37.000 182.795 ;
        RECT 36.730 178.540 36.990 178.860 ;
        RECT 36.270 175.820 36.530 176.140 ;
        RECT 35.870 175.060 36.470 175.200 ;
        RECT 36.330 174.780 36.470 175.060 ;
        RECT 36.270 174.460 36.530 174.780 ;
        RECT 35.810 172.420 36.070 172.740 ;
        RECT 35.870 170.020 36.010 172.420 ;
        RECT 36.260 172.225 36.540 172.595 ;
        RECT 36.330 170.020 36.470 172.225 ;
        RECT 35.810 169.700 36.070 170.020 ;
        RECT 36.270 169.700 36.530 170.020 ;
        RECT 35.870 167.040 36.010 169.700 ;
        RECT 36.330 167.640 36.470 169.700 ;
        RECT 36.270 167.320 36.530 167.640 ;
        RECT 36.790 167.300 36.930 178.540 ;
        RECT 37.250 173.080 37.390 188.060 ;
        RECT 37.710 187.020 37.850 196.220 ;
        RECT 38.110 193.675 38.370 193.820 ;
        RECT 38.100 193.305 38.380 193.675 ;
        RECT 38.630 192.120 38.770 198.940 ;
        RECT 39.090 197.755 39.230 198.940 ;
        RECT 39.020 197.385 39.300 197.755 ;
        RECT 40.010 196.960 40.150 199.280 ;
        RECT 40.470 197.560 40.610 206.225 ;
        RECT 43.160 205.545 43.440 205.915 ;
        RECT 40.870 205.060 41.130 205.380 ;
        RECT 40.930 203.680 41.070 205.060 ;
        RECT 40.870 203.360 41.130 203.680 ;
        RECT 43.230 203.000 43.370 205.545 ;
        RECT 45.930 205.400 46.190 205.720 ;
        RECT 45.000 204.865 45.280 205.235 ;
        RECT 45.070 203.680 45.210 204.865 ;
        RECT 45.010 203.360 45.270 203.680 ;
        RECT 45.990 203.000 46.130 205.400 ;
        RECT 46.910 203.680 47.050 206.760 ;
        RECT 91.460 206.225 91.740 206.595 ;
        RECT 54.210 205.740 54.470 206.060 ;
        RECT 84.110 205.740 84.370 206.060 ;
        RECT 88.710 205.740 88.970 206.060 ;
        RECT 46.850 203.360 47.110 203.680 ;
        RECT 50.530 203.250 50.790 203.340 ;
        RECT 50.130 203.110 50.790 203.250 ;
        RECT 43.170 202.680 43.430 203.000 ;
        RECT 45.930 202.680 46.190 203.000 ;
        RECT 49.610 202.680 49.870 203.000 ;
        RECT 42.250 202.515 42.510 202.660 ;
        RECT 42.240 202.145 42.520 202.515 ;
        RECT 43.630 202.000 43.890 202.320 ;
        RECT 40.870 199.620 41.130 199.940 ;
        RECT 41.790 199.620 42.050 199.940 ;
        RECT 42.710 199.795 42.970 199.940 ;
        RECT 40.410 197.240 40.670 197.560 ;
        RECT 39.030 196.560 39.290 196.880 ;
        RECT 40.010 196.820 40.610 196.960 ;
        RECT 38.110 191.800 38.370 192.120 ;
        RECT 38.570 191.800 38.830 192.120 ;
        RECT 37.650 186.700 37.910 187.020 ;
        RECT 38.170 186.340 38.310 191.800 ;
        RECT 38.570 188.740 38.830 189.060 ;
        RECT 38.110 186.020 38.370 186.340 ;
        RECT 37.650 181.600 37.910 181.920 ;
        RECT 37.710 180.900 37.850 181.600 ;
        RECT 38.170 180.900 38.310 186.020 ;
        RECT 38.630 181.580 38.770 188.740 ;
        RECT 39.090 183.280 39.230 196.560 ;
        RECT 39.950 196.220 40.210 196.540 ;
        RECT 39.490 195.035 39.750 195.180 ;
        RECT 39.480 194.665 39.760 195.035 ;
        RECT 40.010 194.070 40.150 196.220 ;
        RECT 40.470 194.840 40.610 196.820 ;
        RECT 40.410 194.520 40.670 194.840 ;
        RECT 39.550 193.930 40.150 194.070 ;
        RECT 39.550 190.080 39.690 193.930 ;
        RECT 40.470 192.200 40.610 194.520 ;
        RECT 40.930 194.500 41.070 199.620 ;
        RECT 41.850 198.320 41.990 199.620 ;
        RECT 42.700 199.425 42.980 199.795 ;
        RECT 41.390 198.180 41.990 198.320 ;
        RECT 40.870 194.355 41.130 194.500 ;
        RECT 40.860 193.985 41.140 194.355 ;
        RECT 40.870 192.480 41.130 192.800 ;
        RECT 40.010 192.060 40.610 192.200 ;
        RECT 39.490 189.760 39.750 190.080 ;
        RECT 39.480 188.545 39.760 188.915 ;
        RECT 39.550 186.340 39.690 188.545 ;
        RECT 40.010 187.555 40.150 192.060 ;
        RECT 40.930 189.060 41.070 192.480 ;
        RECT 41.390 191.780 41.530 198.180 ;
        RECT 41.790 197.580 42.050 197.900 ;
        RECT 41.850 194.500 41.990 197.580 ;
        RECT 42.710 197.470 42.970 197.560 ;
        RECT 42.310 197.330 42.970 197.470 ;
        RECT 41.790 194.180 42.050 194.500 ;
        RECT 41.330 191.460 41.590 191.780 ;
        RECT 41.330 189.760 41.590 190.080 ;
        RECT 40.870 188.740 41.130 189.060 ;
        RECT 40.410 188.060 40.670 188.380 ;
        RECT 39.940 187.185 40.220 187.555 ;
        RECT 39.490 186.020 39.750 186.340 ;
        RECT 40.010 183.360 40.150 187.185 ;
        RECT 40.470 184.300 40.610 188.060 ;
        RECT 40.870 184.320 41.130 184.640 ;
        RECT 40.410 183.980 40.670 184.300 ;
        RECT 40.930 183.960 41.070 184.320 ;
        RECT 40.870 183.640 41.130 183.960 ;
        RECT 39.030 182.960 39.290 183.280 ;
        RECT 40.010 183.220 41.070 183.360 ;
        RECT 39.020 182.425 39.300 182.795 ;
        RECT 40.400 182.425 40.680 182.795 ;
        RECT 38.570 181.260 38.830 181.580 ;
        RECT 37.650 180.580 37.910 180.900 ;
        RECT 38.110 180.580 38.370 180.900 ;
        RECT 37.650 178.035 37.910 178.180 ;
        RECT 37.640 177.665 37.920 178.035 ;
        RECT 37.650 177.180 37.910 177.500 ;
        RECT 37.190 172.760 37.450 173.080 ;
        RECT 37.190 172.080 37.450 172.400 ;
        RECT 35.870 166.900 36.470 167.040 ;
        RECT 36.730 166.980 36.990 167.300 ;
        RECT 36.330 166.680 36.470 166.900 ;
        RECT 35.810 166.300 36.070 166.620 ;
        RECT 36.330 166.540 36.930 166.680 ;
        RECT 35.870 163.900 36.010 166.300 ;
        RECT 36.270 164.260 36.530 164.580 ;
        RECT 35.810 163.580 36.070 163.900 ;
        RECT 36.330 162.200 36.470 164.260 ;
        RECT 36.270 161.880 36.530 162.200 ;
        RECT 36.790 161.600 36.930 166.540 ;
        RECT 36.330 161.460 36.930 161.600 ;
        RECT 36.330 159.140 36.470 161.460 ;
        RECT 37.250 160.920 37.390 172.080 ;
        RECT 37.710 162.200 37.850 177.180 ;
        RECT 38.170 175.460 38.310 180.580 ;
        RECT 38.570 177.520 38.830 177.840 ;
        RECT 38.110 175.140 38.370 175.460 ;
        RECT 38.170 172.740 38.310 175.140 ;
        RECT 38.110 172.420 38.370 172.740 ;
        RECT 38.110 170.720 38.370 171.040 ;
        RECT 38.170 167.300 38.310 170.720 ;
        RECT 38.110 166.980 38.370 167.300 ;
        RECT 38.630 165.510 38.770 177.520 ;
        RECT 39.090 166.620 39.230 182.425 ;
        RECT 40.470 181.580 40.610 182.425 ;
        RECT 40.410 181.260 40.670 181.580 ;
        RECT 39.950 180.920 40.210 181.240 ;
        RECT 39.490 178.880 39.750 179.200 ;
        RECT 39.030 166.300 39.290 166.620 ;
        RECT 39.030 165.510 39.290 165.600 ;
        RECT 38.630 165.370 39.290 165.510 ;
        RECT 39.030 165.280 39.290 165.370 ;
        RECT 38.110 164.600 38.370 164.920 ;
        RECT 39.030 164.600 39.290 164.920 ;
        RECT 38.170 164.240 38.310 164.600 ;
        RECT 38.110 163.920 38.370 164.240 ;
        RECT 39.090 162.880 39.230 164.600 ;
        RECT 39.550 163.755 39.690 178.880 ;
        RECT 40.010 178.715 40.150 180.920 ;
        RECT 40.410 178.880 40.670 179.200 ;
        RECT 39.940 178.345 40.220 178.715 ;
        RECT 40.470 178.180 40.610 178.880 ;
        RECT 40.930 178.180 41.070 183.220 ;
        RECT 39.940 177.665 40.220 178.035 ;
        RECT 40.410 177.860 40.670 178.180 ;
        RECT 40.870 177.860 41.130 178.180 ;
        RECT 39.950 177.520 40.210 177.665 ;
        RECT 41.390 177.500 41.530 189.760 ;
        RECT 41.850 187.360 41.990 194.180 ;
        RECT 42.310 192.800 42.450 197.330 ;
        RECT 42.710 197.240 42.970 197.330 ;
        RECT 43.170 197.240 43.430 197.560 ;
        RECT 43.230 194.240 43.370 197.240 ;
        RECT 42.770 194.100 43.370 194.240 ;
        RECT 42.250 192.480 42.510 192.800 ;
        RECT 42.250 191.800 42.510 192.120 ;
        RECT 41.790 187.040 42.050 187.360 ;
        RECT 42.310 184.640 42.450 191.800 ;
        RECT 42.770 189.060 42.910 194.100 ;
        RECT 43.170 193.500 43.430 193.820 ;
        RECT 43.230 192.800 43.370 193.500 ;
        RECT 43.170 192.480 43.430 192.800 ;
        RECT 43.690 189.480 43.830 202.000 ;
        RECT 47.510 201.125 49.390 201.495 ;
        RECT 47.310 200.300 47.570 200.620 ;
        RECT 47.370 199.940 47.510 200.300 ;
        RECT 44.090 199.620 44.350 199.940 ;
        RECT 47.310 199.620 47.570 199.940 ;
        RECT 49.150 199.620 49.410 199.940 ;
        RECT 49.670 199.795 49.810 202.680 ;
        RECT 50.130 201.980 50.270 203.110 ;
        RECT 50.530 203.020 50.790 203.110 ;
        RECT 51.450 202.680 51.710 203.000 ;
        RECT 50.070 201.660 50.330 201.980 ;
        RECT 50.530 201.660 50.790 201.980 ;
        RECT 50.990 201.660 51.250 201.980 ;
        RECT 50.590 200.475 50.730 201.660 ;
        RECT 50.520 200.105 50.800 200.475 ;
        RECT 44.150 196.880 44.290 199.620 ;
        RECT 45.010 198.940 45.270 199.260 ;
        RECT 49.210 199.170 49.350 199.620 ;
        RECT 49.600 199.425 49.880 199.795 ;
        RECT 50.070 199.280 50.330 199.600 ;
        RECT 49.210 199.030 49.810 199.170 ;
        RECT 44.550 197.075 44.810 197.220 ;
        RECT 44.090 196.560 44.350 196.880 ;
        RECT 44.540 196.705 44.820 197.075 ;
        RECT 44.080 194.665 44.360 195.035 ;
        RECT 44.150 194.160 44.290 194.665 ;
        RECT 44.090 193.840 44.350 194.160 ;
        RECT 44.550 193.840 44.810 194.160 ;
        RECT 44.610 191.440 44.750 193.840 ;
        RECT 44.550 191.120 44.810 191.440 ;
        RECT 43.230 189.340 43.830 189.480 ;
        RECT 44.090 189.420 44.350 189.740 ;
        RECT 42.710 188.740 42.970 189.060 ;
        RECT 42.250 184.320 42.510 184.640 ;
        RECT 41.790 181.600 42.050 181.920 ;
        RECT 41.330 177.355 41.590 177.500 ;
        RECT 41.320 176.985 41.600 177.355 ;
        RECT 40.860 175.625 41.140 175.995 ;
        RECT 39.950 174.460 40.210 174.780 ;
        RECT 40.010 172.060 40.150 174.460 ;
        RECT 40.410 172.420 40.670 172.740 ;
        RECT 39.950 171.740 40.210 172.060 ;
        RECT 39.480 163.385 39.760 163.755 ;
        RECT 39.030 162.560 39.290 162.880 ;
        RECT 39.490 162.560 39.750 162.880 ;
        RECT 37.650 161.880 37.910 162.200 ;
        RECT 39.030 161.880 39.290 162.200 ;
        RECT 36.790 160.780 37.390 160.920 ;
        RECT 36.270 158.820 36.530 159.140 ;
        RECT 36.790 157.440 36.930 160.780 ;
        RECT 38.560 159.985 38.840 160.355 ;
        RECT 39.090 160.160 39.230 161.880 ;
        RECT 38.100 159.305 38.380 159.675 ;
        RECT 38.630 159.480 38.770 159.985 ;
        RECT 39.030 159.840 39.290 160.160 ;
        RECT 37.650 158.820 37.910 159.140 ;
        RECT 37.190 158.140 37.450 158.460 ;
        RECT 36.730 157.120 36.990 157.440 ;
        RECT 35.810 156.440 36.070 156.760 ;
        RECT 34.890 156.100 35.150 156.420 ;
        RECT 35.350 156.100 35.610 156.420 ;
        RECT 32.130 155.760 32.390 156.080 ;
        RECT 31.670 154.400 31.930 154.720 ;
        RECT 32.190 153.020 32.330 155.760 ;
        RECT 32.510 154.885 34.390 155.255 ;
        RECT 33.050 154.400 33.310 154.720 ;
        RECT 31.270 152.740 31.870 152.880 ;
        RECT 31.210 149.980 31.470 150.300 ;
        RECT 31.270 146.560 31.410 149.980 ;
        RECT 31.730 148.940 31.870 152.740 ;
        RECT 32.130 152.700 32.390 153.020 ;
        RECT 32.190 150.980 32.330 152.700 ;
        RECT 32.130 150.660 32.390 150.980 ;
        RECT 33.110 150.210 33.250 154.400 ;
        RECT 32.190 150.070 33.250 150.210 ;
        RECT 31.670 148.620 31.930 148.940 ;
        RECT 31.210 146.240 31.470 146.560 ;
        RECT 32.190 145.540 32.330 150.070 ;
        RECT 32.510 149.445 34.390 149.815 ;
        RECT 33.970 147.260 34.230 147.580 ;
        RECT 34.030 145.880 34.170 147.260 ;
        RECT 34.950 146.560 35.090 156.100 ;
        RECT 35.870 154.720 36.010 156.440 ;
        RECT 37.250 156.420 37.390 158.140 ;
        RECT 36.270 156.100 36.530 156.420 ;
        RECT 37.190 156.100 37.450 156.420 ;
        RECT 35.810 154.400 36.070 154.720 ;
        RECT 36.330 154.120 36.470 156.100 ;
        RECT 35.870 154.040 36.470 154.120 ;
        RECT 37.190 154.060 37.450 154.380 ;
        RECT 35.810 153.980 36.470 154.040 ;
        RECT 35.810 153.720 36.070 153.980 ;
        RECT 36.270 152.880 36.530 153.020 ;
        RECT 35.870 152.740 36.530 152.880 ;
        RECT 35.870 150.980 36.010 152.740 ;
        RECT 36.270 152.700 36.530 152.740 ;
        RECT 37.250 151.320 37.390 154.060 ;
        RECT 37.710 154.040 37.850 158.820 ;
        RECT 38.170 156.760 38.310 159.305 ;
        RECT 38.570 159.160 38.830 159.480 ;
        RECT 39.030 159.390 39.290 159.480 ;
        RECT 39.550 159.390 39.690 162.560 ;
        RECT 40.010 159.480 40.150 171.740 ;
        RECT 40.470 169.340 40.610 172.420 ;
        RECT 40.930 171.040 41.070 175.625 ;
        RECT 41.330 171.740 41.590 172.060 ;
        RECT 40.870 170.720 41.130 171.040 ;
        RECT 40.410 169.020 40.670 169.340 ;
        RECT 40.470 164.580 40.610 169.020 ;
        RECT 40.870 168.230 41.130 168.320 ;
        RECT 41.390 168.230 41.530 171.740 ;
        RECT 40.870 168.090 41.530 168.230 ;
        RECT 40.870 168.000 41.130 168.090 ;
        RECT 41.330 167.550 41.590 167.640 ;
        RECT 40.930 167.410 41.590 167.550 ;
        RECT 40.410 164.260 40.670 164.580 ;
        RECT 40.400 163.385 40.680 163.755 ;
        RECT 39.030 159.250 39.690 159.390 ;
        RECT 39.030 159.160 39.290 159.250 ;
        RECT 39.950 159.160 40.210 159.480 ;
        RECT 38.110 156.440 38.370 156.760 ;
        RECT 39.950 156.100 40.210 156.420 ;
        RECT 38.110 155.650 38.370 155.740 ;
        RECT 38.110 155.510 38.770 155.650 ;
        RECT 40.010 155.595 40.150 156.100 ;
        RECT 38.110 155.420 38.370 155.510 ;
        RECT 37.650 153.720 37.910 154.040 ;
        RECT 37.190 151.000 37.450 151.320 ;
        RECT 35.810 150.660 36.070 150.980 ;
        RECT 36.270 150.660 36.530 150.980 ;
        RECT 36.330 148.260 36.470 150.660 ;
        RECT 36.270 147.940 36.530 148.260 ;
        RECT 34.890 146.240 35.150 146.560 ;
        RECT 37.250 145.880 37.390 151.000 ;
        RECT 37.710 148.260 37.850 153.720 ;
        RECT 38.110 150.660 38.370 150.980 ;
        RECT 37.650 147.940 37.910 148.260 ;
        RECT 33.970 145.560 34.230 145.880 ;
        RECT 34.890 145.560 35.150 145.880 ;
        RECT 37.190 145.560 37.450 145.880 ;
        RECT 31.670 145.220 31.930 145.540 ;
        RECT 32.130 145.220 32.390 145.540 ;
        RECT 31.210 141.820 31.470 142.140 ;
        RECT 31.270 134.660 31.410 141.820 ;
        RECT 31.730 140.100 31.870 145.220 ;
        RECT 32.190 143.840 32.330 145.220 ;
        RECT 32.510 144.005 34.390 144.375 ;
        RECT 32.130 143.520 32.390 143.840 ;
        RECT 32.190 140.440 32.330 143.520 ;
        RECT 33.050 141.820 33.310 142.140 ;
        RECT 32.590 140.460 32.850 140.780 ;
        RECT 32.130 140.120 32.390 140.440 ;
        RECT 31.670 139.780 31.930 140.100 ;
        RECT 32.650 139.840 32.790 140.460 ;
        RECT 33.110 140.100 33.250 141.820 ;
        RECT 34.950 140.780 35.090 145.560 ;
        RECT 37.650 144.540 37.910 144.860 ;
        RECT 36.270 143.520 36.530 143.840 ;
        RECT 34.890 140.460 35.150 140.780 ;
        RECT 32.190 139.700 32.790 139.840 ;
        RECT 33.050 139.780 33.310 140.100 ;
        RECT 31.670 137.400 31.930 137.720 ;
        RECT 31.210 134.340 31.470 134.660 ;
        RECT 31.210 131.960 31.470 132.280 ;
        RECT 29.370 126.520 29.630 126.840 ;
        RECT 30.290 126.520 30.550 126.840 ;
        RECT 30.750 126.520 31.010 126.840 ;
        RECT 27.530 124.480 27.790 124.800 ;
        RECT 29.430 123.780 29.570 126.520 ;
        RECT 29.370 123.460 29.630 123.780 ;
        RECT 31.270 108.580 31.410 131.960 ;
        RECT 31.730 124.800 31.870 137.400 ;
        RECT 32.190 135.195 32.330 139.700 ;
        RECT 32.510 138.565 34.390 138.935 ;
        RECT 35.810 137.740 36.070 138.060 ;
        RECT 34.430 136.380 34.690 136.700 ;
        RECT 34.490 135.340 34.630 136.380 ;
        RECT 32.120 134.825 32.400 135.195 ;
        RECT 34.430 135.020 34.690 135.340 ;
        RECT 32.130 134.680 32.390 134.825 ;
        RECT 35.350 134.680 35.610 135.000 ;
        RECT 32.510 133.125 34.390 133.495 ;
        RECT 33.970 132.640 34.230 132.960 ;
        RECT 32.130 132.300 32.390 132.620 ;
        RECT 31.670 124.480 31.930 124.800 ;
        RECT 32.190 124.120 32.330 132.300 ;
        RECT 34.030 129.220 34.170 132.640 ;
        RECT 35.410 129.560 35.550 134.680 ;
        RECT 35.350 129.240 35.610 129.560 ;
        RECT 33.970 128.900 34.230 129.220 ;
        RECT 32.510 127.685 34.390 128.055 ;
        RECT 35.870 126.160 36.010 137.740 ;
        RECT 36.330 127.520 36.470 143.520 ;
        RECT 36.730 142.500 36.990 142.820 ;
        RECT 36.790 129.900 36.930 142.500 ;
        RECT 37.710 141.120 37.850 144.540 ;
        RECT 37.650 140.800 37.910 141.120 ;
        RECT 37.190 140.460 37.450 140.780 ;
        RECT 36.730 129.580 36.990 129.900 ;
        RECT 36.270 127.200 36.530 127.520 ;
        RECT 37.250 127.180 37.390 140.460 ;
        RECT 37.650 138.080 37.910 138.400 ;
        RECT 37.710 130.240 37.850 138.080 ;
        RECT 38.170 136.700 38.310 150.660 ;
        RECT 38.630 140.780 38.770 155.510 ;
        RECT 39.940 155.225 40.220 155.595 ;
        RECT 39.490 154.400 39.750 154.720 ;
        RECT 39.030 153.380 39.290 153.700 ;
        RECT 39.090 145.200 39.230 153.380 ;
        RECT 39.550 153.020 39.690 154.400 ;
        RECT 39.490 152.700 39.750 153.020 ;
        RECT 39.950 150.550 40.210 150.640 ;
        RECT 40.470 150.550 40.610 163.385 ;
        RECT 40.930 156.760 41.070 167.410 ;
        RECT 41.330 167.320 41.590 167.410 ;
        RECT 41.330 164.940 41.590 165.260 ;
        RECT 41.850 165.000 41.990 181.600 ;
        RECT 42.250 177.860 42.510 178.180 ;
        RECT 42.310 173.760 42.450 177.860 ;
        RECT 42.710 177.180 42.970 177.500 ;
        RECT 42.250 173.440 42.510 173.760 ;
        RECT 42.250 172.080 42.510 172.400 ;
        RECT 42.310 167.040 42.450 172.080 ;
        RECT 42.770 171.040 42.910 177.180 ;
        RECT 43.230 176.140 43.370 189.340 ;
        RECT 43.630 186.020 43.890 186.340 ;
        RECT 43.690 180.900 43.830 186.020 ;
        RECT 44.150 184.155 44.290 189.420 ;
        RECT 44.540 189.225 44.820 189.595 ;
        RECT 44.610 186.250 44.750 189.225 ;
        RECT 45.070 189.060 45.210 198.940 ;
        RECT 46.390 197.240 46.650 197.560 ;
        RECT 45.930 196.900 46.190 197.220 ;
        RECT 45.470 196.220 45.730 196.540 ;
        RECT 45.530 191.635 45.670 196.220 ;
        RECT 45.460 191.265 45.740 191.635 ;
        RECT 45.470 190.780 45.730 191.100 ;
        RECT 45.010 188.740 45.270 189.060 ;
        RECT 45.530 187.020 45.670 190.780 ;
        RECT 45.990 187.020 46.130 196.900 ;
        RECT 45.470 186.700 45.730 187.020 ;
        RECT 45.930 186.700 46.190 187.020 ;
        RECT 44.610 186.110 45.670 186.250 ;
        RECT 44.550 185.340 44.810 185.660 ;
        RECT 44.080 183.785 44.360 184.155 ;
        RECT 44.610 181.920 44.750 185.340 ;
        RECT 44.550 181.600 44.810 181.920 ;
        RECT 43.630 180.580 43.890 180.900 ;
        RECT 45.010 180.580 45.270 180.900 ;
        RECT 43.630 177.860 43.890 178.180 ;
        RECT 44.550 178.090 44.810 178.180 ;
        RECT 44.150 177.950 44.810 178.090 ;
        RECT 43.170 175.820 43.430 176.140 ;
        RECT 43.690 175.200 43.830 177.860 ;
        RECT 43.230 175.060 43.830 175.200 ;
        RECT 43.230 174.780 43.370 175.060 ;
        RECT 43.170 174.460 43.430 174.780 ;
        RECT 42.710 170.720 42.970 171.040 ;
        RECT 42.710 169.020 42.970 169.340 ;
        RECT 42.770 167.640 42.910 169.020 ;
        RECT 42.710 167.320 42.970 167.640 ;
        RECT 42.310 166.900 42.910 167.040 ;
        RECT 42.250 166.300 42.510 166.620 ;
        RECT 42.310 165.600 42.450 166.300 ;
        RECT 42.250 165.280 42.510 165.600 ;
        RECT 40.870 156.440 41.130 156.760 ;
        RECT 41.390 156.420 41.530 164.940 ;
        RECT 41.850 164.860 42.450 165.000 ;
        RECT 41.790 162.560 42.050 162.880 ;
        RECT 41.850 159.480 41.990 162.560 ;
        RECT 42.310 161.520 42.450 164.860 ;
        RECT 42.250 161.200 42.510 161.520 ;
        RECT 42.250 159.675 42.510 159.820 ;
        RECT 41.790 159.160 42.050 159.480 ;
        RECT 42.240 159.305 42.520 159.675 ;
        RECT 41.790 157.120 42.050 157.440 ;
        RECT 41.330 156.100 41.590 156.420 ;
        RECT 40.870 152.700 41.130 153.020 ;
        RECT 39.950 150.410 40.610 150.550 ;
        RECT 39.950 150.320 40.210 150.410 ;
        RECT 40.930 149.280 41.070 152.700 ;
        RECT 41.850 149.280 41.990 157.120 ;
        RECT 42.770 156.840 42.910 166.900 ;
        RECT 43.230 160.355 43.370 174.460 ;
        RECT 43.620 174.265 43.900 174.635 ;
        RECT 43.160 159.985 43.440 160.355 ;
        RECT 43.690 158.460 43.830 174.265 ;
        RECT 44.150 167.980 44.290 177.950 ;
        RECT 44.550 177.860 44.810 177.950 ;
        RECT 44.550 177.180 44.810 177.500 ;
        RECT 44.090 167.660 44.350 167.980 ;
        RECT 44.610 167.300 44.750 177.180 ;
        RECT 44.550 166.980 44.810 167.300 ;
        RECT 44.610 166.620 44.750 166.980 ;
        RECT 44.550 166.300 44.810 166.620 ;
        RECT 45.070 165.260 45.210 180.580 ;
        RECT 45.530 169.680 45.670 186.110 ;
        RECT 45.990 183.620 46.130 186.700 ;
        RECT 46.450 184.640 46.590 197.240 ;
        RECT 46.850 196.220 47.110 196.540 ;
        RECT 46.910 192.460 47.050 196.220 ;
        RECT 47.510 195.685 49.390 196.055 ;
        RECT 46.850 192.140 47.110 192.460 ;
        RECT 49.670 192.370 49.810 199.030 ;
        RECT 50.130 194.355 50.270 199.280 ;
        RECT 50.060 193.985 50.340 194.355 ;
        RECT 51.050 194.160 51.190 201.660 ;
        RECT 51.510 199.940 51.650 202.680 ;
        RECT 54.270 202.320 54.410 205.740 ;
        RECT 56.970 204.720 57.230 205.040 ;
        RECT 68.930 204.720 69.190 205.040 ;
        RECT 81.810 204.720 82.070 205.040 ;
        RECT 56.040 203.505 56.320 203.875 ;
        RECT 56.110 203.000 56.250 203.505 ;
        RECT 57.030 203.000 57.170 204.720 ;
        RECT 68.990 204.440 69.130 204.720 ;
        RECT 68.990 204.300 70.050 204.440 ;
        RECT 61.560 203.505 61.840 203.875 ;
        RECT 62.510 203.845 64.390 204.215 ;
        RECT 63.410 203.590 63.670 203.680 ;
        RECT 61.570 203.360 61.830 203.505 ;
        RECT 63.410 203.450 64.990 203.590 ;
        RECT 63.410 203.360 63.670 203.450 ;
        RECT 57.890 203.020 58.150 203.340 ;
        RECT 54.670 202.680 54.930 203.000 ;
        RECT 56.050 202.680 56.310 203.000 ;
        RECT 56.970 202.680 57.230 203.000 ;
        RECT 52.830 202.230 53.090 202.320 ;
        RECT 52.830 202.090 53.490 202.230 ;
        RECT 52.830 202.000 53.090 202.090 ;
        RECT 51.450 199.620 51.710 199.940 ;
        RECT 51.910 199.620 52.170 199.940 ;
        RECT 51.450 197.920 51.710 198.240 ;
        RECT 51.510 195.520 51.650 197.920 ;
        RECT 51.450 195.200 51.710 195.520 ;
        RECT 51.440 194.665 51.720 195.035 ;
        RECT 50.990 193.840 51.250 194.160 ;
        RECT 50.520 193.305 50.800 193.675 ;
        RECT 50.070 192.370 50.330 192.460 ;
        RECT 49.670 192.230 50.330 192.370 ;
        RECT 50.070 192.140 50.330 192.230 ;
        RECT 46.850 191.460 47.110 191.780 ;
        RECT 46.910 186.250 47.050 191.460 ;
        RECT 47.510 190.245 49.390 190.615 ;
        RECT 48.690 189.080 48.950 189.400 ;
        RECT 48.750 188.630 48.890 189.080 ;
        RECT 49.150 188.630 49.410 188.720 ;
        RECT 48.750 188.490 49.410 188.630 ;
        RECT 49.150 188.400 49.410 188.490 ;
        RECT 47.770 186.250 48.030 186.340 ;
        RECT 46.910 186.110 48.030 186.250 ;
        RECT 46.390 184.320 46.650 184.640 ;
        RECT 45.930 183.300 46.190 183.620 ;
        RECT 46.450 179.200 46.590 184.320 ;
        RECT 46.910 183.960 47.050 186.110 ;
        RECT 47.770 186.020 48.030 186.110 ;
        RECT 50.130 186.000 50.270 192.140 ;
        RECT 50.590 189.400 50.730 193.305 ;
        RECT 51.510 192.800 51.650 194.665 ;
        RECT 51.450 192.480 51.710 192.800 ;
        RECT 51.450 190.780 51.710 191.100 ;
        RECT 50.530 189.080 50.790 189.400 ;
        RECT 50.530 188.400 50.790 188.720 ;
        RECT 49.610 185.680 49.870 186.000 ;
        RECT 50.070 185.680 50.330 186.000 ;
        RECT 47.510 184.805 49.390 185.175 ;
        RECT 46.850 183.640 47.110 183.960 ;
        RECT 47.770 182.850 48.030 182.940 ;
        RECT 47.370 182.710 48.030 182.850 ;
        RECT 47.370 181.240 47.510 182.710 ;
        RECT 47.770 182.620 48.030 182.710 ;
        RECT 49.670 181.920 49.810 185.680 ;
        RECT 50.060 183.785 50.340 184.155 ;
        RECT 49.610 181.600 49.870 181.920 ;
        RECT 47.310 180.920 47.570 181.240 ;
        RECT 48.230 180.920 48.490 181.240 ;
        RECT 49.610 180.920 49.870 181.240 ;
        RECT 48.290 180.640 48.430 180.920 ;
        RECT 46.910 180.500 48.430 180.640 ;
        RECT 46.390 178.880 46.650 179.200 ;
        RECT 46.910 178.715 47.050 180.500 ;
        RECT 47.510 179.365 49.390 179.735 ;
        RECT 46.840 178.600 47.120 178.715 ;
        RECT 45.930 178.200 46.190 178.520 ;
        RECT 46.450 178.460 47.120 178.600 ;
        RECT 45.990 176.140 46.130 178.200 ;
        RECT 45.930 175.820 46.190 176.140 ;
        RECT 46.450 171.800 46.590 178.460 ;
        RECT 46.840 178.345 47.120 178.460 ;
        RECT 46.850 177.180 47.110 177.500 ;
        RECT 45.990 171.660 46.590 171.800 ;
        RECT 46.910 171.800 47.050 177.180 ;
        RECT 47.510 173.925 49.390 174.295 ;
        RECT 47.300 172.905 47.580 173.275 ;
        RECT 47.370 172.740 47.510 172.905 ;
        RECT 47.310 172.420 47.570 172.740 ;
        RECT 46.910 171.660 47.510 171.800 ;
        RECT 45.470 169.360 45.730 169.680 ;
        RECT 45.010 164.940 45.270 165.260 ;
        RECT 44.090 164.600 44.350 164.920 ;
        RECT 44.150 161.180 44.290 164.600 ;
        RECT 45.010 163.920 45.270 164.240 ;
        RECT 44.540 161.345 44.820 161.715 ;
        RECT 44.090 160.860 44.350 161.180 ;
        RECT 44.150 159.480 44.290 160.860 ;
        RECT 44.610 159.675 44.750 161.345 ;
        RECT 44.090 159.160 44.350 159.480 ;
        RECT 44.540 159.305 44.820 159.675 ;
        RECT 44.550 159.160 44.810 159.305 ;
        RECT 43.630 158.140 43.890 158.460 ;
        RECT 44.540 157.945 44.820 158.315 ;
        RECT 44.610 157.440 44.750 157.945 ;
        RECT 44.090 157.120 44.350 157.440 ;
        RECT 44.550 157.120 44.810 157.440 ;
        RECT 42.770 156.700 43.370 156.840 ;
        RECT 42.710 156.100 42.970 156.420 ;
        RECT 42.250 153.720 42.510 154.040 ;
        RECT 40.870 148.960 41.130 149.280 ;
        RECT 41.790 148.960 42.050 149.280 ;
        RECT 39.950 148.620 40.210 148.940 ;
        RECT 40.010 146.560 40.150 148.620 ;
        RECT 40.410 147.260 40.670 147.580 ;
        RECT 39.950 146.240 40.210 146.560 ;
        RECT 39.030 144.880 39.290 145.200 ;
        RECT 40.470 142.820 40.610 147.260 ;
        RECT 40.410 142.500 40.670 142.820 ;
        RECT 38.570 140.460 38.830 140.780 ;
        RECT 40.470 140.100 40.610 142.500 ;
        RECT 42.310 141.120 42.450 153.720 ;
        RECT 42.770 153.360 42.910 156.100 ;
        RECT 43.230 154.720 43.370 156.700 ;
        RECT 43.630 156.440 43.890 156.760 ;
        RECT 43.690 156.275 43.830 156.440 ;
        RECT 43.620 155.905 43.900 156.275 ;
        RECT 43.630 155.420 43.890 155.740 ;
        RECT 43.170 154.400 43.430 154.720 ;
        RECT 42.710 153.040 42.970 153.360 ;
        RECT 43.230 152.880 43.370 154.400 ;
        RECT 42.770 152.740 43.370 152.880 ;
        RECT 42.770 151.320 42.910 152.740 ;
        RECT 42.710 151.000 42.970 151.320 ;
        RECT 42.710 144.880 42.970 145.200 ;
        RECT 42.250 140.800 42.510 141.120 ;
        RECT 42.250 140.120 42.510 140.440 ;
        RECT 40.410 139.780 40.670 140.100 ;
        RECT 40.470 137.380 40.610 139.780 ;
        RECT 40.410 137.060 40.670 137.380 ;
        RECT 40.870 137.060 41.130 137.380 ;
        RECT 38.110 136.380 38.370 136.700 ;
        RECT 40.470 134.660 40.610 137.060 ;
        RECT 38.110 134.340 38.370 134.660 ;
        RECT 38.570 134.340 38.830 134.660 ;
        RECT 40.410 134.340 40.670 134.660 ;
        RECT 38.170 132.960 38.310 134.340 ;
        RECT 38.110 132.640 38.370 132.960 ;
        RECT 38.630 132.475 38.770 134.340 ;
        RECT 38.560 132.105 38.840 132.475 ;
        RECT 40.470 131.940 40.610 134.340 ;
        RECT 38.570 131.620 38.830 131.940 ;
        RECT 40.410 131.620 40.670 131.940 ;
        RECT 38.110 130.940 38.370 131.260 ;
        RECT 37.650 129.920 37.910 130.240 ;
        RECT 38.170 129.220 38.310 130.940 ;
        RECT 38.110 128.900 38.370 129.220 ;
        RECT 37.190 126.860 37.450 127.180 ;
        RECT 35.810 125.840 36.070 126.160 ;
        RECT 35.350 125.500 35.610 125.820 ;
        RECT 32.130 123.800 32.390 124.120 ;
        RECT 34.890 122.780 35.150 123.100 ;
        RECT 32.510 122.245 34.390 122.615 ;
        RECT 34.950 121.740 35.090 122.780 ;
        RECT 35.410 122.080 35.550 125.500 ;
        RECT 38.630 124.800 38.770 131.620 ;
        RECT 39.030 128.560 39.290 128.880 ;
        RECT 39.490 128.560 39.750 128.880 ;
        RECT 39.090 127.520 39.230 128.560 ;
        RECT 39.030 127.200 39.290 127.520 ;
        RECT 39.550 124.800 39.690 128.560 ;
        RECT 40.470 126.500 40.610 131.620 ;
        RECT 40.930 129.900 41.070 137.060 ;
        RECT 42.310 136.700 42.450 140.120 ;
        RECT 42.250 136.380 42.510 136.700 ;
        RECT 41.780 134.825 42.060 135.195 ;
        RECT 41.330 134.340 41.590 134.660 ;
        RECT 41.390 129.900 41.530 134.340 ;
        RECT 41.850 131.940 41.990 134.825 ;
        RECT 42.310 132.960 42.450 136.380 ;
        RECT 42.770 135.680 42.910 144.880 ;
        RECT 43.690 142.140 43.830 155.420 ;
        RECT 44.150 154.720 44.290 157.120 ;
        RECT 44.550 156.440 44.810 156.760 ;
        RECT 44.090 154.400 44.350 154.720 ;
        RECT 44.090 153.720 44.350 154.040 ;
        RECT 44.150 144.860 44.290 153.720 ;
        RECT 44.090 144.540 44.350 144.860 ;
        RECT 44.610 142.560 44.750 156.440 ;
        RECT 45.070 154.380 45.210 163.920 ;
        RECT 45.470 161.540 45.730 161.860 ;
        RECT 45.530 159.820 45.670 161.540 ;
        RECT 45.990 160.160 46.130 171.660 ;
        RECT 46.390 170.720 46.650 171.040 ;
        RECT 46.450 161.035 46.590 170.720 ;
        RECT 46.840 170.185 47.120 170.555 ;
        RECT 46.850 170.040 47.110 170.185 ;
        RECT 47.370 169.760 47.510 171.660 ;
        RECT 49.670 170.555 49.810 180.920 ;
        RECT 49.600 170.185 49.880 170.555 ;
        RECT 46.910 169.620 47.510 169.760 ;
        RECT 46.910 167.040 47.050 169.620 ;
        RECT 49.610 169.020 49.870 169.340 ;
        RECT 47.510 168.485 49.390 168.855 ;
        RECT 49.670 167.640 49.810 169.020 ;
        RECT 49.610 167.320 49.870 167.640 ;
        RECT 46.910 166.900 49.810 167.040 ;
        RECT 49.150 164.320 49.410 164.580 ;
        RECT 48.290 164.260 49.410 164.320 ;
        RECT 48.290 164.240 49.350 164.260 ;
        RECT 48.230 164.180 49.350 164.240 ;
        RECT 48.230 163.920 48.490 164.180 ;
        RECT 46.850 163.580 47.110 163.900 ;
        RECT 46.910 162.450 47.050 163.580 ;
        RECT 47.510 163.045 49.390 163.415 ;
        RECT 46.910 162.310 48.430 162.450 ;
        RECT 49.670 162.395 49.810 166.900 ;
        RECT 50.130 164.435 50.270 183.785 ;
        RECT 50.590 180.900 50.730 188.400 ;
        RECT 50.990 188.060 51.250 188.380 ;
        RECT 51.050 182.940 51.190 188.060 ;
        RECT 51.510 187.360 51.650 190.780 ;
        RECT 51.970 190.080 52.110 199.620 ;
        RECT 52.830 198.940 53.090 199.260 ;
        RECT 52.370 196.900 52.630 197.220 ;
        RECT 52.430 192.800 52.570 196.900 ;
        RECT 52.890 195.520 53.030 198.940 ;
        RECT 52.830 195.200 53.090 195.520 ;
        RECT 52.370 192.480 52.630 192.800 ;
        RECT 53.350 192.315 53.490 202.090 ;
        RECT 54.210 202.000 54.470 202.320 ;
        RECT 53.750 199.280 54.010 199.600 ;
        RECT 53.810 197.220 53.950 199.280 ;
        RECT 53.750 196.900 54.010 197.220 ;
        RECT 53.810 194.160 53.950 196.900 ;
        RECT 54.210 196.220 54.470 196.540 ;
        RECT 53.750 193.840 54.010 194.160 ;
        RECT 53.280 191.945 53.560 192.315 ;
        RECT 53.810 191.440 53.950 193.840 ;
        RECT 54.270 192.800 54.410 196.220 ;
        RECT 54.210 192.480 54.470 192.800 ;
        RECT 52.370 191.120 52.630 191.440 ;
        RECT 53.750 191.120 54.010 191.440 ;
        RECT 51.910 189.760 52.170 190.080 ;
        RECT 51.450 187.040 51.710 187.360 ;
        RECT 52.430 183.280 52.570 191.120 ;
        RECT 52.830 188.800 53.090 189.060 ;
        RECT 53.810 188.800 53.950 191.120 ;
        RECT 52.830 188.740 53.950 188.800 ;
        RECT 52.890 188.660 53.950 188.740 ;
        RECT 52.830 185.340 53.090 185.660 ;
        RECT 52.890 183.960 53.030 185.340 ;
        RECT 52.830 183.640 53.090 183.960 ;
        RECT 53.810 183.360 53.950 188.660 ;
        RECT 54.730 186.875 54.870 202.680 ;
        RECT 56.510 202.000 56.770 202.320 ;
        RECT 56.570 200.280 56.710 202.000 ;
        RECT 57.430 201.660 57.690 201.980 ;
        RECT 56.970 200.640 57.230 200.960 ;
        RECT 55.590 199.960 55.850 200.280 ;
        RECT 56.510 199.960 56.770 200.280 ;
        RECT 55.650 199.260 55.790 199.960 ;
        RECT 55.590 198.940 55.850 199.260 ;
        RECT 55.130 197.920 55.390 198.240 ;
        RECT 55.190 192.800 55.330 197.920 ;
        RECT 55.590 197.580 55.850 197.900 ;
        RECT 55.130 192.480 55.390 192.800 ;
        RECT 55.190 191.100 55.330 192.480 ;
        RECT 55.130 190.780 55.390 191.100 ;
        RECT 55.650 189.060 55.790 197.580 ;
        RECT 57.030 194.160 57.170 200.640 ;
        RECT 57.490 199.600 57.630 201.660 ;
        RECT 57.950 200.475 58.090 203.020 ;
        RECT 61.110 202.680 61.370 203.000 ;
        RECT 58.810 202.000 59.070 202.320 ;
        RECT 58.350 201.660 58.610 201.980 ;
        RECT 57.880 200.105 58.160 200.475 ;
        RECT 57.430 199.280 57.690 199.600 ;
        RECT 58.410 197.900 58.550 201.660 ;
        RECT 58.870 201.180 59.010 202.000 ;
        RECT 58.870 201.040 59.470 201.180 ;
        RECT 59.330 198.240 59.470 201.040 ;
        RECT 58.810 197.920 59.070 198.240 ;
        RECT 59.270 197.920 59.530 198.240 ;
        RECT 58.350 197.580 58.610 197.900 ;
        RECT 57.430 194.520 57.690 194.840 ;
        RECT 56.970 193.840 57.230 194.160 ;
        RECT 57.490 192.880 57.630 194.520 ;
        RECT 58.870 193.820 59.010 197.920 ;
        RECT 58.810 193.500 59.070 193.820 ;
        RECT 56.570 192.740 57.630 192.880 ;
        RECT 56.570 192.460 56.710 192.740 ;
        RECT 56.510 192.140 56.770 192.460 ;
        RECT 56.510 191.460 56.770 191.780 ;
        RECT 58.350 191.460 58.610 191.780 ;
        RECT 56.570 189.400 56.710 191.460 ;
        RECT 56.050 189.080 56.310 189.400 ;
        RECT 56.510 189.080 56.770 189.400 ;
        RECT 55.590 188.740 55.850 189.060 ;
        RECT 55.130 188.060 55.390 188.380 ;
        RECT 54.660 186.505 54.940 186.875 ;
        RECT 54.670 186.020 54.930 186.340 ;
        RECT 54.210 185.680 54.470 186.000 ;
        RECT 54.270 184.040 54.410 185.680 ;
        RECT 54.730 184.640 54.870 186.020 ;
        RECT 54.670 184.320 54.930 184.640 ;
        RECT 54.270 183.900 54.870 184.040 ;
        RECT 54.210 183.360 54.470 183.620 ;
        RECT 53.810 183.300 54.470 183.360 ;
        RECT 52.370 182.960 52.630 183.280 ;
        RECT 53.810 183.220 54.410 183.300 ;
        RECT 50.990 182.620 51.250 182.940 ;
        RECT 51.440 182.425 51.720 182.795 ;
        RECT 50.530 180.580 50.790 180.900 ;
        RECT 50.590 179.200 50.730 180.580 ;
        RECT 50.530 178.880 50.790 179.200 ;
        RECT 50.530 175.140 50.790 175.460 ;
        RECT 50.590 172.400 50.730 175.140 ;
        RECT 51.510 172.400 51.650 182.425 ;
        RECT 52.370 180.580 52.630 180.900 ;
        RECT 52.430 176.480 52.570 180.580 ;
        RECT 53.810 180.220 53.950 183.220 ;
        RECT 53.750 179.900 54.010 180.220 ;
        RECT 53.810 178.180 53.950 179.900 ;
        RECT 53.750 177.860 54.010 178.180 ;
        RECT 52.830 177.180 53.090 177.500 ;
        RECT 52.890 176.560 53.030 177.180 ;
        RECT 52.370 176.160 52.630 176.480 ;
        RECT 52.890 176.420 53.490 176.560 ;
        RECT 52.830 173.440 53.090 173.760 ;
        RECT 50.530 172.080 50.790 172.400 ;
        RECT 51.450 172.080 51.710 172.400 ;
        RECT 51.450 170.040 51.710 170.360 ;
        RECT 51.510 168.320 51.650 170.040 ;
        RECT 51.450 168.000 51.710 168.320 ;
        RECT 52.890 167.300 53.030 173.440 ;
        RECT 53.350 171.040 53.490 176.420 ;
        RECT 53.810 173.080 53.950 177.860 ;
        RECT 54.730 175.800 54.870 183.900 ;
        RECT 54.670 175.480 54.930 175.800 ;
        RECT 54.210 174.800 54.470 175.120 ;
        RECT 53.750 172.760 54.010 173.080 ;
        RECT 53.290 170.720 53.550 171.040 ;
        RECT 53.750 169.700 54.010 170.020 ;
        RECT 53.290 167.660 53.550 167.980 ;
        RECT 52.830 166.980 53.090 167.300 ;
        RECT 50.530 166.640 50.790 166.960 ;
        RECT 50.590 165.600 50.730 166.640 ;
        RECT 51.450 166.300 51.710 166.620 ;
        RECT 52.370 166.300 52.630 166.620 ;
        RECT 50.530 165.280 50.790 165.600 ;
        RECT 51.510 164.920 51.650 166.300 ;
        RECT 52.430 165.260 52.570 166.300 ;
        RECT 52.370 164.940 52.630 165.260 ;
        RECT 51.450 164.600 51.710 164.920 ;
        RECT 50.060 164.065 50.340 164.435 ;
        RECT 51.910 164.260 52.170 164.580 ;
        RECT 50.530 163.580 50.790 163.900 ;
        RECT 51.450 163.810 51.710 163.900 ;
        RECT 51.050 163.670 51.710 163.810 ;
        RECT 48.290 161.860 48.430 162.310 ;
        RECT 49.600 162.025 49.880 162.395 ;
        RECT 48.230 161.540 48.490 161.860 ;
        RECT 49.610 161.715 49.870 161.860 ;
        RECT 49.600 161.345 49.880 161.715 ;
        RECT 46.380 160.665 46.660 161.035 ;
        RECT 49.610 160.860 49.870 161.180 ;
        RECT 45.930 160.070 46.190 160.160 ;
        RECT 45.930 159.930 46.590 160.070 ;
        RECT 45.930 159.840 46.190 159.930 ;
        RECT 45.470 159.500 45.730 159.820 ;
        RECT 45.930 159.160 46.190 159.480 ;
        RECT 45.990 156.420 46.130 159.160 ;
        RECT 46.450 156.955 46.590 159.930 ;
        RECT 48.230 159.840 48.490 160.160 ;
        RECT 46.840 159.305 47.120 159.675 ;
        RECT 48.290 159.480 48.430 159.840 ;
        RECT 46.850 159.160 47.110 159.305 ;
        RECT 48.230 159.160 48.490 159.480 ;
        RECT 46.380 156.585 46.660 156.955 ;
        RECT 45.930 156.100 46.190 156.420 ;
        RECT 46.390 156.330 46.650 156.420 ;
        RECT 46.910 156.330 47.050 159.160 ;
        RECT 47.510 157.605 49.390 157.975 ;
        RECT 47.760 156.585 48.040 156.955 ;
        RECT 47.830 156.420 47.970 156.585 ;
        RECT 46.390 156.190 47.050 156.330 ;
        RECT 46.390 156.100 46.650 156.190 ;
        RECT 47.770 156.100 48.030 156.420 ;
        RECT 46.840 154.545 47.120 154.915 ;
        RECT 45.010 154.060 45.270 154.380 ;
        RECT 46.390 154.060 46.650 154.380 ;
        RECT 45.470 153.720 45.730 154.040 ;
        RECT 45.010 153.380 45.270 153.700 ;
        RECT 44.150 142.420 44.750 142.560 ;
        RECT 43.630 141.820 43.890 142.140 ;
        RECT 43.170 139.440 43.430 139.760 ;
        RECT 42.710 135.360 42.970 135.680 ;
        RECT 42.710 134.000 42.970 134.320 ;
        RECT 42.250 132.640 42.510 132.960 ;
        RECT 41.790 131.620 42.050 131.940 ;
        RECT 42.770 129.900 42.910 134.000 ;
        RECT 40.870 129.580 41.130 129.900 ;
        RECT 41.330 129.580 41.590 129.900 ;
        RECT 42.710 129.580 42.970 129.900 ;
        RECT 43.230 128.540 43.370 139.440 ;
        RECT 43.630 138.080 43.890 138.400 ;
        RECT 43.170 128.220 43.430 128.540 ;
        RECT 43.690 127.520 43.830 138.080 ;
        RECT 44.150 134.910 44.290 142.420 ;
        RECT 44.550 141.820 44.810 142.140 ;
        RECT 44.610 140.010 44.750 141.820 ;
        RECT 45.070 140.520 45.210 153.380 ;
        RECT 45.530 147.920 45.670 153.720 ;
        RECT 45.930 152.700 46.190 153.020 ;
        RECT 45.990 150.300 46.130 152.700 ;
        RECT 46.450 152.000 46.590 154.060 ;
        RECT 46.910 154.040 47.050 154.545 ;
        RECT 49.670 154.040 49.810 160.860 ;
        RECT 50.060 159.305 50.340 159.675 ;
        RECT 50.130 156.420 50.270 159.305 ;
        RECT 50.070 156.100 50.330 156.420 ;
        RECT 46.850 153.720 47.110 154.040 ;
        RECT 49.610 153.720 49.870 154.040 ;
        RECT 50.060 153.865 50.340 154.235 ;
        RECT 50.070 153.720 50.330 153.865 ;
        RECT 49.600 153.185 49.880 153.555 ;
        RECT 46.850 152.700 47.110 153.020 ;
        RECT 46.390 151.680 46.650 152.000 ;
        RECT 46.380 151.145 46.660 151.515 ;
        RECT 46.450 150.980 46.590 151.145 ;
        RECT 46.390 150.660 46.650 150.980 ;
        RECT 45.930 149.980 46.190 150.300 ;
        RECT 46.910 148.000 47.050 152.700 ;
        RECT 47.510 152.165 49.390 152.535 ;
        RECT 49.670 150.980 49.810 153.185 ;
        RECT 49.610 150.660 49.870 150.980 ;
        RECT 45.470 147.600 45.730 147.920 ;
        RECT 45.990 147.860 47.050 148.000 ;
        RECT 49.610 147.940 49.870 148.260 ;
        RECT 45.990 141.880 46.130 147.860 ;
        RECT 46.850 147.260 47.110 147.580 ;
        RECT 46.910 145.880 47.050 147.260 ;
        RECT 47.510 146.725 49.390 147.095 ;
        RECT 46.850 145.560 47.110 145.880 ;
        RECT 45.990 141.740 46.590 141.880 ;
        RECT 46.850 141.820 47.110 142.140 ;
        RECT 45.070 140.380 45.670 140.520 ;
        RECT 44.610 139.870 45.210 140.010 ;
        RECT 44.550 134.910 44.810 135.000 ;
        RECT 44.150 134.770 44.810 134.910 ;
        RECT 44.550 134.680 44.810 134.770 ;
        RECT 45.070 134.400 45.210 139.870 ;
        RECT 45.530 135.680 45.670 140.380 ;
        RECT 45.470 135.360 45.730 135.680 ;
        RECT 44.150 134.260 45.210 134.400 ;
        RECT 43.630 127.200 43.890 127.520 ;
        RECT 40.870 126.860 41.130 127.180 ;
        RECT 40.410 126.180 40.670 126.500 ;
        RECT 40.410 125.500 40.670 125.820 ;
        RECT 38.570 124.480 38.830 124.800 ;
        RECT 39.490 124.480 39.750 124.800 ;
        RECT 35.350 121.760 35.610 122.080 ;
        RECT 34.890 121.420 35.150 121.740 ;
        RECT 35.810 120.740 36.070 121.060 ;
        RECT 35.870 108.580 36.010 120.740 ;
        RECT 40.470 108.580 40.610 125.500 ;
        RECT 40.930 123.100 41.070 126.860 ;
        RECT 41.330 126.180 41.590 126.500 ;
        RECT 41.390 123.440 41.530 126.180 ;
        RECT 44.150 124.800 44.290 134.260 ;
        RECT 45.530 132.960 45.670 135.360 ;
        RECT 45.470 132.640 45.730 132.960 ;
        RECT 44.550 130.940 44.810 131.260 ;
        RECT 44.610 129.560 44.750 130.940 ;
        RECT 44.550 129.240 44.810 129.560 ;
        RECT 45.010 128.900 45.270 129.220 ;
        RECT 44.090 124.480 44.350 124.800 ;
        RECT 41.330 123.120 41.590 123.440 ;
        RECT 40.870 122.780 41.130 123.100 ;
        RECT 41.390 121.060 41.530 123.120 ;
        RECT 41.330 120.740 41.590 121.060 ;
        RECT 45.070 108.580 45.210 128.900 ;
        RECT 46.450 121.740 46.590 141.740 ;
        RECT 46.910 140.440 47.050 141.820 ;
        RECT 47.510 141.285 49.390 141.655 ;
        RECT 46.850 140.120 47.110 140.440 ;
        RECT 49.150 140.010 49.410 140.100 ;
        RECT 49.670 140.010 49.810 147.940 ;
        RECT 50.590 147.580 50.730 163.580 ;
        RECT 51.050 159.560 51.190 163.670 ;
        RECT 51.450 163.580 51.710 163.670 ;
        RECT 51.050 159.420 51.650 159.560 ;
        RECT 50.990 158.820 51.250 159.140 ;
        RECT 51.050 157.440 51.190 158.820 ;
        RECT 50.990 157.120 51.250 157.440 ;
        RECT 50.990 156.440 51.250 156.760 ;
        RECT 51.050 154.720 51.190 156.440 ;
        RECT 50.990 154.400 51.250 154.720 ;
        RECT 50.980 153.865 51.260 154.235 ;
        RECT 51.050 152.000 51.190 153.865 ;
        RECT 50.990 151.680 51.250 152.000 ;
        RECT 51.510 148.600 51.650 159.420 ;
        RECT 51.970 154.040 52.110 164.260 ;
        RECT 52.430 161.860 52.570 164.940 ;
        RECT 52.890 161.860 53.030 166.980 ;
        RECT 53.350 164.920 53.490 167.660 ;
        RECT 53.810 164.920 53.950 169.700 ;
        RECT 54.270 165.260 54.410 174.800 ;
        RECT 54.670 174.460 54.930 174.780 ;
        RECT 54.730 171.040 54.870 174.460 ;
        RECT 54.670 170.720 54.930 171.040 ;
        RECT 54.730 170.360 54.870 170.720 ;
        RECT 54.670 170.040 54.930 170.360 ;
        RECT 54.670 169.360 54.930 169.680 ;
        RECT 54.730 167.640 54.870 169.360 ;
        RECT 54.670 167.320 54.930 167.640 ;
        RECT 54.670 166.640 54.930 166.960 ;
        RECT 54.210 164.940 54.470 165.260 ;
        RECT 53.290 164.600 53.550 164.920 ;
        RECT 53.750 164.600 54.010 164.920 ;
        RECT 53.350 164.320 53.490 164.600 ;
        RECT 54.210 164.320 54.470 164.580 ;
        RECT 53.350 164.260 54.470 164.320 ;
        RECT 53.350 164.180 54.410 164.260 ;
        RECT 54.730 163.810 54.870 166.640 ;
        RECT 54.270 163.670 54.870 163.810 ;
        RECT 52.370 161.540 52.630 161.860 ;
        RECT 52.830 161.540 53.090 161.860 ;
        RECT 53.750 161.540 54.010 161.860 ;
        RECT 52.830 158.140 53.090 158.460 ;
        RECT 52.360 156.585 52.640 156.955 ;
        RECT 52.430 156.420 52.570 156.585 ;
        RECT 52.370 156.100 52.630 156.420 ;
        RECT 51.910 153.720 52.170 154.040 ;
        RECT 52.890 152.930 53.030 158.140 ;
        RECT 53.290 155.420 53.550 155.740 ;
        RECT 51.970 152.790 53.030 152.930 ;
        RECT 51.450 148.280 51.710 148.600 ;
        RECT 51.970 148.260 52.110 152.790 ;
        RECT 52.370 149.980 52.630 150.300 ;
        RECT 51.910 147.940 52.170 148.260 ;
        RECT 50.530 147.260 50.790 147.580 ;
        RECT 51.910 147.260 52.170 147.580 ;
        RECT 50.530 145.560 50.790 145.880 ;
        RECT 50.070 144.880 50.330 145.200 ;
        RECT 50.130 143.160 50.270 144.880 ;
        RECT 50.070 142.840 50.330 143.160 ;
        RECT 50.130 140.440 50.270 142.840 ;
        RECT 50.070 140.120 50.330 140.440 ;
        RECT 49.150 139.955 49.810 140.010 ;
        RECT 49.140 139.870 49.810 139.955 ;
        RECT 49.140 139.585 49.420 139.870 ;
        RECT 49.610 139.100 49.870 139.420 ;
        RECT 47.510 135.845 49.390 136.215 ;
        RECT 49.670 135.680 49.810 139.100 ;
        RECT 50.130 137.380 50.270 140.120 ;
        RECT 50.070 137.060 50.330 137.380 ;
        RECT 49.610 135.360 49.870 135.680 ;
        RECT 50.070 134.680 50.330 135.000 ;
        RECT 46.850 133.660 47.110 133.980 ;
        RECT 46.910 132.960 47.050 133.660 ;
        RECT 50.130 132.960 50.270 134.680 ;
        RECT 46.850 132.640 47.110 132.960 ;
        RECT 50.070 132.640 50.330 132.960 ;
        RECT 50.590 132.280 50.730 145.560 ;
        RECT 51.450 143.520 51.710 143.840 ;
        RECT 50.990 137.060 51.250 137.380 ;
        RECT 50.530 131.960 50.790 132.280 ;
        RECT 47.510 130.405 49.390 130.775 ;
        RECT 51.050 130.240 51.190 137.060 ;
        RECT 51.510 132.960 51.650 143.520 ;
        RECT 51.450 132.640 51.710 132.960 ;
        RECT 50.990 129.920 51.250 130.240 ;
        RECT 50.990 128.560 51.250 128.880 ;
        RECT 50.530 126.180 50.790 126.500 ;
        RECT 47.510 124.965 49.390 125.335 ;
        RECT 50.590 124.120 50.730 126.180 ;
        RECT 50.530 123.800 50.790 124.120 ;
        RECT 47.310 123.460 47.570 123.780 ;
        RECT 47.370 122.080 47.510 123.460 ;
        RECT 49.610 123.120 49.870 123.440 ;
        RECT 47.310 121.760 47.570 122.080 ;
        RECT 46.390 121.420 46.650 121.740 ;
        RECT 47.510 119.525 49.390 119.895 ;
        RECT 49.670 108.580 49.810 123.120 ;
        RECT 50.590 121.060 50.730 123.800 ;
        RECT 51.050 122.080 51.190 128.560 ;
        RECT 50.990 121.760 51.250 122.080 ;
        RECT 51.970 121.400 52.110 147.260 ;
        RECT 52.430 126.160 52.570 149.980 ;
        RECT 53.350 149.280 53.490 155.420 ;
        RECT 53.810 151.515 53.950 161.540 ;
        RECT 54.270 153.700 54.410 163.670 ;
        RECT 54.670 160.860 54.930 161.180 ;
        RECT 54.730 159.820 54.870 160.860 ;
        RECT 54.670 159.500 54.930 159.820 ;
        RECT 54.670 154.400 54.930 154.720 ;
        RECT 54.210 153.380 54.470 153.700 ;
        RECT 53.740 151.145 54.020 151.515 ;
        RECT 54.730 151.320 54.870 154.400 ;
        RECT 54.670 151.000 54.930 151.320 ;
        RECT 53.750 150.660 54.010 150.980 ;
        RECT 52.830 148.960 53.090 149.280 ;
        RECT 53.290 148.960 53.550 149.280 ;
        RECT 52.890 128.880 53.030 148.960 ;
        RECT 53.810 148.795 53.950 150.660 ;
        RECT 55.190 149.190 55.330 188.060 ;
        RECT 55.650 180.470 55.790 188.740 ;
        RECT 56.110 181.920 56.250 189.080 ;
        RECT 58.410 187.360 58.550 191.460 ;
        RECT 58.870 188.380 59.010 193.500 ;
        RECT 61.170 191.100 61.310 202.680 ;
        RECT 61.630 201.980 61.770 203.360 ;
        RECT 64.850 203.000 64.990 203.450 ;
        RECT 68.990 203.000 69.130 204.300 ;
        RECT 69.910 203.680 70.050 204.300 ;
        RECT 69.390 203.360 69.650 203.680 ;
        RECT 69.850 203.360 70.110 203.680 ;
        RECT 69.450 203.000 69.590 203.360 ;
        RECT 81.870 203.340 82.010 204.720 ;
        RECT 81.810 203.020 82.070 203.340 ;
        RECT 63.410 202.680 63.670 203.000 ;
        RECT 64.790 202.680 65.050 203.000 ;
        RECT 65.710 202.680 65.970 203.000 ;
        RECT 68.930 202.910 69.190 203.000 ;
        RECT 68.530 202.770 69.190 202.910 ;
        RECT 63.470 202.400 63.610 202.680 ;
        RECT 63.470 202.260 64.070 202.400 ;
        RECT 64.330 202.340 64.590 202.660 ;
        RECT 65.250 202.340 65.510 202.660 ;
        RECT 61.570 201.660 61.830 201.980 ;
        RECT 63.930 199.600 64.070 202.260 ;
        RECT 64.390 200.620 64.530 202.340 ;
        RECT 64.790 202.000 65.050 202.320 ;
        RECT 64.330 200.300 64.590 200.620 ;
        RECT 63.870 199.280 64.130 199.600 ;
        RECT 61.560 198.745 61.840 199.115 ;
        RECT 61.630 191.780 61.770 198.745 ;
        RECT 62.510 198.405 64.390 198.775 ;
        RECT 64.850 197.900 64.990 202.000 ;
        RECT 64.790 197.580 65.050 197.900 ;
        RECT 63.870 196.560 64.130 196.880 ;
        RECT 64.320 196.705 64.600 197.075 ;
        RECT 64.790 196.900 65.050 197.220 ;
        RECT 62.940 195.430 63.220 195.715 ;
        RECT 62.090 195.345 63.220 195.430 ;
        RECT 62.090 195.290 63.210 195.345 ;
        RECT 61.570 191.460 61.830 191.780 ;
        RECT 61.110 190.780 61.370 191.100 ;
        RECT 60.190 188.740 60.450 189.060 ;
        RECT 61.110 188.740 61.370 189.060 ;
        RECT 58.810 188.060 59.070 188.380 ;
        RECT 58.350 187.040 58.610 187.360 ;
        RECT 56.510 183.475 56.770 183.620 ;
        RECT 56.500 183.105 56.780 183.475 ;
        RECT 56.050 181.600 56.310 181.920 ;
        RECT 57.430 180.580 57.690 180.900 ;
        RECT 56.050 180.470 56.310 180.560 ;
        RECT 55.650 180.330 56.310 180.470 ;
        RECT 55.650 179.200 55.790 180.330 ;
        RECT 56.050 180.240 56.310 180.330 ;
        RECT 55.590 178.880 55.850 179.200 ;
        RECT 57.490 177.840 57.630 180.580 ;
        RECT 58.870 178.520 59.010 188.060 ;
        RECT 59.720 187.185 60.000 187.555 ;
        RECT 59.730 187.040 59.990 187.185 ;
        RECT 60.250 184.640 60.390 188.740 ;
        RECT 61.170 186.680 61.310 188.740 ;
        RECT 60.650 186.360 60.910 186.680 ;
        RECT 61.110 186.360 61.370 186.680 ;
        RECT 60.190 184.320 60.450 184.640 ;
        RECT 60.710 183.960 60.850 186.360 ;
        RECT 60.650 183.640 60.910 183.960 ;
        RECT 61.170 183.360 61.310 186.360 ;
        RECT 62.090 186.195 62.230 195.290 ;
        RECT 62.950 195.200 63.210 195.290 ;
        RECT 63.930 194.500 64.070 196.560 ;
        RECT 64.390 196.540 64.530 196.705 ;
        RECT 64.330 196.220 64.590 196.540 ;
        RECT 64.850 194.500 64.990 196.900 ;
        RECT 65.310 195.520 65.450 202.340 ;
        RECT 65.770 201.980 65.910 202.680 ;
        RECT 67.550 202.000 67.810 202.320 ;
        RECT 65.710 201.660 65.970 201.980 ;
        RECT 67.090 201.660 67.350 201.980 ;
        RECT 65.250 195.200 65.510 195.520 ;
        RECT 65.770 195.035 65.910 201.660 ;
        RECT 66.170 199.960 66.430 200.280 ;
        RECT 66.230 196.880 66.370 199.960 ;
        RECT 66.630 199.280 66.890 199.600 ;
        RECT 66.690 197.220 66.830 199.280 ;
        RECT 66.630 196.900 66.890 197.220 ;
        RECT 66.170 196.560 66.430 196.880 ;
        RECT 66.230 195.520 66.370 196.560 ;
        RECT 66.170 195.200 66.430 195.520 ;
        RECT 65.700 194.665 65.980 195.035 ;
        RECT 63.870 194.180 64.130 194.500 ;
        RECT 64.790 194.180 65.050 194.500 ;
        RECT 62.510 192.965 64.390 193.335 ;
        RECT 63.410 191.120 63.670 191.440 ;
        RECT 63.470 189.060 63.610 191.120 ;
        RECT 64.850 189.740 64.990 194.180 ;
        RECT 65.250 193.500 65.510 193.820 ;
        RECT 65.310 192.460 65.450 193.500 ;
        RECT 65.250 192.140 65.510 192.460 ;
        RECT 64.790 189.420 65.050 189.740 ;
        RECT 66.230 189.400 66.370 195.200 ;
        RECT 66.170 189.080 66.430 189.400 ;
        RECT 66.690 189.310 66.830 196.900 ;
        RECT 67.150 192.800 67.290 201.660 ;
        RECT 67.090 192.480 67.350 192.800 ;
        RECT 67.610 192.120 67.750 202.000 ;
        RECT 68.010 199.960 68.270 200.280 ;
        RECT 68.070 198.240 68.210 199.960 ;
        RECT 68.010 197.920 68.270 198.240 ;
        RECT 67.550 191.800 67.810 192.120 ;
        RECT 68.070 191.100 68.210 197.920 ;
        RECT 68.530 197.560 68.670 202.770 ;
        RECT 68.930 202.680 69.190 202.770 ;
        RECT 69.390 202.910 69.650 203.000 ;
        RECT 69.390 202.770 70.510 202.910 ;
        RECT 69.390 202.680 69.650 202.770 ;
        RECT 69.390 198.940 69.650 199.260 ;
        RECT 69.850 198.940 70.110 199.260 ;
        RECT 68.470 197.240 68.730 197.560 ;
        RECT 68.930 197.240 69.190 197.560 ;
        RECT 68.460 194.920 68.740 195.035 ;
        RECT 68.990 194.920 69.130 197.240 ;
        RECT 69.450 195.520 69.590 198.940 ;
        RECT 69.390 195.200 69.650 195.520 ;
        RECT 68.460 194.780 69.130 194.920 ;
        RECT 68.460 194.665 68.740 194.780 ;
        RECT 68.470 194.520 68.730 194.665 ;
        RECT 69.450 192.460 69.590 195.200 ;
        RECT 68.930 192.140 69.190 192.460 ;
        RECT 69.390 192.140 69.650 192.460 ;
        RECT 68.010 190.780 68.270 191.100 ;
        RECT 68.470 190.780 68.730 191.100 ;
        RECT 66.690 189.170 67.290 189.310 ;
        RECT 63.410 188.740 63.670 189.060 ;
        RECT 66.170 188.400 66.430 188.720 ;
        RECT 66.630 188.400 66.890 188.720 ;
        RECT 65.710 188.060 65.970 188.380 ;
        RECT 62.510 187.525 64.390 187.895 ;
        RECT 64.330 187.040 64.590 187.360 ;
        RECT 62.020 185.825 62.300 186.195 ;
        RECT 60.710 183.220 61.310 183.360 ;
        RECT 59.260 181.065 59.540 181.435 ;
        RECT 58.810 178.200 59.070 178.520 ;
        RECT 57.430 177.520 57.690 177.840 ;
        RECT 57.890 177.180 58.150 177.500 ;
        RECT 56.510 175.480 56.770 175.800 ;
        RECT 56.050 174.460 56.310 174.780 ;
        RECT 55.590 171.740 55.850 172.060 ;
        RECT 55.650 170.020 55.790 171.740 ;
        RECT 56.110 170.700 56.250 174.460 ;
        RECT 56.570 173.760 56.710 175.480 ;
        RECT 56.510 173.440 56.770 173.760 ;
        RECT 56.050 170.380 56.310 170.700 ;
        RECT 55.590 169.700 55.850 170.020 ;
        RECT 57.430 169.020 57.690 169.340 ;
        RECT 57.490 167.300 57.630 169.020 ;
        RECT 55.590 166.980 55.850 167.300 ;
        RECT 57.430 166.980 57.690 167.300 ;
        RECT 55.650 166.620 55.790 166.980 ;
        RECT 55.590 166.300 55.850 166.620 ;
        RECT 55.650 164.920 55.790 166.300 ;
        RECT 56.970 165.280 57.230 165.600 ;
        RECT 55.590 164.600 55.850 164.920 ;
        RECT 57.030 161.180 57.170 165.280 ;
        RECT 56.970 160.860 57.230 161.180 ;
        RECT 57.430 160.860 57.690 161.180 ;
        RECT 55.590 158.820 55.850 159.140 ;
        RECT 55.650 156.760 55.790 158.820 ;
        RECT 55.590 156.440 55.850 156.760 ;
        RECT 56.050 155.420 56.310 155.740 ;
        RECT 57.490 155.595 57.630 160.860 ;
        RECT 57.950 156.275 58.090 177.180 ;
        RECT 59.330 167.835 59.470 181.065 ;
        RECT 60.710 178.180 60.850 183.220 ;
        RECT 61.110 178.540 61.370 178.860 ;
        RECT 61.170 178.180 61.310 178.540 ;
        RECT 60.650 177.860 60.910 178.180 ;
        RECT 61.110 177.860 61.370 178.180 ;
        RECT 60.190 177.180 60.450 177.500 ;
        RECT 61.170 177.355 61.310 177.860 ;
        RECT 62.090 177.410 62.230 185.825 ;
        RECT 64.390 182.940 64.530 187.040 ;
        RECT 65.250 186.360 65.510 186.680 ;
        RECT 64.790 183.640 65.050 183.960 ;
        RECT 64.330 182.620 64.590 182.940 ;
        RECT 62.510 182.085 64.390 182.455 ;
        RECT 64.850 181.920 64.990 183.640 ;
        RECT 64.790 181.600 65.050 181.920 ;
        RECT 63.400 181.065 63.680 181.435 ;
        RECT 63.470 179.200 63.610 181.065 ;
        RECT 65.310 180.900 65.450 186.360 ;
        RECT 65.770 181.580 65.910 188.060 ;
        RECT 66.230 183.475 66.370 188.400 ;
        RECT 66.160 183.105 66.440 183.475 ;
        RECT 66.230 181.920 66.370 183.105 ;
        RECT 66.170 181.600 66.430 181.920 ;
        RECT 65.710 181.260 65.970 181.580 ;
        RECT 65.250 180.580 65.510 180.900 ;
        RECT 63.410 178.880 63.670 179.200 ;
        RECT 63.870 178.880 64.130 179.200 ;
        RECT 63.470 178.180 63.610 178.880 ;
        RECT 63.930 178.180 64.070 178.880 ;
        RECT 63.410 177.860 63.670 178.180 ;
        RECT 63.870 177.860 64.130 178.180 ;
        RECT 62.490 177.410 62.750 177.500 ;
        RECT 59.720 168.145 60.000 168.515 ;
        RECT 59.790 167.980 59.930 168.145 ;
        RECT 59.260 167.465 59.540 167.835 ;
        RECT 59.730 167.660 59.990 167.980 ;
        RECT 59.270 167.155 59.530 167.300 ;
        RECT 59.260 166.785 59.540 167.155 ;
        RECT 59.330 165.260 59.470 166.785 ;
        RECT 59.270 164.940 59.530 165.260 ;
        RECT 58.350 163.580 58.610 163.900 ;
        RECT 59.730 163.580 59.990 163.900 ;
        RECT 57.880 155.905 58.160 156.275 ;
        RECT 56.110 151.660 56.250 155.420 ;
        RECT 57.420 155.225 57.700 155.595 ;
        RECT 56.510 153.380 56.770 153.700 ;
        RECT 56.050 151.340 56.310 151.660 ;
        RECT 55.590 149.980 55.850 150.300 ;
        RECT 54.270 149.050 55.330 149.190 ;
        RECT 53.740 148.425 54.020 148.795 ;
        RECT 53.750 148.280 54.010 148.425 ;
        RECT 53.290 147.940 53.550 148.260 ;
        RECT 53.350 145.880 53.490 147.940 ;
        RECT 53.290 145.560 53.550 145.880 ;
        RECT 53.290 144.880 53.550 145.200 ;
        RECT 53.350 136.700 53.490 144.880 ;
        RECT 53.750 144.540 54.010 144.860 ;
        RECT 53.810 143.500 53.950 144.540 ;
        RECT 53.750 143.180 54.010 143.500 ;
        RECT 54.270 140.440 54.410 149.050 ;
        RECT 55.650 148.600 55.790 149.980 ;
        RECT 55.590 148.510 55.850 148.600 ;
        RECT 54.730 148.370 55.850 148.510 ;
        RECT 54.730 145.540 54.870 148.370 ;
        RECT 55.590 148.280 55.850 148.370 ;
        RECT 54.670 145.220 54.930 145.540 ;
        RECT 56.050 143.070 56.310 143.160 ;
        RECT 56.570 143.070 56.710 153.380 ;
        RECT 56.970 152.700 57.230 153.020 ;
        RECT 57.030 147.580 57.170 152.700 ;
        RECT 57.890 150.320 58.150 150.640 ;
        RECT 57.950 149.475 58.090 150.320 ;
        RECT 57.880 149.105 58.160 149.475 ;
        RECT 57.420 148.425 57.700 148.795 ;
        RECT 57.950 148.600 58.090 149.105 ;
        RECT 57.430 148.280 57.690 148.425 ;
        RECT 57.890 148.280 58.150 148.600 ;
        RECT 56.970 147.260 57.230 147.580 ;
        RECT 57.490 145.540 57.630 148.280 ;
        RECT 57.950 145.880 58.090 148.280 ;
        RECT 57.890 145.560 58.150 145.880 ;
        RECT 57.430 145.220 57.690 145.540 ;
        RECT 56.970 144.540 57.230 144.860 ;
        RECT 57.430 144.540 57.690 144.860 ;
        RECT 57.890 144.540 58.150 144.860 ;
        RECT 57.030 143.500 57.170 144.540 ;
        RECT 56.970 143.180 57.230 143.500 ;
        RECT 56.050 142.930 56.710 143.070 ;
        RECT 56.050 142.840 56.310 142.930 ;
        RECT 56.570 141.120 56.710 142.930 ;
        RECT 56.510 140.800 56.770 141.120 ;
        RECT 54.210 140.120 54.470 140.440 ;
        RECT 53.290 136.380 53.550 136.700 ;
        RECT 56.570 135.000 56.710 140.800 ;
        RECT 56.510 134.680 56.770 135.000 ;
        RECT 56.050 134.340 56.310 134.660 ;
        RECT 54.210 134.000 54.470 134.320 ;
        RECT 53.740 132.105 54.020 132.475 ;
        RECT 53.810 129.220 53.950 132.105 ;
        RECT 53.750 128.900 54.010 129.220 ;
        RECT 52.830 128.560 53.090 128.880 ;
        RECT 53.810 126.840 53.950 128.900 ;
        RECT 54.270 127.520 54.410 134.000 ;
        RECT 55.590 133.720 55.850 133.980 ;
        RECT 55.190 133.660 55.850 133.720 ;
        RECT 55.190 133.580 55.790 133.660 ;
        RECT 54.670 132.300 54.930 132.620 ;
        RECT 54.730 130.240 54.870 132.300 ;
        RECT 54.670 129.920 54.930 130.240 ;
        RECT 54.210 127.200 54.470 127.520 ;
        RECT 55.190 126.840 55.330 133.580 ;
        RECT 55.590 130.940 55.850 131.260 ;
        RECT 55.650 129.220 55.790 130.940 ;
        RECT 56.110 130.240 56.250 134.340 ;
        RECT 56.570 131.940 56.710 134.680 ;
        RECT 57.490 134.320 57.630 144.540 ;
        RECT 57.950 140.100 58.090 144.540 ;
        RECT 57.890 139.780 58.150 140.100 ;
        RECT 57.890 136.380 58.150 136.700 ;
        RECT 57.430 134.000 57.690 134.320 ;
        RECT 57.950 132.870 58.090 136.380 ;
        RECT 58.410 134.660 58.550 163.580 ;
        RECT 59.790 161.860 59.930 163.580 ;
        RECT 58.810 161.540 59.070 161.860 ;
        RECT 59.270 161.540 59.530 161.860 ;
        RECT 59.730 161.540 59.990 161.860 ;
        RECT 58.870 157.100 59.010 161.540 ;
        RECT 59.330 159.820 59.470 161.540 ;
        RECT 59.790 160.160 59.930 161.540 ;
        RECT 59.730 159.840 59.990 160.160 ;
        RECT 59.270 159.675 59.530 159.820 ;
        RECT 59.260 159.305 59.540 159.675 ;
        RECT 60.250 159.560 60.390 177.180 ;
        RECT 61.100 176.985 61.380 177.355 ;
        RECT 62.090 177.270 62.750 177.410 ;
        RECT 62.490 177.180 62.750 177.270 ;
        RECT 65.710 177.180 65.970 177.500 ;
        RECT 60.640 176.305 60.920 176.675 ;
        RECT 62.510 176.645 64.390 177.015 ;
        RECT 60.710 174.780 60.850 176.305 ;
        RECT 64.790 175.820 65.050 176.140 ;
        RECT 61.570 175.140 61.830 175.460 ;
        RECT 60.650 174.460 60.910 174.780 ;
        RECT 60.710 173.080 60.850 174.460 ;
        RECT 60.650 172.760 60.910 173.080 ;
        RECT 60.650 171.740 60.910 172.060 ;
        RECT 60.710 170.270 60.850 171.740 ;
        RECT 61.110 170.270 61.370 170.360 ;
        RECT 60.710 170.130 61.370 170.270 ;
        RECT 60.710 167.980 60.850 170.130 ;
        RECT 61.110 170.040 61.370 170.130 ;
        RECT 60.650 167.660 60.910 167.980 ;
        RECT 61.110 167.660 61.370 167.980 ;
        RECT 61.170 167.040 61.310 167.660 ;
        RECT 61.630 167.640 61.770 175.140 ;
        RECT 62.510 171.205 64.390 171.575 ;
        RECT 63.860 168.145 64.140 168.515 ;
        RECT 64.850 168.320 64.990 175.820 ;
        RECT 65.770 175.200 65.910 177.180 ;
        RECT 65.310 175.060 65.910 175.200 ;
        RECT 61.570 167.320 61.830 167.640 ;
        RECT 63.930 167.300 64.070 168.145 ;
        RECT 64.790 168.000 65.050 168.320 ;
        RECT 62.950 167.155 63.210 167.300 ;
        RECT 59.790 159.420 60.390 159.560 ;
        RECT 60.710 166.900 61.310 167.040 ;
        RECT 58.810 156.780 59.070 157.100 ;
        RECT 59.790 152.880 59.930 159.420 ;
        RECT 60.190 156.100 60.450 156.420 ;
        RECT 60.250 155.595 60.390 156.100 ;
        RECT 60.180 155.225 60.460 155.595 ;
        RECT 59.790 152.740 60.390 152.880 ;
        RECT 59.270 150.660 59.530 150.980 ;
        RECT 59.330 148.600 59.470 150.660 ;
        RECT 59.270 148.280 59.530 148.600 ;
        RECT 59.270 147.600 59.530 147.920 ;
        RECT 59.330 143.840 59.470 147.600 ;
        RECT 59.270 143.520 59.530 143.840 ;
        RECT 59.270 141.820 59.530 142.140 ;
        RECT 59.330 137.720 59.470 141.820 ;
        RECT 59.730 140.800 59.990 141.120 ;
        RECT 59.270 137.400 59.530 137.720 ;
        RECT 58.350 134.340 58.610 134.660 ;
        RECT 58.350 132.870 58.610 132.960 ;
        RECT 57.950 132.730 58.610 132.870 ;
        RECT 58.350 132.640 58.610 132.730 ;
        RECT 56.510 131.680 56.770 131.940 ;
        RECT 56.510 131.620 57.630 131.680 ;
        RECT 56.570 131.540 57.630 131.620 ;
        RECT 56.050 129.920 56.310 130.240 ;
        RECT 57.490 129.560 57.630 131.540 ;
        RECT 58.410 129.560 58.550 132.640 ;
        RECT 59.790 130.240 59.930 140.800 ;
        RECT 60.250 135.000 60.390 152.740 ;
        RECT 60.710 140.100 60.850 166.900 ;
        RECT 62.940 166.785 63.220 167.155 ;
        RECT 63.870 166.980 64.130 167.300 ;
        RECT 62.510 165.765 64.390 166.135 ;
        RECT 61.570 164.940 61.830 165.260 ;
        RECT 61.630 162.540 61.770 164.940 ;
        RECT 64.790 164.260 65.050 164.580 ;
        RECT 64.320 162.705 64.600 163.075 ;
        RECT 64.330 162.560 64.590 162.705 ;
        RECT 61.570 162.220 61.830 162.540 ;
        RECT 61.110 161.715 61.370 161.860 ;
        RECT 61.100 161.345 61.380 161.715 ;
        RECT 62.510 160.325 64.390 160.695 ;
        RECT 64.850 160.160 64.990 164.260 ;
        RECT 64.790 159.840 65.050 160.160 ;
        RECT 65.310 158.995 65.450 175.060 ;
        RECT 65.710 174.460 65.970 174.780 ;
        RECT 65.770 169.340 65.910 174.460 ;
        RECT 65.710 169.020 65.970 169.340 ;
        RECT 65.710 168.000 65.970 168.320 ;
        RECT 65.770 167.300 65.910 168.000 ;
        RECT 65.710 166.980 65.970 167.300 ;
        RECT 65.240 158.625 65.520 158.995 ;
        RECT 66.170 158.820 66.430 159.140 ;
        RECT 63.870 158.140 64.130 158.460 ;
        RECT 63.930 156.760 64.070 158.140 ;
        RECT 66.230 157.440 66.370 158.820 ;
        RECT 66.170 157.120 66.430 157.440 ;
        RECT 63.870 156.670 64.130 156.760 ;
        RECT 63.870 156.530 64.990 156.670 ;
        RECT 63.870 156.440 64.130 156.530 ;
        RECT 62.030 155.760 62.290 156.080 ;
        RECT 61.110 155.420 61.370 155.740 ;
        RECT 61.170 154.040 61.310 155.420 ;
        RECT 62.090 154.720 62.230 155.760 ;
        RECT 62.510 154.885 64.390 155.255 ;
        RECT 62.030 154.400 62.290 154.720 ;
        RECT 61.110 153.720 61.370 154.040 ;
        RECT 62.030 152.700 62.290 153.020 ;
        RECT 62.090 151.320 62.230 152.700 ;
        RECT 62.030 151.000 62.290 151.320 ;
        RECT 61.560 149.105 61.840 149.475 ;
        RECT 62.510 149.445 64.390 149.815 ;
        RECT 61.570 148.960 61.830 149.105 ;
        RECT 61.110 148.620 61.370 148.940 ;
        RECT 61.170 143.160 61.310 148.620 ;
        RECT 61.560 148.425 61.840 148.795 ;
        RECT 62.490 148.510 62.750 148.600 ;
        RECT 61.570 148.280 61.830 148.425 ;
        RECT 62.090 148.370 62.750 148.510 ;
        RECT 62.090 143.840 62.230 148.370 ;
        RECT 62.490 148.280 62.750 148.370 ;
        RECT 63.410 148.280 63.670 148.600 ;
        RECT 63.470 147.920 63.610 148.280 ;
        RECT 64.850 148.260 64.990 156.530 ;
        RECT 65.710 155.420 65.970 155.740 ;
        RECT 65.770 150.300 65.910 155.420 ;
        RECT 66.170 150.660 66.430 150.980 ;
        RECT 65.710 149.980 65.970 150.300 ;
        RECT 65.770 149.280 65.910 149.980 ;
        RECT 65.710 148.960 65.970 149.280 ;
        RECT 66.230 148.260 66.370 150.660 ;
        RECT 66.690 148.940 66.830 188.400 ;
        RECT 67.150 181.580 67.290 189.170 ;
        RECT 68.010 188.060 68.270 188.380 ;
        RECT 67.550 183.640 67.810 183.960 ;
        RECT 67.610 182.940 67.750 183.640 ;
        RECT 68.070 182.940 68.210 188.060 ;
        RECT 68.530 187.360 68.670 190.780 ;
        RECT 68.470 187.040 68.730 187.360 ;
        RECT 68.990 186.680 69.130 192.140 ;
        RECT 69.910 190.160 70.050 198.940 ;
        RECT 70.370 197.560 70.510 202.770 ;
        RECT 71.230 202.680 71.490 203.000 ;
        RECT 75.370 202.680 75.630 203.000 ;
        RECT 70.770 202.000 71.030 202.320 ;
        RECT 70.830 198.240 70.970 202.000 ;
        RECT 71.290 201.180 71.430 202.680 ;
        RECT 73.070 202.340 73.330 202.660 ;
        RECT 71.290 201.040 72.350 201.180 ;
        RECT 70.770 197.920 71.030 198.240 ;
        RECT 70.310 197.240 70.570 197.560 ;
        RECT 70.370 193.820 70.510 197.240 ;
        RECT 70.310 193.500 70.570 193.820 ;
        RECT 69.450 190.020 70.050 190.160 ;
        RECT 69.450 188.380 69.590 190.020 ;
        RECT 69.850 189.420 70.110 189.740 ;
        RECT 69.390 188.060 69.650 188.380 ;
        RECT 69.910 187.360 70.050 189.420 ;
        RECT 70.370 188.720 70.510 193.500 ;
        RECT 70.830 192.800 70.970 197.920 ;
        RECT 72.210 197.220 72.350 201.040 ;
        RECT 73.130 197.560 73.270 202.340 ;
        RECT 75.430 200.960 75.570 202.680 ;
        RECT 75.830 202.000 76.090 202.320 ;
        RECT 74.910 200.640 75.170 200.960 ;
        RECT 75.370 200.640 75.630 200.960 ;
        RECT 73.530 197.920 73.790 198.240 ;
        RECT 73.070 197.240 73.330 197.560 ;
        RECT 71.230 196.900 71.490 197.220 ;
        RECT 72.150 196.900 72.410 197.220 ;
        RECT 71.290 195.180 71.430 196.900 ;
        RECT 71.230 194.860 71.490 195.180 ;
        RECT 72.210 194.500 72.350 196.900 ;
        RECT 73.130 194.840 73.270 197.240 ;
        RECT 73.590 197.075 73.730 197.920 ;
        RECT 74.970 197.130 75.110 200.640 ;
        RECT 75.890 198.435 76.030 202.000 ;
        RECT 80.890 201.660 81.150 201.980 ;
        RECT 76.280 200.785 76.560 201.155 ;
        RECT 77.510 201.125 79.390 201.495 ;
        RECT 75.820 198.065 76.100 198.435 ;
        RECT 75.830 197.240 76.090 197.560 ;
        RECT 75.370 197.130 75.630 197.220 ;
        RECT 73.520 196.705 73.800 197.075 ;
        RECT 74.970 196.990 75.630 197.130 ;
        RECT 75.370 196.900 75.630 196.990 ;
        RECT 74.450 196.220 74.710 196.540 ;
        RECT 73.070 194.520 73.330 194.840 ;
        RECT 72.150 194.180 72.410 194.500 ;
        RECT 72.150 193.500 72.410 193.820 ;
        RECT 70.770 192.710 71.030 192.800 ;
        RECT 70.770 192.570 71.890 192.710 ;
        RECT 70.770 192.480 71.030 192.570 ;
        RECT 71.750 192.120 71.890 192.570 ;
        RECT 71.230 191.800 71.490 192.120 ;
        RECT 71.690 191.800 71.950 192.120 ;
        RECT 71.290 189.595 71.430 191.800 ;
        RECT 71.220 189.480 71.500 189.595 ;
        RECT 71.220 189.340 71.890 189.480 ;
        RECT 71.220 189.225 71.500 189.340 ;
        RECT 71.230 188.740 71.490 189.060 ;
        RECT 70.310 188.400 70.570 188.720 ;
        RECT 69.390 187.040 69.650 187.360 ;
        RECT 69.850 187.040 70.110 187.360 ;
        RECT 68.470 186.360 68.730 186.680 ;
        RECT 68.930 186.360 69.190 186.680 ;
        RECT 68.530 186.080 68.670 186.360 ;
        RECT 68.530 185.940 69.130 186.080 ;
        RECT 68.470 183.980 68.730 184.300 ;
        RECT 67.550 182.620 67.810 182.940 ;
        RECT 68.010 182.620 68.270 182.940 ;
        RECT 67.090 181.260 67.350 181.580 ;
        RECT 67.090 180.580 67.350 180.900 ;
        RECT 67.150 180.220 67.290 180.580 ;
        RECT 67.090 179.900 67.350 180.220 ;
        RECT 67.150 175.460 67.290 179.900 ;
        RECT 67.610 178.180 67.750 182.620 ;
        RECT 68.070 181.435 68.210 182.620 ;
        RECT 68.000 181.065 68.280 181.435 ;
        RECT 68.000 180.385 68.280 180.755 ;
        RECT 68.070 178.180 68.210 180.385 ;
        RECT 68.530 178.180 68.670 183.980 ;
        RECT 67.550 177.860 67.810 178.180 ;
        RECT 68.010 177.860 68.270 178.180 ;
        RECT 68.470 178.035 68.730 178.180 ;
        RECT 68.460 177.665 68.740 178.035 ;
        RECT 68.990 175.800 69.130 185.940 ;
        RECT 68.930 175.480 69.190 175.800 ;
        RECT 67.090 175.140 67.350 175.460 ;
        RECT 68.470 175.140 68.730 175.460 ;
        RECT 68.010 174.460 68.270 174.780 ;
        RECT 67.090 172.760 67.350 173.080 ;
        RECT 67.150 169.680 67.290 172.760 ;
        RECT 67.090 169.360 67.350 169.680 ;
        RECT 67.150 168.320 67.290 169.360 ;
        RECT 67.550 169.020 67.810 169.340 ;
        RECT 67.610 168.320 67.750 169.020 ;
        RECT 67.090 168.000 67.350 168.320 ;
        RECT 67.550 168.000 67.810 168.320 ;
        RECT 67.540 167.465 67.820 167.835 ;
        RECT 67.550 167.320 67.810 167.465 ;
        RECT 67.080 166.785 67.360 167.155 ;
        RECT 67.090 166.640 67.350 166.785 ;
        RECT 67.090 164.260 67.350 164.580 ;
        RECT 67.150 161.860 67.290 164.260 ;
        RECT 67.090 161.540 67.350 161.860 ;
        RECT 67.090 158.480 67.350 158.800 ;
        RECT 67.150 157.440 67.290 158.480 ;
        RECT 67.090 157.120 67.350 157.440 ;
        RECT 67.610 156.420 67.750 167.320 ;
        RECT 68.070 165.115 68.210 174.460 ;
        RECT 68.000 164.745 68.280 165.115 ;
        RECT 68.530 164.920 68.670 175.140 ;
        RECT 68.930 173.440 69.190 173.760 ;
        RECT 68.990 170.360 69.130 173.440 ;
        RECT 68.930 170.040 69.190 170.360 ;
        RECT 68.070 162.200 68.210 164.745 ;
        RECT 68.470 164.600 68.730 164.920 ;
        RECT 68.010 161.880 68.270 162.200 ;
        RECT 68.010 161.200 68.270 161.520 ;
        RECT 67.550 156.100 67.810 156.420 ;
        RECT 67.090 155.420 67.350 155.740 ;
        RECT 67.150 154.380 67.290 155.420 ;
        RECT 67.090 154.060 67.350 154.380 ;
        RECT 67.610 152.000 67.750 156.100 ;
        RECT 67.550 151.680 67.810 152.000 ;
        RECT 66.630 148.620 66.890 148.940 ;
        RECT 64.790 148.170 65.050 148.260 ;
        RECT 64.790 148.030 65.450 148.170 ;
        RECT 64.790 147.940 65.050 148.030 ;
        RECT 63.410 147.600 63.670 147.920 ;
        RECT 63.470 146.220 63.610 147.600 ;
        RECT 63.410 145.900 63.670 146.220 ;
        RECT 65.310 145.880 65.450 148.030 ;
        RECT 66.170 147.940 66.430 148.260 ;
        RECT 65.250 145.560 65.510 145.880 ;
        RECT 66.230 145.200 66.370 147.940 ;
        RECT 66.630 145.450 66.890 145.540 ;
        RECT 67.610 145.450 67.750 151.680 ;
        RECT 66.630 145.310 67.750 145.450 ;
        RECT 66.630 145.220 66.890 145.310 ;
        RECT 66.170 144.880 66.430 145.200 ;
        RECT 65.250 144.540 65.510 144.860 ;
        RECT 65.710 144.540 65.970 144.860 ;
        RECT 66.690 144.600 66.830 145.220 ;
        RECT 62.510 144.005 64.390 144.375 ;
        RECT 62.030 143.520 62.290 143.840 ;
        RECT 65.310 143.500 65.450 144.540 ;
        RECT 65.770 143.840 65.910 144.540 ;
        RECT 66.230 144.460 66.830 144.600 ;
        RECT 67.090 144.540 67.350 144.860 ;
        RECT 65.710 143.520 65.970 143.840 ;
        RECT 63.870 143.180 64.130 143.500 ;
        RECT 65.250 143.180 65.510 143.500 ;
        RECT 61.110 142.840 61.370 143.160 ;
        RECT 60.650 139.780 60.910 140.100 ;
        RECT 61.170 138.400 61.310 142.840 ;
        RECT 63.930 139.420 64.070 143.180 ;
        RECT 64.330 142.500 64.590 142.820 ;
        RECT 64.390 140.440 64.530 142.500 ;
        RECT 64.330 140.120 64.590 140.440 ;
        RECT 65.770 140.100 65.910 143.520 ;
        RECT 65.710 139.780 65.970 140.100 ;
        RECT 62.030 139.100 62.290 139.420 ;
        RECT 63.870 139.100 64.130 139.420 ;
        RECT 64.790 139.100 65.050 139.420 ;
        RECT 65.710 139.160 65.970 139.420 ;
        RECT 66.230 139.160 66.370 144.460 ;
        RECT 66.630 140.460 66.890 140.780 ;
        RECT 65.710 139.100 66.370 139.160 ;
        RECT 61.110 138.080 61.370 138.400 ;
        RECT 60.650 136.380 60.910 136.700 ;
        RECT 60.190 134.680 60.450 135.000 ;
        RECT 60.710 132.280 60.850 136.380 ;
        RECT 61.170 132.960 61.310 138.080 ;
        RECT 62.090 134.320 62.230 139.100 ;
        RECT 62.510 138.565 64.390 138.935 ;
        RECT 64.850 135.680 64.990 139.100 ;
        RECT 65.770 139.020 66.370 139.100 ;
        RECT 65.250 137.740 65.510 138.060 ;
        RECT 64.790 135.360 65.050 135.680 ;
        RECT 62.030 134.000 62.290 134.320 ;
        RECT 62.510 133.125 64.390 133.495 ;
        RECT 64.850 132.960 64.990 135.360 ;
        RECT 61.110 132.640 61.370 132.960 ;
        RECT 64.790 132.640 65.050 132.960 ;
        RECT 60.650 131.960 60.910 132.280 ;
        RECT 65.310 130.240 65.450 137.740 ;
        RECT 59.730 129.920 59.990 130.240 ;
        RECT 65.250 129.920 65.510 130.240 ;
        RECT 57.430 129.240 57.690 129.560 ;
        RECT 58.350 129.240 58.610 129.560 ;
        RECT 55.590 128.900 55.850 129.220 ;
        RECT 53.750 126.520 54.010 126.840 ;
        RECT 55.130 126.520 55.390 126.840 ;
        RECT 57.490 126.500 57.630 129.240 ;
        RECT 65.770 129.220 65.910 139.020 ;
        RECT 65.710 128.900 65.970 129.220 ;
        RECT 57.890 128.220 58.150 128.540 ;
        RECT 57.950 127.180 58.090 128.220 ;
        RECT 62.510 127.685 64.390 128.055 ;
        RECT 58.810 127.200 59.070 127.520 ;
        RECT 57.890 126.860 58.150 127.180 ;
        RECT 57.430 126.180 57.690 126.500 ;
        RECT 52.370 125.840 52.630 126.160 ;
        RECT 56.050 125.500 56.310 125.820 ;
        RECT 56.110 124.120 56.250 125.500 ;
        RECT 53.750 123.800 54.010 124.120 ;
        RECT 56.050 123.800 56.310 124.120 ;
        RECT 53.810 123.520 53.950 123.800 ;
        RECT 53.810 123.380 54.410 123.520 ;
        RECT 53.290 122.780 53.550 123.100 ;
        RECT 53.350 122.080 53.490 122.780 ;
        RECT 53.290 121.760 53.550 122.080 ;
        RECT 51.910 121.080 52.170 121.400 ;
        RECT 50.530 120.740 50.790 121.060 ;
        RECT 54.270 108.580 54.410 123.380 ;
        RECT 56.050 123.120 56.310 123.440 ;
        RECT 56.110 122.080 56.250 123.120 ;
        RECT 56.050 121.760 56.310 122.080 ;
        RECT 58.870 108.580 59.010 127.200 ;
        RECT 60.650 126.860 60.910 127.180 ;
        RECT 60.710 122.080 60.850 126.860 ;
        RECT 66.690 126.840 66.830 140.460 ;
        RECT 67.150 140.440 67.290 144.540 ;
        RECT 67.090 140.120 67.350 140.440 ;
        RECT 67.150 131.600 67.290 140.120 ;
        RECT 68.070 137.800 68.210 161.200 ;
        RECT 68.990 152.880 69.130 170.040 ;
        RECT 69.450 162.880 69.590 187.040 ;
        RECT 69.910 180.640 70.050 187.040 ;
        RECT 70.370 186.760 70.510 188.400 ;
        RECT 71.290 187.360 71.430 188.740 ;
        RECT 71.230 187.040 71.490 187.360 ;
        RECT 70.770 186.760 71.030 187.020 ;
        RECT 70.370 186.700 71.030 186.760 ;
        RECT 70.370 186.620 70.970 186.700 ;
        RECT 70.370 186.340 70.510 186.620 ;
        RECT 70.310 186.020 70.570 186.340 ;
        RECT 70.370 181.240 70.510 186.020 ;
        RECT 71.290 186.000 71.430 187.040 ;
        RECT 71.230 185.680 71.490 186.000 ;
        RECT 70.770 184.155 71.030 184.300 ;
        RECT 70.760 183.785 71.040 184.155 ;
        RECT 70.770 182.960 71.030 183.280 ;
        RECT 70.830 182.115 70.970 182.960 ;
        RECT 70.760 181.745 71.040 182.115 ;
        RECT 71.290 181.580 71.430 185.680 ;
        RECT 71.230 181.260 71.490 181.580 ;
        RECT 70.310 180.920 70.570 181.240 ;
        RECT 70.770 180.640 71.030 180.900 ;
        RECT 69.910 180.580 71.030 180.640 ;
        RECT 69.910 180.500 70.970 180.580 ;
        RECT 71.230 179.900 71.490 180.220 ;
        RECT 71.750 180.075 71.890 189.340 ;
        RECT 69.850 177.180 70.110 177.500 ;
        RECT 70.770 177.180 71.030 177.500 ;
        RECT 69.910 165.600 70.050 177.180 ;
        RECT 70.830 175.880 70.970 177.180 ;
        RECT 70.370 175.800 70.970 175.880 ;
        RECT 70.310 175.740 70.970 175.800 ;
        RECT 71.290 175.880 71.430 179.900 ;
        RECT 71.680 179.705 71.960 180.075 ;
        RECT 71.690 178.880 71.950 179.200 ;
        RECT 71.750 178.520 71.890 178.880 ;
        RECT 71.690 178.200 71.950 178.520 ;
        RECT 71.690 177.520 71.950 177.840 ;
        RECT 71.750 176.480 71.890 177.520 ;
        RECT 71.690 176.160 71.950 176.480 ;
        RECT 71.290 175.800 71.890 175.880 ;
        RECT 71.290 175.740 71.950 175.800 ;
        RECT 70.310 175.480 70.570 175.740 ;
        RECT 70.830 170.700 70.970 175.740 ;
        RECT 71.690 175.480 71.950 175.740 ;
        RECT 70.770 170.610 71.030 170.700 ;
        RECT 70.770 170.470 71.430 170.610 ;
        RECT 70.770 170.380 71.030 170.470 ;
        RECT 70.760 169.505 71.040 169.875 ;
        RECT 70.300 168.145 70.580 168.515 ;
        RECT 70.370 167.980 70.510 168.145 ;
        RECT 70.310 167.660 70.570 167.980 ;
        RECT 70.370 167.300 70.510 167.660 ;
        RECT 70.310 166.980 70.570 167.300 ;
        RECT 70.830 165.795 70.970 169.505 ;
        RECT 69.850 165.280 70.110 165.600 ;
        RECT 70.760 165.425 71.040 165.795 ;
        RECT 70.770 164.940 71.030 165.260 ;
        RECT 70.830 163.810 70.970 164.940 ;
        RECT 71.290 164.920 71.430 170.470 ;
        RECT 71.690 166.980 71.950 167.300 ;
        RECT 71.750 164.920 71.890 166.980 ;
        RECT 71.230 164.600 71.490 164.920 ;
        RECT 71.690 164.600 71.950 164.920 ;
        RECT 71.220 164.065 71.500 164.435 ;
        RECT 71.230 163.920 71.490 164.065 ;
        RECT 70.600 163.670 70.970 163.810 ;
        RECT 70.600 162.960 70.740 163.670 ;
        RECT 69.390 162.560 69.650 162.880 ;
        RECT 70.600 162.820 70.970 162.960 ;
        RECT 70.830 162.790 70.970 162.820 ;
        RECT 70.830 162.650 71.430 162.790 ;
        RECT 69.450 159.480 69.590 162.560 ;
        RECT 70.310 162.220 70.570 162.540 ;
        RECT 69.390 159.390 69.650 159.480 ;
        RECT 69.390 159.250 70.050 159.390 ;
        RECT 69.390 159.160 69.650 159.250 ;
        RECT 69.390 158.140 69.650 158.460 ;
        RECT 69.450 154.380 69.590 158.140 ;
        RECT 69.910 156.420 70.050 159.250 ;
        RECT 69.850 156.100 70.110 156.420 ;
        RECT 69.850 155.650 70.110 155.740 ;
        RECT 70.370 155.650 70.510 162.220 ;
        RECT 70.760 162.025 71.040 162.395 ;
        RECT 70.770 161.880 71.030 162.025 ;
        RECT 70.770 161.200 71.030 161.520 ;
        RECT 70.830 160.355 70.970 161.200 ;
        RECT 70.760 159.985 71.040 160.355 ;
        RECT 69.850 155.510 70.510 155.650 ;
        RECT 69.850 155.420 70.110 155.510 ;
        RECT 69.390 154.060 69.650 154.380 ;
        RECT 69.910 152.880 70.050 155.420 ;
        RECT 70.770 153.380 71.030 153.700 ;
        RECT 68.530 152.740 69.130 152.880 ;
        RECT 69.450 152.740 70.050 152.880 ;
        RECT 68.530 141.030 68.670 152.740 ;
        RECT 69.450 145.540 69.590 152.740 ;
        RECT 70.830 150.980 70.970 153.380 ;
        RECT 70.770 150.660 71.030 150.980 ;
        RECT 69.850 148.620 70.110 148.940 ;
        RECT 70.770 148.620 71.030 148.940 ;
        RECT 69.910 145.540 70.050 148.620 ;
        RECT 70.830 147.580 70.970 148.620 ;
        RECT 71.290 148.600 71.430 162.650 ;
        RECT 71.750 162.200 71.890 164.600 ;
        RECT 71.690 161.880 71.950 162.200 ;
        RECT 72.210 161.860 72.350 193.500 ;
        RECT 72.610 191.800 72.870 192.120 ;
        RECT 73.070 191.800 73.330 192.120 ;
        RECT 73.530 191.800 73.790 192.120 ;
        RECT 72.670 186.000 72.810 191.800 ;
        RECT 73.130 189.740 73.270 191.800 ;
        RECT 73.070 189.420 73.330 189.740 ;
        RECT 73.590 188.380 73.730 191.800 ;
        RECT 73.530 188.060 73.790 188.380 ;
        RECT 72.610 185.680 72.870 186.000 ;
        RECT 73.060 185.825 73.340 186.195 ;
        RECT 72.670 181.580 72.810 185.680 ;
        RECT 73.130 183.280 73.270 185.825 ;
        RECT 73.530 185.680 73.790 186.000 ;
        RECT 73.070 182.960 73.330 183.280 ;
        RECT 72.610 181.260 72.870 181.580 ;
        RECT 73.070 180.240 73.330 180.560 ;
        RECT 72.600 179.705 72.880 180.075 ;
        RECT 72.670 178.600 72.810 179.705 ;
        RECT 73.130 179.200 73.270 180.240 ;
        RECT 73.070 178.880 73.330 179.200 ;
        RECT 72.670 178.460 73.270 178.600 ;
        RECT 72.610 177.860 72.870 178.180 ;
        RECT 72.670 175.800 72.810 177.860 ;
        RECT 72.610 175.480 72.870 175.800 ;
        RECT 73.130 173.760 73.270 178.460 ;
        RECT 73.070 173.670 73.330 173.760 ;
        RECT 72.670 173.530 73.330 173.670 ;
        RECT 72.670 169.875 72.810 173.530 ;
        RECT 73.070 173.440 73.330 173.530 ;
        RECT 73.070 172.420 73.330 172.740 ;
        RECT 73.130 170.360 73.270 172.420 ;
        RECT 73.070 170.040 73.330 170.360 ;
        RECT 72.600 169.505 72.880 169.875 ;
        RECT 73.130 169.680 73.270 170.040 ;
        RECT 73.070 169.360 73.330 169.680 ;
        RECT 73.070 167.320 73.330 167.640 ;
        RECT 72.610 166.640 72.870 166.960 ;
        RECT 72.150 161.600 72.410 161.860 ;
        RECT 71.750 161.540 72.410 161.600 ;
        RECT 71.750 161.460 72.350 161.540 ;
        RECT 71.750 159.480 71.890 161.460 ;
        RECT 72.150 160.860 72.410 161.180 ;
        RECT 72.210 159.820 72.350 160.860 ;
        RECT 72.150 159.500 72.410 159.820 ;
        RECT 71.690 159.160 71.950 159.480 ;
        RECT 71.750 156.080 71.890 159.160 ;
        RECT 71.690 155.760 71.950 156.080 ;
        RECT 72.670 154.040 72.810 166.640 ;
        RECT 73.130 156.420 73.270 167.320 ;
        RECT 73.590 165.795 73.730 185.680 ;
        RECT 74.510 181.240 74.650 196.220 ;
        RECT 75.890 193.820 76.030 197.240 ;
        RECT 76.350 197.075 76.490 200.785 ;
        RECT 80.950 199.600 81.090 201.660 ;
        RECT 84.170 200.280 84.310 205.740 ;
        RECT 88.770 205.040 88.910 205.740 ;
        RECT 88.710 204.720 88.970 205.040 ;
        RECT 89.170 204.720 89.430 205.040 ;
        RECT 84.570 203.020 84.830 203.340 ;
        RECT 83.650 199.960 83.910 200.280 ;
        RECT 84.110 199.960 84.370 200.280 ;
        RECT 80.890 199.280 81.150 199.600 ;
        RECT 82.730 199.280 82.990 199.600 ;
        RECT 83.180 199.425 83.460 199.795 ;
        RECT 82.790 198.240 82.930 199.280 ;
        RECT 82.730 197.920 82.990 198.240 ;
        RECT 79.970 197.240 80.230 197.560 ;
        RECT 76.280 196.705 76.560 197.075 ;
        RECT 76.750 196.900 77.010 197.220 ;
        RECT 76.290 196.220 76.550 196.540 ;
        RECT 74.910 193.500 75.170 193.820 ;
        RECT 75.830 193.500 76.090 193.820 ;
        RECT 74.970 191.780 75.110 193.500 ;
        RECT 74.910 191.460 75.170 191.780 ;
        RECT 74.970 189.060 75.110 191.460 ;
        RECT 74.910 188.740 75.170 189.060 ;
        RECT 74.910 187.040 75.170 187.360 ;
        RECT 74.970 186.875 75.110 187.040 ;
        RECT 74.900 186.505 75.180 186.875 ;
        RECT 75.370 186.020 75.630 186.340 ;
        RECT 75.830 186.020 76.090 186.340 ;
        RECT 74.900 184.465 75.180 184.835 ;
        RECT 74.910 184.320 75.170 184.465 ;
        RECT 74.910 183.640 75.170 183.960 ;
        RECT 74.450 180.920 74.710 181.240 ;
        RECT 73.990 179.900 74.250 180.220 ;
        RECT 74.050 177.840 74.190 179.900 ;
        RECT 74.510 178.180 74.650 180.920 ;
        RECT 74.970 180.220 75.110 183.640 ;
        RECT 75.430 183.620 75.570 186.020 ;
        RECT 75.890 183.620 76.030 186.020 ;
        RECT 75.370 183.300 75.630 183.620 ;
        RECT 75.830 183.300 76.090 183.620 ;
        RECT 75.370 181.600 75.630 181.920 ;
        RECT 74.910 179.900 75.170 180.220 ;
        RECT 74.910 178.880 75.170 179.200 ;
        RECT 74.970 178.715 75.110 178.880 ;
        RECT 74.900 178.345 75.180 178.715 ;
        RECT 74.450 177.860 74.710 178.180 ;
        RECT 73.990 177.520 74.250 177.840 ;
        RECT 74.450 175.820 74.710 176.140 ;
        RECT 74.970 175.995 75.110 178.345 ;
        RECT 73.990 175.480 74.250 175.800 ;
        RECT 74.050 172.740 74.190 175.480 ;
        RECT 73.990 172.420 74.250 172.740 ;
        RECT 73.990 170.380 74.250 170.700 ;
        RECT 74.050 167.300 74.190 170.380 ;
        RECT 73.990 166.980 74.250 167.300 ;
        RECT 73.990 166.300 74.250 166.620 ;
        RECT 73.520 165.425 73.800 165.795 ;
        RECT 73.530 165.170 73.790 165.260 ;
        RECT 74.050 165.170 74.190 166.300 ;
        RECT 73.530 165.030 74.190 165.170 ;
        RECT 73.530 164.940 73.790 165.030 ;
        RECT 74.510 162.540 74.650 175.820 ;
        RECT 74.900 175.625 75.180 175.995 ;
        RECT 75.430 175.200 75.570 181.600 ;
        RECT 75.890 181.240 76.030 183.300 ;
        RECT 75.830 180.920 76.090 181.240 ;
        RECT 75.890 178.520 76.030 180.920 ;
        RECT 75.830 178.200 76.090 178.520 ;
        RECT 76.350 178.180 76.490 196.220 ;
        RECT 76.810 187.020 76.950 196.900 ;
        RECT 79.510 196.220 79.770 196.540 ;
        RECT 80.030 196.395 80.170 197.240 ;
        RECT 77.510 195.685 79.390 196.055 ;
        RECT 79.570 194.840 79.710 196.220 ;
        RECT 79.960 196.025 80.240 196.395 ;
        RECT 79.510 194.520 79.770 194.840 ;
        RECT 80.030 192.880 80.170 196.025 ;
        RECT 83.250 195.520 83.390 199.425 ;
        RECT 83.710 198.240 83.850 199.960 ;
        RECT 84.100 199.425 84.380 199.795 ;
        RECT 83.650 197.920 83.910 198.240 ;
        RECT 84.170 197.640 84.310 199.425 ;
        RECT 84.630 199.260 84.770 203.020 ;
        RECT 89.230 203.000 89.370 204.720 ;
        RECT 91.530 203.340 91.670 206.225 ;
        RECT 94.690 205.400 94.950 205.720 ;
        RECT 92.510 203.845 94.390 204.215 ;
        RECT 91.930 203.360 92.190 203.680 ;
        RECT 91.470 203.020 91.730 203.340 ;
        RECT 86.870 202.680 87.130 203.000 ;
        RECT 89.170 202.680 89.430 203.000 ;
        RECT 85.020 200.105 85.300 200.475 ;
        RECT 84.570 198.940 84.830 199.260 ;
        RECT 83.710 197.500 84.310 197.640 ;
        RECT 84.630 197.560 84.770 198.940 ;
        RECT 85.090 197.560 85.230 200.105 ;
        RECT 86.930 199.795 87.070 202.680 ;
        RECT 88.310 200.220 90.290 200.360 ;
        RECT 88.310 199.940 88.450 200.220 ;
        RECT 86.860 199.425 87.140 199.795 ;
        RECT 88.250 199.620 88.510 199.940 ;
        RECT 86.870 198.940 87.130 199.260 ;
        RECT 87.790 199.170 88.050 199.260 ;
        RECT 87.790 199.030 88.450 199.170 ;
        RECT 87.790 198.940 88.050 199.030 ;
        RECT 83.190 195.200 83.450 195.520 ;
        RECT 83.710 195.180 83.850 197.500 ;
        RECT 84.570 197.240 84.830 197.560 ;
        RECT 85.030 197.240 85.290 197.560 ;
        RECT 84.110 196.900 84.370 197.220 ;
        RECT 84.170 195.520 84.310 196.900 ;
        RECT 84.110 195.200 84.370 195.520 ;
        RECT 83.650 194.860 83.910 195.180 ;
        RECT 83.710 194.500 83.850 194.860 ;
        RECT 84.630 194.840 84.770 197.240 ;
        RECT 86.930 197.220 87.070 198.940 ;
        RECT 86.870 196.900 87.130 197.220 ;
        RECT 86.930 194.840 87.070 196.900 ;
        RECT 84.570 194.520 84.830 194.840 ;
        RECT 85.950 194.520 86.210 194.840 ;
        RECT 86.870 194.520 87.130 194.840 ;
        RECT 83.650 194.180 83.910 194.500 ;
        RECT 84.110 194.180 84.370 194.500 ;
        RECT 80.430 193.500 80.690 193.820 ;
        RECT 79.570 192.740 80.170 192.880 ;
        RECT 77.510 190.245 79.390 190.615 ;
        RECT 78.130 188.740 78.390 189.060 ;
        RECT 77.210 187.040 77.470 187.360 ;
        RECT 76.750 186.700 77.010 187.020 ;
        RECT 77.270 186.250 77.410 187.040 ;
        RECT 76.810 186.110 77.410 186.250 ;
        RECT 76.810 184.300 76.950 186.110 ;
        RECT 78.190 185.660 78.330 188.740 ;
        RECT 78.130 185.340 78.390 185.660 ;
        RECT 77.510 184.805 79.390 185.175 ;
        RECT 79.570 184.640 79.710 192.740 ;
        RECT 80.490 191.100 80.630 193.500 ;
        RECT 80.430 190.780 80.690 191.100 ;
        RECT 80.490 188.380 80.630 190.780 ;
        RECT 80.430 188.290 80.690 188.380 ;
        RECT 80.030 188.150 80.690 188.290 ;
        RECT 80.030 186.680 80.170 188.150 ;
        RECT 80.430 188.060 80.690 188.150 ;
        RECT 79.970 186.360 80.230 186.680 ;
        RECT 80.430 186.360 80.690 186.680 ;
        RECT 79.510 184.320 79.770 184.640 ;
        RECT 80.490 184.300 80.630 186.360 ;
        RECT 81.350 185.340 81.610 185.660 ;
        RECT 76.750 183.980 77.010 184.300 ;
        RECT 77.210 183.980 77.470 184.300 ;
        RECT 80.430 183.980 80.690 184.300 ;
        RECT 77.270 183.620 77.410 183.980 ;
        RECT 80.490 183.620 80.630 183.980 ;
        RECT 77.210 183.300 77.470 183.620 ;
        RECT 78.130 183.300 78.390 183.620 ;
        RECT 80.430 183.300 80.690 183.620 ;
        RECT 77.210 182.850 77.470 182.940 ;
        RECT 78.190 182.850 78.330 183.300 ;
        RECT 77.210 182.710 78.330 182.850 ;
        RECT 77.210 182.620 77.470 182.710 ;
        RECT 78.190 181.435 78.330 182.710 ;
        RECT 79.970 182.620 80.230 182.940 ;
        RECT 78.120 181.065 78.400 181.435 ;
        RECT 79.510 180.920 79.770 181.240 ;
        RECT 76.750 180.580 77.010 180.900 ;
        RECT 76.290 177.860 76.550 178.180 ;
        RECT 75.430 175.060 76.030 175.200 ;
        RECT 75.370 174.460 75.630 174.780 ;
        RECT 74.910 172.080 75.170 172.400 ;
        RECT 74.970 171.040 75.110 172.080 ;
        RECT 75.430 172.060 75.570 174.460 ;
        RECT 75.370 171.740 75.630 172.060 ;
        RECT 74.910 170.720 75.170 171.040 ;
        RECT 75.370 170.040 75.630 170.360 ;
        RECT 74.910 169.020 75.170 169.340 ;
        RECT 74.970 166.620 75.110 169.020 ;
        RECT 74.910 166.300 75.170 166.620 ;
        RECT 74.970 164.920 75.110 166.300 ;
        RECT 75.430 164.920 75.570 170.040 ;
        RECT 75.890 167.980 76.030 175.060 ;
        RECT 76.810 170.020 76.950 180.580 ;
        RECT 77.510 179.365 79.390 179.735 ;
        RECT 77.510 173.925 79.390 174.295 ;
        RECT 77.670 173.100 77.930 173.420 ;
        RECT 77.730 171.040 77.870 173.100 ;
        RECT 79.570 171.040 79.710 180.920 ;
        RECT 80.030 171.800 80.170 182.620 ;
        RECT 80.490 178.860 80.630 183.300 ;
        RECT 81.410 181.580 81.550 185.340 ;
        RECT 84.170 183.280 84.310 194.180 ;
        RECT 86.010 193.820 86.150 194.520 ;
        RECT 87.790 194.180 88.050 194.500 ;
        RECT 88.310 194.410 88.450 199.030 ;
        RECT 88.710 198.940 88.970 199.260 ;
        RECT 88.770 197.900 88.910 198.940 ;
        RECT 88.710 197.580 88.970 197.900 ;
        RECT 90.150 195.520 90.290 200.220 ;
        RECT 91.010 200.190 91.270 200.280 ;
        RECT 91.010 200.050 91.670 200.190 ;
        RECT 91.010 199.960 91.270 200.050 ;
        RECT 91.000 198.065 91.280 198.435 ;
        RECT 91.530 198.240 91.670 200.050 ;
        RECT 91.070 197.900 91.210 198.065 ;
        RECT 91.470 197.920 91.730 198.240 ;
        RECT 91.010 197.580 91.270 197.900 ;
        RECT 91.990 197.560 92.130 203.360 ;
        RECT 94.750 202.400 94.890 205.400 ;
        RECT 95.150 205.060 95.410 205.380 ;
        RECT 95.210 203.340 95.350 205.060 ;
        RECT 96.070 204.380 96.330 204.700 ;
        RECT 96.130 203.680 96.270 204.380 ;
        RECT 96.070 203.360 96.330 203.680 ;
        RECT 95.150 203.020 95.410 203.340 ;
        RECT 97.450 202.680 97.710 203.000 ;
        RECT 94.750 202.260 95.350 202.400 ;
        RECT 96.530 202.340 96.790 202.660 ;
        RECT 96.990 202.340 97.250 202.660 ;
        RECT 92.510 198.405 94.390 198.775 ;
        RECT 95.210 198.240 95.350 202.260 ;
        RECT 96.070 200.300 96.330 200.620 ;
        RECT 95.600 199.425 95.880 199.795 ;
        RECT 95.150 197.920 95.410 198.240 ;
        RECT 95.670 197.900 95.810 199.425 ;
        RECT 95.610 197.580 95.870 197.900 ;
        RECT 91.930 197.240 92.190 197.560 ;
        RECT 91.470 196.560 91.730 196.880 ;
        RECT 94.690 196.560 94.950 196.880 ;
        RECT 90.090 195.200 90.350 195.520 ;
        RECT 89.160 194.665 89.440 195.035 ;
        RECT 91.010 194.860 91.270 195.180 ;
        RECT 88.710 194.410 88.970 194.500 ;
        RECT 88.310 194.270 88.970 194.410 ;
        RECT 88.710 194.180 88.970 194.270 ;
        RECT 85.950 193.500 86.210 193.820 ;
        RECT 85.490 191.800 85.750 192.120 ;
        RECT 85.030 188.060 85.290 188.380 ;
        RECT 85.090 187.360 85.230 188.060 ;
        RECT 85.030 187.040 85.290 187.360 ;
        RECT 85.030 186.020 85.290 186.340 ;
        RECT 84.570 183.300 84.830 183.620 ;
        RECT 84.110 182.960 84.370 183.280 ;
        RECT 81.350 181.260 81.610 181.580 ;
        RECT 82.720 181.065 83.000 181.435 ;
        RECT 84.630 181.240 84.770 183.300 ;
        RECT 85.090 182.940 85.230 186.020 ;
        RECT 85.550 183.960 85.690 191.800 ;
        RECT 86.010 189.400 86.150 193.500 ;
        RECT 87.850 192.460 87.990 194.180 ;
        RECT 87.790 192.140 88.050 192.460 ;
        RECT 86.870 190.780 87.130 191.100 ;
        RECT 85.950 189.080 86.210 189.400 ;
        RECT 85.950 186.700 86.210 187.020 ;
        RECT 86.010 184.300 86.150 186.700 ;
        RECT 85.950 183.980 86.210 184.300 ;
        RECT 85.490 183.640 85.750 183.960 ;
        RECT 85.030 182.620 85.290 182.940 ;
        RECT 86.410 182.620 86.670 182.940 ;
        RECT 85.090 181.240 85.230 182.620 ;
        RECT 82.730 180.920 82.990 181.065 ;
        RECT 84.570 180.920 84.830 181.240 ;
        RECT 85.030 180.920 85.290 181.240 ;
        RECT 81.350 180.580 81.610 180.900 ;
        RECT 80.430 178.540 80.690 178.860 ;
        RECT 80.430 177.180 80.690 177.500 ;
        RECT 80.490 172.400 80.630 177.180 ;
        RECT 80.890 175.820 81.150 176.140 ;
        RECT 80.430 172.080 80.690 172.400 ;
        RECT 80.030 171.660 80.630 171.800 ;
        RECT 77.670 170.720 77.930 171.040 ;
        RECT 79.510 170.950 79.770 171.040 ;
        RECT 79.510 170.810 80.170 170.950 ;
        RECT 79.510 170.720 79.770 170.810 ;
        RECT 79.510 170.040 79.770 170.360 ;
        RECT 76.750 169.700 77.010 170.020 ;
        RECT 76.810 168.230 76.950 169.700 ;
        RECT 77.510 168.485 79.390 168.855 ;
        RECT 76.810 168.090 78.790 168.230 ;
        RECT 75.830 167.660 76.090 167.980 ;
        RECT 74.910 164.600 75.170 164.920 ;
        RECT 75.370 164.600 75.630 164.920 ;
        RECT 74.450 162.220 74.710 162.540 ;
        RECT 74.970 161.600 75.110 164.600 ;
        RECT 75.430 162.200 75.570 164.600 ;
        RECT 75.890 162.200 76.030 167.660 ;
        RECT 77.210 166.640 77.470 166.960 ;
        RECT 76.750 166.300 77.010 166.620 ;
        RECT 76.280 165.425 76.560 165.795 ;
        RECT 75.370 161.880 75.630 162.200 ;
        RECT 75.830 161.880 76.090 162.200 ;
        RECT 74.970 161.520 75.570 161.600 ;
        RECT 74.970 161.460 75.630 161.520 ;
        RECT 75.370 161.200 75.630 161.460 ;
        RECT 74.910 160.860 75.170 161.180 ;
        RECT 76.350 160.920 76.490 165.425 ;
        RECT 76.810 165.260 76.950 166.300 ;
        RECT 76.750 164.940 77.010 165.260 ;
        RECT 77.270 164.920 77.410 166.640 ;
        RECT 78.650 166.530 78.790 168.090 ;
        RECT 79.050 166.530 79.310 166.620 ;
        RECT 78.650 166.390 79.310 166.530 ;
        RECT 77.660 165.425 77.940 165.795 ;
        RECT 77.730 164.920 77.870 165.425 ;
        RECT 77.210 164.600 77.470 164.920 ;
        RECT 77.670 164.600 77.930 164.920 ;
        RECT 78.650 164.580 78.790 166.390 ;
        RECT 79.050 166.300 79.310 166.390 ;
        RECT 79.570 165.260 79.710 170.040 ;
        RECT 80.030 167.640 80.170 170.810 ;
        RECT 79.970 167.320 80.230 167.640 ;
        RECT 79.510 164.940 79.770 165.260 ;
        RECT 79.970 164.600 80.230 164.920 ;
        RECT 76.740 164.065 77.020 164.435 ;
        RECT 78.590 164.260 78.850 164.580 ;
        RECT 74.450 157.120 74.710 157.440 ;
        RECT 73.070 156.100 73.330 156.420 ;
        RECT 74.510 156.275 74.650 157.120 ;
        RECT 74.440 155.905 74.720 156.275 ;
        RECT 72.610 153.720 72.870 154.040 ;
        RECT 71.690 152.700 71.950 153.020 ;
        RECT 73.990 152.700 74.250 153.020 ;
        RECT 71.230 148.280 71.490 148.600 ;
        RECT 70.310 147.260 70.570 147.580 ;
        RECT 70.770 147.260 71.030 147.580 ;
        RECT 69.390 145.220 69.650 145.540 ;
        RECT 69.850 145.220 70.110 145.540 ;
        RECT 68.530 140.890 69.130 141.030 ;
        RECT 68.460 140.265 68.740 140.635 ;
        RECT 68.530 140.100 68.670 140.265 ;
        RECT 68.470 139.780 68.730 140.100 ;
        RECT 68.070 137.660 68.670 137.800 ;
        RECT 68.010 137.060 68.270 137.380 ;
        RECT 68.070 132.960 68.210 137.060 ;
        RECT 68.010 132.640 68.270 132.960 ;
        RECT 68.530 132.475 68.670 137.660 ;
        RECT 68.460 132.105 68.740 132.475 ;
        RECT 68.990 131.940 69.130 140.890 ;
        RECT 68.930 131.620 69.190 131.940 ;
        RECT 67.090 131.280 67.350 131.600 ;
        RECT 68.990 130.240 69.130 131.620 ;
        RECT 68.930 129.920 69.190 130.240 ;
        RECT 66.630 126.520 66.890 126.840 ;
        RECT 61.110 126.180 61.370 126.500 ;
        RECT 64.790 126.180 65.050 126.500 ;
        RECT 61.170 124.120 61.310 126.180 ;
        RECT 61.110 123.800 61.370 124.120 ;
        RECT 62.030 123.120 62.290 123.440 ;
        RECT 60.650 121.760 60.910 122.080 ;
        RECT 26.600 106.580 26.880 108.580 ;
        RECT 31.200 106.580 31.480 108.580 ;
        RECT 35.800 106.580 36.080 108.580 ;
        RECT 40.400 106.580 40.680 108.580 ;
        RECT 45.000 106.580 45.280 108.580 ;
        RECT 49.600 106.580 49.880 108.580 ;
        RECT 54.200 106.580 54.480 108.580 ;
        RECT 58.800 106.580 59.080 108.580 ;
        RECT 62.090 108.560 62.230 123.120 ;
        RECT 62.510 122.245 64.390 122.615 ;
        RECT 64.850 121.400 64.990 126.180 ;
        RECT 67.550 125.500 67.810 125.820 ;
        RECT 68.930 125.500 69.190 125.820 ;
        RECT 67.610 124.120 67.750 125.500 ;
        RECT 67.550 123.800 67.810 124.120 ;
        RECT 65.710 123.120 65.970 123.440 ;
        RECT 65.770 122.080 65.910 123.120 ;
        RECT 65.710 121.760 65.970 122.080 ;
        RECT 68.990 121.740 69.130 125.500 ;
        RECT 69.450 122.080 69.590 145.220 ;
        RECT 70.370 144.770 70.510 147.260 ;
        RECT 70.830 146.560 70.970 147.260 ;
        RECT 70.770 146.240 71.030 146.560 ;
        RECT 70.770 144.880 71.030 145.200 ;
        RECT 69.910 144.630 70.510 144.770 ;
        RECT 69.910 136.700 70.050 144.630 ;
        RECT 70.830 141.120 70.970 144.880 ;
        RECT 70.770 140.800 71.030 141.120 ;
        RECT 69.850 136.380 70.110 136.700 ;
        RECT 70.310 136.380 70.570 136.700 ;
        RECT 69.910 129.560 70.050 136.380 ;
        RECT 70.370 135.000 70.510 136.380 ;
        RECT 70.310 134.680 70.570 135.000 ;
        RECT 69.850 129.240 70.110 129.560 ;
        RECT 71.750 129.220 71.890 152.700 ;
        RECT 72.610 151.680 72.870 152.000 ;
        RECT 72.670 150.980 72.810 151.680 ;
        RECT 72.150 150.660 72.410 150.980 ;
        RECT 72.610 150.660 72.870 150.980 ;
        RECT 72.210 142.820 72.350 150.660 ;
        RECT 73.530 150.320 73.790 150.640 ;
        RECT 73.590 148.940 73.730 150.320 ;
        RECT 73.530 148.620 73.790 148.940 ;
        RECT 73.070 147.260 73.330 147.580 ;
        RECT 72.150 142.500 72.410 142.820 ;
        RECT 72.210 137.380 72.350 142.500 ;
        RECT 72.150 137.060 72.410 137.380 ;
        RECT 72.210 135.000 72.350 137.060 ;
        RECT 72.150 134.680 72.410 135.000 ;
        RECT 71.690 128.900 71.950 129.220 ;
        RECT 73.130 126.840 73.270 147.260 ;
        RECT 73.530 144.540 73.790 144.860 ;
        RECT 73.590 143.160 73.730 144.540 ;
        RECT 73.530 142.840 73.790 143.160 ;
        RECT 74.050 142.480 74.190 152.700 ;
        RECT 74.450 150.660 74.710 150.980 ;
        RECT 74.510 147.920 74.650 150.660 ;
        RECT 74.450 147.600 74.710 147.920 ;
        RECT 74.450 146.240 74.710 146.560 ;
        RECT 73.990 142.160 74.250 142.480 ;
        RECT 73.990 139.100 74.250 139.420 ;
        RECT 74.050 137.720 74.190 139.100 ;
        RECT 74.510 138.400 74.650 146.240 ;
        RECT 74.970 145.540 75.110 160.860 ;
        RECT 75.430 160.780 76.490 160.920 ;
        RECT 75.430 153.700 75.570 160.780 ;
        RECT 76.290 158.480 76.550 158.800 ;
        RECT 75.820 156.585 76.100 156.955 ;
        RECT 76.350 156.760 76.490 158.480 ;
        RECT 76.810 156.840 76.950 164.065 ;
        RECT 77.510 163.045 79.390 163.415 ;
        RECT 80.030 162.200 80.170 164.600 ;
        RECT 79.970 161.880 80.230 162.200 ;
        RECT 78.590 161.200 78.850 161.520 ;
        RECT 78.650 159.820 78.790 161.200 ;
        RECT 78.590 159.730 78.850 159.820 ;
        RECT 78.590 159.590 79.710 159.730 ;
        RECT 78.590 159.500 78.850 159.590 ;
        RECT 77.510 157.605 79.390 157.975 ;
        RECT 75.830 156.440 76.090 156.585 ;
        RECT 76.290 156.440 76.550 156.760 ;
        RECT 76.810 156.700 78.790 156.840 ;
        RECT 76.350 154.040 76.490 156.440 ;
        RECT 78.650 156.420 78.790 156.700 ;
        RECT 79.570 156.420 79.710 159.590 ;
        RECT 77.670 156.100 77.930 156.420 ;
        RECT 78.590 156.100 78.850 156.420 ;
        RECT 79.510 156.100 79.770 156.420 ;
        RECT 76.290 153.720 76.550 154.040 ;
        RECT 76.750 153.950 77.010 154.040 ;
        RECT 77.730 153.950 77.870 156.100 ;
        RECT 78.650 154.040 78.790 156.100 ;
        RECT 80.490 156.080 80.630 171.660 ;
        RECT 80.950 171.040 81.090 175.820 ;
        RECT 80.890 170.720 81.150 171.040 ;
        RECT 80.890 169.360 81.150 169.680 ;
        RECT 80.950 167.155 81.090 169.360 ;
        RECT 80.880 166.785 81.160 167.155 ;
        RECT 80.950 164.920 81.090 166.785 ;
        RECT 80.890 164.600 81.150 164.920 ;
        RECT 80.890 160.860 81.150 161.180 ;
        RECT 80.950 159.820 81.090 160.860 ;
        RECT 80.890 159.500 81.150 159.820 ;
        RECT 80.890 157.120 81.150 157.440 ;
        RECT 80.430 155.760 80.690 156.080 ;
        RECT 79.510 155.420 79.770 155.740 ;
        RECT 76.750 153.810 77.870 153.950 ;
        RECT 76.750 153.720 77.010 153.810 ;
        RECT 78.590 153.720 78.850 154.040 ;
        RECT 75.370 153.380 75.630 153.700 ;
        RECT 76.350 152.880 76.490 153.720 ;
        RECT 75.890 152.740 76.490 152.880 ;
        RECT 75.890 148.680 76.030 152.740 ;
        RECT 76.810 151.910 76.950 153.720 ;
        RECT 77.510 152.165 79.390 152.535 ;
        RECT 76.810 151.770 77.410 151.910 ;
        RECT 77.270 149.280 77.410 151.770 ;
        RECT 77.210 148.960 77.470 149.280 ;
        RECT 75.890 148.600 76.950 148.680 ;
        RECT 77.270 148.600 77.410 148.960 ;
        RECT 75.890 148.540 77.010 148.600 ;
        RECT 76.750 148.280 77.010 148.540 ;
        RECT 77.210 148.280 77.470 148.600 ;
        RECT 77.670 148.280 77.930 148.600 ;
        RECT 75.830 147.260 76.090 147.580 ;
        RECT 75.360 145.705 75.640 146.075 ;
        RECT 75.370 145.560 75.630 145.705 ;
        RECT 74.910 145.220 75.170 145.540 ;
        RECT 75.370 144.880 75.630 145.200 ;
        RECT 75.430 143.920 75.570 144.880 ;
        RECT 74.970 143.780 75.570 143.920 ;
        RECT 74.970 141.120 75.110 143.780 ;
        RECT 75.370 143.180 75.630 143.500 ;
        RECT 74.910 140.800 75.170 141.120 ;
        RECT 74.450 138.080 74.710 138.400 ;
        RECT 73.990 137.400 74.250 137.720 ;
        RECT 74.970 137.380 75.110 140.800 ;
        RECT 75.430 137.720 75.570 143.180 ;
        RECT 75.890 138.060 76.030 147.260 ;
        RECT 76.810 145.880 76.950 148.280 ;
        RECT 77.730 147.580 77.870 148.280 ;
        RECT 77.670 147.260 77.930 147.580 ;
        RECT 77.510 146.725 79.390 147.095 ;
        RECT 76.750 145.560 77.010 145.880 ;
        RECT 77.670 145.450 77.930 145.540 ;
        RECT 77.670 145.310 78.330 145.450 ;
        RECT 77.670 145.220 77.930 145.310 ;
        RECT 77.670 144.540 77.930 144.860 ;
        RECT 76.750 142.840 77.010 143.160 ;
        RECT 76.810 140.440 76.950 142.840 ;
        RECT 77.730 142.140 77.870 144.540 ;
        RECT 78.190 142.820 78.330 145.310 ;
        RECT 78.130 142.500 78.390 142.820 ;
        RECT 77.670 141.820 77.930 142.140 ;
        RECT 77.510 141.285 79.390 141.655 ;
        RECT 76.750 140.120 77.010 140.440 ;
        RECT 75.830 137.740 76.090 138.060 ;
        RECT 75.370 137.400 75.630 137.720 ;
        RECT 74.910 137.060 75.170 137.380 ;
        RECT 75.430 135.680 75.570 137.400 ;
        RECT 75.370 135.360 75.630 135.680 ;
        RECT 76.810 135.000 76.950 140.120 ;
        RECT 79.570 139.840 79.710 155.420 ;
        RECT 79.970 153.720 80.230 154.040 ;
        RECT 80.030 148.600 80.170 153.720 ;
        RECT 79.970 148.280 80.230 148.600 ;
        RECT 80.030 146.220 80.170 148.280 ;
        RECT 80.430 147.940 80.690 148.260 ;
        RECT 79.970 145.900 80.230 146.220 ;
        RECT 80.030 145.540 80.170 145.900 ;
        RECT 80.490 145.880 80.630 147.940 ;
        RECT 80.430 145.560 80.690 145.880 ;
        RECT 79.970 145.220 80.230 145.540 ;
        RECT 79.970 144.540 80.230 144.860 ;
        RECT 80.030 143.840 80.170 144.540 ;
        RECT 79.970 143.520 80.230 143.840 ;
        RECT 80.030 140.440 80.170 143.520 ;
        RECT 79.970 140.120 80.230 140.440 ;
        RECT 79.570 139.700 80.630 139.840 ;
        RECT 78.130 137.400 78.390 137.720 ;
        RECT 78.190 137.040 78.330 137.400 ;
        RECT 78.130 136.720 78.390 137.040 ;
        RECT 77.510 135.845 79.390 136.215 ;
        RECT 76.750 134.680 77.010 135.000 ;
        RECT 73.990 134.000 74.250 134.320 ;
        RECT 74.050 132.960 74.190 134.000 ;
        RECT 73.990 132.640 74.250 132.960 ;
        RECT 76.290 132.190 76.550 132.280 ;
        RECT 76.810 132.190 76.950 134.680 ;
        RECT 79.510 133.660 79.770 133.980 ;
        RECT 76.290 132.050 76.950 132.190 ;
        RECT 76.290 131.960 76.550 132.050 ;
        RECT 75.830 131.620 76.090 131.940 ;
        RECT 74.910 130.940 75.170 131.260 ;
        RECT 73.070 126.520 73.330 126.840 ;
        RECT 70.310 125.500 70.570 125.820 ;
        RECT 73.990 125.500 74.250 125.820 ;
        RECT 69.390 121.760 69.650 122.080 ;
        RECT 68.930 121.420 69.190 121.740 ;
        RECT 64.790 121.080 65.050 121.400 ;
        RECT 70.370 121.060 70.510 125.500 ;
        RECT 72.610 123.120 72.870 123.440 ;
        RECT 67.550 120.800 67.810 121.060 ;
        RECT 67.550 120.740 68.210 120.800 ;
        RECT 70.310 120.740 70.570 121.060 ;
        RECT 67.610 120.660 68.210 120.740 ;
        RECT 63.010 109.100 63.610 109.240 ;
        RECT 63.010 108.560 63.150 109.100 ;
        RECT 63.470 108.580 63.610 109.100 ;
        RECT 68.070 108.580 68.210 120.660 ;
        RECT 72.670 108.580 72.810 123.120 ;
        RECT 74.050 121.740 74.190 125.500 ;
        RECT 73.990 121.420 74.250 121.740 ;
        RECT 74.970 121.400 75.110 130.940 ;
        RECT 75.890 129.900 76.030 131.620 ;
        RECT 75.830 129.580 76.090 129.900 ;
        RECT 75.370 128.560 75.630 128.880 ;
        RECT 75.430 124.120 75.570 128.560 ;
        RECT 75.830 128.220 76.090 128.540 ;
        RECT 75.890 127.180 76.030 128.220 ;
        RECT 75.830 126.860 76.090 127.180 ;
        RECT 76.350 126.500 76.490 131.960 ;
        RECT 77.510 130.405 79.390 130.775 ;
        RECT 79.570 129.560 79.710 133.660 ;
        RECT 79.960 132.105 80.240 132.475 ;
        RECT 79.510 129.240 79.770 129.560 ;
        RECT 80.030 129.220 80.170 132.105 ;
        RECT 80.490 129.900 80.630 139.700 ;
        RECT 80.950 138.310 81.090 157.120 ;
        RECT 81.410 149.190 81.550 180.580 ;
        RECT 81.810 180.240 82.070 180.560 ;
        RECT 81.870 176.390 82.010 180.240 ;
        RECT 82.730 179.900 82.990 180.220 ;
        RECT 82.270 176.390 82.530 176.480 ;
        RECT 81.870 176.250 82.530 176.390 ;
        RECT 81.870 175.460 82.010 176.250 ;
        RECT 82.270 176.160 82.530 176.250 ;
        RECT 81.810 175.140 82.070 175.460 ;
        RECT 81.870 168.320 82.010 175.140 ;
        RECT 82.270 172.760 82.530 173.080 ;
        RECT 82.330 168.320 82.470 172.760 ;
        RECT 81.810 168.000 82.070 168.320 ;
        RECT 82.270 168.000 82.530 168.320 ;
        RECT 82.270 160.860 82.530 161.180 ;
        RECT 81.810 155.420 82.070 155.740 ;
        RECT 81.870 153.020 82.010 155.420 ;
        RECT 82.330 154.380 82.470 160.860 ;
        RECT 82.790 157.100 82.930 179.900 ;
        RECT 85.090 179.200 85.230 180.920 ;
        RECT 85.030 178.880 85.290 179.200 ;
        RECT 85.090 175.800 85.230 178.880 ;
        RECT 85.950 177.520 86.210 177.840 ;
        RECT 86.010 176.140 86.150 177.520 ;
        RECT 85.950 175.820 86.210 176.140 ;
        RECT 85.030 175.480 85.290 175.800 ;
        RECT 84.570 174.460 84.830 174.780 ;
        RECT 83.190 173.440 83.450 173.760 ;
        RECT 83.250 170.360 83.390 173.440 ;
        RECT 83.190 170.270 83.450 170.360 ;
        RECT 83.190 170.130 83.850 170.270 ;
        RECT 83.190 170.040 83.450 170.130 ;
        RECT 83.190 166.980 83.450 167.300 ;
        RECT 83.250 165.600 83.390 166.980 ;
        RECT 83.710 165.795 83.850 170.130 ;
        RECT 83.190 165.280 83.450 165.600 ;
        RECT 83.640 165.425 83.920 165.795 ;
        RECT 83.710 164.920 83.850 165.425 ;
        RECT 83.650 164.600 83.910 164.920 ;
        RECT 84.630 162.880 84.770 174.460 ;
        RECT 85.090 173.080 85.230 175.480 ;
        RECT 86.010 175.315 86.150 175.820 ;
        RECT 85.940 174.945 86.220 175.315 ;
        RECT 85.030 172.760 85.290 173.080 ;
        RECT 85.090 167.300 85.230 172.760 ;
        RECT 86.470 172.400 86.610 182.620 ;
        RECT 86.930 181.580 87.070 190.780 ;
        RECT 87.790 189.420 88.050 189.740 ;
        RECT 87.330 183.300 87.590 183.620 ;
        RECT 86.870 181.260 87.130 181.580 ;
        RECT 87.390 180.810 87.530 183.300 ;
        RECT 86.930 180.670 87.530 180.810 ;
        RECT 86.930 178.180 87.070 180.670 ;
        RECT 86.870 177.860 87.130 178.180 ;
        RECT 86.930 175.120 87.070 177.860 ;
        RECT 87.850 175.460 87.990 189.420 ;
        RECT 88.250 188.740 88.510 189.060 ;
        RECT 88.310 181.920 88.450 188.740 ;
        RECT 88.770 187.555 88.910 194.180 ;
        RECT 89.230 190.080 89.370 194.665 ;
        RECT 91.070 192.200 91.210 194.860 ;
        RECT 91.530 194.500 91.670 196.560 ;
        RECT 94.220 195.345 94.500 195.715 ;
        RECT 94.290 194.500 94.430 195.345 ;
        RECT 91.470 194.180 91.730 194.500 ;
        RECT 94.230 194.180 94.490 194.500 ;
        RECT 91.470 193.500 91.730 193.820 ;
        RECT 91.530 192.710 91.670 193.500 ;
        RECT 92.510 192.965 94.390 193.335 ;
        RECT 91.530 192.570 92.590 192.710 ;
        RECT 91.070 192.120 91.670 192.200 ;
        RECT 91.070 192.060 91.730 192.120 ;
        RECT 90.090 190.780 90.350 191.100 ;
        RECT 90.550 190.780 90.810 191.100 ;
        RECT 90.150 190.080 90.290 190.780 ;
        RECT 89.170 189.760 89.430 190.080 ;
        RECT 90.090 189.760 90.350 190.080 ;
        RECT 89.630 189.420 89.890 189.740 ;
        RECT 89.160 188.545 89.440 188.915 ;
        RECT 89.170 188.400 89.430 188.545 ;
        RECT 88.700 187.185 88.980 187.555 ;
        RECT 89.690 187.360 89.830 189.420 ;
        RECT 90.090 188.060 90.350 188.380 ;
        RECT 89.630 187.040 89.890 187.360 ;
        RECT 90.150 186.680 90.290 188.060 ;
        RECT 90.610 187.020 90.750 190.780 ;
        RECT 90.550 186.700 90.810 187.020 ;
        RECT 90.090 186.360 90.350 186.680 ;
        RECT 91.070 186.340 91.210 192.060 ;
        RECT 91.470 191.800 91.730 192.060 ;
        RECT 92.450 191.780 92.590 192.570 ;
        RECT 92.390 191.460 92.650 191.780 ;
        RECT 91.930 191.120 92.190 191.440 ;
        RECT 91.990 189.740 92.130 191.120 ;
        RECT 91.930 189.420 92.190 189.740 ;
        RECT 92.380 189.225 92.660 189.595 ;
        RECT 91.470 188.740 91.730 189.060 ;
        RECT 92.450 188.970 92.590 189.225 ;
        RECT 91.990 188.830 92.590 188.970 ;
        RECT 90.540 185.825 90.820 186.195 ;
        RECT 91.010 186.020 91.270 186.340 ;
        RECT 90.090 185.340 90.350 185.660 ;
        RECT 88.700 183.785 88.980 184.155 ;
        RECT 88.770 183.620 88.910 183.785 ;
        RECT 88.710 183.300 88.970 183.620 ;
        RECT 89.170 182.960 89.430 183.280 ;
        RECT 89.230 182.115 89.370 182.960 ;
        RECT 88.250 181.600 88.510 181.920 ;
        RECT 89.160 181.745 89.440 182.115 ;
        RECT 88.250 179.900 88.510 180.220 ;
        RECT 87.790 175.140 88.050 175.460 ;
        RECT 86.870 174.800 87.130 175.120 ;
        RECT 86.930 173.760 87.070 174.800 ;
        RECT 88.310 174.520 88.450 179.900 ;
        RECT 88.710 175.480 88.970 175.800 ;
        RECT 87.850 174.380 88.450 174.520 ;
        RECT 86.870 173.440 87.130 173.760 ;
        RECT 86.410 172.080 86.670 172.400 ;
        RECT 85.950 171.740 86.210 172.060 ;
        RECT 86.010 171.040 86.150 171.740 ;
        RECT 85.950 170.720 86.210 171.040 ;
        RECT 85.490 170.380 85.750 170.700 ;
        RECT 85.030 166.980 85.290 167.300 ;
        RECT 85.550 165.600 85.690 170.380 ;
        RECT 86.870 169.020 87.130 169.340 ;
        RECT 86.930 167.300 87.070 169.020 ;
        RECT 86.870 166.980 87.130 167.300 ;
        RECT 85.490 165.280 85.750 165.600 ;
        RECT 85.490 164.600 85.750 164.920 ;
        RECT 85.950 164.600 86.210 164.920 ;
        RECT 84.570 162.560 84.830 162.880 ;
        RECT 83.190 161.880 83.450 162.200 ;
        RECT 84.110 161.880 84.370 162.200 ;
        RECT 83.250 161.715 83.390 161.880 ;
        RECT 83.180 161.345 83.460 161.715 ;
        RECT 83.650 160.860 83.910 161.180 ;
        RECT 83.710 157.440 83.850 160.860 ;
        RECT 84.170 159.140 84.310 161.880 ;
        RECT 85.550 161.860 85.690 164.600 ;
        RECT 86.010 162.880 86.150 164.600 ;
        RECT 87.330 163.920 87.590 164.240 ;
        RECT 87.390 163.755 87.530 163.920 ;
        RECT 87.320 163.385 87.600 163.755 ;
        RECT 85.950 162.560 86.210 162.880 ;
        RECT 84.570 161.540 84.830 161.860 ;
        RECT 85.490 161.540 85.750 161.860 ;
        RECT 84.110 158.820 84.370 159.140 ;
        RECT 83.650 157.120 83.910 157.440 ;
        RECT 82.730 156.780 82.990 157.100 ;
        RECT 84.170 156.760 84.310 158.820 ;
        RECT 84.110 156.440 84.370 156.760 ;
        RECT 82.270 154.060 82.530 154.380 ;
        RECT 81.810 152.700 82.070 153.020 ;
        RECT 81.870 151.320 82.010 152.700 ;
        RECT 84.170 151.320 84.310 156.440 ;
        RECT 84.630 151.660 84.770 161.540 ;
        RECT 85.490 158.820 85.750 159.140 ;
        RECT 87.330 158.820 87.590 159.140 ;
        RECT 85.550 154.720 85.690 158.820 ;
        RECT 86.410 155.420 86.670 155.740 ;
        RECT 85.490 154.400 85.750 154.720 ;
        RECT 86.470 154.040 86.610 155.420 ;
        RECT 86.410 153.720 86.670 154.040 ;
        RECT 85.950 153.380 86.210 153.700 ;
        RECT 86.870 153.380 87.130 153.700 ;
        RECT 86.010 152.000 86.150 153.380 ;
        RECT 85.950 151.680 86.210 152.000 ;
        RECT 84.570 151.340 84.830 151.660 ;
        RECT 81.810 151.000 82.070 151.320 ;
        RECT 84.110 151.000 84.370 151.320 ;
        RECT 82.270 149.980 82.530 150.300 ;
        RECT 83.650 149.980 83.910 150.300 ;
        RECT 81.810 149.190 82.070 149.280 ;
        RECT 81.410 149.050 82.070 149.190 ;
        RECT 81.810 148.960 82.070 149.050 ;
        RECT 82.330 147.580 82.470 149.980 ;
        RECT 83.710 148.940 83.850 149.980 ;
        RECT 83.650 148.620 83.910 148.940 ;
        RECT 82.270 147.260 82.530 147.580 ;
        RECT 82.330 145.880 82.470 147.260 ;
        RECT 84.170 146.220 84.310 151.000 ;
        RECT 84.630 150.980 84.770 151.340 ;
        RECT 84.570 150.660 84.830 150.980 ;
        RECT 85.030 150.660 85.290 150.980 ;
        RECT 85.090 146.560 85.230 150.660 ;
        RECT 85.950 149.980 86.210 150.300 ;
        RECT 86.410 149.980 86.670 150.300 ;
        RECT 86.010 148.600 86.150 149.980 ;
        RECT 85.950 148.280 86.210 148.600 ;
        RECT 86.470 147.580 86.610 149.980 ;
        RECT 86.410 147.260 86.670 147.580 ;
        RECT 85.030 146.240 85.290 146.560 ;
        RECT 84.110 145.900 84.370 146.220 ;
        RECT 85.490 145.960 85.750 146.220 ;
        RECT 85.090 145.900 85.750 145.960 ;
        RECT 82.270 145.560 82.530 145.880 ;
        RECT 85.090 145.820 85.690 145.900 ;
        RECT 86.470 145.880 86.610 147.260 ;
        RECT 85.090 145.450 85.230 145.820 ;
        RECT 86.410 145.560 86.670 145.880 ;
        RECT 84.170 145.310 85.230 145.450 ;
        RECT 81.810 144.880 82.070 145.200 ;
        RECT 81.870 143.840 82.010 144.880 ;
        RECT 81.810 143.520 82.070 143.840 ;
        RECT 82.270 142.840 82.530 143.160 ;
        RECT 81.350 138.310 81.610 138.400 ;
        RECT 80.950 138.170 81.610 138.310 ;
        RECT 81.350 138.080 81.610 138.170 ;
        RECT 82.330 137.720 82.470 142.840 ;
        RECT 83.650 141.820 83.910 142.140 ;
        RECT 82.730 140.120 82.990 140.440 ;
        RECT 82.790 137.800 82.930 140.120 ;
        RECT 83.190 139.440 83.450 139.760 ;
        RECT 83.250 138.400 83.390 139.440 ;
        RECT 83.190 138.080 83.450 138.400 ;
        RECT 82.790 137.720 83.390 137.800 ;
        RECT 82.270 137.400 82.530 137.720 ;
        RECT 82.790 137.660 83.450 137.720 ;
        RECT 83.190 137.400 83.450 137.660 ;
        RECT 83.190 136.720 83.450 137.040 ;
        RECT 83.250 133.980 83.390 136.720 ;
        RECT 83.190 133.660 83.450 133.980 ;
        RECT 83.250 132.960 83.390 133.660 ;
        RECT 83.190 132.640 83.450 132.960 ;
        RECT 80.430 129.580 80.690 129.900 ;
        RECT 79.970 128.900 80.230 129.220 ;
        RECT 83.710 126.840 83.850 141.820 ;
        RECT 84.170 141.120 84.310 145.310 ;
        RECT 85.950 144.540 86.210 144.860 ;
        RECT 84.110 140.800 84.370 141.120 ;
        RECT 84.170 137.040 84.310 140.800 ;
        RECT 86.010 140.440 86.150 144.540 ;
        RECT 86.930 142.820 87.070 153.380 ;
        RECT 87.390 148.260 87.530 158.820 ;
        RECT 87.850 158.460 87.990 174.380 ;
        RECT 88.240 167.465 88.520 167.835 ;
        RECT 88.310 164.920 88.450 167.465 ;
        RECT 88.250 164.600 88.510 164.920 ;
        RECT 88.770 164.320 88.910 175.480 ;
        RECT 89.170 169.700 89.430 170.020 ;
        RECT 89.230 167.980 89.370 169.700 ;
        RECT 89.170 167.660 89.430 167.980 ;
        RECT 89.170 167.155 89.430 167.300 ;
        RECT 89.160 166.785 89.440 167.155 ;
        RECT 89.630 164.600 89.890 164.920 ;
        RECT 88.310 164.180 88.910 164.320 ;
        RECT 88.310 160.160 88.450 164.180 ;
        RECT 88.710 163.580 88.970 163.900 ;
        RECT 89.170 163.580 89.430 163.900 ;
        RECT 88.250 159.840 88.510 160.160 ;
        RECT 88.770 159.820 88.910 163.580 ;
        RECT 88.710 159.500 88.970 159.820 ;
        RECT 88.700 158.625 88.980 158.995 ;
        RECT 87.790 158.140 88.050 158.460 ;
        RECT 88.770 156.420 88.910 158.625 ;
        RECT 88.710 156.100 88.970 156.420 ;
        RECT 87.790 155.420 88.050 155.740 ;
        RECT 87.850 149.280 87.990 155.420 ;
        RECT 88.710 150.660 88.970 150.980 ;
        RECT 87.790 148.960 88.050 149.280 ;
        RECT 87.330 147.940 87.590 148.260 ;
        RECT 87.390 143.840 87.530 147.940 ;
        RECT 87.330 143.520 87.590 143.840 ;
        RECT 86.870 142.500 87.130 142.820 ;
        RECT 86.930 140.440 87.070 142.500 ;
        RECT 85.950 140.120 86.210 140.440 ;
        RECT 86.870 140.120 87.130 140.440 ;
        RECT 88.770 138.400 88.910 150.660 ;
        RECT 89.230 142.480 89.370 163.580 ;
        RECT 89.690 158.460 89.830 164.600 ;
        RECT 89.630 158.140 89.890 158.460 ;
        RECT 89.630 157.120 89.890 157.440 ;
        RECT 89.690 145.880 89.830 157.120 ;
        RECT 90.150 156.420 90.290 185.340 ;
        RECT 90.610 183.620 90.750 185.825 ;
        RECT 90.550 183.300 90.810 183.620 ;
        RECT 90.550 182.620 90.810 182.940 ;
        RECT 90.090 156.100 90.350 156.420 ;
        RECT 90.610 154.040 90.750 182.620 ;
        RECT 91.530 174.780 91.670 188.740 ;
        RECT 91.990 187.360 92.130 188.830 ;
        RECT 92.510 187.525 94.390 187.895 ;
        RECT 91.930 187.040 92.190 187.360 ;
        RECT 93.770 186.360 94.030 186.680 ;
        RECT 93.830 186.195 93.970 186.360 ;
        RECT 93.760 185.825 94.040 186.195 ;
        RECT 94.230 186.020 94.490 186.340 ;
        RECT 94.290 183.280 94.430 186.020 ;
        RECT 94.750 186.000 94.890 196.560 ;
        RECT 95.150 194.860 95.410 195.180 ;
        RECT 94.690 185.680 94.950 186.000 ;
        RECT 94.230 182.960 94.490 183.280 ;
        RECT 94.690 182.960 94.950 183.280 ;
        RECT 92.510 182.085 94.390 182.455 ;
        RECT 94.230 181.490 94.490 181.580 ;
        RECT 94.750 181.490 94.890 182.960 ;
        RECT 94.230 181.350 94.890 181.490 ;
        RECT 94.230 181.260 94.490 181.350 ;
        RECT 94.690 180.240 94.950 180.560 ;
        RECT 94.750 179.200 94.890 180.240 ;
        RECT 94.690 178.880 94.950 179.200 ;
        RECT 92.510 176.645 94.390 177.015 ;
        RECT 94.750 176.140 94.890 178.880 ;
        RECT 94.690 175.820 94.950 176.140 ;
        RECT 91.470 174.460 91.730 174.780 ;
        RECT 94.750 172.740 94.890 175.820 ;
        RECT 91.530 172.340 92.590 172.480 ;
        RECT 94.690 172.420 94.950 172.740 ;
        RECT 91.530 170.020 91.670 172.340 ;
        RECT 92.450 172.060 92.590 172.340 ;
        RECT 91.930 171.740 92.190 172.060 ;
        RECT 92.390 171.740 92.650 172.060 ;
        RECT 91.990 171.040 92.130 171.740 ;
        RECT 92.510 171.205 94.390 171.575 ;
        RECT 91.930 170.720 92.190 171.040 ;
        RECT 91.470 169.700 91.730 170.020 ;
        RECT 91.530 167.640 91.670 169.700 ;
        RECT 91.470 167.320 91.730 167.640 ;
        RECT 91.990 167.300 92.130 170.720 ;
        RECT 93.310 170.380 93.570 170.700 ;
        RECT 93.370 168.320 93.510 170.380 ;
        RECT 94.750 170.360 94.890 172.420 ;
        RECT 94.690 170.040 94.950 170.360 ;
        RECT 93.310 168.000 93.570 168.320 ;
        RECT 94.690 168.000 94.950 168.320 ;
        RECT 91.930 166.980 92.190 167.300 ;
        RECT 91.010 166.680 91.270 166.960 ;
        RECT 91.010 166.640 91.670 166.680 ;
        RECT 91.070 166.540 91.670 166.640 ;
        RECT 91.530 165.115 91.670 166.540 ;
        RECT 91.460 164.745 91.740 165.115 ;
        RECT 91.990 164.830 92.130 166.980 ;
        RECT 92.510 165.765 94.390 166.135 ;
        RECT 92.850 165.280 93.110 165.600 ;
        RECT 92.390 164.830 92.650 164.920 ;
        RECT 91.470 164.600 91.730 164.745 ;
        RECT 91.990 164.690 92.650 164.830 ;
        RECT 92.390 164.600 92.650 164.690 ;
        RECT 92.910 164.580 93.050 165.280 ;
        RECT 94.220 164.745 94.500 165.115 ;
        RECT 94.750 165.000 94.890 168.000 ;
        RECT 95.210 165.600 95.350 194.860 ;
        RECT 95.610 194.180 95.870 194.500 ;
        RECT 95.670 193.675 95.810 194.180 ;
        RECT 95.600 193.305 95.880 193.675 ;
        RECT 95.670 186.680 95.810 193.305 ;
        RECT 96.130 186.680 96.270 200.300 ;
        RECT 96.590 196.450 96.730 202.340 ;
        RECT 97.050 200.960 97.190 202.340 ;
        RECT 96.990 200.640 97.250 200.960 ;
        RECT 97.510 198.240 97.650 202.680 ;
        RECT 98.820 202.145 99.100 202.515 ;
        RECT 99.290 202.340 99.550 202.660 ;
        RECT 97.910 199.280 98.170 199.600 ;
        RECT 96.990 197.920 97.250 198.240 ;
        RECT 97.450 197.920 97.710 198.240 ;
        RECT 97.050 197.220 97.190 197.920 ;
        RECT 96.990 196.900 97.250 197.220 ;
        RECT 96.590 196.310 97.650 196.450 ;
        RECT 96.530 194.180 96.790 194.500 ;
        RECT 97.510 194.410 97.650 196.310 ;
        RECT 97.970 195.180 98.110 199.280 ;
        RECT 98.370 198.940 98.630 199.260 ;
        RECT 97.910 194.860 98.170 195.180 ;
        RECT 97.510 194.270 98.110 194.410 ;
        RECT 96.590 186.680 96.730 194.180 ;
        RECT 96.990 193.500 97.250 193.820 ;
        RECT 97.050 192.800 97.190 193.500 ;
        RECT 96.990 192.480 97.250 192.800 ;
        RECT 97.970 192.200 98.110 194.270 ;
        RECT 97.510 192.060 98.110 192.200 ;
        RECT 97.510 191.780 97.650 192.060 ;
        RECT 98.430 191.780 98.570 198.940 ;
        RECT 98.890 197.900 99.030 202.145 ;
        RECT 99.350 198.150 99.490 202.340 ;
        RECT 99.810 200.280 99.950 206.760 ;
        RECT 101.120 205.545 101.400 205.915 ;
        RECT 111.250 205.740 111.510 206.060 ;
        RECT 100.210 203.360 100.470 203.680 ;
        RECT 99.750 199.960 100.010 200.280 ;
        RECT 99.350 198.010 99.950 198.150 ;
        RECT 98.830 197.580 99.090 197.900 ;
        RECT 99.810 197.220 99.950 198.010 ;
        RECT 100.270 197.560 100.410 203.360 ;
        RECT 100.670 202.000 100.930 202.320 ;
        RECT 100.210 197.240 100.470 197.560 ;
        RECT 98.830 196.900 99.090 197.220 ;
        RECT 99.750 196.900 100.010 197.220 ;
        RECT 98.890 194.160 99.030 196.900 ;
        RECT 99.750 196.220 100.010 196.540 ;
        RECT 99.810 194.840 99.950 196.220 ;
        RECT 100.730 195.520 100.870 202.000 ;
        RECT 101.190 195.520 101.330 205.545 ;
        RECT 105.260 204.865 105.540 205.235 ;
        RECT 105.330 199.940 105.470 204.865 ;
        RECT 107.110 204.720 107.370 205.040 ;
        RECT 105.270 199.620 105.530 199.940 ;
        RECT 106.650 199.620 106.910 199.940 ;
        RECT 104.340 196.705 104.620 197.075 ;
        RECT 105.270 196.900 105.530 197.220 ;
        RECT 101.590 196.395 101.850 196.540 ;
        RECT 101.580 196.025 101.860 196.395 ;
        RECT 100.670 195.200 100.930 195.520 ;
        RECT 101.130 195.200 101.390 195.520 ;
        RECT 99.750 194.520 100.010 194.840 ;
        RECT 98.830 193.840 99.090 194.160 ;
        RECT 99.810 193.820 99.950 194.520 ;
        RECT 100.210 193.840 100.470 194.160 ;
        RECT 101.120 193.985 101.400 194.355 ;
        RECT 102.510 194.180 102.770 194.500 ;
        RECT 99.750 193.500 100.010 193.820 ;
        RECT 98.830 191.800 99.090 192.120 ;
        RECT 96.980 191.265 97.260 191.635 ;
        RECT 97.450 191.460 97.710 191.780 ;
        RECT 97.910 191.460 98.170 191.780 ;
        RECT 98.370 191.460 98.630 191.780 ;
        RECT 97.050 189.400 97.190 191.265 ;
        RECT 97.450 190.780 97.710 191.100 ;
        RECT 96.990 189.080 97.250 189.400 ;
        RECT 95.610 186.360 95.870 186.680 ;
        RECT 96.070 186.360 96.330 186.680 ;
        RECT 96.530 186.360 96.790 186.680 ;
        RECT 96.590 184.155 96.730 186.360 ;
        RECT 97.510 186.250 97.650 190.780 ;
        RECT 97.970 187.020 98.110 191.460 ;
        RECT 98.430 189.400 98.570 191.460 ;
        RECT 98.370 189.080 98.630 189.400 ;
        RECT 98.890 188.800 99.030 191.800 ;
        RECT 99.290 191.120 99.550 191.440 ;
        RECT 98.430 188.660 99.030 188.800 ;
        RECT 97.910 186.700 98.170 187.020 ;
        RECT 97.510 186.110 98.110 186.250 ;
        RECT 96.520 183.785 96.800 184.155 ;
        RECT 96.990 183.980 97.250 184.300 ;
        RECT 96.070 183.300 96.330 183.620 ;
        RECT 95.610 180.920 95.870 181.240 ;
        RECT 95.670 177.500 95.810 180.920 ;
        RECT 96.130 180.900 96.270 183.300 ;
        RECT 96.530 182.620 96.790 182.940 ;
        RECT 96.590 181.240 96.730 182.620 ;
        RECT 96.530 180.920 96.790 181.240 ;
        RECT 96.070 180.580 96.330 180.900 ;
        RECT 95.610 177.180 95.870 177.500 ;
        RECT 95.610 175.140 95.870 175.460 ;
        RECT 95.670 172.060 95.810 175.140 ;
        RECT 95.610 171.740 95.870 172.060 ;
        RECT 95.610 170.040 95.870 170.360 ;
        RECT 95.670 166.960 95.810 170.040 ;
        RECT 95.610 166.640 95.870 166.960 ;
        RECT 95.150 165.280 95.410 165.600 ;
        RECT 94.750 164.860 95.810 165.000 ;
        RECT 96.130 164.920 96.270 180.580 ;
        RECT 96.590 176.480 96.730 180.920 ;
        RECT 96.530 176.160 96.790 176.480 ;
        RECT 96.520 175.625 96.800 175.995 ;
        RECT 94.230 164.600 94.490 164.745 ;
        RECT 92.850 164.260 93.110 164.580 ;
        RECT 91.010 163.580 91.270 163.900 ;
        RECT 94.690 163.580 94.950 163.900 ;
        RECT 91.070 154.040 91.210 163.580 ;
        RECT 93.300 162.025 93.580 162.395 ;
        RECT 93.310 161.880 93.570 162.025 ;
        RECT 91.470 160.860 91.730 161.180 ;
        RECT 91.930 160.860 92.190 161.180 ;
        RECT 91.530 159.820 91.670 160.860 ;
        RECT 91.470 159.500 91.730 159.820 ;
        RECT 91.990 159.050 92.130 160.860 ;
        RECT 92.510 160.325 94.390 160.695 ;
        RECT 94.220 159.305 94.500 159.675 ;
        RECT 91.530 158.910 92.130 159.050 ;
        RECT 91.530 156.420 91.670 158.910 ;
        RECT 92.390 158.820 92.650 159.140 ;
        RECT 91.930 157.120 92.190 157.440 ;
        RECT 91.470 156.100 91.730 156.420 ;
        RECT 90.550 153.720 90.810 154.040 ;
        RECT 91.010 153.720 91.270 154.040 ;
        RECT 91.990 153.440 92.130 157.120 ;
        RECT 92.450 155.740 92.590 158.820 ;
        RECT 93.770 156.440 94.030 156.760 ;
        RECT 93.830 156.275 93.970 156.440 ;
        RECT 94.290 156.420 94.430 159.305 ;
        RECT 94.750 158.995 94.890 163.580 ;
        RECT 95.150 161.540 95.410 161.860 ;
        RECT 94.680 158.625 94.960 158.995 ;
        RECT 95.210 157.100 95.350 161.540 ;
        RECT 95.150 156.955 95.410 157.100 ;
        RECT 95.140 156.585 95.420 156.955 ;
        RECT 95.210 156.420 95.350 156.585 ;
        RECT 93.760 155.905 94.040 156.275 ;
        RECT 94.230 156.100 94.490 156.420 ;
        RECT 95.150 156.330 95.410 156.420 ;
        RECT 94.750 156.190 95.410 156.330 ;
        RECT 92.390 155.420 92.650 155.740 ;
        RECT 92.510 154.885 94.390 155.255 ;
        RECT 94.750 154.720 94.890 156.190 ;
        RECT 95.150 156.100 95.410 156.190 ;
        RECT 95.150 155.420 95.410 155.740 ;
        RECT 94.690 154.400 94.950 154.720 ;
        RECT 94.690 153.720 94.950 154.040 ;
        RECT 94.750 153.440 94.890 153.720 ;
        RECT 91.990 153.300 92.590 153.440 ;
        RECT 92.450 153.020 92.590 153.300 ;
        RECT 94.290 153.300 94.890 153.440 ;
        RECT 90.550 152.700 90.810 153.020 ;
        RECT 91.930 152.700 92.190 153.020 ;
        RECT 92.390 152.700 92.650 153.020 ;
        RECT 90.610 152.000 90.750 152.700 ;
        RECT 90.550 151.680 90.810 152.000 ;
        RECT 91.010 151.340 91.270 151.660 ;
        RECT 91.070 147.580 91.210 151.340 ;
        RECT 91.470 150.320 91.730 150.640 ;
        RECT 91.010 147.260 91.270 147.580 ;
        RECT 89.630 145.560 89.890 145.880 ;
        RECT 91.070 145.450 91.210 147.260 ;
        RECT 91.530 146.220 91.670 150.320 ;
        RECT 91.470 145.900 91.730 146.220 ;
        RECT 91.470 145.450 91.730 145.540 ;
        RECT 91.070 145.310 91.730 145.450 ;
        RECT 91.470 145.220 91.730 145.310 ;
        RECT 89.630 144.540 89.890 144.860 ;
        RECT 89.690 143.500 89.830 144.540 ;
        RECT 89.630 143.180 89.890 143.500 ;
        RECT 89.170 142.160 89.430 142.480 ;
        RECT 89.690 141.120 89.830 143.180 ;
        RECT 89.630 140.800 89.890 141.120 ;
        RECT 91.010 139.440 91.270 139.760 ;
        RECT 88.710 138.080 88.970 138.400 ;
        RECT 87.790 137.400 88.050 137.720 ;
        RECT 84.570 137.060 84.830 137.380 ;
        RECT 84.110 136.720 84.370 137.040 ;
        RECT 84.170 135.000 84.310 136.720 ;
        RECT 84.110 134.680 84.370 135.000 ;
        RECT 84.630 134.320 84.770 137.060 ;
        RECT 86.410 136.380 86.670 136.700 ;
        RECT 86.470 134.660 86.610 136.380 ;
        RECT 86.410 134.340 86.670 134.660 ;
        RECT 84.570 134.000 84.830 134.320 ;
        RECT 84.630 132.960 84.770 134.000 ;
        RECT 84.570 132.640 84.830 132.960 ;
        RECT 85.950 132.300 86.210 132.620 ;
        RECT 86.010 130.240 86.150 132.300 ;
        RECT 85.950 129.920 86.210 130.240 ;
        RECT 87.850 129.900 87.990 137.400 ;
        RECT 88.770 137.120 88.910 138.080 ;
        RECT 88.310 136.980 88.910 137.120 ;
        RECT 88.310 135.680 88.450 136.980 ;
        RECT 88.710 136.380 88.970 136.700 ;
        RECT 90.550 136.380 90.810 136.700 ;
        RECT 88.250 135.360 88.510 135.680 ;
        RECT 87.790 129.580 88.050 129.900 ;
        RECT 88.770 129.220 88.910 136.380 ;
        RECT 90.610 134.320 90.750 136.380 ;
        RECT 90.550 134.000 90.810 134.320 ;
        RECT 89.630 131.620 89.890 131.940 ;
        RECT 89.690 130.240 89.830 131.620 ;
        RECT 91.070 130.240 91.210 139.440 ;
        RECT 89.630 129.920 89.890 130.240 ;
        RECT 91.010 129.920 91.270 130.240 ;
        RECT 91.990 129.560 92.130 152.700 ;
        RECT 94.290 150.640 94.430 153.300 ;
        RECT 94.690 152.700 94.950 153.020 ;
        RECT 94.750 151.660 94.890 152.700 ;
        RECT 94.690 151.340 94.950 151.660 ;
        RECT 94.230 150.320 94.490 150.640 ;
        RECT 94.690 149.980 94.950 150.300 ;
        RECT 92.510 149.445 94.390 149.815 ;
        RECT 92.390 148.620 92.650 148.940 ;
        RECT 92.450 146.560 92.590 148.620 ;
        RECT 92.390 146.240 92.650 146.560 ;
        RECT 92.510 144.005 94.390 144.375 ;
        RECT 94.750 143.160 94.890 149.980 ;
        RECT 93.310 142.840 93.570 143.160 ;
        RECT 94.690 142.840 94.950 143.160 ;
        RECT 93.370 140.635 93.510 142.840 ;
        RECT 95.210 142.560 95.350 155.420 ;
        RECT 95.670 150.980 95.810 164.860 ;
        RECT 96.070 164.600 96.330 164.920 ;
        RECT 96.070 161.540 96.330 161.860 ;
        RECT 96.130 161.035 96.270 161.540 ;
        RECT 96.590 161.520 96.730 175.625 ;
        RECT 96.530 161.200 96.790 161.520 ;
        RECT 96.060 160.665 96.340 161.035 ;
        RECT 96.130 159.140 96.270 160.665 ;
        RECT 96.590 159.820 96.730 161.200 ;
        RECT 96.530 159.500 96.790 159.820 ;
        RECT 96.070 158.820 96.330 159.140 ;
        RECT 96.530 158.820 96.790 159.140 ;
        RECT 96.070 155.650 96.330 155.740 ;
        RECT 96.590 155.650 96.730 158.820 ;
        RECT 96.070 155.510 96.730 155.650 ;
        RECT 96.070 155.420 96.330 155.510 ;
        RECT 96.130 153.700 96.270 155.420 ;
        RECT 96.070 153.380 96.330 153.700 ;
        RECT 96.530 153.380 96.790 153.700 ;
        RECT 96.590 151.320 96.730 153.380 ;
        RECT 97.050 151.320 97.190 183.980 ;
        RECT 97.450 183.475 97.710 183.620 ;
        RECT 97.440 183.105 97.720 183.475 ;
        RECT 97.450 180.580 97.710 180.900 ;
        RECT 97.510 175.460 97.650 180.580 ;
        RECT 97.970 178.180 98.110 186.110 ;
        RECT 97.910 177.860 98.170 178.180 ;
        RECT 97.450 175.140 97.710 175.460 ;
        RECT 98.430 171.040 98.570 188.660 ;
        RECT 98.830 186.700 99.090 187.020 ;
        RECT 98.890 184.155 99.030 186.700 ;
        RECT 98.820 183.785 99.100 184.155 ;
        RECT 98.890 179.200 99.030 183.785 ;
        RECT 98.830 178.880 99.090 179.200 ;
        RECT 99.350 173.420 99.490 191.120 ;
        RECT 99.750 188.740 100.010 189.060 ;
        RECT 99.810 176.480 99.950 188.740 ;
        RECT 100.270 188.380 100.410 193.840 ;
        RECT 101.190 188.720 101.330 193.985 ;
        RECT 101.590 191.800 101.850 192.120 ;
        RECT 101.130 188.400 101.390 188.720 ;
        RECT 100.210 188.060 100.470 188.380 ;
        RECT 100.670 188.060 100.930 188.380 ;
        RECT 100.270 187.020 100.410 188.060 ;
        RECT 100.730 187.360 100.870 188.060 ;
        RECT 100.670 187.040 100.930 187.360 ;
        RECT 100.210 186.700 100.470 187.020 ;
        RECT 100.210 186.020 100.470 186.340 ;
        RECT 100.270 184.155 100.410 186.020 ;
        RECT 100.200 183.785 100.480 184.155 ;
        RECT 100.730 183.960 100.870 187.040 ;
        RECT 101.120 186.760 101.400 186.875 ;
        RECT 101.650 186.760 101.790 191.800 ;
        RECT 101.120 186.620 101.790 186.760 ;
        RECT 101.120 186.505 101.400 186.620 ;
        RECT 101.190 186.340 101.330 186.505 ;
        RECT 102.570 186.340 102.710 194.180 ;
        RECT 104.410 192.460 104.550 196.705 ;
        RECT 105.330 195.180 105.470 196.900 ;
        RECT 106.180 195.345 106.460 195.715 ;
        RECT 105.270 194.860 105.530 195.180 ;
        RECT 104.810 194.520 105.070 194.840 ;
        RECT 103.890 192.315 104.150 192.460 ;
        RECT 103.880 191.945 104.160 192.315 ;
        RECT 104.350 192.140 104.610 192.460 ;
        RECT 104.870 186.680 105.010 194.520 ;
        RECT 106.250 194.500 106.390 195.345 ;
        RECT 106.190 194.180 106.450 194.500 ;
        RECT 105.270 193.500 105.530 193.820 ;
        RECT 104.810 186.360 105.070 186.680 ;
        RECT 101.130 186.020 101.390 186.340 ;
        RECT 102.510 186.020 102.770 186.340 ;
        RECT 102.970 186.020 103.230 186.340 ;
        RECT 103.030 184.300 103.170 186.020 ;
        RECT 104.340 185.825 104.620 186.195 ;
        RECT 102.970 183.980 103.230 184.300 ;
        RECT 100.670 183.640 100.930 183.960 ;
        RECT 100.210 183.300 100.470 183.620 ;
        RECT 102.970 183.300 103.230 183.620 ;
        RECT 100.270 177.500 100.410 183.300 ;
        RECT 102.510 182.620 102.770 182.940 ;
        RECT 101.590 181.260 101.850 181.580 ;
        RECT 100.670 180.240 100.930 180.560 ;
        RECT 100.210 177.180 100.470 177.500 ;
        RECT 99.750 176.160 100.010 176.480 ;
        RECT 100.730 175.120 100.870 180.240 ;
        RECT 101.130 179.900 101.390 180.220 ;
        RECT 101.190 175.800 101.330 179.900 ;
        RECT 101.130 175.480 101.390 175.800 ;
        RECT 101.650 175.315 101.790 181.260 ;
        RECT 102.050 176.160 102.310 176.480 ;
        RECT 100.670 174.800 100.930 175.120 ;
        RECT 101.580 174.945 101.860 175.315 ;
        RECT 99.290 173.100 99.550 173.420 ;
        RECT 98.830 172.760 99.090 173.080 ;
        RECT 100.730 172.990 100.870 174.800 ;
        RECT 100.270 172.850 100.870 172.990 ;
        RECT 101.590 172.990 101.850 173.080 ;
        RECT 102.110 172.990 102.250 176.160 ;
        RECT 102.570 175.800 102.710 182.620 ;
        RECT 102.510 175.480 102.770 175.800 ;
        RECT 103.030 173.420 103.170 183.300 ;
        RECT 104.410 180.220 104.550 185.825 ;
        RECT 104.350 180.130 104.610 180.220 ;
        RECT 103.950 179.990 104.610 180.130 ;
        RECT 103.430 178.540 103.690 178.860 ;
        RECT 103.490 173.760 103.630 178.540 ;
        RECT 103.430 173.440 103.690 173.760 ;
        RECT 102.970 173.100 103.230 173.420 ;
        RECT 103.950 173.080 104.090 179.990 ;
        RECT 104.350 179.900 104.610 179.990 ;
        RECT 104.350 177.860 104.610 178.180 ;
        RECT 101.590 172.850 102.250 172.990 ;
        RECT 98.370 170.720 98.630 171.040 ;
        RECT 98.370 170.270 98.630 170.360 ;
        RECT 97.510 170.130 98.630 170.270 ;
        RECT 97.510 168.320 97.650 170.130 ;
        RECT 98.370 170.040 98.630 170.130 ;
        RECT 98.370 169.020 98.630 169.340 ;
        RECT 97.450 168.000 97.710 168.320 ;
        RECT 97.510 167.300 97.650 168.000 ;
        RECT 97.910 167.660 98.170 167.980 ;
        RECT 97.450 166.980 97.710 167.300 ;
        RECT 97.510 165.260 97.650 166.980 ;
        RECT 97.970 165.600 98.110 167.660 ;
        RECT 97.910 165.280 98.170 165.600 ;
        RECT 97.450 164.940 97.710 165.260 ;
        RECT 98.430 164.920 98.570 169.020 ;
        RECT 98.890 167.980 99.030 172.760 ;
        RECT 99.290 172.420 99.550 172.740 ;
        RECT 99.350 170.360 99.490 172.420 ;
        RECT 99.290 170.040 99.550 170.360 ;
        RECT 99.740 170.185 100.020 170.555 ;
        RECT 99.750 170.040 100.010 170.185 ;
        RECT 99.290 169.020 99.550 169.340 ;
        RECT 98.830 167.660 99.090 167.980 ;
        RECT 98.830 166.980 99.090 167.300 ;
        RECT 98.370 164.600 98.630 164.920 ;
        RECT 98.890 164.580 99.030 166.980 ;
        RECT 98.830 164.260 99.090 164.580 ;
        RECT 97.450 163.580 97.710 163.900 ;
        RECT 98.370 163.580 98.630 163.900 ;
        RECT 98.830 163.580 99.090 163.900 ;
        RECT 97.510 158.460 97.650 163.580 ;
        RECT 97.910 160.860 98.170 161.180 ;
        RECT 97.970 159.480 98.110 160.860 ;
        RECT 97.910 159.160 98.170 159.480 ;
        RECT 97.450 158.140 97.710 158.460 ;
        RECT 97.970 157.100 98.110 159.160 ;
        RECT 97.440 156.585 97.720 156.955 ;
        RECT 97.910 156.780 98.170 157.100 ;
        RECT 97.510 156.420 97.650 156.585 ;
        RECT 97.970 156.420 98.110 156.780 ;
        RECT 97.450 156.100 97.710 156.420 ;
        RECT 97.910 156.100 98.170 156.420 ;
        RECT 97.510 154.720 97.650 156.100 ;
        RECT 97.910 155.420 98.170 155.740 ;
        RECT 97.450 154.400 97.710 154.720 ;
        RECT 97.450 151.680 97.710 152.000 ;
        RECT 96.530 151.000 96.790 151.320 ;
        RECT 96.990 151.000 97.250 151.320 ;
        RECT 95.610 150.660 95.870 150.980 ;
        RECT 96.530 149.980 96.790 150.300 ;
        RECT 96.070 148.280 96.330 148.600 ;
        RECT 95.610 145.220 95.870 145.540 ;
        RECT 94.750 142.420 95.350 142.560 ;
        RECT 93.300 140.265 93.580 140.635 ;
        RECT 92.510 138.565 94.390 138.935 ;
        RECT 92.510 133.125 94.390 133.495 ;
        RECT 91.930 129.240 92.190 129.560 ;
        RECT 94.750 129.220 94.890 142.420 ;
        RECT 95.150 141.820 95.410 142.140 ;
        RECT 95.210 140.440 95.350 141.820 ;
        RECT 95.150 140.120 95.410 140.440 ;
        RECT 95.670 137.720 95.810 145.220 ;
        RECT 96.130 143.840 96.270 148.280 ;
        RECT 96.070 143.520 96.330 143.840 ;
        RECT 96.070 142.500 96.330 142.820 ;
        RECT 96.130 140.440 96.270 142.500 ;
        RECT 96.070 140.120 96.330 140.440 ;
        RECT 95.610 137.400 95.870 137.720 ;
        RECT 96.130 137.380 96.270 140.120 ;
        RECT 96.070 137.060 96.330 137.380 ;
        RECT 95.610 136.380 95.870 136.700 ;
        RECT 95.150 134.340 95.410 134.660 ;
        RECT 95.210 132.960 95.350 134.340 ;
        RECT 95.150 132.640 95.410 132.960 ;
        RECT 95.670 132.280 95.810 136.380 ;
        RECT 95.610 131.960 95.870 132.280 ;
        RECT 96.130 131.940 96.270 137.060 ;
        RECT 96.070 131.620 96.330 131.940 ;
        RECT 88.710 128.900 88.970 129.220 ;
        RECT 94.690 128.900 94.950 129.220 ;
        RECT 86.870 128.560 87.130 128.880 ;
        RECT 84.110 126.860 84.370 127.180 ;
        RECT 83.650 126.520 83.910 126.840 ;
        RECT 76.290 126.180 76.550 126.500 ;
        RECT 76.750 126.180 77.010 126.500 ;
        RECT 76.350 124.800 76.490 126.180 ;
        RECT 76.290 124.480 76.550 124.800 ;
        RECT 75.370 123.800 75.630 124.120 ;
        RECT 76.350 123.520 76.490 124.480 ;
        RECT 76.810 124.200 76.950 126.180 ;
        RECT 77.510 124.965 79.390 125.335 ;
        RECT 84.170 124.800 84.310 126.860 ;
        RECT 84.110 124.480 84.370 124.800 ;
        RECT 76.810 124.060 77.410 124.200 ;
        RECT 76.350 123.380 76.950 123.520 ;
        RECT 76.810 121.400 76.950 123.380 ;
        RECT 74.910 121.080 75.170 121.400 ;
        RECT 76.750 121.080 77.010 121.400 ;
        RECT 77.270 120.800 77.410 124.060 ;
        RECT 86.930 123.780 87.070 128.560 ;
        RECT 91.470 128.220 91.730 128.540 ;
        RECT 95.150 128.220 95.410 128.540 ;
        RECT 96.070 128.220 96.330 128.540 ;
        RECT 91.530 127.180 91.670 128.220 ;
        RECT 92.510 127.685 94.390 128.055 ;
        RECT 95.210 127.180 95.350 128.220 ;
        RECT 91.470 126.860 91.730 127.180 ;
        RECT 95.150 126.860 95.410 127.180 ;
        RECT 91.010 125.840 91.270 126.160 ;
        RECT 87.330 125.500 87.590 125.820 ;
        RECT 87.390 124.120 87.530 125.500 ;
        RECT 87.330 123.800 87.590 124.120 ;
        RECT 86.870 123.520 87.130 123.780 ;
        RECT 86.870 123.460 87.530 123.520 ;
        RECT 86.930 123.380 87.530 123.460 ;
        RECT 86.410 122.780 86.670 123.100 ;
        RECT 86.870 122.780 87.130 123.100 ;
        RECT 86.470 121.740 86.610 122.780 ;
        RECT 86.410 121.420 86.670 121.740 ;
        RECT 76.810 120.660 77.410 120.800 ;
        RECT 81.810 120.740 82.070 121.060 ;
        RECT 86.930 120.800 87.070 122.780 ;
        RECT 87.390 121.400 87.530 123.380 ;
        RECT 88.250 123.120 88.510 123.440 ;
        RECT 88.310 122.080 88.450 123.120 ;
        RECT 88.250 121.760 88.510 122.080 ;
        RECT 87.330 121.080 87.590 121.400 ;
        RECT 76.810 118.760 76.950 120.660 ;
        RECT 77.510 119.525 79.390 119.895 ;
        RECT 76.810 118.620 77.410 118.760 ;
        RECT 77.270 108.580 77.410 118.620 ;
        RECT 81.870 108.580 82.010 120.740 ;
        RECT 86.470 120.660 87.070 120.800 ;
        RECT 86.470 108.580 86.610 120.660 ;
        RECT 91.070 108.580 91.210 125.840 ;
        RECT 92.510 122.245 94.390 122.615 ;
        RECT 96.130 121.740 96.270 128.220 ;
        RECT 96.590 126.500 96.730 149.980 ;
        RECT 96.990 147.940 97.250 148.260 ;
        RECT 97.050 140.440 97.190 147.940 ;
        RECT 97.510 146.560 97.650 151.680 ;
        RECT 97.970 150.980 98.110 155.420 ;
        RECT 97.910 150.660 98.170 150.980 ;
        RECT 97.450 146.240 97.710 146.560 ;
        RECT 98.430 145.880 98.570 163.580 ;
        RECT 98.890 162.880 99.030 163.580 ;
        RECT 98.830 162.560 99.090 162.880 ;
        RECT 98.890 161.860 99.030 162.560 ;
        RECT 98.830 161.540 99.090 161.860 ;
        RECT 99.350 159.675 99.490 169.020 ;
        RECT 99.810 167.980 99.950 170.040 ;
        RECT 100.270 170.020 100.410 172.850 ;
        RECT 101.590 172.760 101.850 172.850 ;
        RECT 103.890 172.760 104.150 173.080 ;
        RECT 100.670 172.080 100.930 172.400 ;
        RECT 100.210 169.700 100.470 170.020 ;
        RECT 99.750 167.660 100.010 167.980 ;
        RECT 100.270 167.300 100.410 169.700 ;
        RECT 100.210 166.980 100.470 167.300 ;
        RECT 100.210 166.300 100.470 166.620 ;
        RECT 100.270 164.920 100.410 166.300 ;
        RECT 99.750 164.600 100.010 164.920 ;
        RECT 100.210 164.600 100.470 164.920 ;
        RECT 99.810 162.880 99.950 164.600 ;
        RECT 99.750 162.560 100.010 162.880 ;
        RECT 100.210 162.110 100.470 162.200 ;
        RECT 99.810 161.970 100.470 162.110 ;
        RECT 99.280 159.305 99.560 159.675 ;
        RECT 99.810 159.050 99.950 161.970 ;
        RECT 100.210 161.880 100.470 161.970 ;
        RECT 100.210 159.160 100.470 159.480 ;
        RECT 99.350 158.910 99.950 159.050 ;
        RECT 99.350 156.420 99.490 158.910 ;
        RECT 99.750 157.120 100.010 157.440 ;
        RECT 99.290 156.275 99.550 156.420 ;
        RECT 99.280 155.905 99.560 156.275 ;
        RECT 98.830 155.420 99.090 155.740 ;
        RECT 98.890 154.040 99.030 155.420 ;
        RECT 99.290 154.630 99.550 154.720 ;
        RECT 99.810 154.630 99.950 157.120 ;
        RECT 100.270 156.955 100.410 159.160 ;
        RECT 100.200 156.585 100.480 156.955 ;
        RECT 100.270 156.420 100.410 156.585 ;
        RECT 100.210 156.100 100.470 156.420 ;
        RECT 99.290 154.490 99.950 154.630 ;
        RECT 99.290 154.400 99.550 154.490 ;
        RECT 98.830 153.720 99.090 154.040 ;
        RECT 98.890 153.020 99.030 153.720 ;
        RECT 99.290 153.380 99.550 153.700 ;
        RECT 98.830 152.700 99.090 153.020 ;
        RECT 99.350 151.660 99.490 153.380 ;
        RECT 100.730 152.000 100.870 172.080 ;
        RECT 101.650 170.020 101.790 172.760 ;
        RECT 104.410 172.480 104.550 177.860 ;
        RECT 104.810 177.180 105.070 177.500 ;
        RECT 103.950 172.340 104.550 172.480 ;
        RECT 102.050 170.720 102.310 171.040 ;
        RECT 102.110 170.360 102.250 170.720 ;
        RECT 102.050 170.040 102.310 170.360 ;
        RECT 102.510 170.040 102.770 170.360 ;
        RECT 103.420 170.185 103.700 170.555 ;
        RECT 103.430 170.040 103.690 170.185 ;
        RECT 101.590 169.700 101.850 170.020 ;
        RECT 102.110 169.340 102.250 170.040 ;
        RECT 102.050 169.020 102.310 169.340 ;
        RECT 102.570 168.320 102.710 170.040 ;
        RECT 102.510 168.000 102.770 168.320 ;
        RECT 102.970 166.980 103.230 167.300 ;
        RECT 101.590 166.640 101.850 166.960 ;
        RECT 101.650 159.480 101.790 166.640 ;
        RECT 102.050 166.300 102.310 166.620 ;
        RECT 102.110 163.900 102.250 166.300 ;
        RECT 102.050 163.580 102.310 163.900 ;
        RECT 102.050 161.880 102.310 162.200 ;
        RECT 102.500 162.025 102.780 162.395 ;
        RECT 101.590 159.160 101.850 159.480 ;
        RECT 102.110 159.140 102.250 161.880 ;
        RECT 102.570 161.520 102.710 162.025 ;
        RECT 102.510 161.200 102.770 161.520 ;
        RECT 102.510 159.500 102.770 159.820 ;
        RECT 102.050 158.820 102.310 159.140 ;
        RECT 101.130 158.140 101.390 158.460 ;
        RECT 100.670 151.680 100.930 152.000 ;
        RECT 99.290 151.340 99.550 151.660 ;
        RECT 100.200 151.145 100.480 151.515 ;
        RECT 100.270 150.980 100.410 151.145 ;
        RECT 99.290 150.660 99.550 150.980 ;
        RECT 99.750 150.660 100.010 150.980 ;
        RECT 100.210 150.660 100.470 150.980 ;
        RECT 98.830 147.260 99.090 147.580 ;
        RECT 98.370 145.560 98.630 145.880 ;
        RECT 97.450 144.540 97.710 144.860 ;
        RECT 97.510 142.820 97.650 144.540 ;
        RECT 97.450 142.500 97.710 142.820 ;
        RECT 96.990 140.120 97.250 140.440 ;
        RECT 97.050 135.000 97.190 140.120 ;
        RECT 98.370 138.080 98.630 138.400 ;
        RECT 97.910 137.400 98.170 137.720 ;
        RECT 97.970 135.680 98.110 137.400 ;
        RECT 97.910 135.360 98.170 135.680 ;
        RECT 96.990 134.680 97.250 135.000 ;
        RECT 97.050 132.620 97.190 134.680 ;
        RECT 98.430 132.960 98.570 138.080 ;
        RECT 98.890 134.320 99.030 147.260 ;
        RECT 99.350 146.220 99.490 150.660 ;
        RECT 99.290 145.900 99.550 146.220 ;
        RECT 99.810 145.960 99.950 150.660 ;
        RECT 99.350 145.540 99.490 145.900 ;
        RECT 99.810 145.820 100.410 145.960 ;
        RECT 99.290 145.220 99.550 145.540 ;
        RECT 99.750 144.880 100.010 145.200 ;
        RECT 99.810 143.840 99.950 144.880 ;
        RECT 99.750 143.520 100.010 143.840 ;
        RECT 99.290 142.840 99.550 143.160 ;
        RECT 99.350 140.440 99.490 142.840 ;
        RECT 99.290 140.120 99.550 140.440 ;
        RECT 99.290 139.100 99.550 139.420 ;
        RECT 98.830 134.000 99.090 134.320 ;
        RECT 98.370 132.640 98.630 132.960 ;
        RECT 96.990 132.300 97.250 132.620 ;
        RECT 97.050 129.900 97.190 132.300 ;
        RECT 98.360 132.105 98.640 132.475 ;
        RECT 96.990 129.580 97.250 129.900 ;
        RECT 97.050 127.180 97.190 129.580 ;
        RECT 98.430 129.220 98.570 132.105 ;
        RECT 99.350 131.940 99.490 139.100 ;
        RECT 100.270 138.400 100.410 145.820 ;
        RECT 100.670 145.560 100.930 145.880 ;
        RECT 100.730 143.500 100.870 145.560 ;
        RECT 100.670 143.180 100.930 143.500 ;
        RECT 100.210 138.080 100.470 138.400 ;
        RECT 99.750 136.380 100.010 136.700 ;
        RECT 99.810 132.280 99.950 136.380 ;
        RECT 99.750 131.960 100.010 132.280 ;
        RECT 99.290 131.620 99.550 131.940 ;
        RECT 98.370 128.900 98.630 129.220 ;
        RECT 98.830 128.560 99.090 128.880 ;
        RECT 96.990 126.860 97.250 127.180 ;
        RECT 97.910 126.520 98.170 126.840 ;
        RECT 96.530 126.180 96.790 126.500 ;
        RECT 97.970 124.120 98.110 126.520 ;
        RECT 98.370 125.500 98.630 125.820 ;
        RECT 97.910 123.800 98.170 124.120 ;
        RECT 97.970 123.100 98.110 123.800 ;
        RECT 97.910 122.780 98.170 123.100 ;
        RECT 96.070 121.420 96.330 121.740 ;
        RECT 97.970 121.060 98.110 122.780 ;
        RECT 98.430 121.740 98.570 125.500 ;
        RECT 98.890 124.120 99.030 128.560 ;
        RECT 99.290 128.220 99.550 128.540 ;
        RECT 100.670 128.220 100.930 128.540 ;
        RECT 99.350 127.520 99.490 128.220 ;
        RECT 99.290 127.200 99.550 127.520 ;
        RECT 98.830 123.800 99.090 124.120 ;
        RECT 100.730 123.440 100.870 128.220 ;
        RECT 101.190 124.800 101.330 158.140 ;
        RECT 101.590 155.420 101.850 155.740 ;
        RECT 101.650 154.380 101.790 155.420 ;
        RECT 101.590 154.060 101.850 154.380 ;
        RECT 102.110 151.320 102.250 158.820 ;
        RECT 102.570 156.420 102.710 159.500 ;
        RECT 102.510 156.100 102.770 156.420 ;
        RECT 102.050 151.000 102.310 151.320 ;
        RECT 102.510 149.980 102.770 150.300 ;
        RECT 102.570 149.280 102.710 149.980 ;
        RECT 102.510 148.960 102.770 149.280 ;
        RECT 103.030 147.920 103.170 166.980 ;
        RECT 103.430 161.035 103.690 161.180 ;
        RECT 103.420 160.665 103.700 161.035 ;
        RECT 103.430 152.700 103.690 153.020 ;
        RECT 103.490 150.980 103.630 152.700 ;
        RECT 103.430 150.660 103.690 150.980 ;
        RECT 102.970 147.600 103.230 147.920 ;
        RECT 103.030 145.540 103.170 147.600 ;
        RECT 103.950 146.220 104.090 172.340 ;
        RECT 104.870 172.060 105.010 177.180 ;
        RECT 105.330 175.880 105.470 193.500 ;
        RECT 106.250 190.080 106.390 194.180 ;
        RECT 106.190 189.760 106.450 190.080 ;
        RECT 105.730 189.080 105.990 189.400 ;
        RECT 105.790 180.900 105.930 189.080 ;
        RECT 106.710 186.000 106.850 199.620 ;
        RECT 107.170 199.260 107.310 204.720 ;
        RECT 108.030 203.195 108.290 203.340 ;
        RECT 108.020 202.825 108.300 203.195 ;
        RECT 110.330 202.340 110.590 202.660 ;
        RECT 107.510 201.125 109.390 201.495 ;
        RECT 107.110 198.940 107.370 199.260 ;
        RECT 107.170 194.410 107.310 198.940 ;
        RECT 108.950 197.755 109.210 197.900 ;
        RECT 108.940 197.385 109.220 197.755 ;
        RECT 110.390 197.560 110.530 202.340 ;
        RECT 110.790 199.115 111.050 199.260 ;
        RECT 110.780 198.745 111.060 199.115 ;
        RECT 111.310 198.240 111.450 205.740 ;
        RECT 111.250 197.920 111.510 198.240 ;
        RECT 110.330 197.240 110.590 197.560 ;
        RECT 111.710 197.240 111.970 197.560 ;
        RECT 107.510 195.685 109.390 196.055 ;
        RECT 109.400 194.665 109.680 195.035 ;
        RECT 109.470 194.500 109.610 194.665 ;
        RECT 108.030 194.410 108.290 194.500 ;
        RECT 107.170 194.270 108.290 194.410 ;
        RECT 108.030 194.180 108.290 194.270 ;
        RECT 109.410 194.180 109.670 194.500 ;
        RECT 107.110 193.675 107.370 193.820 ;
        RECT 107.100 193.305 107.380 193.675 ;
        RECT 108.950 193.500 109.210 193.820 ;
        RECT 107.170 187.360 107.310 193.305 ;
        RECT 109.010 192.800 109.150 193.500 ;
        RECT 108.950 192.480 109.210 192.800 ;
        RECT 109.870 190.780 110.130 191.100 ;
        RECT 107.510 190.245 109.390 190.615 ;
        RECT 109.930 189.480 110.070 190.780 ;
        RECT 109.470 189.340 110.070 189.480 ;
        RECT 110.390 189.400 110.530 197.240 ;
        RECT 111.250 196.900 111.510 197.220 ;
        RECT 111.310 195.520 111.450 196.900 ;
        RECT 111.250 195.200 111.510 195.520 ;
        RECT 111.770 194.500 111.910 197.240 ;
        RECT 111.710 194.180 111.970 194.500 ;
        RECT 110.790 189.760 111.050 190.080 ;
        RECT 109.470 188.915 109.610 189.340 ;
        RECT 110.330 189.080 110.590 189.400 ;
        RECT 108.030 188.400 108.290 188.720 ;
        RECT 109.400 188.545 109.680 188.915 ;
        RECT 109.870 188.740 110.130 189.060 ;
        RECT 108.090 187.555 108.230 188.400 ;
        RECT 107.110 187.040 107.370 187.360 ;
        RECT 108.020 187.185 108.300 187.555 ;
        RECT 109.470 186.680 109.610 188.545 ;
        RECT 107.570 186.360 107.830 186.680 ;
        RECT 109.410 186.360 109.670 186.680 ;
        RECT 107.630 186.195 107.770 186.360 ;
        RECT 106.650 185.680 106.910 186.000 ;
        RECT 107.560 185.825 107.840 186.195 ;
        RECT 107.110 185.340 107.370 185.660 ;
        RECT 106.190 183.300 106.450 183.620 ;
        RECT 105.730 180.580 105.990 180.900 ;
        RECT 106.250 176.480 106.390 183.300 ;
        RECT 107.170 181.920 107.310 185.340 ;
        RECT 107.510 184.805 109.390 185.175 ;
        RECT 109.930 184.640 110.070 188.740 ;
        RECT 110.330 188.060 110.590 188.380 ;
        RECT 109.870 184.320 110.130 184.640 ;
        RECT 107.110 181.600 107.370 181.920 ;
        RECT 106.650 181.260 106.910 181.580 ;
        RECT 106.190 176.160 106.450 176.480 ;
        RECT 105.330 175.740 106.390 175.880 ;
        RECT 105.730 174.460 105.990 174.780 ;
        RECT 105.790 173.760 105.930 174.460 ;
        RECT 105.730 173.440 105.990 173.760 ;
        RECT 104.350 171.740 104.610 172.060 ;
        RECT 104.810 171.740 105.070 172.060 ;
        RECT 104.410 171.040 104.550 171.740 ;
        RECT 104.350 170.720 104.610 171.040 ;
        RECT 105.720 170.185 106.000 170.555 ;
        RECT 104.810 163.580 105.070 163.900 ;
        RECT 105.790 163.810 105.930 170.185 ;
        RECT 106.250 164.580 106.390 175.740 ;
        RECT 106.710 170.555 106.850 181.260 ;
        RECT 107.170 176.480 107.310 181.600 ;
        RECT 107.510 179.365 109.390 179.735 ;
        RECT 110.390 178.600 110.530 188.060 ;
        RECT 110.850 186.680 110.990 189.760 ;
        RECT 110.790 186.360 111.050 186.680 ;
        RECT 110.790 182.620 111.050 182.940 ;
        RECT 109.470 178.520 110.530 178.600 ;
        RECT 109.410 178.460 110.530 178.520 ;
        RECT 109.410 178.200 109.670 178.460 ;
        RECT 109.870 177.520 110.130 177.840 ;
        RECT 107.110 176.160 107.370 176.480 ;
        RECT 107.110 174.460 107.370 174.780 ;
        RECT 106.640 170.185 106.920 170.555 ;
        RECT 106.650 169.360 106.910 169.680 ;
        RECT 106.710 168.320 106.850 169.360 ;
        RECT 106.650 168.000 106.910 168.320 ;
        RECT 107.170 167.720 107.310 174.460 ;
        RECT 107.510 173.925 109.390 174.295 ;
        RECT 108.490 171.740 108.750 172.060 ;
        RECT 108.550 170.360 108.690 171.740 ;
        RECT 108.490 170.040 108.750 170.360 ;
        RECT 109.410 170.040 109.670 170.360 ;
        RECT 109.470 169.680 109.610 170.040 ;
        RECT 109.410 169.360 109.670 169.680 ;
        RECT 107.510 168.485 109.390 168.855 ;
        RECT 106.710 167.580 107.310 167.720 ;
        RECT 106.190 164.260 106.450 164.580 ;
        RECT 105.790 163.670 106.390 163.810 ;
        RECT 104.870 161.860 105.010 163.580 ;
        RECT 105.730 162.560 105.990 162.880 ;
        RECT 104.810 161.540 105.070 161.860 ;
        RECT 104.870 159.480 105.010 161.540 ;
        RECT 104.810 159.160 105.070 159.480 ;
        RECT 104.350 158.820 104.610 159.140 ;
        RECT 104.410 157.440 104.550 158.820 ;
        RECT 104.350 157.120 104.610 157.440 ;
        RECT 104.810 148.620 105.070 148.940 ;
        RECT 104.870 146.560 105.010 148.620 ;
        RECT 104.810 146.240 105.070 146.560 ;
        RECT 103.890 145.900 104.150 146.220 ;
        RECT 102.050 145.220 102.310 145.540 ;
        RECT 102.970 145.220 103.230 145.540 ;
        RECT 104.350 145.220 104.610 145.540 ;
        RECT 101.590 144.540 101.850 144.860 ;
        RECT 101.650 142.480 101.790 144.540 ;
        RECT 101.590 142.160 101.850 142.480 ;
        RECT 102.110 139.760 102.250 145.220 ;
        RECT 103.430 144.540 103.690 144.860 ;
        RECT 103.490 143.500 103.630 144.540 ;
        RECT 103.430 143.180 103.690 143.500 ;
        RECT 102.050 139.440 102.310 139.760 ;
        RECT 101.590 139.100 101.850 139.420 ;
        RECT 101.650 136.700 101.790 139.100 ;
        RECT 103.430 137.740 103.690 138.060 ;
        RECT 101.590 136.380 101.850 136.700 ;
        RECT 103.490 132.960 103.630 137.740 ;
        RECT 104.410 133.980 104.550 145.220 ;
        RECT 105.790 144.860 105.930 162.560 ;
        RECT 106.250 149.280 106.390 163.670 ;
        RECT 106.190 148.960 106.450 149.280 ;
        RECT 106.710 146.220 106.850 167.580 ;
        RECT 107.510 163.045 109.390 163.415 ;
        RECT 109.930 162.880 110.070 177.520 ;
        RECT 110.330 175.140 110.590 175.460 ;
        RECT 110.390 173.760 110.530 175.140 ;
        RECT 110.330 173.440 110.590 173.760 ;
        RECT 110.850 172.400 110.990 182.620 ;
        RECT 111.250 180.580 111.510 180.900 ;
        RECT 111.310 178.520 111.450 180.580 ;
        RECT 111.250 178.200 111.510 178.520 ;
        RECT 111.310 173.080 111.450 178.200 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 111.250 172.760 111.510 173.080 ;
        RECT 110.790 172.080 111.050 172.400 ;
        RECT 110.330 171.740 110.590 172.060 ;
        RECT 110.390 165.600 110.530 171.740 ;
        RECT 110.790 170.720 111.050 171.040 ;
        RECT 110.330 165.280 110.590 165.600 ;
        RECT 110.330 164.260 110.590 164.580 ;
        RECT 109.870 162.560 110.130 162.880 ;
        RECT 109.870 161.540 110.130 161.860 ;
        RECT 107.110 160.860 107.370 161.180 ;
        RECT 109.410 160.860 109.670 161.180 ;
        RECT 107.170 159.480 107.310 160.860 ;
        RECT 107.110 159.160 107.370 159.480 ;
        RECT 109.470 158.880 109.610 160.860 ;
        RECT 109.930 160.160 110.070 161.540 ;
        RECT 109.870 159.840 110.130 160.160 ;
        RECT 109.470 158.740 110.070 158.880 ;
        RECT 107.110 158.140 107.370 158.460 ;
        RECT 107.170 156.080 107.310 158.140 ;
        RECT 107.510 157.605 109.390 157.975 ;
        RECT 107.110 155.760 107.370 156.080 ;
        RECT 107.510 152.165 109.390 152.535 ;
        RECT 109.930 150.980 110.070 158.740 ;
        RECT 110.390 156.160 110.530 164.260 ;
        RECT 110.850 161.600 110.990 170.720 ;
        RECT 111.310 167.640 111.450 172.760 ;
        RECT 111.710 172.420 111.970 172.740 ;
        RECT 111.770 171.040 111.910 172.420 ;
        RECT 111.710 170.720 111.970 171.040 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 111.710 169.020 111.970 169.340 ;
        RECT 111.770 167.835 111.910 169.020 ;
        RECT 111.250 167.320 111.510 167.640 ;
        RECT 111.700 167.465 111.980 167.835 ;
        RECT 111.310 164.920 111.450 167.320 ;
        RECT 111.710 166.640 111.970 166.960 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 111.250 164.600 111.510 164.920 ;
        RECT 110.850 161.460 111.450 161.600 ;
        RECT 110.790 160.860 111.050 161.180 ;
        RECT 110.850 156.760 110.990 160.860 ;
        RECT 111.310 159.820 111.450 161.460 ;
        RECT 111.250 159.500 111.510 159.820 ;
        RECT 111.250 158.820 111.510 159.140 ;
        RECT 110.790 156.440 111.050 156.760 ;
        RECT 110.390 156.020 110.990 156.160 ;
        RECT 110.330 155.420 110.590 155.740 ;
        RECT 110.390 153.700 110.530 155.420 ;
        RECT 110.330 153.380 110.590 153.700 ;
        RECT 109.870 150.660 110.130 150.980 ;
        RECT 108.490 149.980 108.750 150.300 ;
        RECT 108.550 148.600 108.690 149.980 ;
        RECT 108.490 148.280 108.750 148.600 ;
        RECT 110.390 148.260 110.530 153.380 ;
        RECT 110.850 152.000 110.990 156.020 ;
        RECT 110.790 151.680 111.050 152.000 ;
        RECT 111.310 151.320 111.450 158.820 ;
        RECT 111.770 151.660 111.910 166.640 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 111.710 151.340 111.970 151.660 ;
        RECT 111.250 151.000 111.510 151.320 ;
        RECT 110.790 150.320 111.050 150.640 ;
        RECT 110.850 148.600 110.990 150.320 ;
        RECT 110.790 148.280 111.050 148.600 ;
        RECT 109.410 148.000 109.670 148.260 ;
        RECT 109.410 147.940 110.070 148.000 ;
        RECT 110.330 147.940 110.590 148.260 ;
        RECT 109.470 147.860 110.070 147.940 ;
        RECT 107.510 146.725 109.390 147.095 ;
        RECT 106.650 145.900 106.910 146.220 ;
        RECT 108.950 145.900 109.210 146.220 ;
        RECT 109.010 145.540 109.150 145.900 ;
        RECT 108.950 145.220 109.210 145.540 ;
        RECT 105.730 144.540 105.990 144.860 ;
        RECT 109.410 144.540 109.670 144.860 ;
        RECT 109.470 143.160 109.610 144.540 ;
        RECT 109.410 142.840 109.670 143.160 ;
        RECT 107.510 141.285 109.390 141.655 ;
        RECT 109.410 139.780 109.670 140.100 ;
        RECT 105.730 139.440 105.990 139.760 ;
        RECT 105.790 135.680 105.930 139.440 ;
        RECT 109.470 138.400 109.610 139.780 ;
        RECT 109.410 138.080 109.670 138.400 ;
        RECT 107.570 137.400 107.830 137.720 ;
        RECT 106.650 137.060 106.910 137.380 ;
        RECT 105.730 135.360 105.990 135.680 ;
        RECT 104.810 134.680 105.070 135.000 ;
        RECT 104.350 133.890 104.610 133.980 ;
        RECT 103.950 133.750 104.610 133.890 ;
        RECT 103.430 132.640 103.690 132.960 ;
        RECT 102.970 132.190 103.230 132.280 ;
        RECT 103.950 132.190 104.090 133.750 ;
        RECT 104.350 133.660 104.610 133.750 ;
        RECT 104.350 132.640 104.610 132.960 ;
        RECT 102.970 132.050 104.090 132.190 ;
        RECT 102.970 131.960 103.230 132.050 ;
        RECT 103.030 130.240 103.170 131.960 ;
        RECT 102.970 129.920 103.230 130.240 ;
        RECT 104.410 128.880 104.550 132.640 ;
        RECT 104.870 132.620 105.010 134.680 ;
        RECT 106.710 134.660 106.850 137.060 ;
        RECT 107.630 136.950 107.770 137.400 ;
        RECT 107.170 136.810 107.770 136.950 ;
        RECT 106.650 134.340 106.910 134.660 ;
        RECT 107.170 132.960 107.310 136.810 ;
        RECT 107.510 135.845 109.390 136.215 ;
        RECT 107.110 132.640 107.370 132.960 ;
        RECT 104.810 132.300 105.070 132.620 ;
        RECT 109.930 132.280 110.070 147.860 ;
        RECT 110.390 142.820 110.530 147.940 ;
        RECT 110.850 146.220 110.990 148.280 ;
        RECT 110.790 145.900 111.050 146.220 ;
        RECT 111.700 145.705 111.980 146.075 ;
        RECT 111.770 145.540 111.910 145.705 ;
        RECT 110.780 145.025 111.060 145.395 ;
        RECT 111.710 145.220 111.970 145.540 ;
        RECT 110.850 144.860 110.990 145.025 ;
        RECT 110.790 144.540 111.050 144.860 ;
        RECT 110.330 142.500 110.590 142.820 ;
        RECT 110.390 140.440 110.530 142.500 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 110.330 140.120 110.590 140.440 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 110.390 137.380 110.530 140.120 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 110.330 137.060 110.590 137.380 ;
        RECT 111.250 134.340 111.510 134.660 ;
        RECT 110.790 133.660 111.050 133.980 ;
        RECT 107.110 131.960 107.370 132.280 ;
        RECT 109.870 131.960 110.130 132.280 ;
        RECT 107.170 131.680 107.310 131.960 ;
        RECT 104.870 131.540 107.310 131.680 ;
        RECT 104.350 128.560 104.610 128.880 ;
        RECT 104.350 127.200 104.610 127.520 ;
        RECT 101.130 124.480 101.390 124.800 ;
        RECT 100.210 123.120 100.470 123.440 ;
        RECT 100.670 123.120 100.930 123.440 ;
        RECT 98.370 121.420 98.630 121.740 ;
        RECT 95.610 120.740 95.870 121.060 ;
        RECT 97.910 120.740 98.170 121.060 ;
        RECT 95.670 108.580 95.810 120.740 ;
        RECT 100.270 108.580 100.410 123.120 ;
        RECT 104.410 120.800 104.550 127.200 ;
        RECT 104.870 121.400 105.010 131.540 ;
        RECT 110.330 131.280 110.590 131.600 ;
        RECT 106.190 130.940 106.450 131.260 ;
        RECT 106.650 130.940 106.910 131.260 ;
        RECT 106.250 130.240 106.390 130.940 ;
        RECT 106.190 129.920 106.450 130.240 ;
        RECT 106.710 128.880 106.850 130.940 ;
        RECT 107.510 130.405 109.390 130.775 ;
        RECT 106.650 128.560 106.910 128.880 ;
        RECT 110.390 128.540 110.530 131.280 ;
        RECT 110.850 130.240 110.990 133.660 ;
        RECT 110.790 129.920 111.050 130.240 ;
        RECT 110.330 128.220 110.590 128.540 ;
        RECT 109.870 126.860 110.130 127.180 ;
        RECT 107.510 124.965 109.390 125.335 ;
        RECT 109.930 124.800 110.070 126.860 ;
        RECT 109.870 124.480 110.130 124.800 ;
        RECT 110.390 123.780 110.530 128.220 ;
        RECT 110.330 123.460 110.590 123.780 ;
        RECT 110.330 122.780 110.590 123.100 ;
        RECT 109.870 121.760 110.130 122.080 ;
        RECT 104.810 121.080 105.070 121.400 ;
        RECT 104.410 120.660 105.010 120.800 ;
        RECT 104.870 108.580 105.010 120.660 ;
        RECT 107.510 119.525 109.390 119.895 ;
        RECT 109.930 118.760 110.070 121.760 ;
        RECT 110.390 121.740 110.530 122.780 ;
        RECT 110.330 121.420 110.590 121.740 ;
        RECT 111.310 120.915 111.450 134.340 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 114.010 128.560 114.270 128.880 ;
        RECT 111.710 123.120 111.970 123.440 ;
        RECT 111.770 121.400 111.910 123.120 ;
        RECT 111.710 121.080 111.970 121.400 ;
        RECT 111.240 120.545 111.520 120.915 ;
        RECT 109.470 118.620 110.070 118.760 ;
        RECT 109.470 108.580 109.610 118.620 ;
        RECT 114.070 108.580 114.210 128.560 ;
        RECT 62.090 108.420 63.150 108.560 ;
        RECT 63.400 106.580 63.680 108.580 ;
        RECT 68.000 106.580 68.280 108.580 ;
        RECT 72.600 106.580 72.880 108.580 ;
        RECT 77.200 106.580 77.480 108.580 ;
        RECT 81.800 106.580 82.080 108.580 ;
        RECT 86.400 106.580 86.680 108.580 ;
        RECT 91.000 106.580 91.280 108.580 ;
        RECT 95.600 106.580 95.880 108.580 ;
        RECT 100.200 106.580 100.480 108.580 ;
        RECT 104.800 106.580 105.080 108.580 ;
        RECT 109.400 106.580 109.680 108.580 ;
        RECT 114.000 106.580 114.280 108.580 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 40.375 206.560 40.705 206.575 ;
        RECT 91.435 206.560 91.765 206.575 ;
        RECT 40.375 206.260 91.765 206.560 ;
        RECT 40.375 206.245 40.705 206.260 ;
        RECT 91.435 206.245 91.765 206.260 ;
        RECT 43.135 205.880 43.465 205.895 ;
        RECT 101.095 205.880 101.425 205.895 ;
        RECT 43.135 205.580 101.425 205.880 ;
        RECT 43.135 205.565 43.465 205.580 ;
        RECT 101.095 205.565 101.425 205.580 ;
        RECT 44.975 205.200 45.305 205.215 ;
        RECT 105.235 205.200 105.565 205.215 ;
        RECT 44.975 204.900 105.565 205.200 ;
        RECT 44.975 204.885 45.305 204.900 ;
        RECT 105.235 204.885 105.565 204.900 ;
        RECT 32.460 203.865 34.440 204.195 ;
        RECT 62.460 203.865 64.440 204.195 ;
        RECT 92.460 203.865 94.440 204.195 ;
        RECT 56.015 203.840 56.345 203.855 ;
        RECT 61.535 203.840 61.865 203.855 ;
        RECT 56.015 203.540 61.865 203.840 ;
        RECT 56.015 203.525 56.345 203.540 ;
        RECT 61.535 203.525 61.865 203.540 ;
        RECT 39.915 203.160 40.245 203.175 ;
        RECT 107.995 203.160 108.325 203.175 ;
        RECT 39.915 202.860 108.325 203.160 ;
        RECT 39.915 202.845 40.245 202.860 ;
        RECT 107.995 202.845 108.325 202.860 ;
        RECT 42.215 202.480 42.545 202.495 ;
        RECT 98.795 202.480 99.125 202.495 ;
        RECT 42.215 202.180 99.125 202.480 ;
        RECT 42.215 202.165 42.545 202.180 ;
        RECT 98.795 202.165 99.125 202.180 ;
        RECT 47.460 201.145 49.440 201.475 ;
        RECT 77.460 201.145 79.440 201.475 ;
        RECT 107.460 201.145 109.440 201.475 ;
        RECT 76.255 201.120 76.585 201.135 ;
        RECT 56.720 200.820 76.585 201.120 ;
        RECT 50.495 200.440 50.825 200.455 ;
        RECT 56.720 200.440 57.020 200.820 ;
        RECT 76.255 200.805 76.585 200.820 ;
        RECT 50.495 200.140 57.020 200.440 ;
        RECT 57.855 200.440 58.185 200.455 ;
        RECT 84.995 200.440 85.325 200.455 ;
        RECT 57.855 200.140 85.325 200.440 ;
        RECT 50.495 200.125 50.825 200.140 ;
        RECT 57.855 200.125 58.185 200.140 ;
        RECT 84.995 200.125 85.325 200.140 ;
        RECT 41.960 199.760 42.340 199.770 ;
        RECT 42.675 199.760 43.005 199.775 ;
        RECT 41.960 199.460 43.005 199.760 ;
        RECT 41.960 199.450 42.340 199.460 ;
        RECT 42.675 199.445 43.005 199.460 ;
        RECT 49.575 199.760 49.905 199.775 ;
        RECT 83.155 199.760 83.485 199.775 ;
        RECT 49.575 199.460 83.485 199.760 ;
        RECT 49.575 199.445 49.905 199.460 ;
        RECT 83.155 199.445 83.485 199.460 ;
        RECT 84.075 199.760 84.405 199.775 ;
        RECT 86.835 199.760 87.165 199.775 ;
        RECT 95.575 199.760 95.905 199.775 ;
        RECT 84.075 199.460 95.905 199.760 ;
        RECT 84.075 199.445 84.405 199.460 ;
        RECT 86.835 199.445 87.165 199.460 ;
        RECT 95.575 199.445 95.905 199.460 ;
        RECT 38.075 199.080 38.405 199.095 ;
        RECT 61.535 199.080 61.865 199.095 ;
        RECT 110.755 199.090 111.085 199.095 ;
        RECT 110.755 199.080 111.340 199.090 ;
        RECT 38.075 198.780 61.865 199.080 ;
        RECT 110.530 198.780 111.340 199.080 ;
        RECT 38.075 198.765 38.405 198.780 ;
        RECT 61.535 198.765 61.865 198.780 ;
        RECT 110.755 198.770 111.340 198.780 ;
        RECT 110.755 198.765 111.085 198.770 ;
        RECT 32.460 198.425 34.440 198.755 ;
        RECT 62.460 198.425 64.440 198.755 ;
        RECT 92.460 198.425 94.440 198.755 ;
        RECT 75.795 198.400 76.125 198.415 ;
        RECT 90.975 198.400 91.305 198.415 ;
        RECT 75.795 198.100 91.305 198.400 ;
        RECT 75.795 198.085 76.125 198.100 ;
        RECT 90.975 198.085 91.305 198.100 ;
        RECT 38.995 197.720 39.325 197.735 ;
        RECT 108.915 197.720 109.245 197.735 ;
        RECT 38.995 197.420 109.245 197.720 ;
        RECT 38.995 197.405 39.325 197.420 ;
        RECT 108.915 197.405 109.245 197.420 ;
        RECT 43.800 197.040 44.180 197.050 ;
        RECT 44.515 197.040 44.845 197.055 ;
        RECT 43.800 196.740 44.845 197.040 ;
        RECT 43.800 196.730 44.180 196.740 ;
        RECT 44.515 196.725 44.845 196.740 ;
        RECT 64.295 197.040 64.625 197.055 ;
        RECT 73.495 197.040 73.825 197.055 ;
        RECT 64.295 196.740 73.825 197.040 ;
        RECT 64.295 196.725 64.625 196.740 ;
        RECT 73.495 196.725 73.825 196.740 ;
        RECT 76.255 197.040 76.585 197.055 ;
        RECT 104.315 197.040 104.645 197.055 ;
        RECT 76.255 196.740 104.645 197.040 ;
        RECT 76.255 196.725 76.585 196.740 ;
        RECT 104.315 196.725 104.645 196.740 ;
        RECT 33.935 196.360 34.265 196.375 ;
        RECT 42.880 196.360 43.260 196.370 ;
        RECT 33.935 196.060 43.260 196.360 ;
        RECT 33.935 196.045 34.265 196.060 ;
        RECT 42.880 196.050 43.260 196.060 ;
        RECT 79.935 196.360 80.265 196.375 ;
        RECT 101.555 196.360 101.885 196.375 ;
        RECT 79.935 196.060 101.885 196.360 ;
        RECT 79.935 196.045 80.265 196.060 ;
        RECT 101.555 196.045 101.885 196.060 ;
        RECT 47.460 195.705 49.440 196.035 ;
        RECT 77.460 195.705 79.440 196.035 ;
        RECT 107.460 195.705 109.440 196.035 ;
        RECT 62.915 195.680 63.245 195.695 ;
        RECT 50.510 195.380 63.245 195.680 ;
        RECT 33.015 195.000 33.345 195.015 ;
        RECT 39.455 195.010 39.785 195.015 ;
        RECT 35.520 195.000 35.900 195.010 ;
        RECT 33.015 194.700 35.900 195.000 ;
        RECT 33.015 194.685 33.345 194.700 ;
        RECT 35.520 194.690 35.900 194.700 ;
        RECT 39.200 195.000 39.785 195.010 ;
        RECT 41.960 195.000 42.340 195.010 ;
        RECT 44.055 195.000 44.385 195.015 ;
        RECT 50.510 195.000 50.810 195.380 ;
        RECT 62.915 195.365 63.245 195.380 ;
        RECT 91.640 195.680 92.020 195.690 ;
        RECT 94.195 195.680 94.525 195.695 ;
        RECT 106.155 195.680 106.485 195.695 ;
        RECT 91.640 195.380 106.485 195.680 ;
        RECT 91.640 195.370 92.020 195.380 ;
        RECT 94.195 195.365 94.525 195.380 ;
        RECT 106.155 195.365 106.485 195.380 ;
        RECT 39.200 194.700 40.010 195.000 ;
        RECT 41.960 194.700 44.385 195.000 ;
        RECT 39.200 194.690 39.785 194.700 ;
        RECT 41.960 194.690 42.340 194.700 ;
        RECT 39.455 194.685 39.785 194.690 ;
        RECT 44.055 194.685 44.385 194.700 ;
        RECT 49.360 194.700 50.810 195.000 ;
        RECT 51.415 195.000 51.745 195.015 ;
        RECT 65.675 195.000 66.005 195.015 ;
        RECT 68.435 195.000 68.765 195.015 ;
        RECT 51.415 194.700 68.765 195.000 ;
        RECT 40.120 194.320 40.500 194.330 ;
        RECT 40.835 194.320 41.165 194.335 ;
        RECT 49.360 194.320 49.660 194.700 ;
        RECT 51.415 194.685 51.745 194.700 ;
        RECT 65.675 194.685 66.005 194.700 ;
        RECT 68.435 194.685 68.765 194.700 ;
        RECT 89.135 195.000 89.465 195.015 ;
        RECT 109.375 195.000 109.705 195.015 ;
        RECT 89.135 194.700 109.705 195.000 ;
        RECT 89.135 194.685 89.465 194.700 ;
        RECT 109.375 194.685 109.705 194.700 ;
        RECT 40.120 194.020 49.660 194.320 ;
        RECT 50.035 194.320 50.365 194.335 ;
        RECT 101.095 194.320 101.425 194.335 ;
        RECT 50.035 194.020 101.425 194.320 ;
        RECT 40.120 194.010 40.500 194.020 ;
        RECT 40.835 194.005 41.165 194.020 ;
        RECT 50.035 194.005 50.365 194.020 ;
        RECT 101.095 194.005 101.425 194.020 ;
        RECT 38.075 193.640 38.405 193.655 ;
        RECT 50.495 193.640 50.825 193.655 ;
        RECT 38.075 193.340 50.825 193.640 ;
        RECT 38.075 193.325 38.405 193.340 ;
        RECT 50.495 193.325 50.825 193.340 ;
        RECT 95.575 193.640 95.905 193.655 ;
        RECT 107.075 193.640 107.405 193.655 ;
        RECT 95.575 193.340 107.405 193.640 ;
        RECT 95.575 193.325 95.905 193.340 ;
        RECT 107.075 193.325 107.405 193.340 ;
        RECT 32.460 192.985 34.440 193.315 ;
        RECT 62.460 192.985 64.440 193.315 ;
        RECT 92.460 192.985 94.440 193.315 ;
        RECT 53.255 192.280 53.585 192.295 ;
        RECT 103.855 192.280 104.185 192.295 ;
        RECT 53.255 191.980 104.185 192.280 ;
        RECT 53.255 191.965 53.585 191.980 ;
        RECT 103.855 191.965 104.185 191.980 ;
        RECT 45.435 191.600 45.765 191.615 ;
        RECT 96.955 191.600 97.285 191.615 ;
        RECT 45.435 191.300 97.285 191.600 ;
        RECT 45.435 191.285 45.765 191.300 ;
        RECT 96.955 191.285 97.285 191.300 ;
        RECT 47.460 190.265 49.440 190.595 ;
        RECT 77.460 190.265 79.440 190.595 ;
        RECT 107.460 190.265 109.440 190.595 ;
        RECT 36.695 189.560 37.025 189.575 ;
        RECT 44.515 189.560 44.845 189.575 ;
        RECT 36.695 189.260 44.845 189.560 ;
        RECT 36.695 189.245 37.025 189.260 ;
        RECT 44.515 189.245 44.845 189.260 ;
        RECT 71.195 189.560 71.525 189.575 ;
        RECT 92.355 189.560 92.685 189.575 ;
        RECT 71.195 189.260 92.685 189.560 ;
        RECT 71.195 189.245 71.525 189.260 ;
        RECT 92.355 189.245 92.685 189.260 ;
        RECT 37.155 188.880 37.485 188.895 ;
        RECT 39.455 188.880 39.785 188.895 ;
        RECT 37.155 188.580 39.785 188.880 ;
        RECT 37.155 188.565 37.485 188.580 ;
        RECT 39.455 188.565 39.785 188.580 ;
        RECT 89.135 188.880 89.465 188.895 ;
        RECT 109.375 188.880 109.705 188.895 ;
        RECT 89.135 188.580 109.705 188.880 ;
        RECT 89.135 188.565 89.465 188.580 ;
        RECT 109.375 188.565 109.705 188.580 ;
        RECT 32.460 187.545 34.440 187.875 ;
        RECT 62.460 187.545 64.440 187.875 ;
        RECT 92.460 187.545 94.440 187.875 ;
        RECT 39.915 187.520 40.245 187.535 ;
        RECT 59.695 187.520 60.025 187.535 ;
        RECT 39.915 187.220 60.025 187.520 ;
        RECT 39.915 187.205 40.245 187.220 ;
        RECT 59.695 187.205 60.025 187.220 ;
        RECT 88.675 187.520 89.005 187.535 ;
        RECT 106.360 187.520 106.740 187.530 ;
        RECT 107.995 187.520 108.325 187.535 ;
        RECT 88.675 187.205 89.220 187.520 ;
        RECT 106.360 187.220 108.325 187.520 ;
        RECT 106.360 187.210 106.740 187.220 ;
        RECT 107.995 187.205 108.325 187.220 ;
        RECT 54.635 186.840 54.965 186.855 ;
        RECT 74.875 186.840 75.205 186.855 ;
        RECT 54.635 186.540 75.205 186.840 ;
        RECT 88.920 186.840 89.220 187.205 ;
        RECT 101.095 186.840 101.425 186.855 ;
        RECT 88.920 186.540 101.425 186.840 ;
        RECT 54.635 186.525 54.965 186.540 ;
        RECT 74.875 186.525 75.205 186.540 ;
        RECT 101.095 186.525 101.425 186.540 ;
        RECT 61.995 186.160 62.325 186.175 ;
        RECT 73.035 186.160 73.365 186.175 ;
        RECT 90.515 186.160 90.845 186.175 ;
        RECT 91.640 186.160 92.020 186.170 ;
        RECT 93.735 186.160 94.065 186.175 ;
        RECT 61.995 185.860 94.065 186.160 ;
        RECT 61.995 185.845 62.325 185.860 ;
        RECT 73.035 185.845 73.365 185.860 ;
        RECT 90.515 185.845 90.845 185.860 ;
        RECT 91.640 185.850 92.020 185.860 ;
        RECT 93.735 185.845 94.065 185.860 ;
        RECT 104.315 186.160 104.645 186.175 ;
        RECT 107.535 186.160 107.865 186.175 ;
        RECT 104.315 185.860 107.865 186.160 ;
        RECT 104.315 185.845 104.645 185.860 ;
        RECT 107.535 185.845 107.865 185.860 ;
        RECT 47.460 184.825 49.440 185.155 ;
        RECT 77.460 184.825 79.440 185.155 ;
        RECT 107.460 184.825 109.440 185.155 ;
        RECT 73.240 184.800 73.620 184.810 ;
        RECT 74.875 184.800 75.205 184.815 ;
        RECT 73.240 184.500 75.205 184.800 ;
        RECT 73.240 184.490 73.620 184.500 ;
        RECT 74.875 184.485 75.205 184.500 ;
        RECT 44.055 184.120 44.385 184.135 ;
        RECT 50.035 184.120 50.365 184.135 ;
        RECT 44.055 183.820 50.365 184.120 ;
        RECT 44.055 183.805 44.385 183.820 ;
        RECT 50.035 183.805 50.365 183.820 ;
        RECT 70.735 184.120 71.065 184.135 ;
        RECT 88.675 184.120 89.005 184.135 ;
        RECT 96.495 184.120 96.825 184.135 ;
        RECT 98.795 184.120 99.125 184.135 ;
        RECT 70.735 183.820 99.125 184.120 ;
        RECT 70.735 183.805 71.065 183.820 ;
        RECT 88.675 183.805 89.005 183.820 ;
        RECT 96.495 183.805 96.825 183.820 ;
        RECT 98.795 183.805 99.125 183.820 ;
        RECT 100.175 183.805 100.505 184.135 ;
        RECT 56.475 183.440 56.805 183.455 ;
        RECT 66.135 183.440 66.465 183.455 ;
        RECT 56.475 183.140 66.465 183.440 ;
        RECT 56.475 183.125 56.805 183.140 ;
        RECT 66.135 183.125 66.465 183.140 ;
        RECT 97.415 183.440 97.745 183.455 ;
        RECT 99.000 183.440 99.380 183.450 ;
        RECT 100.190 183.440 100.490 183.805 ;
        RECT 97.415 183.140 100.490 183.440 ;
        RECT 97.415 183.125 97.745 183.140 ;
        RECT 99.000 183.130 99.380 183.140 ;
        RECT 36.695 182.760 37.025 182.775 ;
        RECT 38.995 182.760 39.325 182.775 ;
        RECT 36.695 182.460 39.325 182.760 ;
        RECT 36.695 182.445 37.025 182.460 ;
        RECT 38.995 182.445 39.325 182.460 ;
        RECT 40.375 182.760 40.705 182.775 ;
        RECT 51.415 182.760 51.745 182.775 ;
        RECT 40.375 182.460 51.745 182.760 ;
        RECT 40.375 182.445 40.705 182.460 ;
        RECT 51.415 182.445 51.745 182.460 ;
        RECT 32.460 182.105 34.440 182.435 ;
        RECT 62.460 182.105 64.440 182.435 ;
        RECT 92.460 182.105 94.440 182.435 ;
        RECT 70.735 182.080 71.065 182.095 ;
        RECT 89.135 182.080 89.465 182.095 ;
        RECT 70.735 181.780 89.465 182.080 ;
        RECT 70.735 181.765 71.065 181.780 ;
        RECT 89.135 181.765 89.465 181.780 ;
        RECT 28.875 181.400 29.205 181.415 ;
        RECT 59.235 181.400 59.565 181.415 ;
        RECT 28.875 181.100 59.565 181.400 ;
        RECT 28.875 181.085 29.205 181.100 ;
        RECT 59.235 181.085 59.565 181.100 ;
        RECT 63.375 181.400 63.705 181.415 ;
        RECT 67.975 181.400 68.305 181.415 ;
        RECT 63.375 181.100 68.305 181.400 ;
        RECT 63.375 181.085 63.705 181.100 ;
        RECT 67.975 181.085 68.305 181.100 ;
        RECT 78.095 181.400 78.425 181.415 ;
        RECT 82.695 181.400 83.025 181.415 ;
        RECT 78.095 181.100 83.025 181.400 ;
        RECT 78.095 181.085 78.425 181.100 ;
        RECT 82.695 181.085 83.025 181.100 ;
        RECT 33.015 180.720 33.345 180.735 ;
        RECT 35.520 180.720 35.900 180.730 ;
        RECT 67.975 180.720 68.305 180.735 ;
        RECT 33.015 180.420 68.305 180.720 ;
        RECT 33.015 180.405 33.345 180.420 ;
        RECT 35.520 180.410 35.900 180.420 ;
        RECT 67.975 180.405 68.305 180.420 ;
        RECT 71.655 180.040 71.985 180.055 ;
        RECT 72.575 180.040 72.905 180.055 ;
        RECT 71.655 179.740 72.905 180.040 ;
        RECT 71.655 179.725 71.985 179.740 ;
        RECT 72.575 179.725 72.905 179.740 ;
        RECT 47.460 179.385 49.440 179.715 ;
        RECT 77.460 179.385 79.440 179.715 ;
        RECT 107.460 179.385 109.440 179.715 ;
        RECT 39.915 178.680 40.245 178.695 ;
        RECT 38.320 178.380 40.245 178.680 ;
        RECT 37.615 178.000 37.945 178.015 ;
        RECT 38.320 178.000 38.620 178.380 ;
        RECT 39.915 178.365 40.245 178.380 ;
        RECT 46.815 178.680 47.145 178.695 ;
        RECT 74.875 178.680 75.205 178.695 ;
        RECT 46.815 178.380 75.205 178.680 ;
        RECT 46.815 178.365 47.145 178.380 ;
        RECT 74.875 178.365 75.205 178.380 ;
        RECT 39.915 178.010 40.245 178.015 ;
        RECT 39.915 178.000 40.500 178.010 ;
        RECT 37.615 177.700 38.620 178.000 ;
        RECT 39.690 177.700 40.500 178.000 ;
        RECT 37.615 177.685 37.945 177.700 ;
        RECT 32.460 176.665 34.440 176.995 ;
        RECT 38.320 176.640 38.620 177.700 ;
        RECT 39.915 177.690 40.500 177.700 ;
        RECT 41.960 178.000 42.340 178.010 ;
        RECT 68.435 178.000 68.765 178.015 ;
        RECT 41.960 177.700 68.765 178.000 ;
        RECT 41.960 177.690 42.340 177.700 ;
        RECT 39.915 177.685 40.245 177.690 ;
        RECT 68.435 177.685 68.765 177.700 ;
        RECT 41.295 177.320 41.625 177.335 ;
        RECT 61.075 177.320 61.405 177.335 ;
        RECT 41.295 177.020 61.405 177.320 ;
        RECT 41.295 177.005 41.625 177.020 ;
        RECT 61.075 177.005 61.405 177.020 ;
        RECT 62.460 176.665 64.440 176.995 ;
        RECT 92.460 176.665 94.440 176.995 ;
        RECT 60.615 176.640 60.945 176.655 ;
        RECT 38.320 176.340 60.945 176.640 ;
        RECT 60.615 176.325 60.945 176.340 ;
        RECT 40.835 175.960 41.165 175.975 ;
        RECT 41.960 175.960 42.340 175.970 ;
        RECT 40.835 175.660 42.340 175.960 ;
        RECT 40.835 175.645 41.165 175.660 ;
        RECT 41.960 175.650 42.340 175.660 ;
        RECT 74.875 175.960 75.205 175.975 ;
        RECT 96.495 175.960 96.825 175.975 ;
        RECT 74.875 175.660 96.825 175.960 ;
        RECT 74.875 175.645 75.205 175.660 ;
        RECT 96.495 175.645 96.825 175.660 ;
        RECT 64.960 175.280 65.340 175.290 ;
        RECT 85.915 175.280 86.245 175.295 ;
        RECT 64.960 174.980 86.245 175.280 ;
        RECT 64.960 174.970 65.340 174.980 ;
        RECT 85.915 174.965 86.245 174.980 ;
        RECT 101.555 175.280 101.885 175.295 ;
        RECT 116.970 175.280 118.970 175.430 ;
        RECT 101.555 174.980 118.970 175.280 ;
        RECT 101.555 174.965 101.885 174.980 ;
        RECT 116.970 174.830 118.970 174.980 ;
        RECT 43.595 174.610 43.925 174.615 ;
        RECT 43.595 174.600 44.180 174.610 ;
        RECT 43.595 174.300 44.380 174.600 ;
        RECT 43.595 174.290 44.180 174.300 ;
        RECT 43.595 174.285 43.925 174.290 ;
        RECT 47.460 173.945 49.440 174.275 ;
        RECT 77.460 173.945 79.440 174.275 ;
        RECT 107.460 173.945 109.440 174.275 ;
        RECT 42.880 173.240 43.260 173.250 ;
        RECT 47.275 173.240 47.605 173.255 ;
        RECT 42.880 172.940 47.605 173.240 ;
        RECT 42.880 172.930 43.260 172.940 ;
        RECT 47.275 172.925 47.605 172.940 ;
        RECT 34.395 172.560 34.725 172.575 ;
        RECT 36.235 172.560 36.565 172.575 ;
        RECT 34.395 172.260 36.565 172.560 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 34.395 172.245 34.725 172.260 ;
        RECT 36.235 172.245 36.565 172.260 ;
        RECT 32.460 171.225 34.440 171.555 ;
        RECT 62.460 171.225 64.440 171.555 ;
        RECT 92.460 171.225 94.440 171.555 ;
        RECT 46.815 170.520 47.145 170.535 ;
        RECT 49.575 170.520 49.905 170.535 ;
        RECT 64.960 170.520 65.340 170.530 ;
        RECT 46.815 170.220 65.340 170.520 ;
        RECT 46.815 170.205 47.145 170.220 ;
        RECT 49.575 170.205 49.905 170.220 ;
        RECT 64.960 170.210 65.340 170.220 ;
        RECT 99.715 170.520 100.045 170.535 ;
        RECT 103.395 170.520 103.725 170.535 ;
        RECT 99.715 170.220 103.725 170.520 ;
        RECT 99.715 170.205 100.045 170.220 ;
        RECT 103.395 170.205 103.725 170.220 ;
        RECT 105.695 170.520 106.025 170.535 ;
        RECT 106.615 170.520 106.945 170.535 ;
        RECT 105.695 170.220 106.945 170.520 ;
        RECT 105.695 170.205 106.025 170.220 ;
        RECT 106.615 170.205 106.945 170.220 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 70.735 169.840 71.065 169.855 ;
        RECT 72.575 169.840 72.905 169.855 ;
        RECT 70.735 169.540 72.905 169.840 ;
        RECT 70.735 169.525 71.065 169.540 ;
        RECT 72.575 169.525 72.905 169.540 ;
        RECT 47.460 168.505 49.440 168.835 ;
        RECT 77.460 168.505 79.440 168.835 ;
        RECT 107.460 168.505 109.440 168.835 ;
        RECT 59.695 168.480 60.025 168.495 ;
        RECT 63.835 168.480 64.165 168.495 ;
        RECT 70.275 168.480 70.605 168.495 ;
        RECT 59.695 168.180 70.605 168.480 ;
        RECT 59.695 168.165 60.025 168.180 ;
        RECT 63.835 168.165 64.165 168.180 ;
        RECT 70.275 168.165 70.605 168.180 ;
        RECT 59.235 167.800 59.565 167.815 ;
        RECT 67.515 167.800 67.845 167.815 ;
        RECT 59.235 167.500 67.845 167.800 ;
        RECT 59.235 167.485 59.565 167.500 ;
        RECT 67.515 167.485 67.845 167.500 ;
        RECT 88.215 167.800 88.545 167.815 ;
        RECT 111.675 167.800 112.005 167.815 ;
        RECT 88.215 167.500 112.005 167.800 ;
        RECT 88.215 167.485 88.545 167.500 ;
        RECT 111.675 167.485 112.005 167.500 ;
        RECT 59.235 167.120 59.565 167.135 ;
        RECT 62.915 167.120 63.245 167.135 ;
        RECT 67.055 167.120 67.385 167.135 ;
        RECT 59.235 166.820 67.385 167.120 ;
        RECT 59.235 166.805 59.565 166.820 ;
        RECT 62.915 166.805 63.245 166.820 ;
        RECT 67.055 166.805 67.385 166.820 ;
        RECT 80.855 167.120 81.185 167.135 ;
        RECT 89.135 167.120 89.465 167.135 ;
        RECT 80.855 166.820 89.465 167.120 ;
        RECT 80.855 166.805 81.185 166.820 ;
        RECT 89.135 166.805 89.465 166.820 ;
        RECT 32.460 165.785 34.440 166.115 ;
        RECT 62.460 165.785 64.440 166.115 ;
        RECT 92.460 165.785 94.440 166.115 ;
        RECT 70.735 165.760 71.065 165.775 ;
        RECT 71.400 165.760 71.780 165.770 ;
        RECT 70.735 165.460 71.780 165.760 ;
        RECT 70.735 165.445 71.065 165.460 ;
        RECT 71.400 165.450 71.780 165.460 ;
        RECT 73.495 165.760 73.825 165.775 ;
        RECT 76.255 165.760 76.585 165.775 ;
        RECT 73.495 165.460 76.585 165.760 ;
        RECT 73.495 165.445 73.825 165.460 ;
        RECT 76.255 165.445 76.585 165.460 ;
        RECT 77.635 165.760 77.965 165.775 ;
        RECT 83.615 165.760 83.945 165.775 ;
        RECT 77.635 165.460 83.945 165.760 ;
        RECT 77.635 165.445 77.965 165.460 ;
        RECT 83.615 165.445 83.945 165.460 ;
        RECT 67.975 165.080 68.305 165.095 ;
        RECT 91.435 165.080 91.765 165.095 ;
        RECT 94.195 165.080 94.525 165.095 ;
        RECT 67.975 164.780 94.525 165.080 ;
        RECT 67.975 164.765 68.305 164.780 ;
        RECT 91.435 164.765 91.765 164.780 ;
        RECT 94.195 164.765 94.525 164.780 ;
        RECT 50.035 164.400 50.365 164.415 ;
        RECT 51.160 164.400 51.540 164.410 ;
        RECT 50.035 164.100 51.540 164.400 ;
        RECT 50.035 164.085 50.365 164.100 ;
        RECT 51.160 164.090 51.540 164.100 ;
        RECT 71.195 164.400 71.525 164.415 ;
        RECT 76.715 164.400 77.045 164.415 ;
        RECT 71.195 164.100 77.045 164.400 ;
        RECT 71.195 164.085 71.525 164.100 ;
        RECT 76.715 164.085 77.045 164.100 ;
        RECT 39.455 163.720 39.785 163.735 ;
        RECT 40.375 163.720 40.705 163.735 ;
        RECT 39.455 163.420 40.705 163.720 ;
        RECT 39.455 163.405 39.785 163.420 ;
        RECT 40.375 163.405 40.705 163.420 ;
        RECT 87.295 163.720 87.625 163.735 ;
        RECT 90.720 163.720 91.100 163.730 ;
        RECT 87.295 163.420 91.100 163.720 ;
        RECT 87.295 163.405 87.625 163.420 ;
        RECT 90.720 163.410 91.100 163.420 ;
        RECT 47.460 163.065 49.440 163.395 ;
        RECT 77.460 163.065 79.440 163.395 ;
        RECT 107.460 163.065 109.440 163.395 ;
        RECT 64.295 163.040 64.625 163.055 ;
        RECT 64.960 163.040 65.340 163.050 ;
        RECT 70.480 163.040 70.860 163.050 ;
        RECT 64.295 162.740 70.860 163.040 ;
        RECT 64.295 162.725 64.625 162.740 ;
        RECT 64.960 162.730 65.340 162.740 ;
        RECT 70.480 162.730 70.860 162.740 ;
        RECT 49.575 162.360 49.905 162.375 ;
        RECT 50.240 162.360 50.620 162.370 ;
        RECT 49.575 162.060 50.620 162.360 ;
        RECT 49.575 162.045 49.905 162.060 ;
        RECT 50.240 162.050 50.620 162.060 ;
        RECT 70.735 162.360 71.065 162.375 ;
        RECT 71.400 162.360 71.780 162.370 ;
        RECT 70.735 162.060 71.780 162.360 ;
        RECT 70.735 162.045 71.065 162.060 ;
        RECT 71.400 162.050 71.780 162.060 ;
        RECT 93.275 162.360 93.605 162.375 ;
        RECT 102.475 162.360 102.805 162.375 ;
        RECT 93.275 162.060 102.805 162.360 ;
        RECT 93.275 162.045 93.605 162.060 ;
        RECT 102.475 162.045 102.805 162.060 ;
        RECT 44.515 161.680 44.845 161.695 ;
        RECT 49.575 161.680 49.905 161.695 ;
        RECT 61.075 161.680 61.405 161.695 ;
        RECT 44.515 161.380 61.405 161.680 ;
        RECT 44.515 161.365 44.845 161.380 ;
        RECT 49.575 161.365 49.905 161.380 ;
        RECT 61.075 161.365 61.405 161.380 ;
        RECT 83.155 161.680 83.485 161.695 ;
        RECT 99.000 161.680 99.380 161.690 ;
        RECT 83.155 161.380 99.380 161.680 ;
        RECT 83.155 161.365 83.485 161.380 ;
        RECT 99.000 161.370 99.380 161.380 ;
        RECT 46.355 161.010 46.685 161.015 ;
        RECT 46.355 161.000 46.940 161.010 ;
        RECT 46.130 160.700 46.940 161.000 ;
        RECT 46.355 160.690 46.940 160.700 ;
        RECT 96.035 161.000 96.365 161.015 ;
        RECT 103.395 161.000 103.725 161.015 ;
        RECT 96.035 160.700 103.725 161.000 ;
        RECT 46.355 160.685 46.685 160.690 ;
        RECT 96.035 160.685 96.365 160.700 ;
        RECT 103.395 160.685 103.725 160.700 ;
        RECT 32.460 160.345 34.440 160.675 ;
        RECT 62.460 160.345 64.440 160.675 ;
        RECT 92.460 160.345 94.440 160.675 ;
        RECT 38.535 160.320 38.865 160.335 ;
        RECT 43.135 160.320 43.465 160.335 ;
        RECT 38.535 160.020 43.465 160.320 ;
        RECT 38.535 160.005 38.865 160.020 ;
        RECT 43.135 160.005 43.465 160.020 ;
        RECT 70.735 160.320 71.065 160.335 ;
        RECT 76.000 160.320 76.380 160.330 ;
        RECT 70.735 160.020 76.380 160.320 ;
        RECT 70.735 160.005 71.065 160.020 ;
        RECT 76.000 160.010 76.380 160.020 ;
        RECT 38.075 159.640 38.405 159.655 ;
        RECT 39.200 159.640 39.580 159.650 ;
        RECT 38.075 159.340 39.580 159.640 ;
        RECT 38.075 159.325 38.405 159.340 ;
        RECT 39.200 159.330 39.580 159.340 ;
        RECT 42.215 159.640 42.545 159.655 ;
        RECT 44.515 159.640 44.845 159.655 ;
        RECT 42.215 159.340 44.845 159.640 ;
        RECT 42.215 159.325 42.545 159.340 ;
        RECT 44.515 159.325 44.845 159.340 ;
        RECT 46.815 159.640 47.145 159.655 ;
        RECT 50.035 159.640 50.365 159.655 ;
        RECT 59.235 159.640 59.565 159.655 ;
        RECT 46.815 159.340 59.565 159.640 ;
        RECT 46.815 159.325 47.145 159.340 ;
        RECT 50.035 159.325 50.365 159.340 ;
        RECT 59.235 159.325 59.565 159.340 ;
        RECT 94.195 159.640 94.525 159.655 ;
        RECT 99.255 159.640 99.585 159.655 ;
        RECT 94.195 159.340 99.585 159.640 ;
        RECT 94.195 159.325 94.525 159.340 ;
        RECT 99.255 159.325 99.585 159.340 ;
        RECT 30.715 158.960 31.045 158.975 ;
        RECT 32.555 158.960 32.885 158.975 ;
        RECT 65.215 158.960 65.545 158.975 ;
        RECT 30.715 158.645 31.260 158.960 ;
        RECT 32.555 158.660 65.545 158.960 ;
        RECT 32.555 158.645 32.885 158.660 ;
        RECT 65.215 158.645 65.545 158.660 ;
        RECT 88.675 158.960 89.005 158.975 ;
        RECT 94.655 158.960 94.985 158.975 ;
        RECT 88.675 158.660 94.985 158.960 ;
        RECT 88.675 158.645 89.005 158.660 ;
        RECT 94.655 158.645 94.985 158.660 ;
        RECT 30.960 156.255 31.260 158.645 ;
        RECT 33.935 158.280 34.265 158.295 ;
        RECT 44.515 158.280 44.845 158.295 ;
        RECT 33.935 157.980 44.845 158.280 ;
        RECT 33.935 157.965 34.265 157.980 ;
        RECT 44.515 157.965 44.845 157.980 ;
        RECT 47.460 157.625 49.440 157.955 ;
        RECT 77.460 157.625 79.440 157.955 ;
        RECT 107.460 157.625 109.440 157.955 ;
        RECT 46.355 156.920 46.685 156.935 ;
        RECT 47.735 156.920 48.065 156.935 ;
        RECT 52.335 156.920 52.665 156.935 ;
        RECT 46.355 156.620 52.665 156.920 ;
        RECT 46.355 156.605 46.685 156.620 ;
        RECT 47.735 156.605 48.065 156.620 ;
        RECT 52.335 156.605 52.665 156.620 ;
        RECT 75.795 156.920 76.125 156.935 ;
        RECT 95.115 156.920 95.445 156.935 ;
        RECT 75.795 156.620 95.445 156.920 ;
        RECT 75.795 156.605 76.125 156.620 ;
        RECT 95.115 156.605 95.445 156.620 ;
        RECT 97.415 156.920 97.745 156.935 ;
        RECT 100.175 156.920 100.505 156.935 ;
        RECT 97.415 156.620 100.505 156.920 ;
        RECT 97.415 156.605 97.745 156.620 ;
        RECT 100.175 156.605 100.505 156.620 ;
        RECT 30.960 155.940 31.505 156.255 ;
        RECT 31.175 155.925 31.505 155.940 ;
        RECT 43.595 156.240 43.925 156.255 ;
        RECT 57.855 156.240 58.185 156.255 ;
        RECT 43.595 155.940 58.185 156.240 ;
        RECT 43.595 155.925 43.925 155.940 ;
        RECT 57.855 155.925 58.185 155.940 ;
        RECT 74.415 156.240 74.745 156.255 ;
        RECT 93.735 156.240 94.065 156.255 ;
        RECT 99.255 156.240 99.585 156.255 ;
        RECT 74.415 155.940 99.585 156.240 ;
        RECT 74.415 155.925 74.745 155.940 ;
        RECT 93.735 155.925 94.065 155.940 ;
        RECT 99.255 155.925 99.585 155.940 ;
        RECT 39.915 155.560 40.245 155.575 ;
        RECT 57.395 155.560 57.725 155.575 ;
        RECT 60.155 155.560 60.485 155.575 ;
        RECT 39.915 155.260 60.485 155.560 ;
        RECT 39.915 155.245 40.245 155.260 ;
        RECT 57.395 155.245 57.725 155.260 ;
        RECT 60.155 155.245 60.485 155.260 ;
        RECT 32.460 154.905 34.440 155.235 ;
        RECT 62.460 154.905 64.440 155.235 ;
        RECT 92.460 154.905 94.440 155.235 ;
        RECT 46.815 154.890 47.145 154.895 ;
        RECT 46.560 154.880 47.145 154.890 ;
        RECT 46.360 154.580 47.145 154.880 ;
        RECT 46.560 154.570 47.145 154.580 ;
        RECT 46.815 154.565 47.145 154.570 ;
        RECT 30.255 154.200 30.585 154.215 ;
        RECT 50.035 154.200 50.365 154.215 ;
        RECT 30.255 153.900 50.365 154.200 ;
        RECT 30.255 153.885 30.585 153.900 ;
        RECT 50.035 153.885 50.365 153.900 ;
        RECT 50.955 154.210 51.285 154.215 ;
        RECT 50.955 154.200 51.540 154.210 ;
        RECT 50.955 153.900 51.740 154.200 ;
        RECT 50.955 153.890 51.540 153.900 ;
        RECT 50.955 153.885 51.285 153.890 ;
        RECT 49.575 153.520 49.905 153.535 ;
        RECT 50.240 153.520 50.620 153.530 ;
        RECT 49.575 153.220 50.620 153.520 ;
        RECT 49.575 153.205 49.905 153.220 ;
        RECT 50.240 153.210 50.620 153.220 ;
        RECT 47.460 152.185 49.440 152.515 ;
        RECT 77.460 152.185 79.440 152.515 ;
        RECT 107.460 152.185 109.440 152.515 ;
        RECT 46.355 151.480 46.685 151.495 ;
        RECT 53.715 151.480 54.045 151.495 ;
        RECT 46.355 151.180 54.045 151.480 ;
        RECT 46.355 151.165 46.685 151.180 ;
        RECT 53.715 151.165 54.045 151.180 ;
        RECT 99.000 151.480 99.380 151.490 ;
        RECT 100.175 151.480 100.505 151.495 ;
        RECT 99.000 151.180 100.505 151.480 ;
        RECT 99.000 151.170 99.380 151.180 ;
        RECT 100.175 151.165 100.505 151.180 ;
        RECT 32.460 149.465 34.440 149.795 ;
        RECT 62.460 149.465 64.440 149.795 ;
        RECT 92.460 149.465 94.440 149.795 ;
        RECT 57.855 149.440 58.185 149.455 ;
        RECT 61.535 149.440 61.865 149.455 ;
        RECT 57.855 149.140 61.865 149.440 ;
        RECT 57.855 149.125 58.185 149.140 ;
        RECT 61.535 149.125 61.865 149.140 ;
        RECT 53.715 148.760 54.045 148.775 ;
        RECT 57.395 148.760 57.725 148.775 ;
        RECT 61.535 148.760 61.865 148.775 ;
        RECT 53.715 148.460 61.865 148.760 ;
        RECT 53.715 148.445 54.045 148.460 ;
        RECT 57.395 148.445 57.725 148.460 ;
        RECT 61.535 148.445 61.865 148.460 ;
        RECT 76.000 148.080 76.380 148.090 ;
        RECT 116.970 148.080 118.970 148.230 ;
        RECT 76.000 147.780 118.970 148.080 ;
        RECT 76.000 147.770 76.380 147.780 ;
        RECT 116.970 147.630 118.970 147.780 ;
        RECT 47.460 146.745 49.440 147.075 ;
        RECT 77.460 146.745 79.440 147.075 ;
        RECT 107.460 146.745 109.440 147.075 ;
        RECT 73.240 146.040 73.620 146.050 ;
        RECT 75.335 146.040 75.665 146.055 ;
        RECT 73.240 145.740 75.665 146.040 ;
        RECT 73.240 145.730 73.620 145.740 ;
        RECT 75.335 145.725 75.665 145.740 ;
        RECT 110.960 146.040 111.340 146.050 ;
        RECT 111.675 146.040 112.005 146.055 ;
        RECT 110.960 145.740 112.005 146.040 ;
        RECT 110.960 145.730 111.340 145.740 ;
        RECT 111.675 145.725 112.005 145.740 ;
        RECT 106.360 145.360 106.740 145.370 ;
        RECT 110.755 145.360 111.085 145.375 ;
        RECT 106.360 145.060 111.085 145.360 ;
        RECT 106.360 145.050 106.740 145.060 ;
        RECT 110.755 145.045 111.085 145.060 ;
        RECT 32.460 144.025 34.440 144.355 ;
        RECT 62.460 144.025 64.440 144.355 ;
        RECT 92.460 144.025 94.440 144.355 ;
        RECT 47.460 141.305 49.440 141.635 ;
        RECT 77.460 141.305 79.440 141.635 ;
        RECT 107.460 141.305 109.440 141.635 ;
        RECT 68.435 140.600 68.765 140.615 ;
        RECT 70.480 140.600 70.860 140.610 ;
        RECT 93.275 140.600 93.605 140.615 ;
        RECT 56.720 140.300 93.605 140.600 ;
        RECT 49.115 139.920 49.445 139.935 ;
        RECT 56.720 139.920 57.020 140.300 ;
        RECT 68.435 140.285 68.765 140.300 ;
        RECT 70.480 140.290 70.860 140.300 ;
        RECT 93.275 140.285 93.605 140.300 ;
        RECT 49.115 139.620 57.020 139.920 ;
        RECT 49.115 139.605 49.445 139.620 ;
        RECT 32.460 138.585 34.440 138.915 ;
        RECT 62.460 138.585 64.440 138.915 ;
        RECT 92.460 138.585 94.440 138.915 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 47.460 135.865 49.440 136.195 ;
        RECT 77.460 135.865 79.440 136.195 ;
        RECT 107.460 135.865 109.440 136.195 ;
        RECT 32.095 135.160 32.425 135.175 ;
        RECT 41.755 135.160 42.085 135.175 ;
        RECT 32.095 134.860 42.085 135.160 ;
        RECT 32.095 134.845 32.425 134.860 ;
        RECT 41.755 134.845 42.085 134.860 ;
        RECT 32.460 133.145 34.440 133.475 ;
        RECT 62.460 133.145 64.440 133.475 ;
        RECT 92.460 133.145 94.440 133.475 ;
        RECT 38.535 132.440 38.865 132.455 ;
        RECT 53.715 132.440 54.045 132.455 ;
        RECT 68.435 132.440 68.765 132.455 ;
        RECT 79.935 132.440 80.265 132.455 ;
        RECT 38.535 132.140 80.265 132.440 ;
        RECT 38.535 132.125 38.865 132.140 ;
        RECT 53.715 132.125 54.045 132.140 ;
        RECT 68.435 132.125 68.765 132.140 ;
        RECT 79.935 132.125 80.265 132.140 ;
        RECT 90.720 132.440 91.100 132.450 ;
        RECT 98.335 132.440 98.665 132.455 ;
        RECT 90.720 132.140 98.665 132.440 ;
        RECT 90.720 132.130 91.100 132.140 ;
        RECT 98.335 132.125 98.665 132.140 ;
        RECT 47.460 130.425 49.440 130.755 ;
        RECT 77.460 130.425 79.440 130.755 ;
        RECT 107.460 130.425 109.440 130.755 ;
        RECT 32.460 127.705 34.440 128.035 ;
        RECT 62.460 127.705 64.440 128.035 ;
        RECT 92.460 127.705 94.440 128.035 ;
        RECT 47.460 124.985 49.440 125.315 ;
        RECT 77.460 124.985 79.440 125.315 ;
        RECT 107.460 124.985 109.440 125.315 ;
        RECT 32.460 122.265 34.440 122.595 ;
        RECT 62.460 122.265 64.440 122.595 ;
        RECT 92.460 122.265 94.440 122.595 ;
        RECT 111.215 120.880 111.545 120.895 ;
        RECT 116.970 120.880 118.970 121.030 ;
        RECT 111.215 120.580 118.970 120.880 ;
        RECT 111.215 120.565 111.545 120.580 ;
        RECT 116.970 120.430 118.970 120.580 ;
        RECT 47.460 119.545 49.440 119.875 ;
        RECT 77.460 119.545 79.440 119.875 ;
        RECT 107.460 119.545 109.440 119.875 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 32.450 119.470 34.450 204.270 ;
        RECT 41.985 199.445 42.315 199.775 ;
        RECT 42.000 195.015 42.300 199.445 ;
        RECT 43.825 196.725 44.155 197.055 ;
        RECT 42.905 196.045 43.235 196.375 ;
        RECT 35.545 194.685 35.875 195.015 ;
        RECT 39.225 194.685 39.555 195.015 ;
        RECT 41.985 194.685 42.315 195.015 ;
        RECT 35.560 180.735 35.860 194.685 ;
        RECT 35.545 180.405 35.875 180.735 ;
        RECT 39.240 159.655 39.540 194.685 ;
        RECT 40.145 194.005 40.475 194.335 ;
        RECT 40.160 178.015 40.460 194.005 ;
        RECT 42.000 178.015 42.300 194.685 ;
        RECT 40.145 177.685 40.475 178.015 ;
        RECT 41.985 177.685 42.315 178.015 ;
        RECT 42.000 175.975 42.300 177.685 ;
        RECT 41.985 175.645 42.315 175.975 ;
        RECT 42.920 173.255 43.220 196.045 ;
        RECT 43.840 174.615 44.140 196.725 ;
        RECT 43.825 174.285 44.155 174.615 ;
        RECT 42.905 172.925 43.235 173.255 ;
        RECT 46.585 160.685 46.915 161.015 ;
        RECT 39.225 159.325 39.555 159.655 ;
        RECT 46.600 154.895 46.900 160.685 ;
        RECT 46.585 154.565 46.915 154.895 ;
        RECT 47.450 119.470 49.450 204.270 ;
        RECT 51.185 164.085 51.515 164.415 ;
        RECT 50.265 162.045 50.595 162.375 ;
        RECT 50.280 153.535 50.580 162.045 ;
        RECT 51.200 154.215 51.500 164.085 ;
        RECT 51.185 153.885 51.515 154.215 ;
        RECT 50.265 153.205 50.595 153.535 ;
        RECT 62.450 119.470 64.450 204.270 ;
        RECT 73.265 184.485 73.595 184.815 ;
        RECT 64.985 174.965 65.315 175.295 ;
        RECT 65.000 170.535 65.300 174.965 ;
        RECT 64.985 170.205 65.315 170.535 ;
        RECT 65.000 163.055 65.300 170.205 ;
        RECT 71.425 165.445 71.755 165.775 ;
        RECT 64.985 162.725 65.315 163.055 ;
        RECT 70.505 162.725 70.835 163.055 ;
        RECT 70.520 140.615 70.820 162.725 ;
        RECT 71.440 162.375 71.740 165.445 ;
        RECT 71.425 162.045 71.755 162.375 ;
        RECT 73.280 146.055 73.580 184.485 ;
        RECT 76.025 160.005 76.355 160.335 ;
        RECT 76.040 148.095 76.340 160.005 ;
        RECT 76.025 147.765 76.355 148.095 ;
        RECT 73.265 145.725 73.595 146.055 ;
        RECT 70.505 140.285 70.835 140.615 ;
        RECT 77.450 119.470 79.450 204.270 ;
        RECT 91.665 195.365 91.995 195.695 ;
        RECT 91.680 186.175 91.980 195.365 ;
        RECT 91.665 185.845 91.995 186.175 ;
        RECT 90.745 163.405 91.075 163.735 ;
        RECT 90.760 132.455 91.060 163.405 ;
        RECT 90.745 132.125 91.075 132.455 ;
        RECT 92.450 119.470 94.450 204.270 ;
        RECT 106.385 187.205 106.715 187.535 ;
        RECT 99.025 183.125 99.355 183.455 ;
        RECT 99.040 161.695 99.340 183.125 ;
        RECT 99.025 161.365 99.355 161.695 ;
        RECT 99.040 151.495 99.340 161.365 ;
        RECT 99.025 151.165 99.355 151.495 ;
        RECT 106.400 145.375 106.700 187.205 ;
        RECT 106.385 145.045 106.715 145.375 ;
        RECT 107.450 119.470 109.450 204.270 ;
        RECT 110.985 198.765 111.315 199.095 ;
        RECT 111.000 146.055 111.300 198.765 ;
        RECT 110.985 145.725 111.315 146.055 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

