VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 1199.802979 ;
    ANTENNADIFFAREA 1170.027222 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 9.435 215.805 9.605 215.995 ;
        RECT 10.870 215.855 10.990 215.965 ;
        RECT 12.655 215.805 12.825 215.995 ;
        RECT 14.495 215.805 14.665 215.995 ;
        RECT 20.015 215.805 20.185 215.995 ;
        RECT 25.535 215.805 25.705 215.995 ;
        RECT 27.375 215.805 27.545 215.995 ;
        RECT 32.895 215.805 33.065 215.995 ;
        RECT 38.415 215.805 38.585 215.995 ;
        RECT 40.255 215.805 40.425 215.995 ;
        RECT 45.775 215.805 45.945 215.995 ;
        RECT 51.295 215.805 51.465 215.995 ;
        RECT 53.135 215.805 53.305 215.995 ;
        RECT 58.655 215.805 58.825 215.995 ;
        RECT 64.175 215.805 64.345 215.995 ;
        RECT 66.015 215.805 66.185 215.995 ;
        RECT 71.535 215.805 71.705 215.995 ;
        RECT 77.055 215.805 77.225 215.995 ;
        RECT 78.895 215.805 79.065 215.995 ;
        RECT 84.415 215.805 84.585 215.995 ;
        RECT 89.935 215.805 90.105 215.995 ;
        RECT 91.775 215.805 91.945 215.995 ;
        RECT 97.295 215.805 97.465 215.995 ;
        RECT 102.815 215.805 102.985 215.995 ;
        RECT 104.655 215.805 104.825 215.995 ;
        RECT 110.175 215.805 110.345 215.995 ;
        RECT 115.695 215.805 115.865 215.995 ;
        RECT 116.670 215.855 116.790 215.965 ;
        RECT 122.135 215.805 122.305 215.995 ;
        RECT 127.655 215.805 127.825 215.995 ;
        RECT 129.035 215.805 129.205 215.995 ;
        RECT 9.295 214.995 10.665 215.805 ;
        RECT 11.135 214.995 12.965 215.805 ;
        RECT 12.985 214.935 13.415 215.720 ;
        RECT 13.435 214.995 14.805 215.805 ;
        RECT 14.815 214.995 20.325 215.805 ;
        RECT 20.335 214.995 25.845 215.805 ;
        RECT 25.865 214.935 26.295 215.720 ;
        RECT 26.315 214.995 27.685 215.805 ;
        RECT 27.695 214.995 33.205 215.805 ;
        RECT 33.215 214.995 38.725 215.805 ;
        RECT 38.745 214.935 39.175 215.720 ;
        RECT 39.195 214.995 40.565 215.805 ;
        RECT 40.575 214.995 46.085 215.805 ;
        RECT 46.095 214.995 51.605 215.805 ;
        RECT 51.625 214.935 52.055 215.720 ;
        RECT 52.075 214.995 53.445 215.805 ;
        RECT 53.455 214.995 58.965 215.805 ;
        RECT 58.975 214.995 64.485 215.805 ;
        RECT 64.505 214.935 64.935 215.720 ;
        RECT 64.955 214.995 66.325 215.805 ;
        RECT 66.335 214.995 71.845 215.805 ;
        RECT 71.855 214.995 77.365 215.805 ;
        RECT 77.385 214.935 77.815 215.720 ;
        RECT 77.835 214.995 79.205 215.805 ;
        RECT 79.215 214.995 84.725 215.805 ;
        RECT 84.735 214.995 90.245 215.805 ;
        RECT 90.265 214.935 90.695 215.720 ;
        RECT 90.715 214.995 92.085 215.805 ;
        RECT 92.095 214.995 97.605 215.805 ;
        RECT 97.615 214.995 103.125 215.805 ;
        RECT 103.145 214.935 103.575 215.720 ;
        RECT 103.595 214.995 104.965 215.805 ;
        RECT 104.975 214.995 110.485 215.805 ;
        RECT 110.495 214.995 116.005 215.805 ;
        RECT 116.025 214.935 116.455 215.720 ;
        RECT 116.935 214.995 122.445 215.805 ;
        RECT 122.455 214.995 127.965 215.805 ;
        RECT 127.975 214.995 129.345 215.805 ;
      LAYER nwell ;
        RECT 9.100 211.775 129.540 214.605 ;
      LAYER pwell ;
        RECT 9.295 210.575 10.665 211.385 ;
        RECT 11.135 210.575 14.805 211.385 ;
        RECT 14.815 210.575 20.325 211.385 ;
        RECT 20.335 210.575 25.845 211.385 ;
        RECT 25.865 210.660 26.295 211.445 ;
        RECT 26.775 210.575 29.525 211.385 ;
        RECT 29.535 210.575 35.045 211.385 ;
        RECT 35.055 210.575 40.565 211.385 ;
        RECT 40.575 210.575 46.085 211.385 ;
        RECT 46.095 210.575 51.605 211.385 ;
        RECT 51.625 210.660 52.055 211.445 ;
        RECT 52.535 210.575 55.285 211.385 ;
        RECT 55.295 210.575 60.805 211.385 ;
        RECT 60.815 210.575 66.325 211.385 ;
        RECT 66.335 210.575 71.845 211.385 ;
        RECT 71.855 210.575 77.365 211.385 ;
        RECT 77.385 210.660 77.815 211.445 ;
        RECT 78.295 210.575 81.045 211.385 ;
        RECT 81.055 210.575 86.565 211.385 ;
        RECT 86.575 210.575 92.085 211.385 ;
        RECT 92.095 210.575 97.605 211.385 ;
        RECT 97.615 210.575 103.125 211.385 ;
        RECT 103.145 210.660 103.575 211.445 ;
        RECT 104.055 210.575 105.885 211.385 ;
        RECT 105.895 210.575 111.405 211.385 ;
        RECT 111.415 210.575 116.925 211.385 ;
        RECT 116.935 210.575 122.445 211.385 ;
        RECT 122.455 210.575 127.965 211.385 ;
        RECT 127.975 210.575 129.345 211.385 ;
        RECT 9.435 210.365 9.605 210.575 ;
        RECT 10.870 210.415 10.990 210.525 ;
        RECT 12.655 210.365 12.825 210.555 ;
        RECT 13.630 210.415 13.750 210.525 ;
        RECT 14.495 210.385 14.665 210.575 ;
        RECT 16.335 210.365 16.505 210.555 ;
        RECT 20.015 210.385 20.185 210.575 ;
        RECT 21.855 210.365 22.025 210.555 ;
        RECT 25.535 210.385 25.705 210.575 ;
        RECT 26.510 210.415 26.630 210.525 ;
        RECT 27.375 210.365 27.545 210.555 ;
        RECT 29.215 210.385 29.385 210.575 ;
        RECT 32.895 210.365 33.065 210.555 ;
        RECT 34.735 210.385 34.905 210.575 ;
        RECT 38.415 210.365 38.585 210.555 ;
        RECT 39.390 210.415 39.510 210.525 ;
        RECT 40.255 210.385 40.425 210.575 ;
        RECT 42.095 210.365 42.265 210.555 ;
        RECT 45.775 210.385 45.945 210.575 ;
        RECT 47.615 210.365 47.785 210.555 ;
        RECT 51.295 210.385 51.465 210.575 ;
        RECT 52.270 210.415 52.390 210.525 ;
        RECT 53.135 210.365 53.305 210.555 ;
        RECT 54.975 210.385 55.145 210.575 ;
        RECT 58.655 210.365 58.825 210.555 ;
        RECT 60.495 210.385 60.665 210.575 ;
        RECT 64.175 210.365 64.345 210.555 ;
        RECT 65.150 210.415 65.270 210.525 ;
        RECT 66.015 210.385 66.185 210.575 ;
        RECT 67.855 210.365 68.025 210.555 ;
        RECT 71.535 210.385 71.705 210.575 ;
        RECT 73.375 210.365 73.545 210.555 ;
        RECT 77.055 210.385 77.225 210.575 ;
        RECT 78.030 210.415 78.150 210.525 ;
        RECT 78.895 210.365 79.065 210.555 ;
        RECT 80.735 210.385 80.905 210.575 ;
        RECT 84.415 210.365 84.585 210.555 ;
        RECT 86.255 210.385 86.425 210.575 ;
        RECT 89.935 210.365 90.105 210.555 ;
        RECT 90.910 210.415 91.030 210.525 ;
        RECT 91.775 210.385 91.945 210.575 ;
        RECT 93.615 210.365 93.785 210.555 ;
        RECT 97.295 210.385 97.465 210.575 ;
        RECT 99.135 210.365 99.305 210.555 ;
        RECT 102.815 210.385 102.985 210.575 ;
        RECT 103.790 210.415 103.910 210.525 ;
        RECT 104.655 210.365 104.825 210.555 ;
        RECT 105.575 210.385 105.745 210.575 ;
        RECT 110.175 210.365 110.345 210.555 ;
        RECT 111.095 210.385 111.265 210.575 ;
        RECT 115.695 210.365 115.865 210.555 ;
        RECT 116.615 210.525 116.785 210.575 ;
        RECT 116.615 210.415 116.790 210.525 ;
        RECT 116.615 210.385 116.785 210.415 ;
        RECT 122.135 210.365 122.305 210.575 ;
        RECT 127.655 210.365 127.825 210.575 ;
        RECT 129.035 210.365 129.205 210.575 ;
        RECT 9.295 209.555 10.665 210.365 ;
        RECT 11.135 209.555 12.965 210.365 ;
        RECT 12.985 209.495 13.415 210.280 ;
        RECT 13.895 209.555 16.645 210.365 ;
        RECT 16.655 209.555 22.165 210.365 ;
        RECT 22.175 209.555 27.685 210.365 ;
        RECT 27.695 209.555 33.205 210.365 ;
        RECT 33.215 209.555 38.725 210.365 ;
        RECT 38.745 209.495 39.175 210.280 ;
        RECT 39.655 209.555 42.405 210.365 ;
        RECT 42.415 209.555 47.925 210.365 ;
        RECT 47.935 209.555 53.445 210.365 ;
        RECT 53.455 209.555 58.965 210.365 ;
        RECT 58.975 209.555 64.485 210.365 ;
        RECT 64.505 209.495 64.935 210.280 ;
        RECT 65.415 209.555 68.165 210.365 ;
        RECT 68.175 209.555 73.685 210.365 ;
        RECT 73.695 209.555 79.205 210.365 ;
        RECT 79.215 209.555 84.725 210.365 ;
        RECT 84.735 209.555 90.245 210.365 ;
        RECT 90.265 209.495 90.695 210.280 ;
        RECT 91.175 209.555 93.925 210.365 ;
        RECT 93.935 209.555 99.445 210.365 ;
        RECT 99.455 209.555 104.965 210.365 ;
        RECT 104.975 209.555 110.485 210.365 ;
        RECT 110.495 209.555 116.005 210.365 ;
        RECT 116.025 209.495 116.455 210.280 ;
        RECT 116.935 209.555 122.445 210.365 ;
        RECT 122.455 209.555 127.965 210.365 ;
        RECT 127.975 209.555 129.345 210.365 ;
      LAYER nwell ;
        RECT 9.100 206.335 129.540 209.165 ;
      LAYER pwell ;
        RECT 9.295 205.135 10.665 205.945 ;
        RECT 11.135 205.135 14.805 205.945 ;
        RECT 14.815 205.135 20.325 205.945 ;
        RECT 20.335 205.135 25.845 205.945 ;
        RECT 25.865 205.220 26.295 206.005 ;
        RECT 26.775 205.135 29.525 205.945 ;
        RECT 29.535 205.135 35.045 205.945 ;
        RECT 35.055 205.135 40.565 205.945 ;
        RECT 40.575 205.135 46.085 205.945 ;
        RECT 46.095 205.135 51.605 205.945 ;
        RECT 51.625 205.220 52.055 206.005 ;
        RECT 52.535 205.135 55.285 205.945 ;
        RECT 55.295 205.135 60.805 205.945 ;
        RECT 60.815 205.135 66.325 205.945 ;
        RECT 66.335 205.135 71.845 205.945 ;
        RECT 71.855 205.135 77.365 205.945 ;
        RECT 77.385 205.220 77.815 206.005 ;
        RECT 78.295 205.135 81.045 205.945 ;
        RECT 81.055 205.135 86.565 205.945 ;
        RECT 86.575 205.135 92.085 205.945 ;
        RECT 92.095 205.135 97.605 205.945 ;
        RECT 97.615 205.135 103.125 205.945 ;
        RECT 103.145 205.220 103.575 206.005 ;
        RECT 104.055 205.135 105.885 205.945 ;
        RECT 105.895 205.135 111.405 205.945 ;
        RECT 111.415 205.135 116.925 205.945 ;
        RECT 116.935 205.135 122.445 205.945 ;
        RECT 122.455 205.135 127.965 205.945 ;
        RECT 127.975 205.135 129.345 205.945 ;
        RECT 9.435 204.925 9.605 205.135 ;
        RECT 10.870 204.975 10.990 205.085 ;
        RECT 12.655 204.925 12.825 205.115 ;
        RECT 13.630 204.975 13.750 205.085 ;
        RECT 14.495 204.945 14.665 205.135 ;
        RECT 16.335 204.925 16.505 205.115 ;
        RECT 20.015 204.945 20.185 205.135 ;
        RECT 21.855 204.925 22.025 205.115 ;
        RECT 25.535 204.945 25.705 205.135 ;
        RECT 26.510 204.975 26.630 205.085 ;
        RECT 27.375 204.925 27.545 205.115 ;
        RECT 29.215 204.945 29.385 205.135 ;
        RECT 32.895 204.925 33.065 205.115 ;
        RECT 34.735 204.945 34.905 205.135 ;
        RECT 38.415 204.925 38.585 205.115 ;
        RECT 39.390 204.975 39.510 205.085 ;
        RECT 40.255 204.945 40.425 205.135 ;
        RECT 42.095 204.925 42.265 205.115 ;
        RECT 45.775 204.945 45.945 205.135 ;
        RECT 47.615 204.925 47.785 205.115 ;
        RECT 51.295 204.945 51.465 205.135 ;
        RECT 52.270 204.975 52.390 205.085 ;
        RECT 53.135 204.925 53.305 205.115 ;
        RECT 54.975 204.945 55.145 205.135 ;
        RECT 58.655 204.925 58.825 205.115 ;
        RECT 60.495 204.945 60.665 205.135 ;
        RECT 64.175 204.925 64.345 205.115 ;
        RECT 65.150 204.975 65.270 205.085 ;
        RECT 66.015 204.945 66.185 205.135 ;
        RECT 67.855 204.925 68.025 205.115 ;
        RECT 71.535 204.945 71.705 205.135 ;
        RECT 73.375 204.925 73.545 205.115 ;
        RECT 77.055 204.945 77.225 205.135 ;
        RECT 78.030 204.975 78.150 205.085 ;
        RECT 78.895 204.925 79.065 205.115 ;
        RECT 80.735 204.945 80.905 205.135 ;
        RECT 84.415 204.925 84.585 205.115 ;
        RECT 86.255 204.945 86.425 205.135 ;
        RECT 89.935 204.925 90.105 205.115 ;
        RECT 90.910 204.975 91.030 205.085 ;
        RECT 91.775 204.945 91.945 205.135 ;
        RECT 93.615 204.925 93.785 205.115 ;
        RECT 97.295 204.945 97.465 205.135 ;
        RECT 99.135 204.925 99.305 205.115 ;
        RECT 102.815 204.945 102.985 205.135 ;
        RECT 103.790 204.975 103.910 205.085 ;
        RECT 104.655 204.925 104.825 205.115 ;
        RECT 105.575 204.945 105.745 205.135 ;
        RECT 110.175 204.925 110.345 205.115 ;
        RECT 111.095 204.945 111.265 205.135 ;
        RECT 115.695 204.925 115.865 205.115 ;
        RECT 116.615 205.085 116.785 205.135 ;
        RECT 116.615 204.975 116.790 205.085 ;
        RECT 116.615 204.945 116.785 204.975 ;
        RECT 122.135 204.925 122.305 205.135 ;
        RECT 127.655 204.925 127.825 205.135 ;
        RECT 129.035 204.925 129.205 205.135 ;
        RECT 9.295 204.115 10.665 204.925 ;
        RECT 11.135 204.115 12.965 204.925 ;
        RECT 12.985 204.055 13.415 204.840 ;
        RECT 13.895 204.115 16.645 204.925 ;
        RECT 16.655 204.115 22.165 204.925 ;
        RECT 22.175 204.115 27.685 204.925 ;
        RECT 27.695 204.115 33.205 204.925 ;
        RECT 33.215 204.115 38.725 204.925 ;
        RECT 38.745 204.055 39.175 204.840 ;
        RECT 39.655 204.115 42.405 204.925 ;
        RECT 42.415 204.115 47.925 204.925 ;
        RECT 47.935 204.115 53.445 204.925 ;
        RECT 53.455 204.115 58.965 204.925 ;
        RECT 58.975 204.115 64.485 204.925 ;
        RECT 64.505 204.055 64.935 204.840 ;
        RECT 65.415 204.115 68.165 204.925 ;
        RECT 68.175 204.115 73.685 204.925 ;
        RECT 73.695 204.115 79.205 204.925 ;
        RECT 79.215 204.115 84.725 204.925 ;
        RECT 84.735 204.115 90.245 204.925 ;
        RECT 90.265 204.055 90.695 204.840 ;
        RECT 91.175 204.115 93.925 204.925 ;
        RECT 93.935 204.115 99.445 204.925 ;
        RECT 99.455 204.115 104.965 204.925 ;
        RECT 104.975 204.115 110.485 204.925 ;
        RECT 110.495 204.115 116.005 204.925 ;
        RECT 116.025 204.055 116.455 204.840 ;
        RECT 116.935 204.115 122.445 204.925 ;
        RECT 122.455 204.115 127.965 204.925 ;
        RECT 127.975 204.115 129.345 204.925 ;
      LAYER nwell ;
        RECT 9.100 200.895 129.540 203.725 ;
      LAYER pwell ;
        RECT 9.295 199.695 10.665 200.505 ;
        RECT 11.135 199.695 14.805 200.505 ;
        RECT 14.815 199.695 20.325 200.505 ;
        RECT 20.335 199.695 25.845 200.505 ;
        RECT 25.865 199.780 26.295 200.565 ;
        RECT 26.775 199.695 29.525 200.505 ;
        RECT 29.535 199.695 35.045 200.505 ;
        RECT 35.055 199.695 40.565 200.505 ;
        RECT 40.575 199.695 46.085 200.505 ;
        RECT 46.095 199.695 51.605 200.505 ;
        RECT 51.625 199.780 52.055 200.565 ;
        RECT 52.535 199.695 55.285 200.505 ;
        RECT 55.295 199.695 60.805 200.505 ;
        RECT 60.815 199.695 66.325 200.505 ;
        RECT 66.335 199.695 71.845 200.505 ;
        RECT 71.855 199.695 77.365 200.505 ;
        RECT 77.385 199.780 77.815 200.565 ;
        RECT 78.295 199.695 81.045 200.505 ;
        RECT 81.055 199.695 86.565 200.505 ;
        RECT 86.575 199.695 92.085 200.505 ;
        RECT 92.095 199.695 97.605 200.505 ;
        RECT 97.615 199.695 103.125 200.505 ;
        RECT 103.145 199.780 103.575 200.565 ;
        RECT 104.055 199.695 105.885 200.505 ;
        RECT 105.895 199.695 111.405 200.505 ;
        RECT 111.415 199.695 116.925 200.505 ;
        RECT 116.935 199.695 122.445 200.505 ;
        RECT 122.455 199.695 127.965 200.505 ;
        RECT 127.975 199.695 129.345 200.505 ;
        RECT 9.435 199.485 9.605 199.695 ;
        RECT 10.870 199.535 10.990 199.645 ;
        RECT 12.655 199.485 12.825 199.675 ;
        RECT 13.630 199.535 13.750 199.645 ;
        RECT 14.495 199.505 14.665 199.695 ;
        RECT 16.335 199.485 16.505 199.675 ;
        RECT 20.015 199.505 20.185 199.695 ;
        RECT 21.855 199.485 22.025 199.675 ;
        RECT 25.535 199.505 25.705 199.695 ;
        RECT 26.510 199.535 26.630 199.645 ;
        RECT 27.375 199.485 27.545 199.675 ;
        RECT 29.215 199.505 29.385 199.695 ;
        RECT 32.895 199.485 33.065 199.675 ;
        RECT 34.735 199.505 34.905 199.695 ;
        RECT 38.415 199.485 38.585 199.675 ;
        RECT 39.795 199.530 39.955 199.640 ;
        RECT 40.255 199.505 40.425 199.695 ;
        RECT 43.475 199.485 43.645 199.675 ;
        RECT 45.775 199.505 45.945 199.695 ;
        RECT 48.995 199.485 49.165 199.675 ;
        RECT 51.295 199.505 51.465 199.695 ;
        RECT 52.270 199.535 52.390 199.645 ;
        RECT 54.515 199.485 54.685 199.675 ;
        RECT 54.975 199.485 55.145 199.695 ;
        RECT 60.495 199.505 60.665 199.695 ;
        RECT 66.015 199.485 66.185 199.695 ;
        RECT 66.530 199.535 66.650 199.645 ;
        RECT 69.695 199.485 69.865 199.675 ;
        RECT 71.535 199.505 71.705 199.695 ;
        RECT 73.375 199.485 73.545 199.675 ;
        RECT 77.055 199.505 77.225 199.695 ;
        RECT 78.030 199.535 78.150 199.645 ;
        RECT 78.895 199.485 79.065 199.675 ;
        RECT 80.735 199.505 80.905 199.695 ;
        RECT 84.415 199.485 84.585 199.675 ;
        RECT 86.255 199.505 86.425 199.695 ;
        RECT 89.935 199.485 90.105 199.675 ;
        RECT 91.775 199.505 91.945 199.695 ;
        RECT 92.235 199.485 92.405 199.675 ;
        RECT 97.295 199.505 97.465 199.695 ;
        RECT 97.755 199.485 97.925 199.675 ;
        RECT 99.135 199.485 99.305 199.675 ;
        RECT 100.055 199.530 100.215 199.640 ;
        RECT 100.515 199.485 100.685 199.675 ;
        RECT 102.815 199.485 102.985 199.695 ;
        RECT 103.790 199.535 103.910 199.645 ;
        RECT 105.575 199.505 105.745 199.695 ;
        RECT 108.335 199.485 108.505 199.675 ;
        RECT 111.095 199.505 111.265 199.695 ;
        RECT 113.855 199.485 114.025 199.675 ;
        RECT 115.235 199.485 115.405 199.675 ;
        RECT 116.615 199.645 116.785 199.695 ;
        RECT 115.750 199.535 115.870 199.645 ;
        RECT 116.615 199.535 116.790 199.645 ;
        RECT 116.615 199.505 116.785 199.535 ;
        RECT 122.135 199.485 122.305 199.695 ;
        RECT 127.655 199.485 127.825 199.695 ;
        RECT 129.035 199.485 129.205 199.695 ;
        RECT 9.295 198.675 10.665 199.485 ;
        RECT 11.135 198.675 12.965 199.485 ;
        RECT 12.985 198.615 13.415 199.400 ;
        RECT 13.895 198.675 16.645 199.485 ;
        RECT 16.655 198.675 22.165 199.485 ;
        RECT 22.175 198.675 27.685 199.485 ;
        RECT 27.695 198.675 33.205 199.485 ;
        RECT 33.215 198.675 38.725 199.485 ;
        RECT 38.745 198.615 39.175 199.400 ;
        RECT 40.115 198.675 43.785 199.485 ;
        RECT 43.795 198.675 49.305 199.485 ;
        RECT 49.315 198.675 54.825 199.485 ;
        RECT 54.835 198.805 64.445 199.485 ;
        RECT 59.345 198.585 60.275 198.805 ;
        RECT 63.105 198.575 64.445 198.805 ;
        RECT 64.505 198.615 64.935 199.400 ;
        RECT 64.965 198.575 66.315 199.485 ;
        RECT 66.795 198.575 69.905 199.485 ;
        RECT 70.015 198.675 73.685 199.485 ;
        RECT 73.695 198.675 79.205 199.485 ;
        RECT 79.215 198.675 84.725 199.485 ;
        RECT 84.735 198.675 90.245 199.485 ;
        RECT 90.265 198.615 90.695 199.400 ;
        RECT 90.715 198.675 92.545 199.485 ;
        RECT 92.555 198.675 98.065 199.485 ;
        RECT 98.085 198.575 99.435 199.485 ;
        RECT 100.375 198.705 101.745 199.485 ;
        RECT 101.755 198.675 103.125 199.485 ;
        RECT 103.135 198.675 108.645 199.485 ;
        RECT 108.655 198.675 114.165 199.485 ;
        RECT 114.185 198.575 115.535 199.485 ;
        RECT 116.025 198.615 116.455 199.400 ;
        RECT 116.935 198.675 122.445 199.485 ;
        RECT 122.455 198.675 127.965 199.485 ;
        RECT 127.975 198.675 129.345 199.485 ;
      LAYER nwell ;
        RECT 9.100 195.455 129.540 198.285 ;
      LAYER pwell ;
        RECT 9.295 194.255 10.665 195.065 ;
        RECT 11.135 194.255 14.805 195.065 ;
        RECT 14.815 194.255 20.325 195.065 ;
        RECT 20.335 194.255 25.845 195.065 ;
        RECT 25.865 194.340 26.295 195.125 ;
        RECT 26.775 194.255 32.285 195.065 ;
        RECT 32.295 194.255 37.805 195.065 ;
        RECT 37.815 194.255 43.325 195.065 ;
        RECT 43.335 194.255 44.705 195.035 ;
        RECT 45.645 194.255 46.995 195.165 ;
        RECT 47.475 194.255 50.225 195.065 ;
        RECT 50.245 194.255 51.595 195.165 ;
        RECT 51.625 194.340 52.055 195.125 ;
        RECT 52.075 194.255 53.905 195.065 ;
        RECT 53.915 194.255 55.285 195.035 ;
        RECT 55.295 194.255 56.665 195.065 ;
        RECT 61.185 194.935 62.115 195.155 ;
        RECT 64.835 194.935 67.045 195.165 ;
        RECT 56.675 194.255 67.045 194.935 ;
        RECT 67.255 194.255 68.625 195.035 ;
        RECT 69.095 194.255 72.765 195.065 ;
        RECT 72.785 194.255 74.135 195.165 ;
        RECT 74.255 194.255 77.365 195.165 ;
        RECT 77.385 194.340 77.815 195.125 ;
        RECT 78.295 194.255 83.805 195.065 ;
        RECT 84.185 195.055 85.105 195.165 ;
        RECT 84.185 194.935 86.520 195.055 ;
        RECT 91.185 194.935 92.105 195.155 ;
        RECT 93.935 194.935 94.855 195.165 ;
        RECT 97.685 194.935 98.615 195.155 ;
        RECT 84.185 194.255 93.465 194.935 ;
        RECT 93.935 194.255 103.125 194.935 ;
        RECT 103.145 194.340 103.575 195.125 ;
        RECT 104.515 194.255 110.025 195.065 ;
        RECT 110.045 194.255 111.395 195.165 ;
        RECT 111.415 194.935 112.335 195.165 ;
        RECT 115.165 194.935 116.095 195.155 ;
        RECT 111.415 194.255 120.605 194.935 ;
        RECT 120.615 194.255 122.445 195.065 ;
        RECT 122.455 194.255 127.965 195.065 ;
        RECT 127.975 194.255 129.345 195.065 ;
        RECT 9.435 194.045 9.605 194.255 ;
        RECT 10.870 194.095 10.990 194.205 ;
        RECT 12.655 194.045 12.825 194.235 ;
        RECT 14.035 194.090 14.195 194.200 ;
        RECT 14.495 194.065 14.665 194.255 ;
        RECT 17.715 194.045 17.885 194.235 ;
        RECT 20.015 194.065 20.185 194.255 ;
        RECT 23.235 194.045 23.405 194.235 ;
        RECT 25.535 194.065 25.705 194.255 ;
        RECT 26.510 194.095 26.630 194.205 ;
        RECT 28.755 194.045 28.925 194.235 ;
        RECT 31.975 194.065 32.145 194.255 ;
        RECT 34.275 194.045 34.445 194.235 ;
        RECT 37.495 194.065 37.665 194.255 ;
        RECT 38.140 194.045 38.310 194.235 ;
        RECT 39.335 194.045 39.505 194.235 ;
        RECT 43.015 194.065 43.185 194.255 ;
        RECT 44.395 194.065 44.565 194.255 ;
        RECT 45.315 194.100 45.475 194.210 ;
        RECT 46.695 194.065 46.865 194.255 ;
        RECT 47.210 194.095 47.330 194.205 ;
        RECT 48.590 194.095 48.710 194.205 ;
        RECT 49.915 194.065 50.085 194.255 ;
        RECT 50.375 194.065 50.545 194.255 ;
        RECT 53.595 194.065 53.765 194.255 ;
        RECT 54.055 194.065 54.225 194.255 ;
        RECT 56.355 194.065 56.525 194.255 ;
        RECT 56.815 194.065 56.985 194.255 ;
        RECT 57.735 194.045 57.905 194.235 ;
        RECT 58.250 194.095 58.370 194.205 ;
        RECT 61.875 194.045 62.045 194.235 ;
        RECT 63.255 194.045 63.425 194.235 ;
        RECT 64.175 194.090 64.335 194.200 ;
        RECT 65.150 194.095 65.270 194.205 ;
        RECT 67.395 194.045 67.565 194.235 ;
        RECT 68.315 194.065 68.485 194.255 ;
        RECT 68.830 194.095 68.950 194.205 ;
        RECT 69.690 194.045 69.860 194.235 ;
        RECT 70.150 194.045 70.320 194.235 ;
        RECT 72.455 194.065 72.625 194.255 ;
        RECT 72.915 194.065 73.085 194.255 ;
        RECT 74.295 194.065 74.465 194.255 ;
        RECT 78.030 194.095 78.150 194.205 ;
        RECT 80.275 194.045 80.445 194.235 ;
        RECT 83.495 194.065 83.665 194.255 ;
        RECT 89.935 194.045 90.105 194.235 ;
        RECT 91.775 194.045 91.945 194.235 ;
        RECT 93.155 194.045 93.325 194.255 ;
        RECT 93.670 194.095 93.790 194.205 ;
        RECT 94.535 194.045 94.705 194.235 ;
        RECT 95.050 194.095 95.170 194.205 ;
        RECT 98.860 194.045 99.030 194.235 ;
        RECT 100.515 194.045 100.685 194.235 ;
        RECT 101.895 194.045 102.065 194.235 ;
        RECT 102.815 194.065 102.985 194.255 ;
        RECT 104.195 194.100 104.355 194.210 ;
        RECT 106.495 194.045 106.665 194.235 ;
        RECT 109.715 194.065 109.885 194.255 ;
        RECT 111.095 194.065 111.265 194.255 ;
        RECT 115.695 194.045 115.865 194.235 ;
        RECT 116.615 194.045 116.785 194.235 ;
        RECT 118.455 194.090 118.615 194.200 ;
        RECT 120.295 194.065 120.465 194.255 ;
        RECT 122.135 194.045 122.305 194.255 ;
        RECT 127.655 194.045 127.825 194.255 ;
        RECT 129.035 194.045 129.205 194.255 ;
        RECT 9.295 193.235 10.665 194.045 ;
        RECT 11.135 193.235 12.965 194.045 ;
        RECT 12.985 193.175 13.415 193.960 ;
        RECT 14.355 193.235 18.025 194.045 ;
        RECT 18.035 193.235 23.545 194.045 ;
        RECT 23.555 193.235 29.065 194.045 ;
        RECT 29.075 193.235 34.585 194.045 ;
        RECT 34.825 193.365 38.725 194.045 ;
        RECT 37.795 193.135 38.725 193.365 ;
        RECT 38.745 193.175 39.175 193.960 ;
        RECT 39.195 193.365 48.385 194.045 ;
        RECT 43.705 193.145 44.635 193.365 ;
        RECT 47.465 193.135 48.385 193.365 ;
        RECT 48.855 193.365 58.045 194.045 ;
        RECT 48.855 193.135 49.775 193.365 ;
        RECT 52.605 193.145 53.535 193.365 ;
        RECT 58.515 193.235 62.185 194.045 ;
        RECT 62.205 193.135 63.555 194.045 ;
        RECT 64.505 193.175 64.935 193.960 ;
        RECT 65.415 193.365 67.705 194.045 ;
        RECT 65.415 193.135 66.335 193.365 ;
        RECT 67.715 193.135 70.005 194.045 ;
        RECT 70.035 193.135 71.385 194.045 ;
        RECT 71.395 193.365 80.585 194.045 ;
        RECT 80.965 193.365 90.245 194.045 ;
        RECT 71.395 193.135 72.315 193.365 ;
        RECT 75.145 193.145 76.075 193.365 ;
        RECT 80.965 193.245 83.300 193.365 ;
        RECT 80.965 193.135 81.885 193.245 ;
        RECT 87.965 193.145 88.885 193.365 ;
        RECT 90.265 193.175 90.695 193.960 ;
        RECT 90.725 193.135 92.075 194.045 ;
        RECT 92.105 193.135 93.455 194.045 ;
        RECT 93.475 193.265 94.845 194.045 ;
        RECT 95.545 193.365 99.445 194.045 ;
        RECT 98.515 193.135 99.445 193.365 ;
        RECT 99.455 193.235 100.825 194.045 ;
        RECT 100.845 193.135 102.195 194.045 ;
        RECT 103.135 193.235 106.805 194.045 ;
        RECT 106.815 193.365 116.005 194.045 ;
        RECT 106.815 193.135 107.735 193.365 ;
        RECT 110.565 193.145 111.495 193.365 ;
        RECT 116.025 193.175 116.455 193.960 ;
        RECT 116.475 193.265 117.845 194.045 ;
        RECT 118.775 193.235 122.445 194.045 ;
        RECT 122.455 193.235 127.965 194.045 ;
        RECT 127.975 193.235 129.345 194.045 ;
      LAYER nwell ;
        RECT 9.100 190.015 129.540 192.845 ;
      LAYER pwell ;
        RECT 9.295 188.815 10.665 189.625 ;
        RECT 11.135 188.815 14.805 189.625 ;
        RECT 14.815 188.815 20.325 189.625 ;
        RECT 20.335 188.815 25.845 189.625 ;
        RECT 25.865 188.900 26.295 189.685 ;
        RECT 26.775 188.815 29.525 189.625 ;
        RECT 29.545 188.815 30.895 189.725 ;
        RECT 31.285 189.615 32.205 189.725 ;
        RECT 31.285 189.495 33.620 189.615 ;
        RECT 38.285 189.495 39.205 189.715 ;
        RECT 31.285 188.815 40.565 189.495 ;
        RECT 40.575 188.815 41.945 189.595 ;
        RECT 42.415 189.495 43.335 189.725 ;
        RECT 46.165 189.495 47.095 189.715 ;
        RECT 42.415 188.815 51.605 189.495 ;
        RECT 51.625 188.900 52.055 189.685 ;
        RECT 52.085 188.815 53.435 189.725 ;
        RECT 53.455 188.815 56.205 189.625 ;
        RECT 56.215 188.815 61.725 189.625 ;
        RECT 62.025 188.815 64.945 189.725 ;
        RECT 64.955 189.525 65.885 189.725 ;
        RECT 67.220 189.525 68.165 189.725 ;
        RECT 64.955 189.045 68.165 189.525 ;
        RECT 65.095 188.845 68.165 189.045 ;
        RECT 9.435 188.605 9.605 188.815 ;
        RECT 10.870 188.655 10.990 188.765 ;
        RECT 12.655 188.605 12.825 188.795 ;
        RECT 14.495 188.605 14.665 188.815 ;
        RECT 20.015 188.605 20.185 188.815 ;
        RECT 20.475 188.605 20.645 188.795 ;
        RECT 25.535 188.625 25.705 188.815 ;
        RECT 26.510 188.655 26.630 188.765 ;
        RECT 29.215 188.625 29.385 188.815 ;
        RECT 29.675 188.625 29.845 188.815 ;
        RECT 30.595 188.605 30.765 188.795 ;
        RECT 31.975 188.605 32.145 188.795 ;
        RECT 33.815 188.605 33.985 188.795 ;
        RECT 37.680 188.605 37.850 188.795 ;
        RECT 38.470 188.655 38.590 188.765 ;
        RECT 39.390 188.655 39.510 188.765 ;
        RECT 40.255 188.625 40.425 188.815 ;
        RECT 41.635 188.625 41.805 188.815 ;
        RECT 42.095 188.765 42.265 188.795 ;
        RECT 42.095 188.655 42.270 188.765 ;
        RECT 42.095 188.605 42.265 188.655 ;
        RECT 47.615 188.605 47.785 188.795 ;
        RECT 48.075 188.605 48.245 188.795 ;
        RECT 51.295 188.625 51.465 188.815 ;
        RECT 52.860 188.605 53.030 188.795 ;
        RECT 53.135 188.625 53.305 188.815 ;
        RECT 55.895 188.625 56.065 188.815 ;
        RECT 58.655 188.605 58.825 188.795 ;
        RECT 61.415 188.625 61.585 188.815 ;
        RECT 64.175 188.605 64.345 188.795 ;
        RECT 64.630 188.625 64.800 188.815 ;
        RECT 65.095 188.625 65.265 188.845 ;
        RECT 67.220 188.815 68.165 188.845 ;
        RECT 68.175 189.525 69.120 189.725 ;
        RECT 70.455 189.525 71.385 189.725 ;
        RECT 68.175 189.045 71.385 189.525 ;
        RECT 72.445 189.495 73.375 189.725 ;
        RECT 68.175 188.845 71.245 189.045 ;
        RECT 68.175 188.815 69.120 188.845 ;
        RECT 65.555 188.650 65.715 188.760 ;
        RECT 69.235 188.605 69.405 188.795 ;
        RECT 71.075 188.605 71.245 188.845 ;
        RECT 71.540 188.815 73.375 189.495 ;
        RECT 73.695 189.495 74.615 189.725 ;
        RECT 73.695 188.815 75.985 189.495 ;
        RECT 75.995 188.815 77.365 189.625 ;
        RECT 77.385 188.900 77.815 189.685 ;
        RECT 77.835 188.815 80.585 189.625 ;
        RECT 80.595 188.815 86.105 189.625 ;
        RECT 89.315 189.495 90.245 189.725 ;
        RECT 86.345 188.815 90.245 189.495 ;
        RECT 90.255 188.815 91.625 189.595 ;
        RECT 92.095 188.815 93.925 189.625 ;
        RECT 98.445 189.495 99.375 189.715 ;
        RECT 102.205 189.495 103.125 189.725 ;
        RECT 93.935 188.815 103.125 189.495 ;
        RECT 103.145 188.900 103.575 189.685 ;
        RECT 103.595 188.815 104.965 189.625 ;
        RECT 104.975 188.815 110.485 189.625 ;
        RECT 113.695 189.495 114.625 189.725 ;
        RECT 110.725 188.815 114.625 189.495 ;
        RECT 114.635 188.815 116.005 189.595 ;
        RECT 116.935 188.815 122.445 189.625 ;
        RECT 122.455 188.815 127.965 189.625 ;
        RECT 127.975 188.815 129.345 189.625 ;
        RECT 71.540 188.795 71.705 188.815 ;
        RECT 71.535 188.625 71.705 188.795 ;
        RECT 75.675 188.625 75.845 188.815 ;
        RECT 77.055 188.625 77.225 188.815 ;
        RECT 80.275 188.605 80.445 188.815 ;
        RECT 81.655 188.605 81.825 188.795 ;
        RECT 85.335 188.605 85.505 188.795 ;
        RECT 85.795 188.625 85.965 188.815 ;
        RECT 89.200 188.605 89.370 188.795 ;
        RECT 89.660 188.625 89.830 188.815 ;
        RECT 89.990 188.655 90.110 188.765 ;
        RECT 91.315 188.625 91.485 188.815 ;
        RECT 91.775 188.765 91.945 188.795 ;
        RECT 91.775 188.655 91.950 188.765 ;
        RECT 91.775 188.605 91.945 188.655 ;
        RECT 93.615 188.625 93.785 188.815 ;
        RECT 94.075 188.625 94.245 188.815 ;
        RECT 95.455 188.605 95.625 188.795 ;
        RECT 100.975 188.605 101.145 188.795 ;
        RECT 102.355 188.605 102.525 188.795 ;
        RECT 103.090 188.605 103.260 188.795 ;
        RECT 104.655 188.625 104.825 188.815 ;
        RECT 109.255 188.605 109.425 188.795 ;
        RECT 110.175 188.625 110.345 188.815 ;
        RECT 113.120 188.605 113.290 188.795 ;
        RECT 113.910 188.655 114.030 188.765 ;
        RECT 114.040 188.625 114.210 188.815 ;
        RECT 115.695 188.605 115.865 188.815 ;
        RECT 116.615 188.765 116.775 188.770 ;
        RECT 116.615 188.660 116.790 188.765 ;
        RECT 116.670 188.655 116.790 188.660 ;
        RECT 122.135 188.605 122.305 188.815 ;
        RECT 127.655 188.605 127.825 188.815 ;
        RECT 129.035 188.605 129.205 188.815 ;
        RECT 9.295 187.795 10.665 188.605 ;
        RECT 11.135 187.795 12.965 188.605 ;
        RECT 12.985 187.735 13.415 188.520 ;
        RECT 13.435 187.795 14.805 188.605 ;
        RECT 14.815 187.795 20.325 188.605 ;
        RECT 20.345 187.695 21.695 188.605 ;
        RECT 21.715 187.925 30.905 188.605 ;
        RECT 21.715 187.695 22.635 187.925 ;
        RECT 25.465 187.705 26.395 187.925 ;
        RECT 30.915 187.825 32.285 188.605 ;
        RECT 32.295 187.795 34.125 188.605 ;
        RECT 34.365 187.925 38.265 188.605 ;
        RECT 37.335 187.695 38.265 187.925 ;
        RECT 38.745 187.735 39.175 188.520 ;
        RECT 39.655 187.795 42.405 188.605 ;
        RECT 42.415 187.795 47.925 188.605 ;
        RECT 47.935 187.825 49.305 188.605 ;
        RECT 49.545 187.925 53.445 188.605 ;
        RECT 52.515 187.695 53.445 187.925 ;
        RECT 53.455 187.795 58.965 188.605 ;
        RECT 58.975 187.795 64.485 188.605 ;
        RECT 64.505 187.735 64.935 188.520 ;
        RECT 65.875 187.795 69.545 188.605 ;
        RECT 69.555 187.925 71.385 188.605 ;
        RECT 71.395 187.925 80.585 188.605 ;
        RECT 69.555 187.695 70.900 187.925 ;
        RECT 71.395 187.695 72.315 187.925 ;
        RECT 75.145 187.705 76.075 187.925 ;
        RECT 80.595 187.795 81.965 188.605 ;
        RECT 81.975 187.795 85.645 188.605 ;
        RECT 85.885 187.925 89.785 188.605 ;
        RECT 88.855 187.695 89.785 187.925 ;
        RECT 90.265 187.735 90.695 188.520 ;
        RECT 90.715 187.795 92.085 188.605 ;
        RECT 92.095 187.795 95.765 188.605 ;
        RECT 95.775 187.795 101.285 188.605 ;
        RECT 101.295 187.825 102.665 188.605 ;
        RECT 102.675 187.925 106.575 188.605 ;
        RECT 102.675 187.695 103.605 187.925 ;
        RECT 106.815 187.795 109.565 188.605 ;
        RECT 109.805 187.925 113.705 188.605 ;
        RECT 112.775 187.695 113.705 187.925 ;
        RECT 114.175 187.795 116.005 188.605 ;
        RECT 116.025 187.735 116.455 188.520 ;
        RECT 116.935 187.795 122.445 188.605 ;
        RECT 122.455 187.795 127.965 188.605 ;
        RECT 127.975 187.795 129.345 188.605 ;
      LAYER nwell ;
        RECT 9.100 184.575 129.540 187.405 ;
      LAYER pwell ;
        RECT 9.295 183.375 10.665 184.185 ;
        RECT 11.135 183.375 14.805 184.185 ;
        RECT 14.815 183.375 20.325 184.185 ;
        RECT 20.335 183.375 25.845 184.185 ;
        RECT 25.865 183.460 26.295 184.245 ;
        RECT 29.515 184.055 30.445 184.285 ;
        RECT 26.545 183.375 30.445 184.055 ;
        RECT 30.455 183.375 34.125 184.185 ;
        RECT 34.135 184.055 35.055 184.285 ;
        RECT 37.885 184.055 38.815 184.275 ;
        RECT 34.135 183.375 43.325 184.055 ;
        RECT 43.795 183.375 46.545 184.185 ;
        RECT 46.555 184.055 47.485 184.285 ;
        RECT 46.555 183.375 50.455 184.055 ;
        RECT 51.625 183.460 52.055 184.245 ;
        RECT 52.545 183.375 53.895 184.285 ;
        RECT 53.915 183.375 55.285 184.185 ;
        RECT 55.295 183.375 60.805 184.185 ;
        RECT 60.815 183.375 66.325 184.185 ;
        RECT 68.175 184.055 69.105 184.285 ;
        RECT 66.335 183.375 68.165 184.055 ;
        RECT 68.175 183.375 71.845 184.055 ;
        RECT 71.855 183.375 73.685 184.185 ;
        RECT 73.695 183.375 75.065 184.155 ;
        RECT 75.085 183.375 76.435 184.285 ;
        RECT 77.385 183.460 77.815 184.245 ;
        RECT 78.295 183.375 81.045 184.185 ;
        RECT 81.055 183.375 86.565 184.185 ;
        RECT 89.775 184.055 90.705 184.285 ;
        RECT 86.805 183.375 90.705 184.055 ;
        RECT 90.715 183.375 92.085 184.185 ;
        RECT 92.095 183.375 95.765 184.185 ;
        RECT 98.975 184.055 99.905 184.285 ;
        RECT 96.005 183.375 99.905 184.055 ;
        RECT 100.375 183.375 103.125 184.185 ;
        RECT 103.145 183.460 103.575 184.245 ;
        RECT 103.595 183.375 105.425 184.185 ;
        RECT 105.435 183.375 110.945 184.185 ;
        RECT 110.955 183.375 116.465 184.185 ;
        RECT 116.485 183.375 117.835 184.285 ;
        RECT 117.865 183.375 119.215 184.285 ;
        RECT 120.155 183.375 121.525 184.155 ;
        RECT 122.455 183.375 127.965 184.185 ;
        RECT 127.975 183.375 129.345 184.185 ;
        RECT 9.435 183.165 9.605 183.375 ;
        RECT 10.870 183.215 10.990 183.325 ;
        RECT 12.655 183.165 12.825 183.355 ;
        RECT 13.630 183.215 13.750 183.325 ;
        RECT 14.495 183.185 14.665 183.375 ;
        RECT 15.415 183.165 15.585 183.355 ;
        RECT 20.015 183.185 20.185 183.375 ;
        RECT 20.935 183.165 21.105 183.355 ;
        RECT 21.395 183.165 21.565 183.355 ;
        RECT 25.535 183.185 25.705 183.375 ;
        RECT 25.995 183.165 26.165 183.355 ;
        RECT 27.375 183.165 27.545 183.355 ;
        RECT 29.860 183.185 30.030 183.375 ;
        RECT 30.135 183.165 30.305 183.355 ;
        RECT 33.815 183.185 33.985 183.375 ;
        RECT 35.655 183.165 35.825 183.355 ;
        RECT 36.115 183.165 36.285 183.355 ;
        RECT 37.495 183.165 37.665 183.355 ;
        RECT 39.610 183.165 39.780 183.355 ;
        RECT 43.015 183.185 43.185 183.375 ;
        RECT 43.530 183.215 43.650 183.325 ;
        RECT 46.235 183.185 46.405 183.375 ;
        RECT 46.970 183.185 47.140 183.375 ;
        RECT 48.995 183.165 49.165 183.355 ;
        RECT 51.295 183.220 51.455 183.330 ;
        RECT 52.270 183.215 52.390 183.325 ;
        RECT 53.595 183.185 53.765 183.375 ;
        RECT 54.975 183.185 55.145 183.375 ;
        RECT 58.195 183.165 58.365 183.355 ;
        RECT 58.710 183.215 58.830 183.325 ;
        RECT 60.495 183.185 60.665 183.375 ;
        RECT 64.175 183.165 64.345 183.355 ;
        RECT 65.555 183.210 65.715 183.320 ;
        RECT 66.015 183.185 66.185 183.375 ;
        RECT 67.395 183.165 67.565 183.355 ;
        RECT 67.855 183.185 68.025 183.375 ;
        RECT 71.535 183.185 71.705 183.375 ;
        RECT 71.995 183.165 72.165 183.355 ;
        RECT 72.915 183.210 73.075 183.320 ;
        RECT 73.375 183.165 73.545 183.375 ;
        RECT 73.835 183.185 74.005 183.375 ;
        RECT 75.675 183.165 75.845 183.355 ;
        RECT 76.135 183.185 76.305 183.375 ;
        RECT 77.055 183.165 77.225 183.355 ;
        RECT 78.030 183.215 78.150 183.325 ;
        RECT 80.735 183.165 80.905 183.375 ;
        RECT 86.255 183.185 86.425 183.375 ;
        RECT 89.935 183.165 90.105 183.355 ;
        RECT 90.120 183.185 90.290 183.375 ;
        RECT 91.775 183.165 91.945 183.375 ;
        RECT 92.290 183.215 92.410 183.325 ;
        RECT 95.455 183.185 95.625 183.375 ;
        RECT 99.320 183.185 99.490 183.375 ;
        RECT 100.110 183.215 100.230 183.325 ;
        RECT 101.435 183.165 101.605 183.355 ;
        RECT 102.355 183.210 102.515 183.320 ;
        RECT 102.815 183.185 102.985 183.375 ;
        RECT 105.115 183.185 105.285 183.375 ;
        RECT 106.035 183.165 106.205 183.355 ;
        RECT 110.635 183.185 110.805 183.375 ;
        RECT 111.555 183.165 111.725 183.355 ;
        RECT 115.420 183.165 115.590 183.355 ;
        RECT 116.155 183.185 116.325 183.375 ;
        RECT 116.615 183.185 116.785 183.375 ;
        RECT 117.995 183.185 118.165 183.375 ;
        RECT 119.835 183.220 119.995 183.330 ;
        RECT 120.295 183.185 120.465 183.375 ;
        RECT 122.135 183.220 122.295 183.330 ;
        RECT 125.355 183.165 125.525 183.355 ;
        RECT 125.870 183.215 125.990 183.325 ;
        RECT 127.655 183.165 127.825 183.375 ;
        RECT 129.035 183.165 129.205 183.375 ;
        RECT 9.295 182.355 10.665 183.165 ;
        RECT 11.135 182.355 12.965 183.165 ;
        RECT 12.985 182.295 13.415 183.080 ;
        RECT 13.895 182.355 15.725 183.165 ;
        RECT 15.735 182.355 21.245 183.165 ;
        RECT 21.265 182.255 22.615 183.165 ;
        RECT 22.635 182.355 26.305 183.165 ;
        RECT 26.315 182.385 27.685 183.165 ;
        RECT 27.695 182.355 30.445 183.165 ;
        RECT 30.455 182.355 35.965 183.165 ;
        RECT 35.985 182.255 37.335 183.165 ;
        RECT 37.355 182.385 38.725 183.165 ;
        RECT 38.745 182.295 39.175 183.080 ;
        RECT 39.195 182.485 43.095 183.165 ;
        RECT 39.195 182.255 40.125 182.485 ;
        RECT 43.795 182.355 49.305 183.165 ;
        RECT 49.315 182.485 58.505 183.165 ;
        RECT 49.315 182.255 50.235 182.485 ;
        RECT 53.065 182.265 53.995 182.485 ;
        RECT 58.975 182.355 64.485 183.165 ;
        RECT 64.505 182.295 64.935 183.080 ;
        RECT 65.875 182.485 67.705 183.165 ;
        RECT 67.725 183.125 68.645 183.165 ;
        RECT 67.715 182.935 68.645 183.125 ;
        RECT 70.735 182.935 72.305 183.165 ;
        RECT 67.715 182.575 72.305 182.935 ;
        RECT 67.725 182.485 72.305 182.575 ;
        RECT 67.725 182.255 70.725 182.485 ;
        RECT 73.245 182.255 74.595 183.165 ;
        RECT 74.625 182.255 75.975 183.165 ;
        RECT 75.995 182.355 77.365 183.165 ;
        RECT 77.375 182.355 81.045 183.165 ;
        RECT 81.055 182.485 90.245 183.165 ;
        RECT 81.055 182.255 81.975 182.485 ;
        RECT 84.805 182.265 85.735 182.485 ;
        RECT 90.265 182.295 90.695 183.080 ;
        RECT 90.715 182.385 92.085 183.165 ;
        RECT 92.555 182.485 101.745 183.165 ;
        RECT 92.555 182.255 93.475 182.485 ;
        RECT 96.305 182.265 97.235 182.485 ;
        RECT 102.675 182.355 106.345 183.165 ;
        RECT 106.355 182.355 111.865 183.165 ;
        RECT 112.105 182.485 116.005 183.165 ;
        RECT 115.075 182.255 116.005 182.485 ;
        RECT 116.025 182.295 116.455 183.080 ;
        RECT 116.475 182.485 125.665 183.165 ;
        RECT 116.475 182.255 117.395 182.485 ;
        RECT 120.225 182.265 121.155 182.485 ;
        RECT 126.135 182.355 127.965 183.165 ;
        RECT 127.975 182.355 129.345 183.165 ;
      LAYER nwell ;
        RECT 9.100 179.135 129.540 181.965 ;
      LAYER pwell ;
        RECT 9.295 177.935 10.665 178.745 ;
        RECT 11.135 177.935 16.645 178.745 ;
        RECT 21.165 178.615 22.095 178.835 ;
        RECT 24.925 178.615 25.845 178.845 ;
        RECT 16.655 177.935 25.845 178.615 ;
        RECT 25.865 178.020 26.295 178.805 ;
        RECT 26.315 178.615 27.245 178.845 ;
        RECT 26.315 177.935 30.215 178.615 ;
        RECT 30.455 177.935 33.930 178.845 ;
        RECT 34.135 177.935 37.610 178.845 ;
        RECT 38.275 177.935 41.945 178.745 ;
        RECT 41.955 177.935 47.465 178.745 ;
        RECT 50.675 178.615 51.605 178.845 ;
        RECT 47.705 177.935 51.605 178.615 ;
        RECT 51.625 178.020 52.055 178.805 ;
        RECT 52.995 177.935 54.365 178.715 ;
        RECT 54.385 177.935 57.125 178.615 ;
        RECT 57.135 177.935 62.645 178.745 ;
        RECT 62.655 177.935 68.165 178.745 ;
        RECT 68.175 178.615 69.095 178.845 ;
        RECT 71.925 178.615 72.855 178.835 ;
        RECT 68.175 177.935 77.365 178.615 ;
        RECT 77.385 178.020 77.815 178.805 ;
        RECT 78.295 177.935 81.045 178.745 ;
        RECT 81.055 177.935 83.795 178.615 ;
        RECT 83.815 177.935 87.485 178.745 ;
        RECT 87.505 177.935 88.855 178.845 ;
        RECT 89.795 177.935 95.305 178.745 ;
        RECT 95.325 177.935 96.675 178.845 ;
        RECT 97.155 177.935 98.985 178.745 ;
        RECT 98.995 177.935 100.365 178.715 ;
        RECT 100.375 177.935 103.125 178.745 ;
        RECT 103.145 178.020 103.575 178.805 ;
        RECT 103.595 177.935 105.425 178.745 ;
        RECT 105.435 177.935 108.910 178.845 ;
        RECT 109.115 177.935 111.865 178.745 ;
        RECT 115.075 178.615 116.005 178.845 ;
        RECT 112.105 177.935 116.005 178.615 ;
        RECT 116.015 178.615 116.935 178.845 ;
        RECT 119.765 178.615 120.695 178.835 ;
        RECT 116.015 177.935 125.205 178.615 ;
        RECT 125.215 177.935 127.965 178.745 ;
        RECT 127.975 177.935 129.345 178.745 ;
        RECT 9.435 177.725 9.605 177.935 ;
        RECT 10.870 177.775 10.990 177.885 ;
        RECT 12.655 177.725 12.825 177.915 ;
        RECT 13.630 177.775 13.750 177.885 ;
        RECT 15.415 177.725 15.585 177.915 ;
        RECT 16.335 177.745 16.505 177.935 ;
        RECT 16.795 177.745 16.965 177.935 ;
        RECT 20.935 177.725 21.105 177.915 ;
        RECT 21.395 177.725 21.565 177.915 ;
        RECT 26.730 177.745 26.900 177.935 ;
        RECT 30.600 177.745 30.770 177.935 ;
        RECT 31.515 177.725 31.685 177.915 ;
        RECT 32.250 177.725 32.420 177.915 ;
        RECT 34.280 177.745 34.450 177.935 ;
        RECT 41.635 177.915 41.805 177.935 ;
        RECT 38.010 177.775 38.130 177.885 ;
        RECT 38.415 177.725 38.585 177.915 ;
        RECT 39.390 177.775 39.510 177.885 ;
        RECT 41.175 177.725 41.345 177.915 ;
        RECT 41.635 177.745 41.810 177.915 ;
        RECT 47.155 177.745 47.325 177.935 ;
        RECT 41.640 177.725 41.810 177.745 ;
        RECT 48.720 177.725 48.890 177.915 ;
        RECT 51.020 177.745 51.190 177.935 ;
        RECT 52.675 177.780 52.835 177.890 ;
        RECT 53.135 177.745 53.305 177.935 ;
        RECT 56.815 177.745 56.985 177.935 ;
        RECT 58.195 177.725 58.365 177.915 ;
        RECT 58.710 177.775 58.830 177.885 ;
        RECT 62.335 177.725 62.505 177.935 ;
        RECT 64.175 177.725 64.345 177.915 ;
        RECT 66.015 177.725 66.185 177.915 ;
        RECT 66.475 177.745 66.645 177.915 ;
        RECT 67.855 177.745 68.025 177.935 ;
        RECT 69.750 177.775 69.870 177.885 ;
        RECT 66.575 177.725 66.645 177.745 ;
        RECT 71.535 177.725 71.705 177.915 ;
        RECT 77.055 177.725 77.225 177.935 ;
        RECT 77.520 177.725 77.690 177.915 ;
        RECT 78.030 177.775 78.150 177.885 ;
        RECT 80.280 177.725 80.450 177.915 ;
        RECT 80.735 177.745 80.905 177.935 ;
        RECT 81.195 177.745 81.365 177.935 ;
        RECT 83.960 177.725 84.130 177.915 ;
        RECT 87.175 177.745 87.345 177.935 ;
        RECT 88.555 177.745 88.725 177.935 ;
        RECT 89.475 177.780 89.635 177.890 ;
        RECT 89.935 177.725 90.105 177.915 ;
        RECT 90.910 177.775 91.030 177.885 ;
        RECT 92.695 177.725 92.865 177.915 ;
        RECT 94.995 177.745 95.165 177.935 ;
        RECT 96.375 177.745 96.545 177.935 ;
        RECT 98.675 177.915 98.845 177.935 ;
        RECT 96.890 177.775 97.010 177.885 ;
        RECT 98.215 177.725 98.385 177.915 ;
        RECT 98.675 177.745 98.850 177.915 ;
        RECT 99.135 177.745 99.305 177.935 ;
        RECT 102.410 177.775 102.530 177.885 ;
        RECT 102.815 177.745 102.985 177.935 ;
        RECT 98.680 177.725 98.850 177.745 ;
        RECT 104.195 177.725 104.365 177.915 ;
        RECT 104.660 177.725 104.830 177.915 ;
        RECT 105.115 177.745 105.285 177.935 ;
        RECT 105.580 177.745 105.750 177.935 ;
        RECT 108.340 177.725 108.510 177.915 ;
        RECT 111.555 177.745 111.725 177.935 ;
        RECT 115.230 177.725 115.400 177.915 ;
        RECT 115.420 177.745 115.590 177.935 ;
        RECT 115.750 177.775 115.870 177.885 ;
        RECT 116.670 177.775 116.790 177.885 ;
        RECT 120.295 177.725 120.465 177.915 ;
        RECT 120.755 177.725 120.925 177.915 ;
        RECT 122.190 177.775 122.310 177.885 ;
        RECT 124.895 177.745 125.065 177.935 ;
        RECT 127.655 177.725 127.825 177.935 ;
        RECT 129.035 177.725 129.205 177.935 ;
        RECT 9.295 176.915 10.665 177.725 ;
        RECT 11.135 176.915 12.965 177.725 ;
        RECT 12.985 176.855 13.415 177.640 ;
        RECT 13.895 176.915 15.725 177.725 ;
        RECT 15.735 176.915 21.245 177.725 ;
        RECT 21.265 176.815 22.615 177.725 ;
        RECT 22.635 177.045 31.825 177.725 ;
        RECT 31.835 177.045 35.735 177.725 ;
        RECT 22.635 176.815 23.555 177.045 ;
        RECT 26.385 176.825 27.315 177.045 ;
        RECT 31.835 176.815 32.765 177.045 ;
        RECT 35.975 176.915 38.725 177.725 ;
        RECT 38.745 176.855 39.175 177.640 ;
        RECT 39.655 176.915 41.485 177.725 ;
        RECT 41.495 176.815 44.970 177.725 ;
        RECT 45.405 177.045 49.305 177.725 ;
        RECT 48.375 176.815 49.305 177.045 ;
        RECT 49.315 177.045 58.505 177.725 ;
        RECT 49.315 176.815 50.235 177.045 ;
        RECT 53.065 176.825 53.995 177.045 ;
        RECT 58.975 176.915 62.645 177.725 ;
        RECT 62.655 177.045 64.485 177.725 ;
        RECT 62.655 176.815 64.000 177.045 ;
        RECT 64.505 176.855 64.935 177.640 ;
        RECT 64.955 176.915 66.325 177.725 ;
        RECT 66.575 177.495 68.845 177.725 ;
        RECT 66.575 176.815 69.330 177.495 ;
        RECT 70.015 176.915 71.845 177.725 ;
        RECT 71.855 176.915 77.365 177.725 ;
        RECT 77.375 176.815 79.985 177.725 ;
        RECT 80.135 176.815 83.610 177.725 ;
        RECT 83.815 176.815 86.425 177.725 ;
        RECT 86.575 176.915 90.245 177.725 ;
        RECT 90.265 176.855 90.695 177.640 ;
        RECT 91.175 176.915 93.005 177.725 ;
        RECT 93.015 176.915 98.525 177.725 ;
        RECT 98.535 176.815 102.010 177.725 ;
        RECT 102.675 176.915 104.505 177.725 ;
        RECT 104.515 176.815 107.990 177.725 ;
        RECT 108.195 176.815 111.670 177.725 ;
        RECT 112.070 176.815 115.545 177.725 ;
        RECT 116.025 176.855 116.455 177.640 ;
        RECT 116.935 176.915 120.605 177.725 ;
        RECT 120.615 176.945 121.985 177.725 ;
        RECT 122.455 176.915 127.965 177.725 ;
        RECT 127.975 176.915 129.345 177.725 ;
      LAYER nwell ;
        RECT 9.100 173.695 129.540 176.525 ;
      LAYER pwell ;
        RECT 9.295 172.495 10.665 173.305 ;
        RECT 11.135 172.495 14.805 173.305 ;
        RECT 14.815 172.495 20.325 173.305 ;
        RECT 20.335 172.495 25.845 173.305 ;
        RECT 25.865 172.580 26.295 173.365 ;
        RECT 26.315 172.495 27.685 173.305 ;
        RECT 27.695 172.495 31.365 173.305 ;
        RECT 31.375 172.495 32.745 173.275 ;
        RECT 32.755 172.495 36.230 173.405 ;
        RECT 36.895 172.495 40.370 173.405 ;
        RECT 40.575 172.495 44.050 173.405 ;
        RECT 44.255 172.495 47.730 173.405 ;
        RECT 47.935 172.495 51.410 173.405 ;
        RECT 51.625 172.580 52.055 173.365 ;
        RECT 52.545 172.495 53.895 173.405 ;
        RECT 54.835 172.495 56.205 173.275 ;
        RECT 56.215 172.495 59.885 173.305 ;
        RECT 59.895 173.175 61.240 173.405 ;
        RECT 61.735 173.175 63.080 173.405 ;
        RECT 59.895 172.495 61.725 173.175 ;
        RECT 61.735 172.495 63.565 173.175 ;
        RECT 63.790 172.725 66.545 173.405 ;
        RECT 64.275 172.495 66.545 172.725 ;
        RECT 9.435 172.285 9.605 172.495 ;
        RECT 10.870 172.335 10.990 172.445 ;
        RECT 12.655 172.285 12.825 172.475 ;
        RECT 13.630 172.335 13.750 172.445 ;
        RECT 14.495 172.305 14.665 172.495 ;
        RECT 16.335 172.285 16.505 172.475 ;
        RECT 20.015 172.305 20.185 172.495 ;
        RECT 21.855 172.285 22.025 172.475 ;
        RECT 25.535 172.305 25.705 172.495 ;
        RECT 27.375 172.285 27.545 172.495 ;
        RECT 31.055 172.305 31.225 172.495 ;
        RECT 32.435 172.305 32.605 172.495 ;
        RECT 32.900 172.475 33.070 172.495 ;
        RECT 32.895 172.305 33.070 172.475 ;
        RECT 36.630 172.335 36.750 172.445 ;
        RECT 37.040 172.305 37.210 172.495 ;
        RECT 32.895 172.285 33.065 172.305 ;
        RECT 38.415 172.285 38.585 172.475 ;
        RECT 39.340 172.285 39.510 172.475 ;
        RECT 40.720 172.305 40.890 172.495 ;
        RECT 43.070 172.335 43.190 172.445 ;
        RECT 44.400 172.305 44.570 172.495 ;
        RECT 45.775 172.285 45.945 172.475 ;
        RECT 46.240 172.285 46.410 172.475 ;
        RECT 48.080 172.305 48.250 172.495 ;
        RECT 51.295 172.285 51.465 172.475 ;
        RECT 52.270 172.335 52.390 172.445 ;
        RECT 53.595 172.305 53.765 172.495 ;
        RECT 54.515 172.340 54.675 172.450 ;
        RECT 54.975 172.305 55.145 172.495 ;
        RECT 56.815 172.285 56.985 172.475 ;
        RECT 59.575 172.305 59.745 172.495 ;
        RECT 61.415 172.305 61.585 172.495 ;
        RECT 62.335 172.285 62.505 172.475 ;
        RECT 62.795 172.285 62.965 172.475 ;
        RECT 63.255 172.305 63.425 172.495 ;
        RECT 66.475 172.475 66.545 172.495 ;
        RECT 67.035 172.725 69.790 173.405 ;
        RECT 67.035 172.495 69.305 172.725 ;
        RECT 70.015 172.495 71.845 173.305 ;
        RECT 71.855 172.495 77.365 173.305 ;
        RECT 77.385 172.580 77.815 173.365 ;
        RECT 78.295 172.495 80.125 173.305 ;
        RECT 80.135 172.495 83.610 173.405 ;
        RECT 83.815 172.495 87.290 173.405 ;
        RECT 87.495 172.495 88.865 173.305 ;
        RECT 88.875 172.495 94.385 173.305 ;
        RECT 94.405 172.495 95.755 173.405 ;
        RECT 95.775 172.495 97.605 173.305 ;
        RECT 97.615 172.495 103.125 173.305 ;
        RECT 103.145 172.580 103.575 173.365 ;
        RECT 104.515 172.495 108.185 173.305 ;
        RECT 108.195 172.495 111.670 173.405 ;
        RECT 111.875 172.495 113.245 173.305 ;
        RECT 113.255 172.495 116.925 173.305 ;
        RECT 116.935 172.495 122.445 173.305 ;
        RECT 122.455 172.495 127.965 173.305 ;
        RECT 127.975 172.495 129.345 173.305 ;
        RECT 67.035 172.475 67.105 172.495 ;
        RECT 66.475 172.305 66.645 172.475 ;
        RECT 66.935 172.305 67.105 172.475 ;
        RECT 69.235 172.285 69.405 172.475 ;
        RECT 69.695 172.285 69.865 172.475 ;
        RECT 71.535 172.305 71.705 172.495 ;
        RECT 74.350 172.335 74.470 172.445 ;
        RECT 77.055 172.305 77.225 172.495 ;
        RECT 78.030 172.335 78.150 172.445 ;
        RECT 79.815 172.285 79.985 172.495 ;
        RECT 80.280 172.285 80.450 172.495 ;
        RECT 83.960 172.305 84.130 172.495 ;
        RECT 84.415 172.330 84.575 172.440 ;
        RECT 88.555 172.305 88.725 172.495 ;
        RECT 89.935 172.285 90.105 172.475 ;
        RECT 90.910 172.335 91.030 172.445 ;
        RECT 91.315 172.285 91.485 172.475 ;
        RECT 94.075 172.305 94.245 172.495 ;
        RECT 94.535 172.305 94.705 172.495 ;
        RECT 97.295 172.305 97.465 172.495 ;
        RECT 101.435 172.285 101.605 172.475 ;
        RECT 101.895 172.285 102.065 172.475 ;
        RECT 102.815 172.305 102.985 172.495 ;
        RECT 103.330 172.335 103.450 172.445 ;
        RECT 104.195 172.340 104.355 172.450 ;
        RECT 107.875 172.305 108.045 172.495 ;
        RECT 108.340 172.305 108.510 172.495 ;
        RECT 108.795 172.285 108.965 172.475 ;
        RECT 110.175 172.285 110.345 172.475 ;
        RECT 112.935 172.305 113.105 172.495 ;
        RECT 115.695 172.285 115.865 172.475 ;
        RECT 116.615 172.445 116.785 172.495 ;
        RECT 116.615 172.335 116.790 172.445 ;
        RECT 116.615 172.305 116.785 172.335 ;
        RECT 117.075 172.285 117.245 172.475 ;
        RECT 118.455 172.285 118.625 172.475 ;
        RECT 119.890 172.335 120.010 172.445 ;
        RECT 122.135 172.305 122.305 172.495 ;
        RECT 122.595 172.285 122.765 172.475 ;
        RECT 124.435 172.285 124.605 172.475 ;
        RECT 124.950 172.335 125.070 172.445 ;
        RECT 127.655 172.285 127.825 172.495 ;
        RECT 129.035 172.285 129.205 172.495 ;
        RECT 9.295 171.475 10.665 172.285 ;
        RECT 11.135 171.475 12.965 172.285 ;
        RECT 12.985 171.415 13.415 172.200 ;
        RECT 13.895 171.475 16.645 172.285 ;
        RECT 16.655 171.475 22.165 172.285 ;
        RECT 22.175 171.475 27.685 172.285 ;
        RECT 27.695 171.475 33.205 172.285 ;
        RECT 33.215 171.475 38.725 172.285 ;
        RECT 38.745 171.415 39.175 172.200 ;
        RECT 39.195 171.375 42.670 172.285 ;
        RECT 43.335 171.475 46.085 172.285 ;
        RECT 46.095 171.375 49.570 172.285 ;
        RECT 49.775 171.475 51.605 172.285 ;
        RECT 51.615 171.475 57.125 172.285 ;
        RECT 57.135 171.475 62.645 172.285 ;
        RECT 62.655 171.605 64.485 172.285 ;
        RECT 63.140 171.375 64.485 171.605 ;
        RECT 64.505 171.415 64.935 172.200 ;
        RECT 64.995 171.375 69.545 172.285 ;
        RECT 69.555 172.055 71.125 172.285 ;
        RECT 73.215 172.245 74.135 172.285 ;
        RECT 73.215 172.055 74.145 172.245 ;
        RECT 69.555 171.695 74.145 172.055 ;
        RECT 69.555 171.605 74.135 171.695 ;
        RECT 71.135 171.375 74.135 171.605 ;
        RECT 74.615 171.475 80.125 172.285 ;
        RECT 80.135 171.375 83.610 172.285 ;
        RECT 84.735 171.475 90.245 172.285 ;
        RECT 90.265 171.415 90.695 172.200 ;
        RECT 91.175 171.605 100.365 172.285 ;
        RECT 95.685 171.385 96.615 171.605 ;
        RECT 99.445 171.375 100.365 171.605 ;
        RECT 100.375 171.475 101.745 172.285 ;
        RECT 101.765 171.375 103.115 172.285 ;
        RECT 103.595 171.475 109.105 172.285 ;
        RECT 109.125 171.375 110.475 172.285 ;
        RECT 110.495 171.475 116.005 172.285 ;
        RECT 116.025 171.415 116.455 172.200 ;
        RECT 116.945 171.375 118.295 172.285 ;
        RECT 118.325 171.375 119.675 172.285 ;
        RECT 120.155 171.475 122.905 172.285 ;
        RECT 122.915 171.605 124.745 172.285 ;
        RECT 125.215 171.475 127.965 172.285 ;
        RECT 127.975 171.475 129.345 172.285 ;
      LAYER nwell ;
        RECT 9.100 168.255 129.540 171.085 ;
      LAYER pwell ;
        RECT 9.295 167.055 10.665 167.865 ;
        RECT 11.135 167.055 14.805 167.865 ;
        RECT 14.815 167.055 20.325 167.865 ;
        RECT 20.335 167.055 25.845 167.865 ;
        RECT 25.865 167.140 26.295 167.925 ;
        RECT 26.775 167.055 28.605 167.865 ;
        RECT 28.615 167.055 34.125 167.865 ;
        RECT 34.135 167.055 39.645 167.865 ;
        RECT 39.665 167.055 41.015 167.965 ;
        RECT 41.955 167.055 45.625 167.865 ;
        RECT 45.635 167.055 48.795 167.965 ;
        RECT 48.855 167.055 51.605 167.865 ;
        RECT 51.625 167.140 52.055 167.925 ;
        RECT 52.075 167.055 53.445 167.865 ;
        RECT 53.455 167.055 58.965 167.865 ;
        RECT 58.975 167.055 64.485 167.865 ;
        RECT 64.505 167.055 65.855 167.965 ;
        RECT 66.360 167.735 67.705 167.965 ;
        RECT 65.875 167.055 67.705 167.735 ;
        RECT 67.955 167.285 70.710 167.965 ;
        RECT 67.955 167.055 70.225 167.285 ;
        RECT 71.855 167.055 77.365 167.865 ;
        RECT 77.385 167.140 77.815 167.925 ;
        RECT 78.295 167.055 81.045 167.865 ;
        RECT 84.255 167.735 85.185 167.965 ;
        RECT 81.285 167.055 85.185 167.735 ;
        RECT 86.125 167.055 87.475 167.965 ;
        RECT 88.415 167.055 92.085 167.865 ;
        RECT 95.295 167.735 96.225 167.965 ;
        RECT 92.325 167.055 96.225 167.735 ;
        RECT 96.695 167.055 98.065 167.835 ;
        RECT 102.195 167.735 103.125 167.965 ;
        RECT 99.225 167.055 103.125 167.735 ;
        RECT 103.145 167.140 103.575 167.925 ;
        RECT 103.595 167.735 104.515 167.965 ;
        RECT 107.345 167.735 108.275 167.955 ;
        RECT 115.995 167.735 116.925 167.965 ;
        RECT 103.595 167.055 112.785 167.735 ;
        RECT 113.025 167.055 116.925 167.735 ;
        RECT 116.935 167.735 117.855 167.965 ;
        RECT 120.685 167.735 121.615 167.955 ;
        RECT 116.935 167.055 126.125 167.735 ;
        RECT 126.135 167.055 127.965 167.865 ;
        RECT 127.975 167.055 129.345 167.865 ;
        RECT 9.435 166.845 9.605 167.055 ;
        RECT 10.870 166.895 10.990 167.005 ;
        RECT 12.655 166.845 12.825 167.035 ;
        RECT 14.495 166.845 14.665 167.055 ;
        RECT 14.955 166.845 15.125 167.035 ;
        RECT 20.015 166.865 20.185 167.055 ;
        RECT 25.075 166.845 25.245 167.035 ;
        RECT 25.535 167.005 25.705 167.055 ;
        RECT 25.535 166.895 25.710 167.005 ;
        RECT 26.510 166.895 26.630 167.005 ;
        RECT 25.535 166.865 25.705 166.895 ;
        RECT 27.375 166.845 27.545 167.035 ;
        RECT 27.835 166.845 28.005 167.035 ;
        RECT 28.295 166.865 28.465 167.055 ;
        RECT 33.815 166.865 33.985 167.055 ;
        RECT 37.955 166.845 38.125 167.035 ;
        RECT 39.335 167.005 39.505 167.055 ;
        RECT 38.470 166.895 38.590 167.005 ;
        RECT 39.335 166.895 39.510 167.005 ;
        RECT 39.335 166.865 39.505 166.895 ;
        RECT 39.795 166.845 39.965 167.035 ;
        RECT 40.715 166.865 40.885 167.055 ;
        RECT 41.635 166.900 41.795 167.010 ;
        RECT 45.315 166.865 45.485 167.055 ;
        RECT 48.535 166.865 48.705 167.055 ;
        RECT 49.050 166.895 49.170 167.005 ;
        RECT 50.375 166.845 50.545 167.035 ;
        RECT 51.295 166.865 51.465 167.055 ;
        RECT 52.215 166.845 52.385 167.035 ;
        RECT 53.135 166.865 53.305 167.055 ;
        RECT 54.970 166.845 55.140 167.035 ;
        RECT 56.355 166.845 56.525 167.035 ;
        RECT 58.655 166.865 58.825 167.055 ;
        RECT 59.110 166.845 59.280 167.035 ;
        RECT 60.495 166.845 60.665 167.035 ;
        RECT 64.175 166.845 64.345 167.055 ;
        RECT 64.635 166.865 64.805 167.055 ;
        RECT 65.150 166.895 65.270 167.005 ;
        RECT 66.015 166.865 66.185 167.055 ;
        RECT 67.955 167.035 68.025 167.055 ;
        RECT 67.855 166.845 68.025 167.035 ;
        RECT 69.695 166.845 69.865 167.035 ;
        RECT 71.535 166.900 71.695 167.010 ;
        RECT 73.375 166.845 73.545 167.035 ;
        RECT 77.055 166.865 77.225 167.055 ;
        RECT 78.030 166.895 78.150 167.005 ;
        RECT 78.895 166.845 79.065 167.035 ;
        RECT 79.355 166.845 79.525 167.035 ;
        RECT 80.735 166.865 80.905 167.055 ;
        RECT 84.600 166.865 84.770 167.055 ;
        RECT 85.795 166.900 85.955 167.010 ;
        RECT 87.175 166.865 87.345 167.055 ;
        RECT 88.095 166.900 88.255 167.010 ;
        RECT 89.935 166.845 90.105 167.035 ;
        RECT 91.775 166.845 91.945 167.055 ;
        RECT 92.290 166.895 92.410 167.005 ;
        RECT 94.995 166.845 95.165 167.035 ;
        RECT 95.455 166.845 95.625 167.035 ;
        RECT 95.640 166.865 95.810 167.055 ;
        RECT 96.430 166.895 96.550 167.005 ;
        RECT 97.755 166.865 97.925 167.055 ;
        RECT 98.675 166.900 98.835 167.010 ;
        RECT 102.540 166.865 102.710 167.055 ;
        RECT 106.035 166.845 106.205 167.035 ;
        RECT 112.475 166.865 112.645 167.055 ;
        RECT 115.235 166.845 115.405 167.035 ;
        RECT 115.750 166.895 115.870 167.005 ;
        RECT 116.340 166.865 116.510 167.055 ;
        RECT 125.355 166.845 125.525 167.035 ;
        RECT 125.815 166.865 125.985 167.055 ;
        RECT 126.735 166.845 126.905 167.035 ;
        RECT 127.655 166.865 127.825 167.055 ;
        RECT 129.035 166.845 129.205 167.055 ;
        RECT 9.295 166.035 10.665 166.845 ;
        RECT 11.135 166.035 12.965 166.845 ;
        RECT 12.985 165.975 13.415 166.760 ;
        RECT 13.435 166.035 14.805 166.845 ;
        RECT 14.815 166.165 24.005 166.845 ;
        RECT 19.325 165.945 20.255 166.165 ;
        RECT 23.085 165.935 24.005 166.165 ;
        RECT 24.025 165.935 25.375 166.845 ;
        RECT 25.855 166.035 27.685 166.845 ;
        RECT 27.705 165.935 29.055 166.845 ;
        RECT 29.075 166.165 38.265 166.845 ;
        RECT 29.075 165.935 29.995 166.165 ;
        RECT 32.825 165.945 33.755 166.165 ;
        RECT 38.745 165.975 39.175 166.760 ;
        RECT 39.655 166.165 48.760 166.845 ;
        RECT 49.325 165.935 50.675 166.845 ;
        RECT 50.695 166.035 52.525 166.845 ;
        RECT 52.675 165.935 55.285 166.845 ;
        RECT 55.295 166.035 56.665 166.845 ;
        RECT 56.815 165.935 59.425 166.845 ;
        RECT 59.435 166.035 60.805 166.845 ;
        RECT 60.815 166.035 64.485 166.845 ;
        RECT 64.505 165.975 64.935 166.760 ;
        RECT 65.415 166.035 68.165 166.845 ;
        RECT 68.175 166.165 70.005 166.845 ;
        RECT 68.175 165.935 69.520 166.165 ;
        RECT 70.015 166.035 73.685 166.845 ;
        RECT 73.695 166.035 79.205 166.845 ;
        RECT 79.215 166.065 80.585 166.845 ;
        RECT 80.965 166.165 90.245 166.845 ;
        RECT 80.965 166.045 83.300 166.165 ;
        RECT 80.965 165.935 81.885 166.045 ;
        RECT 87.965 165.945 88.885 166.165 ;
        RECT 90.265 165.975 90.695 166.760 ;
        RECT 90.715 166.065 92.085 166.845 ;
        RECT 92.555 166.035 95.305 166.845 ;
        RECT 95.315 166.165 104.420 166.845 ;
        RECT 104.515 166.035 106.345 166.845 ;
        RECT 106.355 166.165 115.545 166.845 ;
        RECT 106.355 165.935 107.275 166.165 ;
        RECT 110.105 165.945 111.035 166.165 ;
        RECT 116.025 165.975 116.455 166.760 ;
        RECT 116.475 166.165 125.665 166.845 ;
        RECT 116.475 165.935 117.395 166.165 ;
        RECT 120.225 165.945 121.155 166.165 ;
        RECT 125.675 166.065 127.045 166.845 ;
        RECT 127.975 166.035 129.345 166.845 ;
      LAYER nwell ;
        RECT 9.100 162.815 129.540 165.645 ;
      LAYER pwell ;
        RECT 9.295 161.615 10.665 162.425 ;
        RECT 11.595 161.615 15.265 162.425 ;
        RECT 15.275 161.615 16.645 162.395 ;
        RECT 21.165 162.295 22.095 162.515 ;
        RECT 24.925 162.295 25.845 162.525 ;
        RECT 16.655 161.615 25.845 162.295 ;
        RECT 25.865 161.700 26.295 162.485 ;
        RECT 26.775 162.295 27.705 162.525 ;
        RECT 26.775 161.615 30.675 162.295 ;
        RECT 31.835 161.615 33.205 162.395 ;
        RECT 37.725 162.295 38.655 162.515 ;
        RECT 41.485 162.295 42.405 162.525 ;
        RECT 33.215 161.615 42.405 162.295 ;
        RECT 42.415 162.295 43.335 162.525 ;
        RECT 46.165 162.295 47.095 162.515 ;
        RECT 42.415 161.615 51.605 162.295 ;
        RECT 51.625 161.700 52.055 162.485 ;
        RECT 52.075 161.615 54.825 162.425 ;
        RECT 54.835 161.615 60.345 162.425 ;
        RECT 60.495 161.615 63.105 162.525 ;
        RECT 63.575 161.615 69.085 162.425 ;
        RECT 69.095 161.615 71.815 162.525 ;
        RECT 71.855 161.615 74.595 162.295 ;
        RECT 74.615 161.615 75.985 162.425 ;
        RECT 76.005 161.615 77.355 162.525 ;
        RECT 77.385 161.700 77.815 162.485 ;
        RECT 78.205 162.415 79.125 162.525 ;
        RECT 78.205 162.295 80.540 162.415 ;
        RECT 85.205 162.295 86.125 162.515 ;
        RECT 78.205 161.615 87.485 162.295 ;
        RECT 87.580 161.615 96.685 162.295 ;
        RECT 97.155 161.615 98.985 162.425 ;
        RECT 102.195 162.295 103.125 162.525 ;
        RECT 99.225 161.615 103.125 162.295 ;
        RECT 103.145 161.700 103.575 162.485 ;
        RECT 104.515 161.615 105.885 162.395 ;
        RECT 105.895 161.615 107.265 162.395 ;
        RECT 107.735 161.615 109.565 162.425 ;
        RECT 112.775 162.295 113.705 162.525 ;
        RECT 109.805 161.615 113.705 162.295 ;
        RECT 113.715 161.615 115.085 162.395 ;
        RECT 118.295 162.295 119.225 162.525 ;
        RECT 115.325 161.615 119.225 162.295 ;
        RECT 119.235 161.615 121.065 162.425 ;
        RECT 121.075 161.615 122.445 162.395 ;
        RECT 122.455 161.615 127.965 162.425 ;
        RECT 127.975 161.615 129.345 162.425 ;
        RECT 9.435 161.405 9.605 161.615 ;
        RECT 10.870 161.455 10.990 161.565 ;
        RECT 11.275 161.460 11.435 161.570 ;
        RECT 12.655 161.405 12.825 161.595 ;
        RECT 13.630 161.455 13.750 161.565 ;
        RECT 14.955 161.425 15.125 161.615 ;
        RECT 15.415 161.425 15.585 161.615 ;
        RECT 16.795 161.425 16.965 161.615 ;
        RECT 17.255 161.405 17.425 161.595 ;
        RECT 18.635 161.405 18.805 161.595 ;
        RECT 19.370 161.405 19.540 161.595 ;
        RECT 23.290 161.455 23.410 161.565 ;
        RECT 25.995 161.405 26.165 161.595 ;
        RECT 26.510 161.455 26.630 161.565 ;
        RECT 27.190 161.425 27.360 161.615 ;
        RECT 27.375 161.405 27.545 161.595 ;
        RECT 31.515 161.460 31.675 161.570 ;
        RECT 31.975 161.425 32.145 161.615 ;
        RECT 33.355 161.425 33.525 161.615 ;
        RECT 36.575 161.405 36.745 161.595 ;
        RECT 38.415 161.405 38.585 161.595 ;
        RECT 39.390 161.455 39.510 161.565 ;
        RECT 40.715 161.405 40.885 161.595 ;
        RECT 41.450 161.405 41.620 161.595 ;
        RECT 48.720 161.405 48.890 161.595 ;
        RECT 50.375 161.405 50.545 161.595 ;
        RECT 51.295 161.425 51.465 161.615 ;
        RECT 51.755 161.405 51.925 161.595 ;
        RECT 53.135 161.405 53.305 161.595 ;
        RECT 54.515 161.425 54.685 161.615 ;
        RECT 58.655 161.405 58.825 161.595 ;
        RECT 60.035 161.425 60.205 161.615 ;
        RECT 62.790 161.425 62.960 161.615 ;
        RECT 63.310 161.455 63.430 161.565 ;
        RECT 64.175 161.405 64.345 161.595 ;
        RECT 66.475 161.405 66.645 161.595 ;
        RECT 68.775 161.425 68.945 161.615 ;
        RECT 69.235 161.405 69.405 161.615 ;
        RECT 71.995 161.425 72.165 161.615 ;
        RECT 72.915 161.405 73.085 161.595 ;
        RECT 75.675 161.425 75.845 161.615 ;
        RECT 77.055 161.425 77.225 161.615 ;
        RECT 78.435 161.405 78.605 161.595 ;
        RECT 79.170 161.405 79.340 161.595 ;
        RECT 83.955 161.405 84.125 161.595 ;
        RECT 85.335 161.405 85.505 161.595 ;
        RECT 85.795 161.405 85.965 161.595 ;
        RECT 87.175 161.425 87.345 161.615 ;
        RECT 89.935 161.405 90.105 161.595 ;
        RECT 90.910 161.455 91.030 161.565 ;
        RECT 93.615 161.405 93.785 161.595 ;
        RECT 94.995 161.405 95.165 161.595 ;
        RECT 95.510 161.455 95.630 161.565 ;
        RECT 96.375 161.425 96.545 161.615 ;
        RECT 96.890 161.455 97.010 161.565 ;
        RECT 97.295 161.405 97.465 161.595 ;
        RECT 98.675 161.425 98.845 161.615 ;
        RECT 102.540 161.425 102.710 161.615 ;
        RECT 104.195 161.460 104.355 161.570 ;
        RECT 104.655 161.425 104.825 161.615 ;
        RECT 106.035 161.425 106.205 161.615 ;
        RECT 106.955 161.405 107.125 161.595 ;
        RECT 107.470 161.455 107.590 161.565 ;
        RECT 109.255 161.425 109.425 161.615 ;
        RECT 110.175 161.405 110.345 161.595 ;
        RECT 113.120 161.425 113.290 161.615 ;
        RECT 114.775 161.425 114.945 161.615 ;
        RECT 115.695 161.405 115.865 161.595 ;
        RECT 117.995 161.405 118.165 161.595 ;
        RECT 118.640 161.425 118.810 161.615 ;
        RECT 120.755 161.595 120.925 161.615 ;
        RECT 120.750 161.425 120.925 161.595 ;
        RECT 121.215 161.425 121.385 161.615 ;
        RECT 120.750 161.405 120.920 161.425 ;
        RECT 122.135 161.405 122.305 161.595 ;
        RECT 127.655 161.405 127.825 161.615 ;
        RECT 129.035 161.405 129.205 161.615 ;
        RECT 9.295 160.595 10.665 161.405 ;
        RECT 11.135 160.595 12.965 161.405 ;
        RECT 12.985 160.535 13.415 161.320 ;
        RECT 13.895 160.595 17.565 161.405 ;
        RECT 17.585 160.495 18.935 161.405 ;
        RECT 18.955 160.725 22.855 161.405 ;
        RECT 18.955 160.495 19.885 160.725 ;
        RECT 23.555 160.595 26.305 161.405 ;
        RECT 26.315 160.625 27.685 161.405 ;
        RECT 27.780 160.725 36.885 161.405 ;
        RECT 36.895 160.595 38.725 161.405 ;
        RECT 38.745 160.535 39.175 161.320 ;
        RECT 39.655 160.625 41.025 161.405 ;
        RECT 41.035 160.725 44.935 161.405 ;
        RECT 45.405 160.725 49.305 161.405 ;
        RECT 41.035 160.495 41.965 160.725 ;
        RECT 48.375 160.495 49.305 160.725 ;
        RECT 49.315 160.595 50.685 161.405 ;
        RECT 50.695 160.625 52.065 161.405 ;
        RECT 52.075 160.595 53.445 161.405 ;
        RECT 53.455 160.595 58.965 161.405 ;
        RECT 58.975 160.595 64.485 161.405 ;
        RECT 64.505 160.535 64.935 161.320 ;
        RECT 64.955 160.725 66.785 161.405 ;
        RECT 66.805 160.725 69.545 161.405 ;
        RECT 64.955 160.495 66.300 160.725 ;
        RECT 69.555 160.595 73.225 161.405 ;
        RECT 73.235 160.595 78.745 161.405 ;
        RECT 78.755 160.725 82.655 161.405 ;
        RECT 78.755 160.495 79.685 160.725 ;
        RECT 82.895 160.595 84.265 161.405 ;
        RECT 84.285 160.495 85.635 161.405 ;
        RECT 85.655 160.625 87.025 161.405 ;
        RECT 87.035 160.495 90.195 161.405 ;
        RECT 90.265 160.535 90.695 161.320 ;
        RECT 91.175 160.595 93.925 161.405 ;
        RECT 93.945 160.495 95.295 161.405 ;
        RECT 95.775 160.595 97.605 161.405 ;
        RECT 97.985 160.725 107.265 161.405 ;
        RECT 97.985 160.605 100.320 160.725 ;
        RECT 97.985 160.495 98.905 160.605 ;
        RECT 104.985 160.505 105.905 160.725 ;
        RECT 107.735 160.595 110.485 161.405 ;
        RECT 110.495 160.595 116.005 161.405 ;
        RECT 116.025 160.535 116.455 161.320 ;
        RECT 116.475 160.595 118.305 161.405 ;
        RECT 118.455 160.495 121.065 161.405 ;
        RECT 121.075 160.595 122.445 161.405 ;
        RECT 122.455 160.595 127.965 161.405 ;
        RECT 127.975 160.595 129.345 161.405 ;
      LAYER nwell ;
        RECT 9.100 157.375 129.540 160.205 ;
      LAYER pwell ;
        RECT 9.295 156.175 10.665 156.985 ;
        RECT 11.505 156.975 12.425 157.085 ;
        RECT 11.505 156.855 13.840 156.975 ;
        RECT 18.505 156.855 19.425 157.075 ;
        RECT 11.505 156.175 20.785 156.855 ;
        RECT 20.795 156.175 24.465 156.985 ;
        RECT 24.485 156.175 25.835 157.085 ;
        RECT 25.865 156.260 26.295 157.045 ;
        RECT 29.515 156.855 30.445 157.085 ;
        RECT 34.595 156.855 35.525 157.085 ;
        RECT 26.545 156.175 30.445 156.855 ;
        RECT 31.755 156.175 34.180 156.855 ;
        RECT 34.595 156.175 38.495 156.855 ;
        RECT 38.735 156.175 40.565 156.985 ;
        RECT 40.575 156.175 46.085 156.985 ;
        RECT 46.095 156.175 51.605 156.985 ;
        RECT 51.625 156.260 52.055 157.045 ;
        RECT 52.085 156.175 53.435 157.085 ;
        RECT 53.595 156.175 56.205 157.085 ;
        RECT 56.215 156.855 57.135 157.085 ;
        RECT 59.965 156.855 60.895 157.075 ;
        RECT 56.215 156.175 65.405 156.855 ;
        RECT 65.415 156.175 66.785 156.985 ;
        RECT 66.795 156.855 68.140 157.085 ;
        RECT 69.120 156.855 70.465 157.085 ;
        RECT 70.960 156.855 72.305 157.085 ;
        RECT 66.795 156.175 68.625 156.855 ;
        RECT 68.635 156.175 70.465 156.855 ;
        RECT 70.475 156.175 72.305 156.855 ;
        RECT 72.315 156.175 73.685 156.985 ;
        RECT 73.695 156.175 77.365 156.985 ;
        RECT 77.385 156.260 77.815 157.045 ;
        RECT 78.295 156.175 80.125 156.985 ;
        RECT 80.505 156.975 81.425 157.085 ;
        RECT 80.505 156.855 82.840 156.975 ;
        RECT 87.505 156.855 88.425 157.075 ;
        RECT 90.625 156.975 91.545 157.085 ;
        RECT 90.625 156.855 92.960 156.975 ;
        RECT 97.625 156.855 98.545 157.075 ;
        RECT 80.505 156.175 89.785 156.855 ;
        RECT 90.625 156.175 99.905 156.855 ;
        RECT 99.915 156.175 101.285 156.955 ;
        RECT 101.295 156.175 102.660 156.855 ;
        RECT 103.145 156.260 103.575 157.045 ;
        RECT 103.605 156.175 104.955 157.085 ;
        RECT 105.435 156.175 107.265 156.985 ;
        RECT 107.275 156.175 112.785 156.985 ;
        RECT 112.795 156.175 118.305 156.985 ;
        RECT 118.325 156.175 119.675 157.085 ;
        RECT 119.705 156.175 121.055 157.085 ;
        RECT 121.075 156.175 122.445 156.985 ;
        RECT 122.455 156.175 127.965 156.985 ;
        RECT 127.975 156.175 129.345 156.985 ;
        RECT 9.435 155.965 9.605 156.175 ;
        RECT 10.870 156.015 10.990 156.125 ;
        RECT 12.655 155.965 12.825 156.155 ;
        RECT 14.955 155.965 15.125 156.155 ;
        RECT 16.335 155.965 16.505 156.155 ;
        RECT 18.175 155.965 18.345 156.155 ;
        RECT 19.555 155.965 19.725 156.155 ;
        RECT 20.475 155.985 20.645 156.175 ;
        RECT 22.315 155.965 22.485 156.155 ;
        RECT 24.155 155.985 24.325 156.175 ;
        RECT 24.615 155.985 24.785 156.175 ;
        RECT 29.860 155.985 30.030 156.175 ;
        RECT 31.055 156.020 31.215 156.130 ;
        RECT 31.975 155.965 32.145 156.155 ;
        RECT 32.490 156.015 32.610 156.125 ;
        RECT 34.275 155.965 34.445 156.155 ;
        RECT 34.740 155.965 34.910 156.155 ;
        RECT 35.010 155.985 35.180 156.175 ;
        RECT 38.470 156.015 38.590 156.125 ;
        RECT 39.390 156.015 39.510 156.125 ;
        RECT 40.255 155.985 40.425 156.175 ;
        RECT 44.855 155.965 45.025 156.155 ;
        RECT 45.320 155.965 45.490 156.155 ;
        RECT 45.775 155.985 45.945 156.175 ;
        RECT 49.050 156.015 49.170 156.125 ;
        RECT 51.295 155.985 51.465 156.175 ;
        RECT 51.755 155.965 51.925 156.155 ;
        RECT 52.215 155.985 52.385 156.175 ;
        RECT 55.890 155.985 56.060 156.175 ;
        RECT 61.415 155.965 61.585 156.155 ;
        RECT 61.875 155.965 62.045 156.155 ;
        RECT 64.175 155.965 64.345 156.155 ;
        RECT 65.095 155.985 65.265 156.175 ;
        RECT 66.475 155.965 66.645 156.175 ;
        RECT 68.315 155.965 68.485 156.175 ;
        RECT 68.775 155.985 68.945 156.175 ;
        RECT 70.155 155.965 70.325 156.155 ;
        RECT 70.615 155.985 70.785 156.175 ;
        RECT 71.075 156.010 71.235 156.120 ;
        RECT 73.375 155.985 73.545 156.175 ;
        RECT 77.055 156.155 77.225 156.175 ;
        RECT 76.595 155.965 76.765 156.155 ;
        RECT 77.055 155.985 77.230 156.155 ;
        RECT 78.030 156.015 78.150 156.125 ;
        RECT 79.815 155.985 79.985 156.175 ;
        RECT 81.195 156.010 81.355 156.120 ;
        RECT 77.060 155.965 77.230 155.985 ;
        RECT 85.060 155.965 85.230 156.155 ;
        RECT 86.255 156.010 86.415 156.120 ;
        RECT 89.475 155.985 89.645 156.175 ;
        RECT 89.935 156.125 90.105 156.155 ;
        RECT 89.935 156.015 90.110 156.125 ;
        RECT 90.910 156.015 91.030 156.125 ;
        RECT 89.935 155.965 90.105 156.015 ;
        RECT 93.615 155.965 93.785 156.155 ;
        RECT 97.480 155.965 97.650 156.155 ;
        RECT 98.675 156.010 98.835 156.120 ;
        RECT 99.595 155.985 99.765 156.175 ;
        RECT 100.975 155.985 101.145 156.175 ;
        RECT 102.355 155.965 102.525 156.155 ;
        RECT 102.815 155.985 102.985 156.155 ;
        RECT 104.655 155.985 104.825 156.175 ;
        RECT 105.170 156.015 105.290 156.125 ;
        RECT 106.955 155.985 107.125 156.175 ;
        RECT 107.875 155.965 108.045 156.155 ;
        RECT 108.340 155.965 108.510 156.155 ;
        RECT 112.475 155.985 112.645 156.175 ;
        RECT 112.935 155.965 113.105 156.155 ;
        RECT 113.400 155.965 113.570 156.155 ;
        RECT 116.670 156.015 116.790 156.125 ;
        RECT 117.995 155.985 118.165 156.175 ;
        RECT 118.455 155.985 118.625 156.175 ;
        RECT 119.835 155.985 120.005 156.175 ;
        RECT 122.135 155.985 122.305 156.175 ;
        RECT 125.815 155.965 125.985 156.155 ;
        RECT 127.655 155.965 127.825 156.175 ;
        RECT 129.035 155.965 129.205 156.175 ;
        RECT 9.295 155.155 10.665 155.965 ;
        RECT 11.135 155.155 12.965 155.965 ;
        RECT 12.985 155.095 13.415 155.880 ;
        RECT 13.435 155.155 15.265 155.965 ;
        RECT 15.285 155.055 16.635 155.965 ;
        RECT 16.655 155.155 18.485 155.965 ;
        RECT 18.495 155.185 19.865 155.965 ;
        RECT 19.875 155.155 22.625 155.965 ;
        RECT 23.005 155.285 32.285 155.965 ;
        RECT 23.005 155.165 25.340 155.285 ;
        RECT 23.005 155.055 23.925 155.165 ;
        RECT 30.005 155.065 30.925 155.285 ;
        RECT 32.755 155.155 34.585 155.965 ;
        RECT 34.595 155.055 38.070 155.965 ;
        RECT 38.745 155.095 39.175 155.880 ;
        RECT 39.655 155.155 45.165 155.965 ;
        RECT 45.175 155.055 48.650 155.965 ;
        RECT 49.315 155.155 52.065 155.965 ;
        RECT 52.445 155.285 61.725 155.965 ;
        RECT 52.445 155.165 54.780 155.285 ;
        RECT 52.445 155.055 53.365 155.165 ;
        RECT 59.445 155.065 60.365 155.285 ;
        RECT 61.745 155.055 63.095 155.965 ;
        RECT 63.115 155.155 64.485 155.965 ;
        RECT 64.505 155.095 64.935 155.880 ;
        RECT 64.955 155.155 66.785 155.965 ;
        RECT 66.795 155.285 68.625 155.965 ;
        RECT 68.635 155.285 70.465 155.965 ;
        RECT 66.795 155.055 68.140 155.285 ;
        RECT 68.635 155.055 69.980 155.285 ;
        RECT 71.395 155.155 76.905 155.965 ;
        RECT 76.915 155.055 80.390 155.965 ;
        RECT 81.745 155.285 85.645 155.965 ;
        RECT 84.715 155.055 85.645 155.285 ;
        RECT 86.575 155.155 90.245 155.965 ;
        RECT 90.265 155.095 90.695 155.880 ;
        RECT 91.175 155.155 93.925 155.965 ;
        RECT 94.165 155.285 98.065 155.965 ;
        RECT 97.135 155.055 98.065 155.285 ;
        RECT 98.995 155.155 102.665 155.965 ;
        RECT 102.675 155.155 108.185 155.965 ;
        RECT 108.195 155.055 111.670 155.965 ;
        RECT 111.875 155.155 113.245 155.965 ;
        RECT 113.255 155.055 115.865 155.965 ;
        RECT 116.025 155.095 116.455 155.880 ;
        RECT 116.935 155.285 126.125 155.965 ;
        RECT 116.935 155.055 117.855 155.285 ;
        RECT 120.685 155.065 121.615 155.285 ;
        RECT 126.135 155.155 127.965 155.965 ;
        RECT 127.975 155.155 129.345 155.965 ;
      LAYER nwell ;
        RECT 9.100 151.935 129.540 154.765 ;
      LAYER pwell ;
        RECT 9.295 150.735 10.665 151.545 ;
        RECT 10.675 150.735 16.185 151.545 ;
        RECT 19.395 151.415 20.325 151.645 ;
        RECT 16.425 150.735 20.325 151.415 ;
        RECT 20.335 150.735 25.845 151.545 ;
        RECT 25.865 150.820 26.295 151.605 ;
        RECT 26.775 150.735 29.525 151.545 ;
        RECT 29.535 150.735 30.905 151.515 ;
        RECT 31.375 150.735 34.125 151.545 ;
        RECT 34.330 150.735 37.805 151.645 ;
        RECT 38.010 150.735 41.485 151.645 ;
        RECT 42.610 150.735 46.085 151.645 ;
        RECT 46.095 150.735 51.605 151.545 ;
        RECT 51.625 150.820 52.055 151.605 ;
        RECT 52.075 150.735 53.905 151.545 ;
        RECT 57.115 151.415 58.045 151.645 ;
        RECT 54.145 150.735 58.045 151.415 ;
        RECT 58.055 150.735 59.425 151.515 ;
        RECT 59.895 150.735 62.645 151.545 ;
        RECT 62.655 150.735 64.025 151.515 ;
        RECT 64.495 150.735 67.245 151.545 ;
        RECT 67.740 151.415 69.085 151.645 ;
        RECT 69.580 151.415 70.925 151.645 ;
        RECT 67.255 150.735 69.085 151.415 ;
        RECT 69.095 150.735 70.925 151.415 ;
        RECT 70.935 150.735 73.655 151.645 ;
        RECT 73.890 150.735 77.365 151.645 ;
        RECT 77.385 150.820 77.815 151.605 ;
        RECT 77.835 150.735 81.310 151.645 ;
        RECT 82.435 150.735 86.105 151.545 ;
        RECT 86.115 150.735 91.625 151.545 ;
        RECT 91.635 150.735 97.145 151.545 ;
        RECT 97.155 150.735 100.630 151.645 ;
        RECT 101.295 150.735 103.125 151.545 ;
        RECT 103.145 150.820 103.575 151.605 ;
        RECT 104.055 150.735 105.885 151.545 ;
        RECT 106.090 150.735 109.565 151.645 ;
        RECT 109.770 150.735 113.245 151.645 ;
        RECT 113.255 150.735 116.005 151.545 ;
        RECT 117.765 151.535 118.685 151.645 ;
        RECT 116.015 150.735 117.385 151.515 ;
        RECT 117.765 151.415 120.100 151.535 ;
        RECT 124.765 151.415 125.685 151.635 ;
        RECT 117.765 150.735 127.045 151.415 ;
        RECT 127.975 150.735 129.345 151.545 ;
        RECT 9.435 150.525 9.605 150.735 ;
        RECT 10.870 150.575 10.990 150.685 ;
        RECT 12.655 150.525 12.825 150.715 ;
        RECT 14.495 150.525 14.665 150.715 ;
        RECT 14.955 150.525 15.125 150.715 ;
        RECT 15.875 150.545 16.045 150.735 ;
        RECT 16.610 150.525 16.780 150.715 ;
        RECT 19.740 150.545 19.910 150.735 ;
        RECT 25.535 150.525 25.705 150.735 ;
        RECT 26.510 150.575 26.630 150.685 ;
        RECT 29.215 150.545 29.385 150.735 ;
        RECT 29.675 150.545 29.845 150.735 ;
        RECT 31.055 150.685 31.225 150.715 ;
        RECT 31.055 150.575 31.230 150.685 ;
        RECT 31.055 150.525 31.225 150.575 ;
        RECT 31.520 150.525 31.690 150.715 ;
        RECT 33.815 150.545 33.985 150.735 ;
        RECT 37.490 150.545 37.660 150.735 ;
        RECT 38.410 150.525 38.580 150.715 ;
        RECT 39.795 150.570 39.955 150.680 ;
        RECT 41.170 150.545 41.340 150.735 ;
        RECT 42.095 150.580 42.255 150.690 ;
        RECT 43.475 150.525 43.645 150.715 ;
        RECT 45.770 150.545 45.940 150.735 ;
        RECT 51.295 150.715 51.465 150.735 ;
        RECT 9.295 149.715 10.665 150.525 ;
        RECT 11.135 149.715 12.965 150.525 ;
        RECT 12.985 149.655 13.415 150.440 ;
        RECT 13.445 149.615 14.795 150.525 ;
        RECT 14.815 149.745 16.185 150.525 ;
        RECT 16.195 149.845 20.095 150.525 ;
        RECT 16.195 149.615 17.125 149.845 ;
        RECT 20.335 149.715 25.845 150.525 ;
        RECT 25.855 149.715 31.365 150.525 ;
        RECT 31.375 149.615 34.850 150.525 ;
        RECT 35.250 149.615 38.725 150.525 ;
        RECT 38.745 149.655 39.175 150.440 ;
        RECT 40.115 149.715 43.785 150.525 ;
        RECT 43.795 150.495 44.740 150.525 ;
        RECT 46.230 150.495 46.400 150.715 ;
        RECT 46.555 150.495 47.500 150.525 ;
        RECT 48.990 150.495 49.160 150.715 ;
        RECT 50.835 150.525 51.005 150.715 ;
        RECT 51.295 150.545 51.470 150.715 ;
        RECT 53.595 150.545 53.765 150.735 ;
        RECT 55.435 150.570 55.595 150.680 ;
        RECT 57.460 150.545 57.630 150.735 ;
        RECT 58.195 150.545 58.365 150.735 ;
        RECT 51.300 150.525 51.470 150.545 ;
        RECT 59.115 150.525 59.285 150.715 ;
        RECT 59.630 150.575 59.750 150.685 ;
        RECT 62.335 150.545 62.505 150.735 ;
        RECT 62.795 150.545 62.965 150.735 ;
        RECT 62.980 150.525 63.150 150.715 ;
        RECT 64.230 150.680 64.350 150.685 ;
        RECT 64.175 150.575 64.350 150.680 ;
        RECT 64.175 150.570 64.335 150.575 ;
        RECT 66.475 150.525 66.645 150.715 ;
        RECT 66.935 150.545 67.105 150.735 ;
        RECT 67.395 150.545 67.565 150.735 ;
        RECT 68.315 150.525 68.485 150.715 ;
        RECT 69.235 150.545 69.405 150.735 ;
        RECT 71.075 150.525 71.245 150.735 ;
        RECT 71.535 150.525 71.705 150.715 ;
        RECT 73.430 150.575 73.550 150.685 ;
        RECT 75.215 150.525 75.385 150.715 ;
        RECT 75.675 150.525 75.845 150.715 ;
        RECT 77.050 150.545 77.220 150.735 ;
        RECT 77.980 150.545 78.150 150.735 ;
        RECT 78.440 150.525 78.610 150.715 ;
        RECT 82.115 150.685 82.275 150.690 ;
        RECT 82.115 150.580 82.290 150.685 ;
        RECT 82.170 150.575 82.290 150.580 ;
        RECT 85.795 150.525 85.965 150.735 ;
        RECT 89.660 150.525 89.830 150.715 ;
        RECT 91.315 150.545 91.485 150.735 ;
        RECT 92.235 150.525 92.405 150.715 ;
        RECT 93.615 150.525 93.785 150.715 ;
        RECT 94.130 150.575 94.250 150.685 ;
        RECT 94.535 150.525 94.705 150.715 ;
        RECT 96.835 150.525 97.005 150.735 ;
        RECT 97.300 150.545 97.470 150.735 ;
        RECT 101.030 150.575 101.150 150.685 ;
        RECT 102.355 150.525 102.525 150.715 ;
        RECT 102.815 150.545 102.985 150.735 ;
        RECT 103.790 150.575 103.910 150.685 ;
        RECT 105.575 150.545 105.745 150.735 ;
        RECT 106.030 150.525 106.200 150.715 ;
        RECT 106.500 150.525 106.670 150.715 ;
        RECT 109.250 150.545 109.420 150.735 ;
        RECT 111.555 150.525 111.725 150.715 ;
        RECT 112.930 150.545 113.100 150.735 ;
        RECT 115.420 150.525 115.590 150.715 ;
        RECT 115.695 150.545 115.865 150.735 ;
        RECT 116.155 150.545 116.325 150.735 ;
        RECT 117.075 150.570 117.235 150.680 ;
        RECT 117.810 150.525 117.980 150.715 ;
        RECT 121.675 150.525 121.845 150.715 ;
        RECT 123.975 150.525 124.145 150.715 ;
        RECT 126.735 150.545 126.905 150.735 ;
        RECT 127.655 150.525 127.825 150.715 ;
        RECT 129.035 150.525 129.205 150.735 ;
        RECT 43.795 149.815 46.545 150.495 ;
        RECT 46.555 149.815 49.305 150.495 ;
        RECT 43.795 149.615 44.740 149.815 ;
        RECT 46.555 149.615 47.500 149.815 ;
        RECT 49.315 149.715 51.145 150.525 ;
        RECT 51.155 149.615 54.630 150.525 ;
        RECT 55.755 149.715 59.425 150.525 ;
        RECT 59.665 149.845 63.565 150.525 ;
        RECT 62.635 149.615 63.565 149.845 ;
        RECT 64.505 149.655 64.935 150.440 ;
        RECT 64.955 149.845 66.785 150.525 ;
        RECT 66.795 149.845 68.625 150.525 ;
        RECT 68.645 149.845 71.385 150.525 ;
        RECT 71.395 149.845 73.225 150.525 ;
        RECT 64.955 149.615 66.300 149.845 ;
        RECT 66.795 149.615 68.140 149.845 ;
        RECT 71.880 149.615 73.225 149.845 ;
        RECT 73.695 149.715 75.525 150.525 ;
        RECT 75.535 149.845 78.275 150.525 ;
        RECT 78.295 149.615 81.770 150.525 ;
        RECT 82.435 149.715 86.105 150.525 ;
        RECT 86.345 149.845 90.245 150.525 ;
        RECT 89.315 149.615 90.245 149.845 ;
        RECT 90.265 149.655 90.695 150.440 ;
        RECT 90.715 149.715 92.545 150.525 ;
        RECT 92.565 149.615 93.915 150.525 ;
        RECT 94.395 149.745 95.765 150.525 ;
        RECT 95.775 149.715 97.145 150.525 ;
        RECT 97.155 149.715 102.665 150.525 ;
        RECT 102.870 149.615 106.345 150.525 ;
        RECT 106.355 149.615 109.830 150.525 ;
        RECT 110.035 149.715 111.865 150.525 ;
        RECT 112.105 149.845 116.005 150.525 ;
        RECT 115.075 149.615 116.005 149.845 ;
        RECT 116.025 149.655 116.455 150.440 ;
        RECT 117.395 149.845 121.295 150.525 ;
        RECT 117.395 149.615 118.325 149.845 ;
        RECT 121.535 149.745 122.905 150.525 ;
        RECT 122.915 149.715 124.285 150.525 ;
        RECT 124.295 149.715 127.965 150.525 ;
        RECT 127.975 149.715 129.345 150.525 ;
      LAYER nwell ;
        RECT 9.100 146.495 129.540 149.325 ;
      LAYER pwell ;
        RECT 9.295 145.295 10.665 146.105 ;
        RECT 11.045 146.095 11.965 146.205 ;
        RECT 11.045 145.975 13.380 146.095 ;
        RECT 18.045 145.975 18.965 146.195 ;
        RECT 11.045 145.295 20.325 145.975 ;
        RECT 20.345 145.295 21.695 146.205 ;
        RECT 24.915 145.975 25.845 146.205 ;
        RECT 21.945 145.295 25.845 145.975 ;
        RECT 25.865 145.380 26.295 146.165 ;
        RECT 26.775 145.295 28.145 146.075 ;
        RECT 28.615 145.295 32.285 146.105 ;
        RECT 32.295 146.005 33.240 146.205 ;
        RECT 32.295 145.325 35.045 146.005 ;
        RECT 32.295 145.295 33.240 145.325 ;
        RECT 9.435 145.085 9.605 145.295 ;
        RECT 10.870 145.135 10.990 145.245 ;
        RECT 12.655 145.085 12.825 145.275 ;
        RECT 14.495 145.085 14.665 145.275 ;
        RECT 14.955 145.085 15.125 145.275 ;
        RECT 16.610 145.085 16.780 145.275 ;
        RECT 20.015 145.105 20.185 145.295 ;
        RECT 20.475 145.105 20.645 145.295 ;
        RECT 25.260 145.105 25.430 145.295 ;
        RECT 26.510 145.135 26.630 145.245 ;
        RECT 26.915 145.105 27.085 145.295 ;
        RECT 28.350 145.135 28.470 145.245 ;
        RECT 29.675 145.085 29.845 145.275 ;
        RECT 30.190 145.135 30.310 145.245 ;
        RECT 31.975 145.085 32.145 145.295 ;
        RECT 32.440 145.085 32.610 145.275 ;
        RECT 34.730 145.105 34.900 145.325 ;
        RECT 35.250 145.295 38.725 146.205 ;
        RECT 38.735 145.295 40.565 146.105 ;
        RECT 40.575 145.295 46.085 146.105 ;
        RECT 46.105 145.295 47.455 146.205 ;
        RECT 50.675 145.975 51.605 146.205 ;
        RECT 47.705 145.295 51.605 145.975 ;
        RECT 51.625 145.380 52.055 146.165 ;
        RECT 52.075 145.295 55.550 146.205 ;
        RECT 56.215 145.295 59.885 146.105 ;
        RECT 70.040 145.975 71.385 146.205 ;
        RECT 59.980 145.295 69.085 145.975 ;
        RECT 69.555 145.295 71.385 145.975 ;
        RECT 71.855 145.295 77.365 146.105 ;
        RECT 77.385 145.380 77.815 146.165 ;
        RECT 77.835 146.005 78.780 146.205 ;
        RECT 77.835 145.325 80.585 146.005 ;
        RECT 77.835 145.295 78.780 145.325 ;
        RECT 38.410 145.275 38.580 145.295 ;
        RECT 38.410 145.105 38.585 145.275 ;
        RECT 40.255 145.105 40.425 145.295 ;
        RECT 38.415 145.085 38.585 145.105 ;
        RECT 42.555 145.085 42.725 145.275 ;
        RECT 9.295 144.275 10.665 145.085 ;
        RECT 11.135 144.275 12.965 145.085 ;
        RECT 12.985 144.215 13.415 145.000 ;
        RECT 13.435 144.275 14.805 145.085 ;
        RECT 14.815 144.305 16.185 145.085 ;
        RECT 16.195 144.405 20.095 145.085 ;
        RECT 20.705 144.405 29.985 145.085 ;
        RECT 16.195 144.175 17.125 144.405 ;
        RECT 20.705 144.285 23.040 144.405 ;
        RECT 20.705 144.175 21.625 144.285 ;
        RECT 27.705 144.185 28.625 144.405 ;
        RECT 30.455 144.275 32.285 145.085 ;
        RECT 32.295 144.175 35.770 145.085 ;
        RECT 35.975 144.275 38.725 145.085 ;
        RECT 38.745 144.215 39.175 145.000 ;
        RECT 39.195 144.275 42.865 145.085 ;
        RECT 42.875 145.055 43.820 145.085 ;
        RECT 45.310 145.055 45.480 145.275 ;
        RECT 45.775 145.105 45.945 145.295 ;
        RECT 46.235 145.105 46.405 145.295 ;
        RECT 51.020 145.105 51.190 145.295 ;
        RECT 52.220 145.105 52.390 145.295 ;
        RECT 54.975 145.085 55.145 145.275 ;
        RECT 55.490 145.135 55.610 145.245 ;
        RECT 55.950 145.135 56.070 145.245 ;
        RECT 59.115 145.085 59.285 145.275 ;
        RECT 59.575 145.085 59.745 145.295 ;
        RECT 60.960 145.085 61.130 145.275 ;
        RECT 65.555 145.130 65.715 145.240 ;
        RECT 68.775 145.105 68.945 145.295 ;
        RECT 69.290 145.135 69.410 145.245 ;
        RECT 69.695 145.105 69.865 145.295 ;
        RECT 71.075 145.085 71.245 145.275 ;
        RECT 71.590 145.135 71.710 145.245 ;
        RECT 76.595 145.085 76.765 145.275 ;
        RECT 77.055 145.105 77.225 145.295 ;
        RECT 80.270 145.085 80.440 145.325 ;
        RECT 81.055 145.295 83.805 146.105 ;
        RECT 83.825 145.295 85.175 146.205 ;
        RECT 88.395 145.975 89.325 146.205 ;
        RECT 85.425 145.295 89.325 145.975 ;
        RECT 89.795 145.975 90.715 146.205 ;
        RECT 93.545 145.975 94.475 146.195 ;
        RECT 89.795 145.295 98.985 145.975 ;
        RECT 99.455 145.295 103.125 146.105 ;
        RECT 103.145 145.380 103.575 146.165 ;
        RECT 103.595 146.005 104.540 146.205 ;
        RECT 103.595 145.325 106.345 146.005 ;
        RECT 103.595 145.295 104.540 145.325 ;
        RECT 80.790 145.135 80.910 145.245 ;
        RECT 83.495 145.105 83.665 145.295 ;
        RECT 84.875 145.105 85.045 145.295 ;
        RECT 88.740 145.105 88.910 145.295 ;
        RECT 89.530 145.135 89.650 145.245 ;
        RECT 89.935 145.085 90.105 145.275 ;
        RECT 91.775 145.085 91.945 145.275 ;
        RECT 93.615 145.085 93.785 145.275 ;
        RECT 98.675 145.105 98.845 145.295 ;
        RECT 99.135 145.245 99.305 145.275 ;
        RECT 99.135 145.135 99.310 145.245 ;
        RECT 99.135 145.085 99.305 145.135 ;
        RECT 102.815 145.105 102.985 145.295 ;
        RECT 104.655 145.085 104.825 145.275 ;
        RECT 42.875 144.375 45.625 145.055 ;
        RECT 46.005 144.405 55.285 145.085 ;
        RECT 42.875 144.175 43.820 144.375 ;
        RECT 46.005 144.285 48.340 144.405 ;
        RECT 46.005 144.175 46.925 144.285 ;
        RECT 53.005 144.185 53.925 144.405 ;
        RECT 55.755 144.275 59.425 145.085 ;
        RECT 59.445 144.175 60.795 145.085 ;
        RECT 60.815 144.175 64.290 145.085 ;
        RECT 64.505 144.215 64.935 145.000 ;
        RECT 65.875 144.275 71.385 145.085 ;
        RECT 71.395 144.275 76.905 145.085 ;
        RECT 77.110 144.175 80.585 145.085 ;
        RECT 80.965 144.405 90.245 145.085 ;
        RECT 80.965 144.285 83.300 144.405 ;
        RECT 80.965 144.175 81.885 144.285 ;
        RECT 87.965 144.185 88.885 144.405 ;
        RECT 90.265 144.215 90.695 145.000 ;
        RECT 90.715 144.305 92.085 145.085 ;
        RECT 92.095 144.275 93.925 145.085 ;
        RECT 93.935 144.275 99.445 145.085 ;
        RECT 99.455 144.275 104.965 145.085 ;
        RECT 105.120 145.055 105.290 145.275 ;
        RECT 106.030 145.105 106.200 145.325 ;
        RECT 106.355 145.295 109.830 146.205 ;
        RECT 110.035 145.295 113.510 146.205 ;
        RECT 114.175 145.295 116.925 146.105 ;
        RECT 116.935 145.295 122.445 146.105 ;
        RECT 122.455 145.295 127.965 146.105 ;
        RECT 127.975 145.295 129.345 146.105 ;
        RECT 106.500 145.105 106.670 145.295 ;
        RECT 108.795 145.085 108.965 145.275 ;
        RECT 110.180 145.105 110.350 145.295 ;
        RECT 112.470 145.085 112.640 145.275 ;
        RECT 106.780 145.055 107.725 145.085 ;
        RECT 104.975 144.375 107.725 145.055 ;
        RECT 106.780 144.175 107.725 144.375 ;
        RECT 107.735 144.275 109.105 145.085 ;
        RECT 109.310 144.175 112.785 145.085 ;
        RECT 112.940 145.055 113.110 145.275 ;
        RECT 116.615 145.245 116.785 145.295 ;
        RECT 113.910 145.135 114.030 145.245 ;
        RECT 115.750 145.135 115.870 145.245 ;
        RECT 116.615 145.135 116.790 145.245 ;
        RECT 116.615 145.105 116.785 145.135 ;
        RECT 122.135 145.085 122.305 145.295 ;
        RECT 127.655 145.085 127.825 145.295 ;
        RECT 129.035 145.085 129.205 145.295 ;
        RECT 114.600 145.055 115.545 145.085 ;
        RECT 112.795 144.375 115.545 145.055 ;
        RECT 114.600 144.175 115.545 144.375 ;
        RECT 116.025 144.215 116.455 145.000 ;
        RECT 116.935 144.275 122.445 145.085 ;
        RECT 122.455 144.275 127.965 145.085 ;
        RECT 127.975 144.275 129.345 145.085 ;
      LAYER nwell ;
        RECT 9.100 141.055 129.540 143.885 ;
      LAYER pwell ;
        RECT 9.295 139.855 10.665 140.665 ;
        RECT 10.675 139.855 14.345 140.665 ;
        RECT 15.715 140.535 16.635 140.755 ;
        RECT 22.715 140.655 23.635 140.765 ;
        RECT 21.300 140.535 23.635 140.655 ;
        RECT 14.355 139.855 23.635 140.535 ;
        RECT 24.015 139.855 25.845 140.665 ;
        RECT 25.865 139.940 26.295 140.725 ;
        RECT 26.775 139.855 32.285 140.665 ;
        RECT 32.295 139.855 35.770 140.765 ;
        RECT 35.975 139.855 37.345 140.665 ;
        RECT 37.355 139.855 41.025 140.665 ;
        RECT 41.035 139.855 46.545 140.665 ;
        RECT 46.555 139.855 50.030 140.765 ;
        RECT 50.235 139.855 51.605 140.665 ;
        RECT 51.625 139.940 52.055 140.725 ;
        RECT 52.535 139.855 53.905 140.635 ;
        RECT 53.915 139.855 55.745 140.665 ;
        RECT 55.755 139.855 58.965 140.765 ;
        RECT 60.335 140.535 61.255 140.755 ;
        RECT 67.335 140.655 68.255 140.765 ;
        RECT 65.920 140.535 68.255 140.655 ;
        RECT 58.975 139.855 68.255 140.535 ;
        RECT 68.635 139.855 72.110 140.765 ;
        RECT 72.325 139.855 73.675 140.765 ;
        RECT 73.695 139.855 77.365 140.665 ;
        RECT 77.385 139.940 77.815 140.725 ;
        RECT 77.835 140.565 78.780 140.765 ;
        RECT 77.835 139.885 80.585 140.565 ;
        RECT 77.835 139.855 78.780 139.885 ;
        RECT 9.435 139.645 9.605 139.855 ;
        RECT 10.870 139.695 10.990 139.805 ;
        RECT 12.655 139.645 12.825 139.835 ;
        RECT 13.630 139.695 13.750 139.805 ;
        RECT 14.035 139.665 14.205 139.855 ;
        RECT 14.495 139.665 14.665 139.855 ;
        RECT 17.255 139.645 17.425 139.835 ;
        RECT 17.715 139.645 17.885 139.835 ;
        RECT 21.395 139.645 21.565 139.835 ;
        RECT 25.535 139.665 25.705 139.855 ;
        RECT 26.510 139.695 26.630 139.805 ;
        RECT 26.915 139.645 27.085 139.835 ;
        RECT 9.295 138.835 10.665 139.645 ;
        RECT 11.135 138.835 12.965 139.645 ;
        RECT 12.985 138.775 13.415 139.560 ;
        RECT 13.895 138.835 17.565 139.645 ;
        RECT 17.585 138.735 18.935 139.645 ;
        RECT 18.955 138.835 21.705 139.645 ;
        RECT 21.715 138.835 27.225 139.645 ;
        RECT 27.235 139.615 28.180 139.645 ;
        RECT 29.670 139.615 29.840 139.835 ;
        RECT 31.975 139.665 32.145 139.855 ;
        RECT 32.440 139.835 32.610 139.855 ;
        RECT 32.430 139.665 32.610 139.835 ;
        RECT 29.995 139.615 30.940 139.645 ;
        RECT 32.430 139.615 32.600 139.665 ;
        RECT 32.755 139.615 33.700 139.645 ;
        RECT 35.190 139.615 35.360 139.835 ;
        RECT 35.710 139.695 35.830 139.805 ;
        RECT 37.035 139.665 37.205 139.855 ;
        RECT 38.415 139.645 38.585 139.835 ;
        RECT 39.390 139.695 39.510 139.805 ;
        RECT 40.715 139.665 40.885 139.855 ;
        RECT 42.095 139.645 42.265 139.835 ;
        RECT 46.235 139.665 46.405 139.855 ;
        RECT 46.700 139.665 46.870 139.855 ;
        RECT 47.615 139.645 47.785 139.835 ;
        RECT 48.350 139.645 48.520 139.835 ;
        RECT 51.295 139.665 51.465 139.855 ;
        RECT 52.270 139.695 52.390 139.805 ;
        RECT 52.675 139.665 52.845 139.855 ;
        RECT 54.975 139.645 55.145 139.835 ;
        RECT 55.435 139.665 55.605 139.855 ;
        RECT 55.895 139.665 56.065 139.855 ;
        RECT 59.115 139.665 59.285 139.855 ;
        RECT 60.495 139.645 60.665 139.835 ;
        RECT 60.960 139.645 61.130 139.835 ;
        RECT 65.150 139.695 65.270 139.805 ;
        RECT 67.855 139.645 68.025 139.835 ;
        RECT 68.780 139.665 68.950 139.855 ;
        RECT 73.375 139.665 73.545 139.855 ;
        RECT 77.055 139.665 77.225 139.855 ;
        RECT 77.515 139.645 77.685 139.835 ;
        RECT 78.895 139.645 79.065 139.835 ;
        RECT 79.360 139.645 79.530 139.835 ;
        RECT 80.270 139.665 80.440 139.885 ;
        RECT 81.055 139.855 86.565 140.665 ;
        RECT 86.575 139.855 92.085 140.665 ;
        RECT 92.095 139.855 97.605 140.665 ;
        RECT 97.615 139.855 103.125 140.665 ;
        RECT 103.145 139.940 103.575 140.725 ;
        RECT 103.595 139.855 104.965 140.665 ;
        RECT 104.975 139.855 108.645 140.665 ;
        RECT 108.655 139.855 112.130 140.765 ;
        RECT 112.795 139.855 116.465 140.665 ;
        RECT 116.485 139.855 117.835 140.765 ;
        RECT 121.055 140.535 121.985 140.765 ;
        RECT 118.085 139.855 121.985 140.535 ;
        RECT 122.915 139.855 124.285 140.635 ;
        RECT 124.295 139.855 127.965 140.665 ;
        RECT 127.975 139.855 129.345 140.665 ;
        RECT 80.790 139.695 80.910 139.805 ;
        RECT 83.090 139.695 83.210 139.805 ;
        RECT 86.255 139.665 86.425 139.855 ;
        RECT 88.555 139.645 88.725 139.835 ;
        RECT 89.935 139.645 90.105 139.835 ;
        RECT 90.910 139.695 91.030 139.805 ;
        RECT 91.775 139.665 91.945 139.855 ;
        RECT 96.375 139.645 96.545 139.835 ;
        RECT 97.295 139.665 97.465 139.855 ;
        RECT 27.235 138.935 29.985 139.615 ;
        RECT 29.995 138.935 32.745 139.615 ;
        RECT 32.755 138.935 35.505 139.615 ;
        RECT 27.235 138.735 28.180 138.935 ;
        RECT 29.995 138.735 30.940 138.935 ;
        RECT 32.755 138.735 33.700 138.935 ;
        RECT 35.975 138.835 38.725 139.645 ;
        RECT 38.745 138.775 39.175 139.560 ;
        RECT 39.655 138.835 42.405 139.645 ;
        RECT 42.415 138.835 47.925 139.645 ;
        RECT 47.935 138.965 51.835 139.645 ;
        RECT 47.935 138.735 48.865 138.965 ;
        RECT 52.535 138.835 55.285 139.645 ;
        RECT 55.295 138.835 60.805 139.645 ;
        RECT 60.815 138.735 64.290 139.645 ;
        RECT 64.505 138.775 64.935 139.560 ;
        RECT 65.415 138.835 68.165 139.645 ;
        RECT 68.545 138.965 77.825 139.645 ;
        RECT 68.545 138.845 70.880 138.965 ;
        RECT 68.545 138.735 69.465 138.845 ;
        RECT 75.545 138.745 76.465 138.965 ;
        RECT 77.835 138.835 79.205 139.645 ;
        RECT 79.215 138.735 82.690 139.645 ;
        RECT 83.355 138.835 88.865 139.645 ;
        RECT 88.885 138.735 90.235 139.645 ;
        RECT 90.265 138.775 90.695 139.560 ;
        RECT 91.175 138.835 96.685 139.645 ;
        RECT 96.695 139.615 97.640 139.645 ;
        RECT 99.130 139.615 99.300 139.835 ;
        RECT 99.600 139.645 99.770 139.835 ;
        RECT 102.815 139.665 102.985 139.855 ;
        RECT 103.330 139.695 103.450 139.805 ;
        RECT 104.655 139.665 104.825 139.855 ;
        RECT 96.695 138.935 99.445 139.615 ;
        RECT 96.695 138.735 97.640 138.935 ;
        RECT 99.455 138.735 102.930 139.645 ;
        RECT 103.595 139.615 104.540 139.645 ;
        RECT 106.030 139.615 106.200 139.835 ;
        RECT 106.500 139.645 106.670 139.835 ;
        RECT 108.335 139.665 108.505 139.855 ;
        RECT 108.800 139.665 108.970 139.855 ;
        RECT 111.555 139.645 111.725 139.835 ;
        RECT 112.530 139.695 112.650 139.805 ;
        RECT 115.420 139.645 115.590 139.835 ;
        RECT 116.155 139.665 116.325 139.855 ;
        RECT 116.615 139.645 116.785 139.855 ;
        RECT 121.400 139.665 121.570 139.855 ;
        RECT 122.595 139.700 122.755 139.810 ;
        RECT 123.055 139.665 123.225 139.855 ;
        RECT 127.195 139.645 127.365 139.835 ;
        RECT 127.655 139.805 127.825 139.855 ;
        RECT 127.655 139.695 127.830 139.805 ;
        RECT 127.655 139.665 127.825 139.695 ;
        RECT 129.035 139.645 129.205 139.855 ;
        RECT 103.595 138.935 106.345 139.615 ;
        RECT 103.595 138.735 104.540 138.935 ;
        RECT 106.355 138.735 109.830 139.645 ;
        RECT 110.035 138.835 111.865 139.645 ;
        RECT 112.105 138.965 116.005 139.645 ;
        RECT 115.075 138.735 116.005 138.965 ;
        RECT 116.025 138.775 116.455 139.560 ;
        RECT 116.485 138.735 117.835 139.645 ;
        RECT 118.225 138.965 127.505 139.645 ;
        RECT 118.225 138.845 120.560 138.965 ;
        RECT 118.225 138.735 119.145 138.845 ;
        RECT 125.225 138.745 126.145 138.965 ;
        RECT 127.975 138.835 129.345 139.645 ;
      LAYER nwell ;
        RECT 9.100 135.615 129.540 138.445 ;
      LAYER pwell ;
        RECT 9.295 134.415 10.665 135.225 ;
        RECT 11.135 134.415 14.805 135.225 ;
        RECT 14.815 134.415 20.325 135.225 ;
        RECT 20.335 134.415 25.845 135.225 ;
        RECT 25.865 134.500 26.295 135.285 ;
        RECT 26.775 134.415 28.605 135.225 ;
        RECT 28.615 134.415 34.125 135.225 ;
        RECT 34.135 134.415 39.645 135.225 ;
        RECT 39.665 134.415 41.015 135.325 ;
        RECT 41.405 135.215 42.325 135.325 ;
        RECT 41.405 135.095 43.740 135.215 ;
        RECT 48.405 135.095 49.325 135.315 ;
        RECT 41.405 134.415 50.685 135.095 ;
        RECT 51.625 134.500 52.055 135.285 ;
        RECT 52.995 134.415 58.505 135.225 ;
        RECT 58.515 134.415 64.025 135.225 ;
        RECT 64.035 134.415 67.510 135.325 ;
        RECT 70.915 135.095 71.845 135.325 ;
        RECT 67.945 134.415 71.845 135.095 ;
        RECT 71.855 134.415 73.225 135.225 ;
        RECT 73.235 134.415 74.605 135.195 ;
        RECT 74.615 134.415 77.365 135.225 ;
        RECT 77.385 134.500 77.815 135.285 ;
        RECT 78.755 134.415 84.265 135.225 ;
        RECT 84.645 135.215 85.565 135.325 ;
        RECT 84.645 135.095 86.980 135.215 ;
        RECT 91.645 135.095 92.565 135.315 ;
        RECT 84.645 134.415 93.925 135.095 ;
        RECT 93.935 134.415 97.605 135.225 ;
        RECT 97.615 134.415 103.125 135.225 ;
        RECT 103.145 134.500 103.575 135.285 ;
        RECT 104.055 134.415 106.805 135.225 ;
        RECT 106.815 135.125 107.760 135.325 ;
        RECT 106.815 134.445 109.565 135.125 ;
        RECT 106.815 134.415 107.760 134.445 ;
        RECT 9.435 134.205 9.605 134.415 ;
        RECT 10.870 134.255 10.990 134.365 ;
        RECT 12.655 134.205 12.825 134.395 ;
        RECT 14.495 134.225 14.665 134.415 ;
        RECT 15.875 134.205 16.045 134.395 ;
        RECT 19.740 134.205 19.910 134.395 ;
        RECT 20.015 134.225 20.185 134.415 ;
        RECT 25.535 134.205 25.705 134.415 ;
        RECT 25.995 134.225 26.165 134.395 ;
        RECT 26.510 134.255 26.630 134.365 ;
        RECT 28.295 134.225 28.465 134.415 ;
        RECT 30.595 134.225 30.765 134.395 ;
        RECT 32.950 134.255 33.070 134.365 ;
        RECT 33.815 134.225 33.985 134.415 ;
        RECT 26.015 134.205 26.165 134.225 ;
        RECT 28.315 134.205 28.465 134.225 ;
        RECT 30.615 134.205 30.765 134.225 ;
        RECT 38.415 134.205 38.585 134.395 ;
        RECT 39.335 134.225 39.505 134.415 ;
        RECT 39.795 134.225 39.965 134.415 ;
        RECT 40.715 134.205 40.885 134.395 ;
        RECT 9.295 133.395 10.665 134.205 ;
        RECT 11.135 133.395 12.965 134.205 ;
        RECT 12.985 133.335 13.415 134.120 ;
        RECT 13.435 133.395 16.185 134.205 ;
        RECT 16.425 133.525 20.325 134.205 ;
        RECT 19.395 133.295 20.325 133.525 ;
        RECT 20.335 133.395 25.845 134.205 ;
        RECT 26.015 133.385 27.945 134.205 ;
        RECT 28.315 133.385 30.245 134.205 ;
        RECT 30.615 133.385 32.545 134.205 ;
        RECT 33.215 133.395 38.725 134.205 ;
        RECT 26.995 133.295 27.945 133.385 ;
        RECT 29.295 133.295 30.245 133.385 ;
        RECT 31.595 133.295 32.545 133.385 ;
        RECT 38.745 133.335 39.175 134.120 ;
        RECT 39.195 133.395 41.025 134.205 ;
        RECT 41.035 134.175 41.980 134.205 ;
        RECT 43.470 134.175 43.640 134.395 ;
        RECT 45.315 134.205 45.485 134.395 ;
        RECT 45.780 134.205 45.950 134.395 ;
        RECT 50.375 134.205 50.545 134.415 ;
        RECT 51.295 134.250 51.455 134.370 ;
        RECT 52.675 134.260 52.835 134.370 ;
        RECT 54.975 134.205 55.145 134.395 ;
        RECT 55.435 134.205 55.605 134.395 ;
        RECT 56.815 134.205 56.985 134.395 ;
        RECT 58.195 134.225 58.365 134.415 ;
        RECT 58.655 134.250 58.815 134.360 ;
        RECT 63.715 134.225 63.885 134.415 ;
        RECT 64.180 134.395 64.350 134.415 ;
        RECT 64.175 134.225 64.350 134.395 ;
        RECT 65.150 134.255 65.270 134.365 ;
        RECT 64.175 134.205 64.345 134.225 ;
        RECT 68.775 134.205 68.945 134.395 ;
        RECT 71.260 134.225 71.430 134.415 ;
        RECT 72.915 134.225 73.085 134.415 ;
        RECT 73.375 134.225 73.545 134.415 ;
        RECT 74.295 134.205 74.465 134.395 ;
        RECT 77.055 134.225 77.225 134.415 ;
        RECT 78.435 134.260 78.595 134.370 ;
        RECT 79.815 134.205 79.985 134.395 ;
        RECT 80.280 134.205 80.450 134.395 ;
        RECT 83.955 134.365 84.125 134.415 ;
        RECT 83.955 134.255 84.130 134.365 ;
        RECT 83.955 134.225 84.125 134.255 ;
        RECT 87.820 134.205 87.990 134.395 ;
        RECT 88.610 134.255 88.730 134.365 ;
        RECT 89.015 134.205 89.185 134.395 ;
        RECT 93.615 134.225 93.785 134.415 ;
        RECT 95.915 134.205 96.085 134.395 ;
        RECT 96.375 134.205 96.545 134.395 ;
        RECT 97.295 134.225 97.465 134.415 ;
        RECT 101.160 134.205 101.330 134.395 ;
        RECT 102.355 134.250 102.515 134.360 ;
        RECT 102.815 134.225 102.985 134.415 ;
        RECT 103.790 134.255 103.910 134.365 ;
        RECT 106.495 134.225 106.665 134.415 ;
        RECT 107.875 134.205 108.045 134.395 ;
        RECT 109.250 134.225 109.420 134.445 ;
        RECT 109.575 134.415 111.405 135.225 ;
        RECT 111.415 134.415 116.925 135.225 ;
        RECT 117.305 135.215 118.225 135.325 ;
        RECT 117.305 135.095 119.640 135.215 ;
        RECT 124.305 135.095 125.225 135.315 ;
        RECT 117.305 134.415 126.585 135.095 ;
        RECT 126.595 134.415 127.965 135.225 ;
        RECT 127.975 134.415 129.345 135.225 ;
        RECT 111.095 134.225 111.265 134.415 ;
        RECT 111.740 134.205 111.910 134.395 ;
        RECT 112.475 134.205 112.645 134.395 ;
        RECT 113.910 134.255 114.030 134.365 ;
        RECT 115.695 134.205 115.865 134.395 ;
        RECT 116.615 134.365 116.785 134.415 ;
        RECT 116.615 134.255 116.790 134.365 ;
        RECT 116.615 134.225 116.785 134.255 ;
        RECT 122.135 134.205 122.305 134.395 ;
        RECT 122.595 134.205 122.765 134.395 ;
        RECT 124.030 134.255 124.150 134.365 ;
        RECT 126.275 134.225 126.445 134.415 ;
        RECT 127.655 134.205 127.825 134.415 ;
        RECT 129.035 134.205 129.205 134.415 ;
        RECT 41.035 133.495 43.785 134.175 ;
        RECT 41.035 133.295 41.980 133.495 ;
        RECT 43.795 133.395 45.625 134.205 ;
        RECT 45.635 133.295 49.110 134.205 ;
        RECT 49.315 133.425 50.685 134.205 ;
        RECT 51.615 133.395 55.285 134.205 ;
        RECT 55.305 133.295 56.655 134.205 ;
        RECT 56.675 133.425 58.045 134.205 ;
        RECT 58.975 133.395 64.485 134.205 ;
        RECT 64.505 133.335 64.935 134.120 ;
        RECT 65.415 133.395 69.085 134.205 ;
        RECT 69.095 133.395 74.605 134.205 ;
        RECT 74.615 133.395 80.125 134.205 ;
        RECT 80.135 133.295 83.610 134.205 ;
        RECT 84.505 133.525 88.405 134.205 ;
        RECT 87.475 133.295 88.405 133.525 ;
        RECT 88.875 133.425 90.245 134.205 ;
        RECT 90.265 133.335 90.695 134.120 ;
        RECT 90.715 133.395 96.225 134.205 ;
        RECT 96.245 133.295 97.595 134.205 ;
        RECT 97.845 133.525 101.745 134.205 ;
        RECT 100.815 133.295 101.745 133.525 ;
        RECT 102.675 133.395 108.185 134.205 ;
        RECT 108.425 133.525 112.325 134.205 ;
        RECT 111.395 133.295 112.325 133.525 ;
        RECT 112.335 133.425 113.705 134.205 ;
        RECT 114.175 133.395 116.005 134.205 ;
        RECT 116.025 133.335 116.455 134.120 ;
        RECT 116.935 133.395 122.445 134.205 ;
        RECT 122.455 133.425 123.825 134.205 ;
        RECT 124.295 133.395 127.965 134.205 ;
        RECT 127.975 133.395 129.345 134.205 ;
      LAYER nwell ;
        RECT 9.100 130.175 129.540 133.005 ;
      LAYER pwell ;
        RECT 9.295 128.975 10.665 129.785 ;
        RECT 11.965 129.775 12.885 129.885 ;
        RECT 11.965 129.655 14.300 129.775 ;
        RECT 18.965 129.655 19.885 129.875 ;
        RECT 11.965 128.975 21.245 129.655 ;
        RECT 21.255 128.975 22.625 129.755 ;
        RECT 23.095 128.975 24.465 129.755 ;
        RECT 24.475 128.975 25.845 129.785 ;
        RECT 25.865 129.060 26.295 129.845 ;
        RECT 33.435 129.795 34.385 129.885 ;
        RECT 27.235 128.975 30.905 129.785 ;
        RECT 30.915 128.975 32.285 129.755 ;
        RECT 32.455 128.975 34.385 129.795 ;
        RECT 34.595 128.975 36.425 129.785 ;
        RECT 36.435 129.685 37.380 129.885 ;
        RECT 39.195 129.685 40.140 129.885 ;
        RECT 36.435 129.005 39.185 129.685 ;
        RECT 39.195 129.005 41.945 129.685 ;
        RECT 36.435 128.975 37.380 129.005 ;
        RECT 9.435 128.765 9.605 128.975 ;
        RECT 11.275 128.810 11.435 128.930 ;
        RECT 12.655 128.765 12.825 128.955 ;
        RECT 20.935 128.785 21.105 128.975 ;
        RECT 22.315 128.785 22.485 128.975 ;
        RECT 22.775 128.925 22.945 128.955 ;
        RECT 22.775 128.815 22.950 128.925 ;
        RECT 22.775 128.765 22.945 128.815 ;
        RECT 24.155 128.785 24.325 128.975 ;
        RECT 25.535 128.785 25.705 128.975 ;
        RECT 26.640 128.765 26.810 128.955 ;
        RECT 26.915 128.820 27.075 128.930 ;
        RECT 30.595 128.785 30.765 128.975 ;
        RECT 31.055 128.785 31.225 128.975 ;
        RECT 32.455 128.955 32.605 128.975 ;
        RECT 32.435 128.785 32.605 128.955 ;
        RECT 36.115 128.765 36.285 128.975 ;
        RECT 36.630 128.815 36.750 128.925 ;
        RECT 38.415 128.765 38.585 128.955 ;
        RECT 38.870 128.785 39.040 129.005 ;
        RECT 39.195 128.975 40.140 129.005 ;
        RECT 39.795 128.810 39.955 128.920 ;
        RECT 41.630 128.785 41.800 129.005 ;
        RECT 41.955 128.975 43.785 129.785 ;
        RECT 43.795 128.975 47.270 129.885 ;
        RECT 50.675 129.655 51.605 129.885 ;
        RECT 47.705 128.975 51.605 129.655 ;
        RECT 51.625 129.060 52.055 129.845 ;
        RECT 52.445 129.775 53.365 129.885 ;
        RECT 52.445 129.655 54.780 129.775 ;
        RECT 59.445 129.655 60.365 129.875 ;
        RECT 52.445 128.975 61.725 129.655 ;
        RECT 62.195 128.975 65.865 129.785 ;
        RECT 69.075 129.655 70.005 129.885 ;
        RECT 66.105 128.975 70.005 129.655 ;
        RECT 70.475 128.975 71.845 129.755 ;
        RECT 71.855 128.975 74.605 129.785 ;
        RECT 74.615 129.685 75.560 129.885 ;
        RECT 74.615 129.005 77.365 129.685 ;
        RECT 77.385 129.060 77.815 129.845 ;
        RECT 74.615 128.975 75.560 129.005 ;
        RECT 43.475 128.785 43.645 128.975 ;
        RECT 43.940 128.785 44.110 128.975 ;
        RECT 45.315 128.765 45.485 128.955 ;
        RECT 47.615 128.785 47.785 128.955 ;
        RECT 47.615 128.765 47.765 128.785 ;
        RECT 48.080 128.765 48.250 128.955 ;
        RECT 51.020 128.785 51.190 128.975 ;
        RECT 51.810 128.815 51.930 128.925 ;
        RECT 53.595 128.765 53.765 128.955 ;
        RECT 57.460 128.765 57.630 128.955 ;
        RECT 59.115 128.765 59.285 128.955 ;
        RECT 61.415 128.785 61.585 128.975 ;
        RECT 61.930 128.815 62.050 128.925 ;
        RECT 62.795 128.765 62.965 128.955 ;
        RECT 63.255 128.765 63.425 128.955 ;
        RECT 65.150 128.815 65.270 128.925 ;
        RECT 65.555 128.785 65.725 128.975 ;
        RECT 69.420 128.785 69.590 128.975 ;
        RECT 70.210 128.815 70.330 128.925 ;
        RECT 70.615 128.785 70.785 128.975 ;
        RECT 74.295 128.785 74.465 128.975 ;
        RECT 74.755 128.765 74.925 128.955 ;
        RECT 77.050 128.785 77.220 129.005 ;
        RECT 77.835 128.975 79.665 129.785 ;
        RECT 79.675 128.975 83.150 129.885 ;
        RECT 83.355 128.975 85.185 129.785 ;
        RECT 88.395 129.655 89.325 129.885 ;
        RECT 85.425 128.975 89.325 129.655 ;
        RECT 89.335 128.975 90.705 129.755 ;
        RECT 90.715 128.975 93.465 129.785 ;
        RECT 93.845 129.775 94.765 129.885 ;
        RECT 93.845 129.655 96.180 129.775 ;
        RECT 100.845 129.655 101.765 129.875 ;
        RECT 93.845 128.975 103.125 129.655 ;
        RECT 103.145 129.060 103.575 129.845 ;
        RECT 104.055 128.975 105.885 129.785 ;
        RECT 106.265 129.775 107.185 129.885 ;
        RECT 106.265 129.655 108.600 129.775 ;
        RECT 113.265 129.655 114.185 129.875 ;
        RECT 106.265 128.975 115.545 129.655 ;
        RECT 115.555 128.975 116.925 129.785 ;
        RECT 116.935 128.975 122.445 129.785 ;
        RECT 122.455 128.975 127.965 129.785 ;
        RECT 127.975 128.975 129.345 129.785 ;
        RECT 77.515 128.765 77.685 128.955 ;
        RECT 79.355 128.785 79.525 128.975 ;
        RECT 79.820 128.785 79.990 128.975 ;
        RECT 9.295 127.955 10.665 128.765 ;
        RECT 11.605 127.855 12.955 128.765 ;
        RECT 12.985 127.895 13.415 128.680 ;
        RECT 13.805 128.085 23.085 128.765 ;
        RECT 23.325 128.085 27.225 128.765 ;
        RECT 27.320 128.085 36.425 128.765 ;
        RECT 13.805 127.965 16.140 128.085 ;
        RECT 13.805 127.855 14.725 127.965 ;
        RECT 20.805 127.865 21.725 128.085 ;
        RECT 26.295 127.855 27.225 128.085 ;
        RECT 36.895 127.955 38.725 128.765 ;
        RECT 38.745 127.895 39.175 128.680 ;
        RECT 40.115 127.955 45.625 128.765 ;
        RECT 45.835 127.945 47.765 128.765 ;
        RECT 45.835 127.855 46.785 127.945 ;
        RECT 47.935 127.855 51.410 128.765 ;
        RECT 52.075 127.955 53.905 128.765 ;
        RECT 54.145 128.085 58.045 128.765 ;
        RECT 57.115 127.855 58.045 128.085 ;
        RECT 58.055 127.955 59.425 128.765 ;
        RECT 59.435 127.955 63.105 128.765 ;
        RECT 63.125 127.855 64.475 128.765 ;
        RECT 64.505 127.895 64.935 128.680 ;
        RECT 65.785 128.085 75.065 128.765 ;
        RECT 65.785 127.965 68.120 128.085 ;
        RECT 65.785 127.855 66.705 127.965 ;
        RECT 72.785 127.865 73.705 128.085 ;
        RECT 75.075 127.955 77.825 128.765 ;
        RECT 77.835 128.735 78.780 128.765 ;
        RECT 80.270 128.735 80.440 128.955 ;
        RECT 84.875 128.785 85.045 128.975 ;
        RECT 88.740 128.785 88.910 128.975 ;
        RECT 89.935 128.765 90.105 128.955 ;
        RECT 90.395 128.785 90.565 128.975 ;
        RECT 91.775 128.765 91.945 128.955 ;
        RECT 93.155 128.765 93.325 128.975 ;
        RECT 96.835 128.765 97.005 128.955 ;
        RECT 97.295 128.785 97.465 128.955 ;
        RECT 100.055 128.810 100.215 128.920 ;
        RECT 97.315 128.765 97.465 128.785 ;
        RECT 101.435 128.765 101.605 128.955 ;
        RECT 101.950 128.815 102.070 128.925 ;
        RECT 102.815 128.785 102.985 128.975 ;
        RECT 103.735 128.925 103.905 128.955 ;
        RECT 103.735 128.815 103.910 128.925 ;
        RECT 103.735 128.765 103.905 128.815 ;
        RECT 104.195 128.785 104.365 128.955 ;
        RECT 105.575 128.785 105.745 128.975 ;
        RECT 106.955 128.810 107.115 128.920 ;
        RECT 104.215 128.765 104.365 128.785 ;
        RECT 107.415 128.765 107.585 128.955 ;
        RECT 110.635 128.785 110.805 128.955 ;
        RECT 111.555 128.810 111.715 128.920 ;
        RECT 112.015 128.785 112.185 128.955 ;
        RECT 115.235 128.785 115.405 128.975 ;
        RECT 110.635 128.765 110.785 128.785 ;
        RECT 77.835 128.055 80.585 128.735 ;
        RECT 80.965 128.085 90.245 128.765 ;
        RECT 77.835 127.855 78.780 128.055 ;
        RECT 80.965 127.965 83.300 128.085 ;
        RECT 80.965 127.855 81.885 127.965 ;
        RECT 87.965 127.865 88.885 128.085 ;
        RECT 90.265 127.895 90.695 128.680 ;
        RECT 90.725 127.855 92.075 128.765 ;
        RECT 92.095 127.955 93.465 128.765 ;
        RECT 93.475 127.955 97.145 128.765 ;
        RECT 97.315 127.945 99.245 128.765 ;
        RECT 100.375 127.985 101.745 128.765 ;
        RECT 102.215 127.955 104.045 128.765 ;
        RECT 104.215 127.945 106.145 128.765 ;
        RECT 98.295 127.855 99.245 127.945 ;
        RECT 105.195 127.855 106.145 127.945 ;
        RECT 107.285 127.855 108.635 128.765 ;
        RECT 108.855 127.945 110.785 128.765 ;
        RECT 112.035 128.765 112.185 128.785 ;
        RECT 115.695 128.765 115.865 128.955 ;
        RECT 116.615 128.925 116.785 128.975 ;
        RECT 116.615 128.815 116.790 128.925 ;
        RECT 116.615 128.785 116.785 128.815 ;
        RECT 122.135 128.765 122.305 128.975 ;
        RECT 127.655 128.765 127.825 128.975 ;
        RECT 129.035 128.765 129.205 128.975 ;
        RECT 112.035 127.945 113.965 128.765 ;
        RECT 114.175 127.955 116.005 128.765 ;
        RECT 108.855 127.855 109.805 127.945 ;
        RECT 113.015 127.855 113.965 127.945 ;
        RECT 116.025 127.895 116.455 128.680 ;
        RECT 116.935 127.955 122.445 128.765 ;
        RECT 122.455 127.955 127.965 128.765 ;
        RECT 127.975 127.955 129.345 128.765 ;
      LAYER nwell ;
        RECT 9.100 124.735 129.540 127.565 ;
      LAYER pwell ;
        RECT 9.295 123.535 10.665 124.345 ;
        RECT 11.595 123.535 15.265 124.345 ;
        RECT 15.285 123.535 16.635 124.445 ;
        RECT 19.855 124.215 20.785 124.445 ;
        RECT 16.885 123.535 20.785 124.215 ;
        RECT 20.795 123.535 24.465 124.345 ;
        RECT 24.485 123.535 25.835 124.445 ;
        RECT 25.865 123.620 26.295 124.405 ;
        RECT 26.685 124.335 27.605 124.445 ;
        RECT 26.685 124.215 29.020 124.335 ;
        RECT 33.685 124.215 34.605 124.435 ;
        RECT 26.685 123.535 35.965 124.215 ;
        RECT 35.975 123.535 37.340 124.215 ;
        RECT 38.745 123.535 40.095 124.445 ;
        RECT 41.035 123.535 50.140 124.215 ;
        RECT 50.235 123.535 51.605 124.345 ;
        RECT 51.625 123.620 52.055 124.405 ;
        RECT 52.535 123.535 58.045 124.345 ;
        RECT 58.055 123.535 59.425 124.315 ;
        RECT 62.635 124.215 63.565 124.445 ;
        RECT 68.375 124.355 69.325 124.445 ;
        RECT 59.665 123.535 63.565 124.215 ;
        RECT 64.495 123.535 66.325 124.215 ;
        RECT 66.335 123.535 68.165 124.215 ;
        RECT 68.375 123.535 70.305 124.355 ;
        RECT 70.475 123.535 71.845 124.345 ;
        RECT 71.855 123.535 77.365 124.345 ;
        RECT 77.385 123.620 77.815 124.405 ;
        RECT 77.835 123.535 80.585 124.345 ;
        RECT 80.595 123.535 89.700 124.215 ;
        RECT 90.255 123.535 93.925 124.345 ;
        RECT 93.935 123.535 103.040 124.215 ;
        RECT 103.145 123.620 103.575 124.405 ;
        RECT 107.015 124.355 107.965 124.445 ;
        RECT 111.155 124.355 112.105 124.445 ;
        RECT 104.055 123.535 106.805 124.345 ;
        RECT 107.015 123.535 108.945 124.355 ;
        RECT 109.115 123.535 110.945 124.345 ;
        RECT 111.155 123.535 113.085 124.355 ;
        RECT 113.255 123.535 116.005 124.345 ;
        RECT 116.025 123.535 117.375 124.445 ;
        RECT 117.765 124.335 118.685 124.445 ;
        RECT 117.765 124.215 120.100 124.335 ;
        RECT 124.765 124.215 125.685 124.435 ;
        RECT 117.765 123.535 127.045 124.215 ;
        RECT 127.975 123.535 129.345 124.345 ;
        RECT 9.435 123.325 9.605 123.535 ;
        RECT 10.870 123.375 10.990 123.485 ;
        RECT 11.275 123.380 11.435 123.490 ;
        RECT 12.655 123.325 12.825 123.515 ;
        RECT 14.955 123.345 15.125 123.535 ;
        RECT 15.415 123.345 15.585 123.535 ;
        RECT 18.635 123.325 18.805 123.515 ;
        RECT 20.200 123.345 20.370 123.535 ;
        RECT 24.155 123.325 24.325 123.535 ;
        RECT 24.615 123.345 24.785 123.535 ;
        RECT 29.675 123.325 29.845 123.515 ;
        RECT 30.135 123.345 30.305 123.515 ;
        RECT 32.435 123.345 32.605 123.515 ;
        RECT 35.655 123.345 35.825 123.535 ;
        RECT 37.495 123.345 37.665 123.515 ;
        RECT 30.155 123.325 30.305 123.345 ;
        RECT 32.455 123.325 32.605 123.345 ;
        RECT 38.140 123.325 38.310 123.515 ;
        RECT 38.415 123.380 38.575 123.490 ;
        RECT 38.875 123.345 39.045 123.535 ;
        RECT 39.390 123.375 39.510 123.485 ;
        RECT 39.795 123.345 39.965 123.515 ;
        RECT 40.715 123.380 40.875 123.490 ;
        RECT 41.175 123.345 41.345 123.535 ;
        RECT 39.815 123.325 39.965 123.345 ;
        RECT 42.095 123.325 42.265 123.515 ;
        RECT 46.695 123.325 46.865 123.515 ;
        RECT 49.915 123.345 50.085 123.515 ;
        RECT 51.295 123.345 51.465 123.535 ;
        RECT 52.270 123.375 52.390 123.485 ;
        RECT 53.595 123.325 53.765 123.515 ;
        RECT 57.735 123.345 57.905 123.535 ;
        RECT 58.195 123.345 58.365 123.535 ;
        RECT 62.980 123.345 63.150 123.535 ;
        RECT 63.255 123.325 63.425 123.515 ;
        RECT 64.175 123.370 64.335 123.490 ;
        RECT 66.015 123.345 66.185 123.535 ;
        RECT 66.475 123.345 66.645 123.535 ;
        RECT 70.155 123.515 70.305 123.535 ;
        RECT 67.395 123.325 67.565 123.515 ;
        RECT 68.775 123.325 68.945 123.515 ;
        RECT 69.235 123.325 69.405 123.515 ;
        RECT 70.155 123.345 70.325 123.515 ;
        RECT 71.535 123.345 71.705 123.535 ;
        RECT 74.295 123.325 74.465 123.515 ;
        RECT 74.755 123.345 74.925 123.515 ;
        RECT 77.055 123.345 77.225 123.535 ;
        RECT 78.895 123.345 79.065 123.515 ;
        RECT 79.410 123.375 79.530 123.485 ;
        RECT 80.275 123.345 80.445 123.535 ;
        RECT 80.735 123.345 80.905 123.535 ;
        RECT 81.655 123.345 81.825 123.515 ;
        RECT 83.955 123.345 84.125 123.515 ;
        RECT 84.470 123.375 84.590 123.485 ;
        RECT 74.775 123.325 74.925 123.345 ;
        RECT 78.895 123.325 79.045 123.345 ;
        RECT 81.655 123.325 81.805 123.345 ;
        RECT 83.955 123.325 84.105 123.345 ;
        RECT 86.255 123.325 86.425 123.515 ;
        RECT 89.475 123.345 89.645 123.515 ;
        RECT 89.990 123.375 90.110 123.485 ;
        RECT 93.155 123.325 93.325 123.515 ;
        RECT 93.615 123.345 93.785 123.535 ;
        RECT 94.075 123.345 94.245 123.535 ;
        RECT 98.675 123.325 98.845 123.515 ;
        RECT 103.790 123.375 103.910 123.485 ;
        RECT 104.195 123.325 104.365 123.515 ;
        RECT 104.655 123.325 104.825 123.515 ;
        RECT 106.090 123.375 106.210 123.485 ;
        RECT 106.495 123.345 106.665 123.535 ;
        RECT 108.795 123.515 108.945 123.535 ;
        RECT 108.795 123.345 108.965 123.515 ;
        RECT 109.900 123.325 110.070 123.515 ;
        RECT 110.635 123.345 110.805 123.535 ;
        RECT 112.935 123.515 113.085 123.535 ;
        RECT 111.555 123.325 111.725 123.515 ;
        RECT 112.935 123.345 113.105 123.515 ;
        RECT 115.420 123.325 115.590 123.515 ;
        RECT 115.695 123.345 115.865 123.535 ;
        RECT 116.155 123.345 116.325 123.535 ;
        RECT 125.815 123.325 125.985 123.515 ;
        RECT 126.735 123.345 126.905 123.535 ;
        RECT 127.195 123.325 127.365 123.515 ;
        RECT 127.655 123.485 127.815 123.490 ;
        RECT 127.655 123.380 127.830 123.485 ;
        RECT 127.710 123.375 127.830 123.380 ;
        RECT 129.035 123.325 129.205 123.535 ;
        RECT 9.295 122.515 10.665 123.325 ;
        RECT 11.135 122.515 12.965 123.325 ;
        RECT 12.985 122.455 13.415 123.240 ;
        RECT 13.435 122.515 18.945 123.325 ;
        RECT 18.955 122.515 24.465 123.325 ;
        RECT 24.475 122.515 29.985 123.325 ;
        RECT 30.155 122.505 32.085 123.325 ;
        RECT 32.455 122.505 34.385 123.325 ;
        RECT 34.825 122.645 38.725 123.325 ;
        RECT 31.135 122.415 32.085 122.505 ;
        RECT 33.435 122.415 34.385 122.505 ;
        RECT 37.795 122.415 38.725 122.645 ;
        RECT 38.745 122.455 39.175 123.240 ;
        RECT 39.815 122.505 41.745 123.325 ;
        RECT 41.955 122.545 43.325 123.325 ;
        RECT 43.335 122.515 47.005 123.325 ;
        RECT 47.395 122.645 49.820 123.325 ;
        RECT 50.235 122.515 53.905 123.325 ;
        RECT 54.285 122.645 63.565 123.325 ;
        RECT 54.285 122.525 56.620 122.645 ;
        RECT 40.795 122.415 41.745 122.505 ;
        RECT 54.285 122.415 55.205 122.525 ;
        RECT 61.285 122.425 62.205 122.645 ;
        RECT 64.505 122.455 64.935 123.240 ;
        RECT 64.965 122.645 67.705 123.325 ;
        RECT 67.715 122.515 69.085 123.325 ;
        RECT 69.095 122.645 71.835 123.325 ;
        RECT 71.855 122.515 74.605 123.325 ;
        RECT 74.775 122.505 76.705 123.325 ;
        RECT 75.755 122.415 76.705 122.505 ;
        RECT 77.115 122.505 79.045 123.325 ;
        RECT 79.875 122.505 81.805 123.325 ;
        RECT 82.175 122.505 84.105 123.325 ;
        RECT 84.735 122.515 86.565 123.325 ;
        RECT 86.955 122.645 89.380 123.325 ;
        RECT 77.115 122.415 78.065 122.505 ;
        RECT 79.875 122.415 80.825 122.505 ;
        RECT 82.175 122.415 83.125 122.505 ;
        RECT 90.265 122.455 90.695 123.240 ;
        RECT 90.715 122.515 93.465 123.325 ;
        RECT 93.475 122.515 98.985 123.325 ;
        RECT 98.995 122.515 104.505 123.325 ;
        RECT 104.525 122.415 105.875 123.325 ;
        RECT 106.585 122.645 110.485 123.325 ;
        RECT 109.555 122.415 110.485 122.645 ;
        RECT 110.495 122.515 111.865 123.325 ;
        RECT 112.105 122.645 116.005 123.325 ;
        RECT 115.075 122.415 116.005 122.645 ;
        RECT 116.025 122.455 116.455 123.240 ;
        RECT 116.845 122.645 126.125 123.325 ;
        RECT 116.845 122.525 119.180 122.645 ;
        RECT 116.845 122.415 117.765 122.525 ;
        RECT 123.845 122.425 124.765 122.645 ;
        RECT 126.135 122.545 127.505 123.325 ;
        RECT 127.975 122.515 129.345 123.325 ;
      LAYER nwell ;
        RECT 9.100 119.295 129.540 122.125 ;
      LAYER pwell ;
        RECT 9.295 118.095 10.665 118.905 ;
        RECT 11.135 118.095 16.645 118.905 ;
        RECT 19.855 118.775 20.785 119.005 ;
        RECT 16.885 118.095 20.785 118.775 ;
        RECT 21.715 118.775 22.645 119.005 ;
        RECT 21.715 118.095 25.615 118.775 ;
        RECT 25.865 118.180 26.295 118.965 ;
        RECT 27.235 118.095 30.905 118.905 ;
        RECT 30.915 118.775 31.845 119.005 ;
        RECT 35.885 118.895 36.805 119.005 ;
        RECT 35.885 118.775 38.220 118.895 ;
        RECT 42.885 118.775 43.805 118.995 ;
        RECT 45.375 118.915 46.325 119.005 ;
        RECT 48.595 118.915 49.545 119.005 ;
        RECT 30.915 118.095 34.815 118.775 ;
        RECT 35.885 118.095 45.165 118.775 ;
        RECT 45.375 118.095 47.305 118.915 ;
        RECT 48.595 118.095 50.525 118.915 ;
        RECT 51.625 118.180 52.055 118.965 ;
        RECT 52.995 118.095 58.505 118.905 ;
        RECT 58.525 118.095 59.875 119.005 ;
        RECT 60.815 118.095 64.485 118.905 ;
        RECT 64.495 118.095 65.865 118.875 ;
        RECT 66.335 118.095 71.845 118.905 ;
        RECT 71.855 118.095 77.365 118.905 ;
        RECT 77.385 118.180 77.815 118.965 ;
        RECT 77.835 118.095 79.205 118.905 ;
        RECT 79.215 118.095 80.585 118.875 ;
        RECT 84.715 118.775 85.645 119.005 ;
        RECT 81.745 118.095 85.645 118.775 ;
        RECT 85.655 118.095 87.025 118.905 ;
        RECT 87.405 118.895 88.325 119.005 ;
        RECT 87.405 118.775 89.740 118.895 ;
        RECT 94.405 118.775 95.325 118.995 ;
        RECT 87.405 118.095 96.685 118.775 ;
        RECT 96.695 118.095 98.065 118.905 ;
        RECT 101.275 118.775 102.205 119.005 ;
        RECT 98.305 118.095 102.205 118.775 ;
        RECT 103.145 118.180 103.575 118.965 ;
        RECT 103.965 118.895 104.885 119.005 ;
        RECT 103.965 118.775 106.300 118.895 ;
        RECT 110.965 118.775 111.885 118.995 ;
        RECT 103.965 118.095 113.245 118.775 ;
        RECT 113.715 118.095 115.545 118.905 ;
        RECT 118.755 118.775 119.685 119.005 ;
        RECT 115.785 118.095 119.685 118.775 ;
        RECT 120.165 118.095 121.515 119.005 ;
        RECT 121.535 118.095 122.905 118.875 ;
        RECT 122.915 118.095 124.285 118.905 ;
        RECT 124.295 118.095 127.965 118.905 ;
        RECT 127.975 118.095 129.345 118.905 ;
        RECT 9.435 117.885 9.605 118.095 ;
        RECT 10.870 117.935 10.990 118.045 ;
        RECT 12.655 117.885 12.825 118.075 ;
        RECT 13.575 117.885 13.745 118.075 ;
        RECT 16.335 117.905 16.505 118.095 ;
        RECT 20.200 117.905 20.370 118.095 ;
        RECT 21.395 117.940 21.555 118.050 ;
        RECT 22.130 117.905 22.300 118.095 ;
        RECT 24.155 117.885 24.325 118.075 ;
        RECT 26.915 117.940 27.075 118.050 ;
        RECT 30.595 117.905 30.765 118.095 ;
        RECT 31.330 117.905 31.500 118.095 ;
        RECT 33.815 117.885 33.985 118.075 ;
        RECT 35.195 118.045 35.365 118.075 ;
        RECT 34.735 117.930 34.895 118.040 ;
        RECT 35.195 117.935 35.370 118.045 ;
        RECT 36.630 117.935 36.750 118.045 ;
        RECT 35.195 117.885 35.365 117.935 ;
        RECT 38.415 117.885 38.585 118.075 ;
        RECT 40.255 117.885 40.425 118.075 ;
        RECT 41.635 117.885 41.805 118.075 ;
        RECT 42.555 117.930 42.715 118.040 ;
        RECT 44.855 117.905 45.025 118.095 ;
        RECT 47.155 118.075 47.305 118.095 ;
        RECT 50.375 118.075 50.525 118.095 ;
        RECT 47.155 117.905 47.325 118.075 ;
        RECT 48.075 117.885 48.245 118.075 ;
        RECT 48.535 117.885 48.705 118.075 ;
        RECT 50.375 117.905 50.545 118.075 ;
        RECT 51.295 117.940 51.455 118.050 ;
        RECT 52.675 117.940 52.835 118.050 ;
        RECT 53.320 117.885 53.490 118.075 ;
        RECT 54.055 117.885 54.225 118.075 ;
        RECT 57.730 117.885 57.900 118.075 ;
        RECT 58.195 117.905 58.365 118.095 ;
        RECT 58.655 117.930 58.815 118.040 ;
        RECT 59.575 117.905 59.745 118.095 ;
        RECT 60.495 117.940 60.655 118.050 ;
        RECT 62.335 117.885 62.505 118.075 ;
        RECT 62.795 117.885 62.965 118.075 ;
        RECT 64.175 118.045 64.345 118.095 ;
        RECT 64.175 117.935 64.350 118.045 ;
        RECT 64.175 117.905 64.345 117.935 ;
        RECT 64.635 117.905 64.805 118.095 ;
        RECT 65.555 117.930 65.715 118.040 ;
        RECT 66.070 117.935 66.190 118.045 ;
        RECT 71.075 117.885 71.245 118.075 ;
        RECT 71.535 117.905 71.705 118.095 ;
        RECT 77.055 117.905 77.225 118.095 ;
        RECT 78.895 117.905 79.065 118.095 ;
        RECT 80.275 117.905 80.445 118.095 ;
        RECT 80.735 117.885 80.905 118.075 ;
        RECT 81.195 117.940 81.355 118.050 ;
        RECT 81.470 117.885 81.640 118.075 ;
        RECT 85.060 117.905 85.230 118.095 ;
        RECT 85.795 117.930 85.955 118.040 ;
        RECT 86.715 117.905 86.885 118.095 ;
        RECT 89.660 117.885 89.830 118.075 ;
        RECT 91.315 117.930 91.475 118.040 ;
        RECT 96.375 117.905 96.545 118.095 ;
        RECT 97.755 117.905 97.925 118.095 ;
        RECT 100.975 117.885 101.145 118.075 ;
        RECT 101.620 117.905 101.790 118.095 ;
        RECT 102.355 117.885 102.525 118.075 ;
        RECT 102.815 117.940 102.975 118.050 ;
        RECT 103.275 117.930 103.435 118.040 ;
        RECT 106.955 117.885 107.125 118.075 ;
        RECT 108.335 117.885 108.505 118.075 ;
        RECT 108.795 117.885 108.965 118.075 ;
        RECT 110.230 117.935 110.350 118.045 ;
        RECT 112.935 117.905 113.105 118.095 ;
        RECT 113.450 117.935 113.570 118.045 ;
        RECT 115.235 117.905 115.405 118.095 ;
        RECT 115.695 117.885 115.865 118.075 ;
        RECT 117.995 117.885 118.165 118.075 ;
        RECT 119.100 117.905 119.270 118.095 ;
        RECT 119.375 117.885 119.545 118.075 ;
        RECT 119.890 117.935 120.010 118.045 ;
        RECT 120.295 117.905 120.465 118.095 ;
        RECT 121.675 117.905 121.845 118.095 ;
        RECT 122.135 117.885 122.305 118.075 ;
        RECT 123.975 117.905 124.145 118.095 ;
        RECT 127.655 117.885 127.825 118.095 ;
        RECT 129.035 117.885 129.205 118.095 ;
        RECT 9.295 117.075 10.665 117.885 ;
        RECT 11.135 117.075 12.965 117.885 ;
        RECT 12.985 117.015 13.415 117.800 ;
        RECT 13.445 116.975 14.795 117.885 ;
        RECT 15.185 117.205 24.465 117.885 ;
        RECT 24.845 117.205 34.125 117.885 ;
        RECT 15.185 117.085 17.520 117.205 ;
        RECT 15.185 116.975 16.105 117.085 ;
        RECT 22.185 116.985 23.105 117.205 ;
        RECT 24.845 117.085 27.180 117.205 ;
        RECT 24.845 116.975 25.765 117.085 ;
        RECT 31.845 116.985 32.765 117.205 ;
        RECT 35.065 116.975 36.415 117.885 ;
        RECT 36.895 117.075 38.725 117.885 ;
        RECT 38.745 117.015 39.175 117.800 ;
        RECT 39.195 117.075 40.565 117.885 ;
        RECT 40.575 117.105 41.945 117.885 ;
        RECT 42.875 117.075 48.385 117.885 ;
        RECT 48.405 116.975 49.755 117.885 ;
        RECT 50.005 117.205 53.905 117.885 ;
        RECT 52.975 116.975 53.905 117.205 ;
        RECT 53.915 117.105 55.285 117.885 ;
        RECT 55.435 116.975 58.045 117.885 ;
        RECT 58.975 117.075 62.645 117.885 ;
        RECT 62.665 116.975 64.015 117.885 ;
        RECT 64.505 117.015 64.935 117.800 ;
        RECT 65.875 117.075 71.385 117.885 ;
        RECT 71.765 117.205 81.045 117.885 ;
        RECT 81.055 117.205 84.955 117.885 ;
        RECT 86.345 117.205 90.245 117.885 ;
        RECT 71.765 117.085 74.100 117.205 ;
        RECT 71.765 116.975 72.685 117.085 ;
        RECT 78.765 116.985 79.685 117.205 ;
        RECT 81.055 116.975 81.985 117.205 ;
        RECT 89.315 116.975 90.245 117.205 ;
        RECT 90.265 117.015 90.695 117.800 ;
        RECT 92.005 117.205 101.285 117.885 ;
        RECT 92.005 117.085 94.340 117.205 ;
        RECT 92.005 116.975 92.925 117.085 ;
        RECT 99.005 116.985 99.925 117.205 ;
        RECT 101.295 117.105 102.665 117.885 ;
        RECT 103.595 117.075 107.265 117.885 ;
        RECT 107.275 117.105 108.645 117.885 ;
        RECT 108.655 117.105 110.025 117.885 ;
        RECT 110.495 117.075 116.005 117.885 ;
        RECT 116.025 117.015 116.455 117.800 ;
        RECT 116.475 117.075 118.305 117.885 ;
        RECT 118.325 116.975 119.675 117.885 ;
        RECT 119.695 117.075 122.445 117.885 ;
        RECT 122.455 117.075 127.965 117.885 ;
        RECT 127.975 117.075 129.345 117.885 ;
      LAYER nwell ;
        RECT 9.100 113.855 129.540 116.685 ;
      LAYER pwell ;
        RECT 9.295 112.655 10.665 113.465 ;
        RECT 11.965 113.455 12.885 113.565 ;
        RECT 11.965 113.335 14.300 113.455 ;
        RECT 18.965 113.335 19.885 113.555 ;
        RECT 11.965 112.655 21.245 113.335 ;
        RECT 21.255 112.655 22.625 113.435 ;
        RECT 23.095 112.655 24.465 113.435 ;
        RECT 24.475 112.655 25.845 113.465 ;
        RECT 25.865 112.740 26.295 113.525 ;
        RECT 26.315 112.655 28.145 113.465 ;
        RECT 28.165 112.655 29.515 113.565 ;
        RECT 32.205 113.455 33.125 113.565 ;
        RECT 30.455 112.655 31.825 113.435 ;
        RECT 32.205 113.335 34.540 113.455 ;
        RECT 39.205 113.335 40.125 113.555 ;
        RECT 41.495 113.335 42.425 113.565 ;
        RECT 32.205 112.655 41.485 113.335 ;
        RECT 41.495 112.655 45.395 113.335 ;
        RECT 46.105 112.655 47.455 113.565 ;
        RECT 50.675 113.335 51.605 113.565 ;
        RECT 47.705 112.655 51.605 113.335 ;
        RECT 51.625 112.740 52.055 113.525 ;
        RECT 52.445 113.455 53.365 113.565 ;
        RECT 52.445 113.335 54.780 113.455 ;
        RECT 59.445 113.335 60.365 113.555 ;
        RECT 62.105 113.455 63.025 113.565 ;
        RECT 62.105 113.335 64.440 113.455 ;
        RECT 69.105 113.335 70.025 113.555 ;
        RECT 52.445 112.655 61.725 113.335 ;
        RECT 62.105 112.655 71.385 113.335 ;
        RECT 71.405 112.655 72.755 113.565 ;
        RECT 75.975 113.335 76.905 113.565 ;
        RECT 73.005 112.655 76.905 113.335 ;
        RECT 77.385 112.740 77.815 113.525 ;
        RECT 77.845 112.655 79.195 113.565 ;
        RECT 79.215 112.655 80.585 113.435 ;
        RECT 80.595 112.655 81.965 113.465 ;
        RECT 83.335 113.335 84.255 113.555 ;
        RECT 90.335 113.455 91.255 113.565 ;
        RECT 88.920 113.335 91.255 113.455 ;
        RECT 81.975 112.655 91.255 113.335 ;
        RECT 91.645 112.655 92.995 113.565 ;
        RECT 93.025 112.655 94.375 113.565 ;
        RECT 94.395 112.655 95.765 113.435 ;
        RECT 95.775 112.655 97.605 113.465 ;
        RECT 97.615 112.655 103.125 113.465 ;
        RECT 103.145 112.740 103.575 113.525 ;
        RECT 107.255 113.335 108.185 113.565 ;
        RECT 104.285 112.655 108.185 113.335 ;
        RECT 108.205 112.655 109.555 113.565 ;
        RECT 113.695 113.335 114.625 113.565 ;
        RECT 110.725 112.655 114.625 113.335 ;
        RECT 115.005 113.455 115.925 113.565 ;
        RECT 115.005 113.335 117.340 113.455 ;
        RECT 122.005 113.335 122.925 113.555 ;
        RECT 115.005 112.655 124.285 113.335 ;
        RECT 124.295 112.655 127.965 113.465 ;
        RECT 127.975 112.655 129.345 113.465 ;
        RECT 9.435 112.445 9.605 112.655 ;
        RECT 10.870 112.495 10.990 112.605 ;
        RECT 11.275 112.500 11.435 112.610 ;
        RECT 12.655 112.445 12.825 112.635 ;
        RECT 13.630 112.495 13.750 112.605 ;
        RECT 15.415 112.445 15.585 112.635 ;
        RECT 16.795 112.445 16.965 112.635 ;
        RECT 18.175 112.445 18.345 112.635 ;
        RECT 20.935 112.465 21.105 112.655 ;
        RECT 21.855 112.445 22.025 112.635 ;
        RECT 22.315 112.465 22.485 112.655 ;
        RECT 22.830 112.495 22.950 112.605 ;
        RECT 24.155 112.465 24.325 112.655 ;
        RECT 25.535 112.465 25.705 112.655 ;
        RECT 27.375 112.445 27.545 112.635 ;
        RECT 27.835 112.465 28.005 112.655 ;
        RECT 29.215 112.465 29.385 112.655 ;
        RECT 30.135 112.500 30.295 112.610 ;
        RECT 30.595 112.465 30.765 112.655 ;
        RECT 32.895 112.445 33.065 112.635 ;
        RECT 38.415 112.445 38.585 112.635 ;
        RECT 39.795 112.490 39.955 112.600 ;
        RECT 41.175 112.465 41.345 112.655 ;
        RECT 41.910 112.465 42.080 112.655 ;
        RECT 45.315 112.445 45.485 112.635 ;
        RECT 45.830 112.495 45.950 112.605 ;
        RECT 46.235 112.465 46.405 112.655 ;
        RECT 51.020 112.465 51.190 112.655 ;
        RECT 54.975 112.445 55.145 112.635 ;
        RECT 58.655 112.445 58.825 112.635 ;
        RECT 61.415 112.465 61.585 112.655 ;
        RECT 64.175 112.445 64.345 112.635 ;
        RECT 65.150 112.495 65.270 112.605 ;
        RECT 67.855 112.445 68.025 112.635 ;
        RECT 71.075 112.465 71.245 112.655 ;
        RECT 71.535 112.465 71.705 112.655 ;
        RECT 76.320 112.465 76.490 112.655 ;
        RECT 77.110 112.495 77.230 112.605 ;
        RECT 77.515 112.445 77.685 112.635 ;
        RECT 78.435 112.490 78.595 112.600 ;
        RECT 78.895 112.465 79.065 112.655 ;
        RECT 80.275 112.465 80.445 112.655 ;
        RECT 81.655 112.465 81.825 112.655 ;
        RECT 82.115 112.465 82.285 112.655 ;
        RECT 83.955 112.445 84.125 112.635 ;
        RECT 85.335 112.445 85.505 112.635 ;
        RECT 86.715 112.445 86.885 112.635 ;
        RECT 87.230 112.495 87.350 112.605 ;
        RECT 89.935 112.445 90.105 112.635 ;
        RECT 92.235 112.445 92.405 112.635 ;
        RECT 92.695 112.465 92.865 112.655 ;
        RECT 93.155 112.465 93.325 112.655 ;
        RECT 94.535 112.465 94.705 112.655 ;
        RECT 97.295 112.465 97.465 112.655 ;
        RECT 97.755 112.445 97.925 112.635 ;
        RECT 102.815 112.465 102.985 112.655 ;
        RECT 103.275 112.445 103.445 112.635 ;
        RECT 103.735 112.605 103.905 112.635 ;
        RECT 103.735 112.495 103.910 112.605 ;
        RECT 103.735 112.445 103.905 112.495 ;
        RECT 107.600 112.465 107.770 112.655 ;
        RECT 109.255 112.465 109.425 112.655 ;
        RECT 110.175 112.500 110.335 112.610 ;
        RECT 114.040 112.465 114.210 112.655 ;
        RECT 115.695 112.445 115.865 112.635 ;
        RECT 118.915 112.445 119.085 112.635 ;
        RECT 119.375 112.445 119.545 112.635 ;
        RECT 122.135 112.445 122.305 112.635 ;
        RECT 123.975 112.465 124.145 112.655 ;
        RECT 127.655 112.445 127.825 112.655 ;
        RECT 129.035 112.445 129.205 112.655 ;
        RECT 9.295 111.635 10.665 112.445 ;
        RECT 11.135 111.635 12.965 112.445 ;
        RECT 12.985 111.575 13.415 112.360 ;
        RECT 13.895 111.635 15.725 112.445 ;
        RECT 15.745 111.535 17.095 112.445 ;
        RECT 17.115 111.635 18.485 112.445 ;
        RECT 18.495 111.635 22.165 112.445 ;
        RECT 22.175 111.635 27.685 112.445 ;
        RECT 27.695 111.635 33.205 112.445 ;
        RECT 33.215 111.635 38.725 112.445 ;
        RECT 38.745 111.575 39.175 112.360 ;
        RECT 40.115 111.635 45.625 112.445 ;
        RECT 46.005 111.765 55.285 112.445 ;
        RECT 46.005 111.645 48.340 111.765 ;
        RECT 46.005 111.535 46.925 111.645 ;
        RECT 53.005 111.545 53.925 111.765 ;
        RECT 55.295 111.635 58.965 112.445 ;
        RECT 58.975 111.635 64.485 112.445 ;
        RECT 64.505 111.575 64.935 112.360 ;
        RECT 65.415 111.635 68.165 112.445 ;
        RECT 68.545 111.765 77.825 112.445 ;
        RECT 68.545 111.645 70.880 111.765 ;
        RECT 68.545 111.535 69.465 111.645 ;
        RECT 75.545 111.545 76.465 111.765 ;
        RECT 78.755 111.635 84.265 112.445 ;
        RECT 84.275 111.665 85.645 112.445 ;
        RECT 85.665 111.535 87.015 112.445 ;
        RECT 87.495 111.635 90.245 112.445 ;
        RECT 90.265 111.575 90.695 112.360 ;
        RECT 90.715 111.635 92.545 112.445 ;
        RECT 92.555 111.635 98.065 112.445 ;
        RECT 98.075 111.635 103.585 112.445 ;
        RECT 103.595 111.765 112.875 112.445 ;
        RECT 104.955 111.545 105.875 111.765 ;
        RECT 110.540 111.645 112.875 111.765 ;
        RECT 111.955 111.535 112.875 111.645 ;
        RECT 113.255 111.635 116.005 112.445 ;
        RECT 116.025 111.575 116.455 112.360 ;
        RECT 116.475 111.635 119.225 112.445 ;
        RECT 119.235 111.665 120.605 112.445 ;
        RECT 120.615 111.635 122.445 112.445 ;
        RECT 122.455 111.635 127.965 112.445 ;
        RECT 127.975 111.635 129.345 112.445 ;
      LAYER nwell ;
        RECT 9.100 108.415 129.540 111.245 ;
      LAYER pwell ;
        RECT 9.295 107.215 10.665 108.025 ;
        RECT 10.675 107.895 11.595 108.125 ;
        RECT 14.425 107.895 15.355 108.115 ;
        RECT 10.675 107.215 19.865 107.895 ;
        RECT 19.875 107.215 21.245 108.025 ;
        RECT 21.255 107.215 22.625 107.995 ;
        RECT 23.095 107.215 25.845 108.025 ;
        RECT 25.865 107.300 26.295 108.085 ;
        RECT 27.235 107.215 28.605 107.995 ;
        RECT 29.535 107.215 35.045 108.025 ;
        RECT 35.055 107.215 40.565 108.025 ;
        RECT 40.575 107.215 46.085 108.025 ;
        RECT 46.095 107.215 51.605 108.025 ;
        RECT 51.625 107.300 52.055 108.085 ;
        RECT 52.075 107.215 53.445 107.995 ;
        RECT 53.455 107.215 55.285 108.025 ;
        RECT 55.295 107.215 60.805 108.025 ;
        RECT 60.815 107.215 66.325 108.025 ;
        RECT 66.335 107.215 71.845 108.025 ;
        RECT 71.855 107.215 77.365 108.025 ;
        RECT 77.385 107.300 77.815 108.085 ;
        RECT 78.295 107.215 80.125 108.025 ;
        RECT 80.135 107.215 82.745 108.125 ;
        RECT 83.815 107.215 87.485 108.025 ;
        RECT 87.495 107.215 93.005 108.025 ;
        RECT 93.015 107.215 98.525 108.025 ;
        RECT 98.535 107.215 99.905 107.995 ;
        RECT 100.375 107.215 103.125 108.025 ;
        RECT 103.145 107.300 103.575 108.085 ;
        RECT 103.595 107.215 104.965 108.025 ;
        RECT 104.975 107.215 110.485 108.025 ;
        RECT 110.495 107.215 116.005 108.025 ;
        RECT 116.015 107.215 121.525 108.025 ;
        RECT 121.535 107.215 122.905 107.995 ;
        RECT 122.915 107.215 124.285 107.995 ;
        RECT 124.295 107.215 127.965 108.025 ;
        RECT 127.975 107.215 129.345 108.025 ;
        RECT 9.435 107.005 9.605 107.215 ;
        RECT 10.870 107.055 10.990 107.165 ;
        RECT 12.655 107.005 12.825 107.195 ;
        RECT 14.035 107.050 14.195 107.160 ;
        RECT 15.415 107.005 15.585 107.195 ;
        RECT 19.555 107.025 19.725 107.215 ;
        RECT 20.935 107.025 21.105 107.215 ;
        RECT 22.315 107.025 22.485 107.215 ;
        RECT 22.830 107.055 22.950 107.165 ;
        RECT 24.615 107.005 24.785 107.195 ;
        RECT 25.130 107.055 25.250 107.165 ;
        RECT 25.535 107.025 25.705 107.215 ;
        RECT 26.915 107.005 27.085 107.195 ;
        RECT 28.295 107.005 28.465 107.215 ;
        RECT 29.215 107.060 29.375 107.170 ;
        RECT 31.055 107.005 31.225 107.195 ;
        RECT 32.435 107.005 32.605 107.195 ;
        RECT 32.950 107.055 33.070 107.165 ;
        RECT 34.735 107.025 34.905 107.215 ;
        RECT 36.575 107.005 36.745 107.195 ;
        RECT 37.955 107.005 38.125 107.195 ;
        RECT 38.470 107.055 38.590 107.165 ;
        RECT 39.795 107.050 39.955 107.160 ;
        RECT 40.255 107.025 40.425 107.215 ;
        RECT 41.175 107.005 41.345 107.195 ;
        RECT 42.555 107.005 42.725 107.195 ;
        RECT 43.070 107.055 43.190 107.165 ;
        RECT 44.855 107.005 45.025 107.195 ;
        RECT 45.315 107.005 45.485 107.195 ;
        RECT 45.775 107.025 45.945 107.215 ;
        RECT 46.750 107.055 46.870 107.165 ;
        RECT 48.535 107.005 48.705 107.195 ;
        RECT 51.295 107.025 51.465 107.215 ;
        RECT 52.215 107.025 52.385 107.215 ;
        RECT 54.055 107.005 54.225 107.195 ;
        RECT 54.975 107.025 55.145 107.215 ;
        RECT 55.435 107.005 55.605 107.195 ;
        RECT 57.275 107.005 57.445 107.195 ;
        RECT 57.735 107.005 57.905 107.195 ;
        RECT 60.495 107.025 60.665 107.215 ;
        RECT 61.410 107.005 61.580 107.195 ;
        RECT 62.795 107.005 62.965 107.195 ;
        RECT 64.175 107.005 64.345 107.195 ;
        RECT 66.015 107.025 66.185 107.215 ;
        RECT 67.395 107.005 67.565 107.195 ;
        RECT 71.535 107.025 71.705 107.215 ;
        RECT 72.915 107.005 73.085 107.195 ;
        RECT 74.295 107.005 74.465 107.195 ;
        RECT 77.055 107.025 77.225 107.215 ;
        RECT 78.030 107.055 78.150 107.165 ;
        RECT 79.815 107.025 79.985 107.215 ;
        RECT 80.280 107.025 80.450 107.215 ;
        RECT 83.495 107.005 83.665 107.195 ;
        RECT 84.415 107.050 84.575 107.160 ;
        RECT 87.175 107.025 87.345 107.215 ;
        RECT 89.935 107.005 90.105 107.195 ;
        RECT 91.315 107.050 91.475 107.160 ;
        RECT 91.775 107.005 91.945 107.195 ;
        RECT 92.695 107.025 92.865 107.215 ;
        RECT 93.210 107.055 93.330 107.165 ;
        RECT 98.215 107.025 98.385 107.215 ;
        RECT 98.675 107.025 98.845 107.215 ;
        RECT 100.110 107.055 100.230 107.165 ;
        RECT 102.355 107.005 102.525 107.195 ;
        RECT 102.815 107.165 102.985 107.215 ;
        RECT 102.815 107.055 102.990 107.165 ;
        RECT 102.815 107.025 102.985 107.055 ;
        RECT 104.655 107.005 104.825 107.215 ;
        RECT 105.115 107.005 105.285 107.195 ;
        RECT 106.955 107.050 107.115 107.160 ;
        RECT 107.415 107.005 107.585 107.195 ;
        RECT 108.795 107.005 108.965 107.195 ;
        RECT 110.175 107.025 110.345 107.215 ;
        RECT 113.395 107.005 113.565 107.195 ;
        RECT 113.855 107.005 114.025 107.195 ;
        RECT 115.695 107.025 115.865 107.215 ;
        RECT 117.075 107.050 117.235 107.160 ;
        RECT 117.535 107.005 117.705 107.195 ;
        RECT 118.915 107.005 119.085 107.195 ;
        RECT 121.215 107.025 121.385 107.215 ;
        RECT 122.595 107.025 122.765 107.215 ;
        RECT 123.975 107.025 124.145 107.215 ;
        RECT 127.655 107.025 127.825 107.215 ;
        RECT 129.035 107.005 129.205 107.215 ;
        RECT 9.295 106.195 10.665 107.005 ;
        RECT 11.135 106.195 12.965 107.005 ;
        RECT 12.985 106.135 13.415 106.920 ;
        RECT 14.365 106.095 15.715 107.005 ;
        RECT 15.735 106.325 24.925 107.005 ;
        RECT 15.735 106.095 16.655 106.325 ;
        RECT 19.485 106.105 20.415 106.325 ;
        RECT 25.395 106.195 27.225 107.005 ;
        RECT 27.235 106.225 28.605 107.005 ;
        RECT 28.615 106.195 31.365 107.005 ;
        RECT 31.375 106.225 32.745 107.005 ;
        RECT 33.215 106.195 36.885 107.005 ;
        RECT 36.895 106.225 38.265 107.005 ;
        RECT 38.745 106.135 39.175 106.920 ;
        RECT 40.125 106.095 41.475 107.005 ;
        RECT 41.495 106.225 42.865 107.005 ;
        RECT 43.335 106.195 45.165 107.005 ;
        RECT 45.175 106.225 46.545 107.005 ;
        RECT 47.015 106.195 48.845 107.005 ;
        RECT 48.855 106.195 54.365 107.005 ;
        RECT 54.375 106.225 55.745 107.005 ;
        RECT 55.755 106.195 57.585 107.005 ;
        RECT 57.595 106.225 58.965 107.005 ;
        RECT 59.115 106.095 61.725 107.005 ;
        RECT 61.735 106.195 63.105 107.005 ;
        RECT 63.115 106.225 64.485 107.005 ;
        RECT 64.505 106.135 64.935 106.920 ;
        RECT 64.955 106.195 67.705 107.005 ;
        RECT 67.715 106.195 73.225 107.005 ;
        RECT 73.245 106.095 74.595 107.005 ;
        RECT 74.615 106.325 83.805 107.005 ;
        RECT 74.615 106.095 75.535 106.325 ;
        RECT 78.365 106.105 79.295 106.325 ;
        RECT 84.735 106.195 90.245 107.005 ;
        RECT 90.265 106.135 90.695 106.920 ;
        RECT 91.635 106.225 93.005 107.005 ;
        RECT 93.475 106.325 102.665 107.005 ;
        RECT 93.475 106.095 94.395 106.325 ;
        RECT 97.225 106.105 98.155 106.325 ;
        RECT 103.135 106.195 104.965 107.005 ;
        RECT 104.975 106.225 106.345 107.005 ;
        RECT 107.285 106.095 108.635 107.005 ;
        RECT 108.655 106.225 110.025 107.005 ;
        RECT 110.035 106.195 113.705 107.005 ;
        RECT 113.715 106.225 115.085 107.005 ;
        RECT 116.025 106.135 116.455 106.920 ;
        RECT 117.405 106.095 118.755 107.005 ;
        RECT 118.775 106.325 127.965 107.005 ;
        RECT 123.285 106.105 124.215 106.325 ;
        RECT 127.045 106.095 127.965 106.325 ;
        RECT 127.975 106.195 129.345 107.005 ;
      LAYER nwell ;
        RECT 9.100 102.975 129.540 105.805 ;
      LAYER pwell ;
        RECT 9.295 101.775 10.665 102.585 ;
        RECT 11.595 101.775 15.265 102.585 ;
        RECT 15.285 101.775 16.635 102.685 ;
        RECT 16.655 102.455 17.575 102.685 ;
        RECT 20.405 102.455 21.335 102.675 ;
        RECT 16.655 101.775 25.845 102.455 ;
        RECT 25.865 101.860 26.295 102.645 ;
        RECT 26.785 101.775 28.135 102.685 ;
        RECT 28.155 101.775 31.825 102.585 ;
        RECT 31.845 101.775 33.195 102.685 ;
        RECT 37.725 102.455 38.655 102.675 ;
        RECT 41.485 102.455 42.405 102.685 ;
        RECT 33.215 101.775 42.405 102.455 ;
        RECT 42.415 102.455 43.335 102.685 ;
        RECT 46.165 102.455 47.095 102.675 ;
        RECT 42.415 101.775 51.605 102.455 ;
        RECT 51.625 101.860 52.055 102.645 ;
        RECT 52.075 101.775 53.905 102.585 ;
        RECT 53.925 101.775 55.275 102.685 ;
        RECT 55.755 101.775 57.585 102.585 ;
        RECT 57.605 101.775 58.955 102.685 ;
        RECT 58.985 101.775 60.335 102.685 ;
        RECT 64.865 102.455 65.795 102.675 ;
        RECT 68.625 102.455 69.545 102.685 ;
        RECT 60.355 101.775 69.545 102.455 ;
        RECT 69.555 101.775 70.925 102.585 ;
        RECT 70.935 101.775 74.605 102.585 ;
        RECT 74.625 101.775 75.975 102.685 ;
        RECT 76.005 101.775 77.355 102.685 ;
        RECT 77.385 101.860 77.815 102.645 ;
        RECT 77.835 101.775 79.205 102.555 ;
        RECT 79.215 101.775 80.585 102.555 ;
        RECT 80.595 101.775 84.265 102.585 ;
        RECT 84.285 101.775 85.635 102.685 ;
        RECT 85.655 101.775 87.025 102.555 ;
        RECT 87.045 101.775 88.395 102.685 ;
        RECT 88.415 102.455 89.335 102.685 ;
        RECT 92.165 102.455 93.095 102.675 ;
        RECT 88.415 101.775 97.605 102.455 ;
        RECT 97.625 101.775 98.975 102.685 ;
        RECT 98.995 101.775 101.745 102.585 ;
        RECT 101.765 101.775 103.115 102.685 ;
        RECT 103.145 101.860 103.575 102.645 ;
        RECT 109.025 102.455 109.955 102.675 ;
        RECT 112.785 102.455 113.705 102.685 ;
        RECT 104.515 101.775 113.705 102.455 ;
        RECT 113.715 101.775 115.545 102.585 ;
        RECT 115.565 101.775 116.915 102.685 ;
        RECT 117.405 101.775 118.755 102.685 ;
        RECT 123.285 102.455 124.215 102.675 ;
        RECT 127.045 102.455 127.965 102.685 ;
        RECT 118.775 101.775 127.965 102.455 ;
        RECT 127.975 101.775 129.345 102.585 ;
        RECT 9.435 101.565 9.605 101.775 ;
        RECT 10.870 101.615 10.990 101.725 ;
        RECT 11.275 101.620 11.435 101.730 ;
        RECT 12.655 101.565 12.825 101.755 ;
        RECT 14.955 101.585 15.125 101.775 ;
        RECT 16.335 101.585 16.505 101.775 ;
        RECT 18.635 101.565 18.805 101.755 ;
        RECT 19.095 101.565 19.265 101.755 ;
        RECT 20.475 101.565 20.645 101.755 ;
        RECT 25.535 101.585 25.705 101.775 ;
        RECT 26.510 101.615 26.630 101.725 ;
        RECT 27.835 101.585 28.005 101.775 ;
        RECT 31.515 101.585 31.685 101.775 ;
        RECT 31.975 101.585 32.145 101.775 ;
        RECT 33.355 101.585 33.525 101.775 ;
        RECT 38.415 101.565 38.585 101.755 ;
        RECT 44.395 101.565 44.565 101.755 ;
        RECT 44.855 101.565 45.025 101.755 ;
        RECT 46.235 101.565 46.405 101.755 ;
        RECT 51.295 101.585 51.465 101.775 ;
        RECT 53.595 101.585 53.765 101.775 ;
        RECT 54.975 101.585 55.145 101.775 ;
        RECT 55.490 101.615 55.610 101.725 ;
        RECT 57.275 101.585 57.445 101.775 ;
        RECT 57.735 101.585 57.905 101.775 ;
        RECT 59.115 101.585 59.285 101.775 ;
        RECT 60.495 101.585 60.665 101.775 ;
        RECT 64.175 101.565 64.345 101.755 ;
        RECT 65.555 101.610 65.715 101.720 ;
        RECT 70.615 101.585 70.785 101.775 ;
        RECT 71.075 101.565 71.245 101.755 ;
        RECT 74.295 101.585 74.465 101.775 ;
        RECT 75.675 101.585 75.845 101.775 ;
        RECT 77.055 101.585 77.225 101.775 ;
        RECT 77.975 101.585 78.145 101.775 ;
        RECT 79.355 101.585 79.525 101.775 ;
        RECT 80.275 101.565 80.445 101.755 ;
        RECT 80.790 101.615 80.910 101.725 ;
        RECT 83.955 101.585 84.125 101.775 ;
        RECT 85.335 101.585 85.505 101.775 ;
        RECT 85.795 101.585 85.965 101.775 ;
        RECT 87.175 101.585 87.345 101.775 ;
        RECT 89.935 101.565 90.105 101.755 ;
        RECT 94.075 101.565 94.245 101.755 ;
        RECT 97.295 101.585 97.465 101.775 ;
        RECT 98.675 101.585 98.845 101.775 ;
        RECT 99.595 101.565 99.765 101.755 ;
        RECT 101.435 101.585 101.605 101.775 ;
        RECT 101.895 101.585 102.065 101.775 ;
        RECT 104.195 101.620 104.355 101.730 ;
        RECT 104.655 101.585 104.825 101.775 ;
        RECT 108.795 101.565 108.965 101.755 ;
        RECT 110.175 101.565 110.345 101.755 ;
        RECT 115.235 101.585 115.405 101.775 ;
        RECT 115.695 101.565 115.865 101.775 ;
        RECT 117.130 101.615 117.250 101.725 ;
        RECT 117.535 101.585 117.705 101.775 ;
        RECT 118.915 101.585 119.085 101.775 ;
        RECT 125.355 101.565 125.525 101.755 ;
        RECT 126.275 101.610 126.435 101.720 ;
        RECT 127.645 101.565 127.815 101.755 ;
        RECT 129.035 101.565 129.205 101.775 ;
        RECT 9.295 100.755 10.665 101.565 ;
        RECT 11.135 100.755 12.965 101.565 ;
        RECT 12.985 100.695 13.415 101.480 ;
        RECT 13.435 100.755 18.945 101.565 ;
        RECT 18.965 100.655 20.315 101.565 ;
        RECT 20.335 100.885 29.525 101.565 ;
        RECT 24.845 100.665 25.775 100.885 ;
        RECT 28.605 100.655 29.525 100.885 ;
        RECT 29.535 100.885 38.725 101.565 ;
        RECT 29.535 100.655 30.455 100.885 ;
        RECT 33.285 100.665 34.215 100.885 ;
        RECT 38.745 100.695 39.175 101.480 ;
        RECT 39.195 100.755 44.705 101.565 ;
        RECT 44.725 100.655 46.075 101.565 ;
        RECT 46.095 100.885 55.285 101.565 ;
        RECT 50.605 100.665 51.535 100.885 ;
        RECT 54.365 100.655 55.285 100.885 ;
        RECT 55.295 100.885 64.485 101.565 ;
        RECT 55.295 100.655 56.215 100.885 ;
        RECT 59.045 100.665 59.975 100.885 ;
        RECT 64.505 100.695 64.935 101.480 ;
        RECT 65.875 100.755 71.385 101.565 ;
        RECT 71.395 100.885 80.585 101.565 ;
        RECT 81.055 100.885 90.245 101.565 ;
        RECT 71.395 100.655 72.315 100.885 ;
        RECT 75.145 100.665 76.075 100.885 ;
        RECT 81.055 100.655 81.975 100.885 ;
        RECT 84.805 100.665 85.735 100.885 ;
        RECT 90.265 100.695 90.695 101.480 ;
        RECT 90.715 100.755 94.385 101.565 ;
        RECT 94.395 100.755 99.905 101.565 ;
        RECT 99.915 100.885 109.105 101.565 ;
        RECT 99.915 100.655 100.835 100.885 ;
        RECT 103.665 100.665 104.595 100.885 ;
        RECT 109.115 100.755 110.485 101.565 ;
        RECT 110.495 100.755 116.005 101.565 ;
        RECT 116.025 100.695 116.455 101.480 ;
        RECT 116.475 100.885 125.665 101.565 ;
        RECT 116.475 100.655 117.395 100.885 ;
        RECT 120.225 100.665 121.155 100.885 ;
        RECT 126.595 100.785 127.965 101.565 ;
        RECT 127.975 100.755 129.345 101.565 ;
      LAYER nwell ;
        RECT 9.100 97.535 129.540 100.365 ;
      LAYER pwell ;
        RECT 9.295 96.335 10.665 97.145 ;
        RECT 11.135 96.335 12.965 97.145 ;
        RECT 12.985 96.420 13.415 97.205 ;
        RECT 13.435 96.335 14.805 97.145 ;
        RECT 14.815 96.335 20.325 97.145 ;
        RECT 20.335 96.335 25.845 97.145 ;
        RECT 25.865 96.420 26.295 97.205 ;
        RECT 26.315 96.335 27.685 97.145 ;
        RECT 27.695 96.335 33.205 97.145 ;
        RECT 33.215 96.335 38.725 97.145 ;
        RECT 38.745 96.420 39.175 97.205 ;
        RECT 39.195 96.335 40.565 97.145 ;
        RECT 40.575 96.335 46.085 97.145 ;
        RECT 46.095 96.335 51.605 97.145 ;
        RECT 51.625 96.420 52.055 97.205 ;
        RECT 52.075 96.335 53.445 97.145 ;
        RECT 53.455 96.335 58.965 97.145 ;
        RECT 58.975 96.335 64.485 97.145 ;
        RECT 64.505 96.420 64.935 97.205 ;
        RECT 64.955 96.335 66.325 97.145 ;
        RECT 66.335 96.335 71.845 97.145 ;
        RECT 71.855 96.335 77.365 97.145 ;
        RECT 77.385 96.420 77.815 97.205 ;
        RECT 77.835 96.335 79.205 97.145 ;
        RECT 79.215 96.335 84.725 97.145 ;
        RECT 84.735 96.335 90.245 97.145 ;
        RECT 90.265 96.420 90.695 97.205 ;
        RECT 90.715 96.335 92.085 97.145 ;
        RECT 92.095 96.335 97.605 97.145 ;
        RECT 97.615 96.335 103.125 97.145 ;
        RECT 103.145 96.420 103.575 97.205 ;
        RECT 103.595 96.335 104.965 97.145 ;
        RECT 104.975 96.335 110.485 97.145 ;
        RECT 110.495 96.335 116.005 97.145 ;
        RECT 116.025 96.420 116.455 97.205 ;
        RECT 116.935 96.335 122.445 97.145 ;
        RECT 122.455 96.335 127.965 97.145 ;
        RECT 127.975 96.335 129.345 97.145 ;
        RECT 9.435 96.145 9.605 96.335 ;
        RECT 10.870 96.175 10.990 96.285 ;
        RECT 12.655 96.145 12.825 96.335 ;
        RECT 14.495 96.145 14.665 96.335 ;
        RECT 20.015 96.145 20.185 96.335 ;
        RECT 25.535 96.145 25.705 96.335 ;
        RECT 27.375 96.145 27.545 96.335 ;
        RECT 32.895 96.145 33.065 96.335 ;
        RECT 38.415 96.145 38.585 96.335 ;
        RECT 40.255 96.145 40.425 96.335 ;
        RECT 45.775 96.145 45.945 96.335 ;
        RECT 51.295 96.145 51.465 96.335 ;
        RECT 53.135 96.145 53.305 96.335 ;
        RECT 58.655 96.145 58.825 96.335 ;
        RECT 64.175 96.145 64.345 96.335 ;
        RECT 66.015 96.145 66.185 96.335 ;
        RECT 71.535 96.145 71.705 96.335 ;
        RECT 77.055 96.145 77.225 96.335 ;
        RECT 78.895 96.145 79.065 96.335 ;
        RECT 84.415 96.145 84.585 96.335 ;
        RECT 89.935 96.145 90.105 96.335 ;
        RECT 91.775 96.145 91.945 96.335 ;
        RECT 97.295 96.145 97.465 96.335 ;
        RECT 102.815 96.145 102.985 96.335 ;
        RECT 104.655 96.145 104.825 96.335 ;
        RECT 110.175 96.145 110.345 96.335 ;
        RECT 115.695 96.145 115.865 96.335 ;
        RECT 116.670 96.175 116.790 96.285 ;
        RECT 122.135 96.145 122.305 96.335 ;
        RECT 127.655 96.145 127.825 96.335 ;
        RECT 129.035 96.145 129.205 96.335 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 9.290 215.825 129.350 215.995 ;
        RECT 9.375 215.075 10.585 215.825 ;
        RECT 9.375 214.535 9.895 215.075 ;
        RECT 11.215 215.055 12.885 215.825 ;
        RECT 13.055 215.100 13.345 215.825 ;
        RECT 13.515 215.075 14.725 215.825 ;
        RECT 14.900 215.280 20.245 215.825 ;
        RECT 20.420 215.280 25.765 215.825 ;
        RECT 10.065 214.365 10.585 214.905 ;
        RECT 9.375 213.275 10.585 214.365 ;
        RECT 11.215 214.365 11.965 214.885 ;
        RECT 12.135 214.535 12.885 215.055 ;
        RECT 11.215 213.275 12.885 214.365 ;
        RECT 13.055 213.275 13.345 214.440 ;
        RECT 13.515 214.365 14.035 214.905 ;
        RECT 14.205 214.535 14.725 215.075 ;
        RECT 13.515 213.275 14.725 214.365 ;
        RECT 16.490 213.710 16.840 214.960 ;
        RECT 18.320 214.450 18.660 215.280 ;
        RECT 22.010 213.710 22.360 214.960 ;
        RECT 23.840 214.450 24.180 215.280 ;
        RECT 25.935 215.100 26.225 215.825 ;
        RECT 26.395 215.075 27.605 215.825 ;
        RECT 27.780 215.280 33.125 215.825 ;
        RECT 33.300 215.280 38.645 215.825 ;
        RECT 14.900 213.275 20.245 213.710 ;
        RECT 20.420 213.275 25.765 213.710 ;
        RECT 25.935 213.275 26.225 214.440 ;
        RECT 26.395 214.365 26.915 214.905 ;
        RECT 27.085 214.535 27.605 215.075 ;
        RECT 26.395 213.275 27.605 214.365 ;
        RECT 29.370 213.710 29.720 214.960 ;
        RECT 31.200 214.450 31.540 215.280 ;
        RECT 34.890 213.710 35.240 214.960 ;
        RECT 36.720 214.450 37.060 215.280 ;
        RECT 38.815 215.100 39.105 215.825 ;
        RECT 39.275 215.075 40.485 215.825 ;
        RECT 40.660 215.280 46.005 215.825 ;
        RECT 46.180 215.280 51.525 215.825 ;
        RECT 27.780 213.275 33.125 213.710 ;
        RECT 33.300 213.275 38.645 213.710 ;
        RECT 38.815 213.275 39.105 214.440 ;
        RECT 39.275 214.365 39.795 214.905 ;
        RECT 39.965 214.535 40.485 215.075 ;
        RECT 39.275 213.275 40.485 214.365 ;
        RECT 42.250 213.710 42.600 214.960 ;
        RECT 44.080 214.450 44.420 215.280 ;
        RECT 47.770 213.710 48.120 214.960 ;
        RECT 49.600 214.450 49.940 215.280 ;
        RECT 51.695 215.100 51.985 215.825 ;
        RECT 52.155 215.075 53.365 215.825 ;
        RECT 53.540 215.280 58.885 215.825 ;
        RECT 59.060 215.280 64.405 215.825 ;
        RECT 40.660 213.275 46.005 213.710 ;
        RECT 46.180 213.275 51.525 213.710 ;
        RECT 51.695 213.275 51.985 214.440 ;
        RECT 52.155 214.365 52.675 214.905 ;
        RECT 52.845 214.535 53.365 215.075 ;
        RECT 52.155 213.275 53.365 214.365 ;
        RECT 55.130 213.710 55.480 214.960 ;
        RECT 56.960 214.450 57.300 215.280 ;
        RECT 60.650 213.710 61.000 214.960 ;
        RECT 62.480 214.450 62.820 215.280 ;
        RECT 64.575 215.100 64.865 215.825 ;
        RECT 65.035 215.075 66.245 215.825 ;
        RECT 66.420 215.280 71.765 215.825 ;
        RECT 71.940 215.280 77.285 215.825 ;
        RECT 53.540 213.275 58.885 213.710 ;
        RECT 59.060 213.275 64.405 213.710 ;
        RECT 64.575 213.275 64.865 214.440 ;
        RECT 65.035 214.365 65.555 214.905 ;
        RECT 65.725 214.535 66.245 215.075 ;
        RECT 65.035 213.275 66.245 214.365 ;
        RECT 68.010 213.710 68.360 214.960 ;
        RECT 69.840 214.450 70.180 215.280 ;
        RECT 73.530 213.710 73.880 214.960 ;
        RECT 75.360 214.450 75.700 215.280 ;
        RECT 77.455 215.100 77.745 215.825 ;
        RECT 77.915 215.075 79.125 215.825 ;
        RECT 79.300 215.280 84.645 215.825 ;
        RECT 84.820 215.280 90.165 215.825 ;
        RECT 66.420 213.275 71.765 213.710 ;
        RECT 71.940 213.275 77.285 213.710 ;
        RECT 77.455 213.275 77.745 214.440 ;
        RECT 77.915 214.365 78.435 214.905 ;
        RECT 78.605 214.535 79.125 215.075 ;
        RECT 77.915 213.275 79.125 214.365 ;
        RECT 80.890 213.710 81.240 214.960 ;
        RECT 82.720 214.450 83.060 215.280 ;
        RECT 86.410 213.710 86.760 214.960 ;
        RECT 88.240 214.450 88.580 215.280 ;
        RECT 90.335 215.100 90.625 215.825 ;
        RECT 90.795 215.075 92.005 215.825 ;
        RECT 92.180 215.280 97.525 215.825 ;
        RECT 97.700 215.280 103.045 215.825 ;
        RECT 79.300 213.275 84.645 213.710 ;
        RECT 84.820 213.275 90.165 213.710 ;
        RECT 90.335 213.275 90.625 214.440 ;
        RECT 90.795 214.365 91.315 214.905 ;
        RECT 91.485 214.535 92.005 215.075 ;
        RECT 90.795 213.275 92.005 214.365 ;
        RECT 93.770 213.710 94.120 214.960 ;
        RECT 95.600 214.450 95.940 215.280 ;
        RECT 99.290 213.710 99.640 214.960 ;
        RECT 101.120 214.450 101.460 215.280 ;
        RECT 103.215 215.100 103.505 215.825 ;
        RECT 103.675 215.075 104.885 215.825 ;
        RECT 105.060 215.280 110.405 215.825 ;
        RECT 110.580 215.280 115.925 215.825 ;
        RECT 92.180 213.275 97.525 213.710 ;
        RECT 97.700 213.275 103.045 213.710 ;
        RECT 103.215 213.275 103.505 214.440 ;
        RECT 103.675 214.365 104.195 214.905 ;
        RECT 104.365 214.535 104.885 215.075 ;
        RECT 103.675 213.275 104.885 214.365 ;
        RECT 106.650 213.710 107.000 214.960 ;
        RECT 108.480 214.450 108.820 215.280 ;
        RECT 112.170 213.710 112.520 214.960 ;
        RECT 114.000 214.450 114.340 215.280 ;
        RECT 116.095 215.100 116.385 215.825 ;
        RECT 117.020 215.280 122.365 215.825 ;
        RECT 122.540 215.280 127.885 215.825 ;
        RECT 105.060 213.275 110.405 213.710 ;
        RECT 110.580 213.275 115.925 213.710 ;
        RECT 116.095 213.275 116.385 214.440 ;
        RECT 118.610 213.710 118.960 214.960 ;
        RECT 120.440 214.450 120.780 215.280 ;
        RECT 124.130 213.710 124.480 214.960 ;
        RECT 125.960 214.450 126.300 215.280 ;
        RECT 128.055 215.075 129.265 215.825 ;
        RECT 128.055 214.365 128.575 214.905 ;
        RECT 128.745 214.535 129.265 215.075 ;
        RECT 117.020 213.275 122.365 213.710 ;
        RECT 122.540 213.275 127.885 213.710 ;
        RECT 128.055 213.275 129.265 214.365 ;
        RECT 9.290 213.105 129.350 213.275 ;
        RECT 9.375 212.015 10.585 213.105 ;
        RECT 9.375 211.305 9.895 211.845 ;
        RECT 10.065 211.475 10.585 212.015 ;
        RECT 11.215 212.015 14.725 213.105 ;
        RECT 14.900 212.670 20.245 213.105 ;
        RECT 20.420 212.670 25.765 213.105 ;
        RECT 11.215 211.495 12.905 212.015 ;
        RECT 13.075 211.325 14.725 211.845 ;
        RECT 16.490 211.420 16.840 212.670 ;
        RECT 9.375 210.555 10.585 211.305 ;
        RECT 11.215 210.555 14.725 211.325 ;
        RECT 18.320 211.100 18.660 211.930 ;
        RECT 22.010 211.420 22.360 212.670 ;
        RECT 25.935 211.940 26.225 213.105 ;
        RECT 26.855 212.015 29.445 213.105 ;
        RECT 29.620 212.670 34.965 213.105 ;
        RECT 35.140 212.670 40.485 213.105 ;
        RECT 40.660 212.670 46.005 213.105 ;
        RECT 46.180 212.670 51.525 213.105 ;
        RECT 23.840 211.100 24.180 211.930 ;
        RECT 26.855 211.495 28.065 212.015 ;
        RECT 28.235 211.325 29.445 211.845 ;
        RECT 31.210 211.420 31.560 212.670 ;
        RECT 14.900 210.555 20.245 211.100 ;
        RECT 20.420 210.555 25.765 211.100 ;
        RECT 25.935 210.555 26.225 211.280 ;
        RECT 26.855 210.555 29.445 211.325 ;
        RECT 33.040 211.100 33.380 211.930 ;
        RECT 36.730 211.420 37.080 212.670 ;
        RECT 38.560 211.100 38.900 211.930 ;
        RECT 42.250 211.420 42.600 212.670 ;
        RECT 44.080 211.100 44.420 211.930 ;
        RECT 47.770 211.420 48.120 212.670 ;
        RECT 51.695 211.940 51.985 213.105 ;
        RECT 52.615 212.015 55.205 213.105 ;
        RECT 55.380 212.670 60.725 213.105 ;
        RECT 60.900 212.670 66.245 213.105 ;
        RECT 66.420 212.670 71.765 213.105 ;
        RECT 71.940 212.670 77.285 213.105 ;
        RECT 49.600 211.100 49.940 211.930 ;
        RECT 52.615 211.495 53.825 212.015 ;
        RECT 53.995 211.325 55.205 211.845 ;
        RECT 56.970 211.420 57.320 212.670 ;
        RECT 29.620 210.555 34.965 211.100 ;
        RECT 35.140 210.555 40.485 211.100 ;
        RECT 40.660 210.555 46.005 211.100 ;
        RECT 46.180 210.555 51.525 211.100 ;
        RECT 51.695 210.555 51.985 211.280 ;
        RECT 52.615 210.555 55.205 211.325 ;
        RECT 58.800 211.100 59.140 211.930 ;
        RECT 62.490 211.420 62.840 212.670 ;
        RECT 64.320 211.100 64.660 211.930 ;
        RECT 68.010 211.420 68.360 212.670 ;
        RECT 69.840 211.100 70.180 211.930 ;
        RECT 73.530 211.420 73.880 212.670 ;
        RECT 77.455 211.940 77.745 213.105 ;
        RECT 78.375 212.015 80.965 213.105 ;
        RECT 81.140 212.670 86.485 213.105 ;
        RECT 86.660 212.670 92.005 213.105 ;
        RECT 92.180 212.670 97.525 213.105 ;
        RECT 97.700 212.670 103.045 213.105 ;
        RECT 75.360 211.100 75.700 211.930 ;
        RECT 78.375 211.495 79.585 212.015 ;
        RECT 79.755 211.325 80.965 211.845 ;
        RECT 82.730 211.420 83.080 212.670 ;
        RECT 55.380 210.555 60.725 211.100 ;
        RECT 60.900 210.555 66.245 211.100 ;
        RECT 66.420 210.555 71.765 211.100 ;
        RECT 71.940 210.555 77.285 211.100 ;
        RECT 77.455 210.555 77.745 211.280 ;
        RECT 78.375 210.555 80.965 211.325 ;
        RECT 84.560 211.100 84.900 211.930 ;
        RECT 88.250 211.420 88.600 212.670 ;
        RECT 90.080 211.100 90.420 211.930 ;
        RECT 93.770 211.420 94.120 212.670 ;
        RECT 95.600 211.100 95.940 211.930 ;
        RECT 99.290 211.420 99.640 212.670 ;
        RECT 103.215 211.940 103.505 213.105 ;
        RECT 104.135 212.015 105.805 213.105 ;
        RECT 105.980 212.670 111.325 213.105 ;
        RECT 111.500 212.670 116.845 213.105 ;
        RECT 117.020 212.670 122.365 213.105 ;
        RECT 122.540 212.670 127.885 213.105 ;
        RECT 101.120 211.100 101.460 211.930 ;
        RECT 104.135 211.495 104.885 212.015 ;
        RECT 105.055 211.325 105.805 211.845 ;
        RECT 107.570 211.420 107.920 212.670 ;
        RECT 81.140 210.555 86.485 211.100 ;
        RECT 86.660 210.555 92.005 211.100 ;
        RECT 92.180 210.555 97.525 211.100 ;
        RECT 97.700 210.555 103.045 211.100 ;
        RECT 103.215 210.555 103.505 211.280 ;
        RECT 104.135 210.555 105.805 211.325 ;
        RECT 109.400 211.100 109.740 211.930 ;
        RECT 113.090 211.420 113.440 212.670 ;
        RECT 114.920 211.100 115.260 211.930 ;
        RECT 118.610 211.420 118.960 212.670 ;
        RECT 120.440 211.100 120.780 211.930 ;
        RECT 124.130 211.420 124.480 212.670 ;
        RECT 128.055 212.015 129.265 213.105 ;
        RECT 125.960 211.100 126.300 211.930 ;
        RECT 128.055 211.475 128.575 212.015 ;
        RECT 128.745 211.305 129.265 211.845 ;
        RECT 105.980 210.555 111.325 211.100 ;
        RECT 111.500 210.555 116.845 211.100 ;
        RECT 117.020 210.555 122.365 211.100 ;
        RECT 122.540 210.555 127.885 211.100 ;
        RECT 128.055 210.555 129.265 211.305 ;
        RECT 9.290 210.385 129.350 210.555 ;
        RECT 9.375 209.635 10.585 210.385 ;
        RECT 9.375 209.095 9.895 209.635 ;
        RECT 11.215 209.615 12.885 210.385 ;
        RECT 13.055 209.660 13.345 210.385 ;
        RECT 13.975 209.615 16.565 210.385 ;
        RECT 16.740 209.840 22.085 210.385 ;
        RECT 22.260 209.840 27.605 210.385 ;
        RECT 27.780 209.840 33.125 210.385 ;
        RECT 33.300 209.840 38.645 210.385 ;
        RECT 10.065 208.925 10.585 209.465 ;
        RECT 9.375 207.835 10.585 208.925 ;
        RECT 11.215 208.925 11.965 209.445 ;
        RECT 12.135 209.095 12.885 209.615 ;
        RECT 11.215 207.835 12.885 208.925 ;
        RECT 13.055 207.835 13.345 209.000 ;
        RECT 13.975 208.925 15.185 209.445 ;
        RECT 15.355 209.095 16.565 209.615 ;
        RECT 13.975 207.835 16.565 208.925 ;
        RECT 18.330 208.270 18.680 209.520 ;
        RECT 20.160 209.010 20.500 209.840 ;
        RECT 23.850 208.270 24.200 209.520 ;
        RECT 25.680 209.010 26.020 209.840 ;
        RECT 29.370 208.270 29.720 209.520 ;
        RECT 31.200 209.010 31.540 209.840 ;
        RECT 34.890 208.270 35.240 209.520 ;
        RECT 36.720 209.010 37.060 209.840 ;
        RECT 38.815 209.660 39.105 210.385 ;
        RECT 39.735 209.615 42.325 210.385 ;
        RECT 42.500 209.840 47.845 210.385 ;
        RECT 48.020 209.840 53.365 210.385 ;
        RECT 53.540 209.840 58.885 210.385 ;
        RECT 59.060 209.840 64.405 210.385 ;
        RECT 16.740 207.835 22.085 208.270 ;
        RECT 22.260 207.835 27.605 208.270 ;
        RECT 27.780 207.835 33.125 208.270 ;
        RECT 33.300 207.835 38.645 208.270 ;
        RECT 38.815 207.835 39.105 209.000 ;
        RECT 39.735 208.925 40.945 209.445 ;
        RECT 41.115 209.095 42.325 209.615 ;
        RECT 39.735 207.835 42.325 208.925 ;
        RECT 44.090 208.270 44.440 209.520 ;
        RECT 45.920 209.010 46.260 209.840 ;
        RECT 49.610 208.270 49.960 209.520 ;
        RECT 51.440 209.010 51.780 209.840 ;
        RECT 55.130 208.270 55.480 209.520 ;
        RECT 56.960 209.010 57.300 209.840 ;
        RECT 60.650 208.270 61.000 209.520 ;
        RECT 62.480 209.010 62.820 209.840 ;
        RECT 64.575 209.660 64.865 210.385 ;
        RECT 65.495 209.615 68.085 210.385 ;
        RECT 68.260 209.840 73.605 210.385 ;
        RECT 73.780 209.840 79.125 210.385 ;
        RECT 79.300 209.840 84.645 210.385 ;
        RECT 84.820 209.840 90.165 210.385 ;
        RECT 42.500 207.835 47.845 208.270 ;
        RECT 48.020 207.835 53.365 208.270 ;
        RECT 53.540 207.835 58.885 208.270 ;
        RECT 59.060 207.835 64.405 208.270 ;
        RECT 64.575 207.835 64.865 209.000 ;
        RECT 65.495 208.925 66.705 209.445 ;
        RECT 66.875 209.095 68.085 209.615 ;
        RECT 65.495 207.835 68.085 208.925 ;
        RECT 69.850 208.270 70.200 209.520 ;
        RECT 71.680 209.010 72.020 209.840 ;
        RECT 75.370 208.270 75.720 209.520 ;
        RECT 77.200 209.010 77.540 209.840 ;
        RECT 80.890 208.270 81.240 209.520 ;
        RECT 82.720 209.010 83.060 209.840 ;
        RECT 86.410 208.270 86.760 209.520 ;
        RECT 88.240 209.010 88.580 209.840 ;
        RECT 90.335 209.660 90.625 210.385 ;
        RECT 91.255 209.615 93.845 210.385 ;
        RECT 94.020 209.840 99.365 210.385 ;
        RECT 99.540 209.840 104.885 210.385 ;
        RECT 105.060 209.840 110.405 210.385 ;
        RECT 110.580 209.840 115.925 210.385 ;
        RECT 68.260 207.835 73.605 208.270 ;
        RECT 73.780 207.835 79.125 208.270 ;
        RECT 79.300 207.835 84.645 208.270 ;
        RECT 84.820 207.835 90.165 208.270 ;
        RECT 90.335 207.835 90.625 209.000 ;
        RECT 91.255 208.925 92.465 209.445 ;
        RECT 92.635 209.095 93.845 209.615 ;
        RECT 91.255 207.835 93.845 208.925 ;
        RECT 95.610 208.270 95.960 209.520 ;
        RECT 97.440 209.010 97.780 209.840 ;
        RECT 101.130 208.270 101.480 209.520 ;
        RECT 102.960 209.010 103.300 209.840 ;
        RECT 106.650 208.270 107.000 209.520 ;
        RECT 108.480 209.010 108.820 209.840 ;
        RECT 112.170 208.270 112.520 209.520 ;
        RECT 114.000 209.010 114.340 209.840 ;
        RECT 116.095 209.660 116.385 210.385 ;
        RECT 117.020 209.840 122.365 210.385 ;
        RECT 122.540 209.840 127.885 210.385 ;
        RECT 94.020 207.835 99.365 208.270 ;
        RECT 99.540 207.835 104.885 208.270 ;
        RECT 105.060 207.835 110.405 208.270 ;
        RECT 110.580 207.835 115.925 208.270 ;
        RECT 116.095 207.835 116.385 209.000 ;
        RECT 118.610 208.270 118.960 209.520 ;
        RECT 120.440 209.010 120.780 209.840 ;
        RECT 124.130 208.270 124.480 209.520 ;
        RECT 125.960 209.010 126.300 209.840 ;
        RECT 128.055 209.635 129.265 210.385 ;
        RECT 128.055 208.925 128.575 209.465 ;
        RECT 128.745 209.095 129.265 209.635 ;
        RECT 117.020 207.835 122.365 208.270 ;
        RECT 122.540 207.835 127.885 208.270 ;
        RECT 128.055 207.835 129.265 208.925 ;
        RECT 9.290 207.665 129.350 207.835 ;
        RECT 9.375 206.575 10.585 207.665 ;
        RECT 9.375 205.865 9.895 206.405 ;
        RECT 10.065 206.035 10.585 206.575 ;
        RECT 11.215 206.575 14.725 207.665 ;
        RECT 14.900 207.230 20.245 207.665 ;
        RECT 20.420 207.230 25.765 207.665 ;
        RECT 11.215 206.055 12.905 206.575 ;
        RECT 13.075 205.885 14.725 206.405 ;
        RECT 16.490 205.980 16.840 207.230 ;
        RECT 9.375 205.115 10.585 205.865 ;
        RECT 11.215 205.115 14.725 205.885 ;
        RECT 18.320 205.660 18.660 206.490 ;
        RECT 22.010 205.980 22.360 207.230 ;
        RECT 25.935 206.500 26.225 207.665 ;
        RECT 26.855 206.575 29.445 207.665 ;
        RECT 29.620 207.230 34.965 207.665 ;
        RECT 35.140 207.230 40.485 207.665 ;
        RECT 40.660 207.230 46.005 207.665 ;
        RECT 46.180 207.230 51.525 207.665 ;
        RECT 23.840 205.660 24.180 206.490 ;
        RECT 26.855 206.055 28.065 206.575 ;
        RECT 28.235 205.885 29.445 206.405 ;
        RECT 31.210 205.980 31.560 207.230 ;
        RECT 14.900 205.115 20.245 205.660 ;
        RECT 20.420 205.115 25.765 205.660 ;
        RECT 25.935 205.115 26.225 205.840 ;
        RECT 26.855 205.115 29.445 205.885 ;
        RECT 33.040 205.660 33.380 206.490 ;
        RECT 36.730 205.980 37.080 207.230 ;
        RECT 38.560 205.660 38.900 206.490 ;
        RECT 42.250 205.980 42.600 207.230 ;
        RECT 44.080 205.660 44.420 206.490 ;
        RECT 47.770 205.980 48.120 207.230 ;
        RECT 51.695 206.500 51.985 207.665 ;
        RECT 52.615 206.575 55.205 207.665 ;
        RECT 55.380 207.230 60.725 207.665 ;
        RECT 60.900 207.230 66.245 207.665 ;
        RECT 66.420 207.230 71.765 207.665 ;
        RECT 71.940 207.230 77.285 207.665 ;
        RECT 49.600 205.660 49.940 206.490 ;
        RECT 52.615 206.055 53.825 206.575 ;
        RECT 53.995 205.885 55.205 206.405 ;
        RECT 56.970 205.980 57.320 207.230 ;
        RECT 29.620 205.115 34.965 205.660 ;
        RECT 35.140 205.115 40.485 205.660 ;
        RECT 40.660 205.115 46.005 205.660 ;
        RECT 46.180 205.115 51.525 205.660 ;
        RECT 51.695 205.115 51.985 205.840 ;
        RECT 52.615 205.115 55.205 205.885 ;
        RECT 58.800 205.660 59.140 206.490 ;
        RECT 62.490 205.980 62.840 207.230 ;
        RECT 64.320 205.660 64.660 206.490 ;
        RECT 68.010 205.980 68.360 207.230 ;
        RECT 69.840 205.660 70.180 206.490 ;
        RECT 73.530 205.980 73.880 207.230 ;
        RECT 77.455 206.500 77.745 207.665 ;
        RECT 78.375 206.575 80.965 207.665 ;
        RECT 81.140 207.230 86.485 207.665 ;
        RECT 86.660 207.230 92.005 207.665 ;
        RECT 92.180 207.230 97.525 207.665 ;
        RECT 97.700 207.230 103.045 207.665 ;
        RECT 75.360 205.660 75.700 206.490 ;
        RECT 78.375 206.055 79.585 206.575 ;
        RECT 79.755 205.885 80.965 206.405 ;
        RECT 82.730 205.980 83.080 207.230 ;
        RECT 55.380 205.115 60.725 205.660 ;
        RECT 60.900 205.115 66.245 205.660 ;
        RECT 66.420 205.115 71.765 205.660 ;
        RECT 71.940 205.115 77.285 205.660 ;
        RECT 77.455 205.115 77.745 205.840 ;
        RECT 78.375 205.115 80.965 205.885 ;
        RECT 84.560 205.660 84.900 206.490 ;
        RECT 88.250 205.980 88.600 207.230 ;
        RECT 90.080 205.660 90.420 206.490 ;
        RECT 93.770 205.980 94.120 207.230 ;
        RECT 95.600 205.660 95.940 206.490 ;
        RECT 99.290 205.980 99.640 207.230 ;
        RECT 103.215 206.500 103.505 207.665 ;
        RECT 104.135 206.575 105.805 207.665 ;
        RECT 105.980 207.230 111.325 207.665 ;
        RECT 111.500 207.230 116.845 207.665 ;
        RECT 117.020 207.230 122.365 207.665 ;
        RECT 122.540 207.230 127.885 207.665 ;
        RECT 101.120 205.660 101.460 206.490 ;
        RECT 104.135 206.055 104.885 206.575 ;
        RECT 105.055 205.885 105.805 206.405 ;
        RECT 107.570 205.980 107.920 207.230 ;
        RECT 81.140 205.115 86.485 205.660 ;
        RECT 86.660 205.115 92.005 205.660 ;
        RECT 92.180 205.115 97.525 205.660 ;
        RECT 97.700 205.115 103.045 205.660 ;
        RECT 103.215 205.115 103.505 205.840 ;
        RECT 104.135 205.115 105.805 205.885 ;
        RECT 109.400 205.660 109.740 206.490 ;
        RECT 113.090 205.980 113.440 207.230 ;
        RECT 114.920 205.660 115.260 206.490 ;
        RECT 118.610 205.980 118.960 207.230 ;
        RECT 120.440 205.660 120.780 206.490 ;
        RECT 124.130 205.980 124.480 207.230 ;
        RECT 128.055 206.575 129.265 207.665 ;
        RECT 125.960 205.660 126.300 206.490 ;
        RECT 128.055 206.035 128.575 206.575 ;
        RECT 128.745 205.865 129.265 206.405 ;
        RECT 105.980 205.115 111.325 205.660 ;
        RECT 111.500 205.115 116.845 205.660 ;
        RECT 117.020 205.115 122.365 205.660 ;
        RECT 122.540 205.115 127.885 205.660 ;
        RECT 128.055 205.115 129.265 205.865 ;
        RECT 9.290 204.945 129.350 205.115 ;
        RECT 9.375 204.195 10.585 204.945 ;
        RECT 9.375 203.655 9.895 204.195 ;
        RECT 11.215 204.175 12.885 204.945 ;
        RECT 13.055 204.220 13.345 204.945 ;
        RECT 13.975 204.175 16.565 204.945 ;
        RECT 16.740 204.400 22.085 204.945 ;
        RECT 22.260 204.400 27.605 204.945 ;
        RECT 27.780 204.400 33.125 204.945 ;
        RECT 33.300 204.400 38.645 204.945 ;
        RECT 10.065 203.485 10.585 204.025 ;
        RECT 9.375 202.395 10.585 203.485 ;
        RECT 11.215 203.485 11.965 204.005 ;
        RECT 12.135 203.655 12.885 204.175 ;
        RECT 11.215 202.395 12.885 203.485 ;
        RECT 13.055 202.395 13.345 203.560 ;
        RECT 13.975 203.485 15.185 204.005 ;
        RECT 15.355 203.655 16.565 204.175 ;
        RECT 13.975 202.395 16.565 203.485 ;
        RECT 18.330 202.830 18.680 204.080 ;
        RECT 20.160 203.570 20.500 204.400 ;
        RECT 23.850 202.830 24.200 204.080 ;
        RECT 25.680 203.570 26.020 204.400 ;
        RECT 29.370 202.830 29.720 204.080 ;
        RECT 31.200 203.570 31.540 204.400 ;
        RECT 34.890 202.830 35.240 204.080 ;
        RECT 36.720 203.570 37.060 204.400 ;
        RECT 38.815 204.220 39.105 204.945 ;
        RECT 39.735 204.175 42.325 204.945 ;
        RECT 42.500 204.400 47.845 204.945 ;
        RECT 48.020 204.400 53.365 204.945 ;
        RECT 53.540 204.400 58.885 204.945 ;
        RECT 59.060 204.400 64.405 204.945 ;
        RECT 16.740 202.395 22.085 202.830 ;
        RECT 22.260 202.395 27.605 202.830 ;
        RECT 27.780 202.395 33.125 202.830 ;
        RECT 33.300 202.395 38.645 202.830 ;
        RECT 38.815 202.395 39.105 203.560 ;
        RECT 39.735 203.485 40.945 204.005 ;
        RECT 41.115 203.655 42.325 204.175 ;
        RECT 39.735 202.395 42.325 203.485 ;
        RECT 44.090 202.830 44.440 204.080 ;
        RECT 45.920 203.570 46.260 204.400 ;
        RECT 49.610 202.830 49.960 204.080 ;
        RECT 51.440 203.570 51.780 204.400 ;
        RECT 55.130 202.830 55.480 204.080 ;
        RECT 56.960 203.570 57.300 204.400 ;
        RECT 60.650 202.830 61.000 204.080 ;
        RECT 62.480 203.570 62.820 204.400 ;
        RECT 64.575 204.220 64.865 204.945 ;
        RECT 65.495 204.175 68.085 204.945 ;
        RECT 68.260 204.400 73.605 204.945 ;
        RECT 73.780 204.400 79.125 204.945 ;
        RECT 79.300 204.400 84.645 204.945 ;
        RECT 84.820 204.400 90.165 204.945 ;
        RECT 42.500 202.395 47.845 202.830 ;
        RECT 48.020 202.395 53.365 202.830 ;
        RECT 53.540 202.395 58.885 202.830 ;
        RECT 59.060 202.395 64.405 202.830 ;
        RECT 64.575 202.395 64.865 203.560 ;
        RECT 65.495 203.485 66.705 204.005 ;
        RECT 66.875 203.655 68.085 204.175 ;
        RECT 65.495 202.395 68.085 203.485 ;
        RECT 69.850 202.830 70.200 204.080 ;
        RECT 71.680 203.570 72.020 204.400 ;
        RECT 75.370 202.830 75.720 204.080 ;
        RECT 77.200 203.570 77.540 204.400 ;
        RECT 80.890 202.830 81.240 204.080 ;
        RECT 82.720 203.570 83.060 204.400 ;
        RECT 86.410 202.830 86.760 204.080 ;
        RECT 88.240 203.570 88.580 204.400 ;
        RECT 90.335 204.220 90.625 204.945 ;
        RECT 91.255 204.175 93.845 204.945 ;
        RECT 94.020 204.400 99.365 204.945 ;
        RECT 99.540 204.400 104.885 204.945 ;
        RECT 105.060 204.400 110.405 204.945 ;
        RECT 110.580 204.400 115.925 204.945 ;
        RECT 68.260 202.395 73.605 202.830 ;
        RECT 73.780 202.395 79.125 202.830 ;
        RECT 79.300 202.395 84.645 202.830 ;
        RECT 84.820 202.395 90.165 202.830 ;
        RECT 90.335 202.395 90.625 203.560 ;
        RECT 91.255 203.485 92.465 204.005 ;
        RECT 92.635 203.655 93.845 204.175 ;
        RECT 91.255 202.395 93.845 203.485 ;
        RECT 95.610 202.830 95.960 204.080 ;
        RECT 97.440 203.570 97.780 204.400 ;
        RECT 101.130 202.830 101.480 204.080 ;
        RECT 102.960 203.570 103.300 204.400 ;
        RECT 106.650 202.830 107.000 204.080 ;
        RECT 108.480 203.570 108.820 204.400 ;
        RECT 112.170 202.830 112.520 204.080 ;
        RECT 114.000 203.570 114.340 204.400 ;
        RECT 116.095 204.220 116.385 204.945 ;
        RECT 117.020 204.400 122.365 204.945 ;
        RECT 122.540 204.400 127.885 204.945 ;
        RECT 94.020 202.395 99.365 202.830 ;
        RECT 99.540 202.395 104.885 202.830 ;
        RECT 105.060 202.395 110.405 202.830 ;
        RECT 110.580 202.395 115.925 202.830 ;
        RECT 116.095 202.395 116.385 203.560 ;
        RECT 118.610 202.830 118.960 204.080 ;
        RECT 120.440 203.570 120.780 204.400 ;
        RECT 124.130 202.830 124.480 204.080 ;
        RECT 125.960 203.570 126.300 204.400 ;
        RECT 128.055 204.195 129.265 204.945 ;
        RECT 128.055 203.485 128.575 204.025 ;
        RECT 128.745 203.655 129.265 204.195 ;
        RECT 117.020 202.395 122.365 202.830 ;
        RECT 122.540 202.395 127.885 202.830 ;
        RECT 128.055 202.395 129.265 203.485 ;
        RECT 9.290 202.225 129.350 202.395 ;
        RECT 9.375 201.135 10.585 202.225 ;
        RECT 9.375 200.425 9.895 200.965 ;
        RECT 10.065 200.595 10.585 201.135 ;
        RECT 11.215 201.135 14.725 202.225 ;
        RECT 14.900 201.790 20.245 202.225 ;
        RECT 20.420 201.790 25.765 202.225 ;
        RECT 11.215 200.615 12.905 201.135 ;
        RECT 13.075 200.445 14.725 200.965 ;
        RECT 16.490 200.540 16.840 201.790 ;
        RECT 9.375 199.675 10.585 200.425 ;
        RECT 11.215 199.675 14.725 200.445 ;
        RECT 18.320 200.220 18.660 201.050 ;
        RECT 22.010 200.540 22.360 201.790 ;
        RECT 25.935 201.060 26.225 202.225 ;
        RECT 26.855 201.135 29.445 202.225 ;
        RECT 29.620 201.790 34.965 202.225 ;
        RECT 35.140 201.790 40.485 202.225 ;
        RECT 40.660 201.790 46.005 202.225 ;
        RECT 46.180 201.790 51.525 202.225 ;
        RECT 23.840 200.220 24.180 201.050 ;
        RECT 26.855 200.615 28.065 201.135 ;
        RECT 28.235 200.445 29.445 200.965 ;
        RECT 31.210 200.540 31.560 201.790 ;
        RECT 14.900 199.675 20.245 200.220 ;
        RECT 20.420 199.675 25.765 200.220 ;
        RECT 25.935 199.675 26.225 200.400 ;
        RECT 26.855 199.675 29.445 200.445 ;
        RECT 33.040 200.220 33.380 201.050 ;
        RECT 36.730 200.540 37.080 201.790 ;
        RECT 38.560 200.220 38.900 201.050 ;
        RECT 42.250 200.540 42.600 201.790 ;
        RECT 44.080 200.220 44.420 201.050 ;
        RECT 47.770 200.540 48.120 201.790 ;
        RECT 51.695 201.060 51.985 202.225 ;
        RECT 52.615 201.135 55.205 202.225 ;
        RECT 55.380 201.790 60.725 202.225 ;
        RECT 60.900 201.790 66.245 202.225 ;
        RECT 66.420 201.790 71.765 202.225 ;
        RECT 71.940 201.790 77.285 202.225 ;
        RECT 49.600 200.220 49.940 201.050 ;
        RECT 52.615 200.615 53.825 201.135 ;
        RECT 53.995 200.445 55.205 200.965 ;
        RECT 56.970 200.540 57.320 201.790 ;
        RECT 29.620 199.675 34.965 200.220 ;
        RECT 35.140 199.675 40.485 200.220 ;
        RECT 40.660 199.675 46.005 200.220 ;
        RECT 46.180 199.675 51.525 200.220 ;
        RECT 51.695 199.675 51.985 200.400 ;
        RECT 52.615 199.675 55.205 200.445 ;
        RECT 58.800 200.220 59.140 201.050 ;
        RECT 62.490 200.540 62.840 201.790 ;
        RECT 64.320 200.220 64.660 201.050 ;
        RECT 68.010 200.540 68.360 201.790 ;
        RECT 69.840 200.220 70.180 201.050 ;
        RECT 73.530 200.540 73.880 201.790 ;
        RECT 77.455 201.060 77.745 202.225 ;
        RECT 78.375 201.135 80.965 202.225 ;
        RECT 81.140 201.790 86.485 202.225 ;
        RECT 86.660 201.790 92.005 202.225 ;
        RECT 92.180 201.790 97.525 202.225 ;
        RECT 97.700 201.790 103.045 202.225 ;
        RECT 75.360 200.220 75.700 201.050 ;
        RECT 78.375 200.615 79.585 201.135 ;
        RECT 79.755 200.445 80.965 200.965 ;
        RECT 82.730 200.540 83.080 201.790 ;
        RECT 55.380 199.675 60.725 200.220 ;
        RECT 60.900 199.675 66.245 200.220 ;
        RECT 66.420 199.675 71.765 200.220 ;
        RECT 71.940 199.675 77.285 200.220 ;
        RECT 77.455 199.675 77.745 200.400 ;
        RECT 78.375 199.675 80.965 200.445 ;
        RECT 84.560 200.220 84.900 201.050 ;
        RECT 88.250 200.540 88.600 201.790 ;
        RECT 90.080 200.220 90.420 201.050 ;
        RECT 93.770 200.540 94.120 201.790 ;
        RECT 95.600 200.220 95.940 201.050 ;
        RECT 99.290 200.540 99.640 201.790 ;
        RECT 103.215 201.060 103.505 202.225 ;
        RECT 104.135 201.135 105.805 202.225 ;
        RECT 105.980 201.790 111.325 202.225 ;
        RECT 111.500 201.790 116.845 202.225 ;
        RECT 117.020 201.790 122.365 202.225 ;
        RECT 122.540 201.790 127.885 202.225 ;
        RECT 101.120 200.220 101.460 201.050 ;
        RECT 104.135 200.615 104.885 201.135 ;
        RECT 105.055 200.445 105.805 200.965 ;
        RECT 107.570 200.540 107.920 201.790 ;
        RECT 81.140 199.675 86.485 200.220 ;
        RECT 86.660 199.675 92.005 200.220 ;
        RECT 92.180 199.675 97.525 200.220 ;
        RECT 97.700 199.675 103.045 200.220 ;
        RECT 103.215 199.675 103.505 200.400 ;
        RECT 104.135 199.675 105.805 200.445 ;
        RECT 109.400 200.220 109.740 201.050 ;
        RECT 113.090 200.540 113.440 201.790 ;
        RECT 114.920 200.220 115.260 201.050 ;
        RECT 118.610 200.540 118.960 201.790 ;
        RECT 120.440 200.220 120.780 201.050 ;
        RECT 124.130 200.540 124.480 201.790 ;
        RECT 128.055 201.135 129.265 202.225 ;
        RECT 125.960 200.220 126.300 201.050 ;
        RECT 128.055 200.595 128.575 201.135 ;
        RECT 128.745 200.425 129.265 200.965 ;
        RECT 105.980 199.675 111.325 200.220 ;
        RECT 111.500 199.675 116.845 200.220 ;
        RECT 117.020 199.675 122.365 200.220 ;
        RECT 122.540 199.675 127.885 200.220 ;
        RECT 128.055 199.675 129.265 200.425 ;
        RECT 9.290 199.505 129.350 199.675 ;
        RECT 9.375 198.755 10.585 199.505 ;
        RECT 9.375 198.215 9.895 198.755 ;
        RECT 11.215 198.735 12.885 199.505 ;
        RECT 13.055 198.780 13.345 199.505 ;
        RECT 13.975 198.735 16.565 199.505 ;
        RECT 16.740 198.960 22.085 199.505 ;
        RECT 22.260 198.960 27.605 199.505 ;
        RECT 27.780 198.960 33.125 199.505 ;
        RECT 33.300 198.960 38.645 199.505 ;
        RECT 10.065 198.045 10.585 198.585 ;
        RECT 9.375 196.955 10.585 198.045 ;
        RECT 11.215 198.045 11.965 198.565 ;
        RECT 12.135 198.215 12.885 198.735 ;
        RECT 11.215 196.955 12.885 198.045 ;
        RECT 13.055 196.955 13.345 198.120 ;
        RECT 13.975 198.045 15.185 198.565 ;
        RECT 15.355 198.215 16.565 198.735 ;
        RECT 13.975 196.955 16.565 198.045 ;
        RECT 18.330 197.390 18.680 198.640 ;
        RECT 20.160 198.130 20.500 198.960 ;
        RECT 23.850 197.390 24.200 198.640 ;
        RECT 25.680 198.130 26.020 198.960 ;
        RECT 29.370 197.390 29.720 198.640 ;
        RECT 31.200 198.130 31.540 198.960 ;
        RECT 34.890 197.390 35.240 198.640 ;
        RECT 36.720 198.130 37.060 198.960 ;
        RECT 38.815 198.780 39.105 199.505 ;
        RECT 40.195 198.735 43.705 199.505 ;
        RECT 43.880 198.960 49.225 199.505 ;
        RECT 49.400 198.960 54.745 199.505 ;
        RECT 16.740 196.955 22.085 197.390 ;
        RECT 22.260 196.955 27.605 197.390 ;
        RECT 27.780 196.955 33.125 197.390 ;
        RECT 33.300 196.955 38.645 197.390 ;
        RECT 38.815 196.955 39.105 198.120 ;
        RECT 40.195 198.045 41.885 198.565 ;
        RECT 42.055 198.215 43.705 198.735 ;
        RECT 40.195 196.955 43.705 198.045 ;
        RECT 45.470 197.390 45.820 198.640 ;
        RECT 47.300 198.130 47.640 198.960 ;
        RECT 50.990 197.390 51.340 198.640 ;
        RECT 52.820 198.130 53.160 198.960 ;
        RECT 54.920 198.955 55.175 199.245 ;
        RECT 55.345 199.125 55.675 199.505 ;
        RECT 54.920 198.785 55.670 198.955 ;
        RECT 54.920 197.965 55.270 198.615 ;
        RECT 55.440 197.795 55.670 198.785 ;
        RECT 54.920 197.625 55.670 197.795 ;
        RECT 43.880 196.955 49.225 197.390 ;
        RECT 49.400 196.955 54.745 197.390 ;
        RECT 54.920 197.125 55.175 197.625 ;
        RECT 55.345 196.955 55.675 197.455 ;
        RECT 55.845 197.125 56.015 199.245 ;
        RECT 56.375 199.145 56.705 199.505 ;
        RECT 56.875 199.115 57.370 199.285 ;
        RECT 57.575 199.115 58.430 199.285 ;
        RECT 56.245 197.925 56.705 198.975 ;
        RECT 56.185 197.140 56.510 197.925 ;
        RECT 56.875 197.755 57.045 199.115 ;
        RECT 57.215 198.205 57.565 198.825 ;
        RECT 57.735 198.605 58.090 198.825 ;
        RECT 57.735 198.015 57.905 198.605 ;
        RECT 58.260 198.405 58.430 199.115 ;
        RECT 59.305 199.045 59.635 199.505 ;
        RECT 59.845 199.145 60.195 199.315 ;
        RECT 58.635 198.575 59.425 198.825 ;
        RECT 59.845 198.755 60.105 199.145 ;
        RECT 60.415 199.055 61.365 199.335 ;
        RECT 61.535 199.065 61.725 199.505 ;
        RECT 61.895 199.125 62.965 199.295 ;
        RECT 59.595 198.405 59.765 198.585 ;
        RECT 56.875 197.585 57.270 197.755 ;
        RECT 57.440 197.625 57.905 198.015 ;
        RECT 58.075 198.235 59.765 198.405 ;
        RECT 57.100 197.455 57.270 197.585 ;
        RECT 58.075 197.455 58.245 198.235 ;
        RECT 59.935 198.065 60.105 198.755 ;
        RECT 58.605 197.895 60.105 198.065 ;
        RECT 60.295 198.095 60.505 198.885 ;
        RECT 60.675 198.265 61.025 198.885 ;
        RECT 61.195 198.275 61.365 199.055 ;
        RECT 61.895 198.895 62.065 199.125 ;
        RECT 61.535 198.725 62.065 198.895 ;
        RECT 61.535 198.445 61.755 198.725 ;
        RECT 62.235 198.555 62.475 198.955 ;
        RECT 61.195 198.105 61.600 198.275 ;
        RECT 61.935 198.185 62.475 198.555 ;
        RECT 62.645 198.770 62.965 199.125 ;
        RECT 63.210 199.045 63.515 199.505 ;
        RECT 63.685 198.795 63.935 199.325 ;
        RECT 62.645 198.595 62.970 198.770 ;
        RECT 62.645 198.295 63.560 198.595 ;
        RECT 62.820 198.265 63.560 198.295 ;
        RECT 60.295 197.935 60.970 198.095 ;
        RECT 61.430 198.015 61.600 198.105 ;
        RECT 60.295 197.925 61.260 197.935 ;
        RECT 59.935 197.755 60.105 197.895 ;
        RECT 56.680 196.955 56.930 197.415 ;
        RECT 57.100 197.125 57.350 197.455 ;
        RECT 57.565 197.125 58.245 197.455 ;
        RECT 58.415 197.555 59.490 197.725 ;
        RECT 59.935 197.585 60.495 197.755 ;
        RECT 60.800 197.635 61.260 197.925 ;
        RECT 61.430 197.845 62.650 198.015 ;
        RECT 58.415 197.215 58.585 197.555 ;
        RECT 58.820 196.955 59.150 197.385 ;
        RECT 59.320 197.215 59.490 197.555 ;
        RECT 59.785 196.955 60.155 197.415 ;
        RECT 60.325 197.125 60.495 197.585 ;
        RECT 61.430 197.465 61.600 197.845 ;
        RECT 62.820 197.675 62.990 198.265 ;
        RECT 63.730 198.145 63.935 198.795 ;
        RECT 64.105 198.750 64.355 199.505 ;
        RECT 64.575 198.780 64.865 199.505 ;
        RECT 65.095 198.685 65.305 199.505 ;
        RECT 65.475 198.705 65.805 199.335 ;
        RECT 60.730 197.125 61.600 197.465 ;
        RECT 62.190 197.505 62.990 197.675 ;
        RECT 61.770 196.955 62.020 197.415 ;
        RECT 62.190 197.215 62.360 197.505 ;
        RECT 62.540 196.955 62.870 197.335 ;
        RECT 63.210 196.955 63.515 198.095 ;
        RECT 63.685 197.265 63.935 198.145 ;
        RECT 64.105 196.955 64.355 198.095 ;
        RECT 64.575 196.955 64.865 198.120 ;
        RECT 65.475 198.105 65.725 198.705 ;
        RECT 65.975 198.685 66.205 199.505 ;
        RECT 66.875 198.765 67.195 199.245 ;
        RECT 67.365 198.935 67.595 199.335 ;
        RECT 67.765 199.115 68.115 199.505 ;
        RECT 67.365 198.855 67.875 198.935 ;
        RECT 68.285 198.855 68.615 199.335 ;
        RECT 67.365 198.765 68.615 198.855 ;
        RECT 65.895 198.265 66.225 198.515 ;
        RECT 65.095 196.955 65.305 198.095 ;
        RECT 65.475 197.125 65.805 198.105 ;
        RECT 65.975 196.955 66.205 198.095 ;
        RECT 66.875 197.835 67.045 198.765 ;
        RECT 67.705 198.685 68.615 198.765 ;
        RECT 68.785 198.685 68.955 199.505 ;
        RECT 69.460 198.765 69.925 199.310 ;
        RECT 67.215 198.175 67.385 198.595 ;
        RECT 67.615 198.345 68.215 198.515 ;
        RECT 67.215 198.005 67.875 198.175 ;
        RECT 66.875 197.635 67.535 197.835 ;
        RECT 67.705 197.805 67.875 198.005 ;
        RECT 68.045 198.145 68.215 198.345 ;
        RECT 68.385 198.315 69.080 198.515 ;
        RECT 69.340 198.145 69.585 198.595 ;
        RECT 68.045 197.975 69.585 198.145 ;
        RECT 69.755 197.805 69.925 198.765 ;
        RECT 70.095 198.735 73.605 199.505 ;
        RECT 73.780 198.960 79.125 199.505 ;
        RECT 79.300 198.960 84.645 199.505 ;
        RECT 84.820 198.960 90.165 199.505 ;
        RECT 67.705 197.635 69.925 197.805 ;
        RECT 70.095 198.045 71.785 198.565 ;
        RECT 71.955 198.215 73.605 198.735 ;
        RECT 67.365 197.465 67.535 197.635 ;
        RECT 66.895 196.955 67.195 197.465 ;
        RECT 67.365 197.295 67.745 197.465 ;
        RECT 68.325 196.955 68.955 197.465 ;
        RECT 69.125 197.125 69.455 197.635 ;
        RECT 69.625 196.955 69.925 197.465 ;
        RECT 70.095 196.955 73.605 198.045 ;
        RECT 75.370 197.390 75.720 198.640 ;
        RECT 77.200 198.130 77.540 198.960 ;
        RECT 80.890 197.390 81.240 198.640 ;
        RECT 82.720 198.130 83.060 198.960 ;
        RECT 86.410 197.390 86.760 198.640 ;
        RECT 88.240 198.130 88.580 198.960 ;
        RECT 90.335 198.780 90.625 199.505 ;
        RECT 90.795 198.735 92.465 199.505 ;
        RECT 92.640 198.960 97.985 199.505 ;
        RECT 73.780 196.955 79.125 197.390 ;
        RECT 79.300 196.955 84.645 197.390 ;
        RECT 84.820 196.955 90.165 197.390 ;
        RECT 90.335 196.955 90.625 198.120 ;
        RECT 90.795 198.045 91.545 198.565 ;
        RECT 91.715 198.215 92.465 198.735 ;
        RECT 90.795 196.955 92.465 198.045 ;
        RECT 94.230 197.390 94.580 198.640 ;
        RECT 96.060 198.130 96.400 198.960 ;
        RECT 98.215 198.685 98.425 199.505 ;
        RECT 98.595 198.705 98.925 199.335 ;
        RECT 98.595 198.105 98.845 198.705 ;
        RECT 99.095 198.685 99.325 199.505 ;
        RECT 100.545 198.955 100.715 199.335 ;
        RECT 100.895 199.125 101.225 199.505 ;
        RECT 100.545 198.785 101.210 198.955 ;
        RECT 101.405 198.830 101.665 199.335 ;
        RECT 99.015 198.265 99.345 198.515 ;
        RECT 100.475 198.235 100.805 198.605 ;
        RECT 101.040 198.530 101.210 198.785 ;
        RECT 101.040 198.200 101.325 198.530 ;
        RECT 92.640 196.955 97.985 197.390 ;
        RECT 98.215 196.955 98.425 198.095 ;
        RECT 98.595 197.125 98.925 198.105 ;
        RECT 99.095 196.955 99.325 198.095 ;
        RECT 101.040 198.055 101.210 198.200 ;
        RECT 100.545 197.885 101.210 198.055 ;
        RECT 101.495 198.030 101.665 198.830 ;
        RECT 101.835 198.755 103.045 199.505 ;
        RECT 103.220 198.960 108.565 199.505 ;
        RECT 108.740 198.960 114.085 199.505 ;
        RECT 100.545 197.125 100.715 197.885 ;
        RECT 100.895 196.955 101.225 197.715 ;
        RECT 101.395 197.125 101.665 198.030 ;
        RECT 101.835 198.045 102.355 198.585 ;
        RECT 102.525 198.215 103.045 198.755 ;
        RECT 101.835 196.955 103.045 198.045 ;
        RECT 104.810 197.390 105.160 198.640 ;
        RECT 106.640 198.130 106.980 198.960 ;
        RECT 110.330 197.390 110.680 198.640 ;
        RECT 112.160 198.130 112.500 198.960 ;
        RECT 114.315 198.685 114.525 199.505 ;
        RECT 114.695 198.705 115.025 199.335 ;
        RECT 114.695 198.105 114.945 198.705 ;
        RECT 115.195 198.685 115.425 199.505 ;
        RECT 116.095 198.780 116.385 199.505 ;
        RECT 117.020 198.960 122.365 199.505 ;
        RECT 122.540 198.960 127.885 199.505 ;
        RECT 115.115 198.265 115.445 198.515 ;
        RECT 103.220 196.955 108.565 197.390 ;
        RECT 108.740 196.955 114.085 197.390 ;
        RECT 114.315 196.955 114.525 198.095 ;
        RECT 114.695 197.125 115.025 198.105 ;
        RECT 115.195 196.955 115.425 198.095 ;
        RECT 116.095 196.955 116.385 198.120 ;
        RECT 118.610 197.390 118.960 198.640 ;
        RECT 120.440 198.130 120.780 198.960 ;
        RECT 124.130 197.390 124.480 198.640 ;
        RECT 125.960 198.130 126.300 198.960 ;
        RECT 128.055 198.755 129.265 199.505 ;
        RECT 128.055 198.045 128.575 198.585 ;
        RECT 128.745 198.215 129.265 198.755 ;
        RECT 117.020 196.955 122.365 197.390 ;
        RECT 122.540 196.955 127.885 197.390 ;
        RECT 128.055 196.955 129.265 198.045 ;
        RECT 9.290 196.785 129.350 196.955 ;
        RECT 9.375 195.695 10.585 196.785 ;
        RECT 9.375 194.985 9.895 195.525 ;
        RECT 10.065 195.155 10.585 195.695 ;
        RECT 11.215 195.695 14.725 196.785 ;
        RECT 14.900 196.350 20.245 196.785 ;
        RECT 20.420 196.350 25.765 196.785 ;
        RECT 11.215 195.175 12.905 195.695 ;
        RECT 13.075 195.005 14.725 195.525 ;
        RECT 16.490 195.100 16.840 196.350 ;
        RECT 9.375 194.235 10.585 194.985 ;
        RECT 11.215 194.235 14.725 195.005 ;
        RECT 18.320 194.780 18.660 195.610 ;
        RECT 22.010 195.100 22.360 196.350 ;
        RECT 25.935 195.620 26.225 196.785 ;
        RECT 26.860 196.350 32.205 196.785 ;
        RECT 32.380 196.350 37.725 196.785 ;
        RECT 37.900 196.350 43.245 196.785 ;
        RECT 23.840 194.780 24.180 195.610 ;
        RECT 28.450 195.100 28.800 196.350 ;
        RECT 14.900 194.235 20.245 194.780 ;
        RECT 20.420 194.235 25.765 194.780 ;
        RECT 25.935 194.235 26.225 194.960 ;
        RECT 30.280 194.780 30.620 195.610 ;
        RECT 33.970 195.100 34.320 196.350 ;
        RECT 35.800 194.780 36.140 195.610 ;
        RECT 39.490 195.100 39.840 196.350 ;
        RECT 43.415 195.710 43.685 196.615 ;
        RECT 43.855 196.025 44.185 196.785 ;
        RECT 44.365 195.855 44.535 196.615 ;
        RECT 41.320 194.780 41.660 195.610 ;
        RECT 43.415 194.910 43.585 195.710 ;
        RECT 43.870 195.685 44.535 195.855 ;
        RECT 43.870 195.540 44.040 195.685 ;
        RECT 45.775 195.645 45.985 196.785 ;
        RECT 43.755 195.210 44.040 195.540 ;
        RECT 46.155 195.635 46.485 196.615 ;
        RECT 46.655 195.645 46.885 196.785 ;
        RECT 47.555 195.695 50.145 196.785 ;
        RECT 43.870 194.955 44.040 195.210 ;
        RECT 44.275 195.135 44.605 195.505 ;
        RECT 26.860 194.235 32.205 194.780 ;
        RECT 32.380 194.235 37.725 194.780 ;
        RECT 37.900 194.235 43.245 194.780 ;
        RECT 43.415 194.405 43.675 194.910 ;
        RECT 43.870 194.785 44.535 194.955 ;
        RECT 43.855 194.235 44.185 194.615 ;
        RECT 44.365 194.405 44.535 194.785 ;
        RECT 45.775 194.235 45.985 195.055 ;
        RECT 46.155 195.035 46.405 195.635 ;
        RECT 46.575 195.225 46.905 195.475 ;
        RECT 47.555 195.175 48.765 195.695 ;
        RECT 50.355 195.645 50.585 196.785 ;
        RECT 50.755 195.635 51.085 196.615 ;
        RECT 51.255 195.645 51.465 196.785 ;
        RECT 46.155 194.405 46.485 195.035 ;
        RECT 46.655 194.235 46.885 195.055 ;
        RECT 48.935 195.005 50.145 195.525 ;
        RECT 50.335 195.225 50.665 195.475 ;
        RECT 47.555 194.235 50.145 195.005 ;
        RECT 50.355 194.235 50.585 195.055 ;
        RECT 50.835 195.035 51.085 195.635 ;
        RECT 51.695 195.620 51.985 196.785 ;
        RECT 52.155 195.695 53.825 196.785 ;
        RECT 54.085 195.855 54.255 196.615 ;
        RECT 54.435 196.025 54.765 196.785 ;
        RECT 52.155 195.175 52.905 195.695 ;
        RECT 54.085 195.685 54.750 195.855 ;
        RECT 54.935 195.710 55.205 196.615 ;
        RECT 54.580 195.540 54.750 195.685 ;
        RECT 50.755 194.405 51.085 195.035 ;
        RECT 51.255 194.235 51.465 195.055 ;
        RECT 53.075 195.005 53.825 195.525 ;
        RECT 54.015 195.135 54.345 195.505 ;
        RECT 54.580 195.210 54.865 195.540 ;
        RECT 51.695 194.235 51.985 194.960 ;
        RECT 52.155 194.235 53.825 195.005 ;
        RECT 54.580 194.955 54.750 195.210 ;
        RECT 54.085 194.785 54.750 194.955 ;
        RECT 55.035 194.910 55.205 195.710 ;
        RECT 55.375 195.695 56.585 196.785 ;
        RECT 56.760 196.115 57.015 196.615 ;
        RECT 57.185 196.285 57.515 196.785 ;
        RECT 56.760 195.945 57.510 196.115 ;
        RECT 55.375 195.155 55.895 195.695 ;
        RECT 56.065 194.985 56.585 195.525 ;
        RECT 56.760 195.125 57.110 195.775 ;
        RECT 54.085 194.405 54.255 194.785 ;
        RECT 54.435 194.235 54.765 194.615 ;
        RECT 54.945 194.405 55.205 194.910 ;
        RECT 55.375 194.235 56.585 194.985 ;
        RECT 57.280 194.955 57.510 195.945 ;
        RECT 56.760 194.785 57.510 194.955 ;
        RECT 56.760 194.495 57.015 194.785 ;
        RECT 57.185 194.235 57.515 194.615 ;
        RECT 57.685 194.495 57.855 196.615 ;
        RECT 58.025 195.815 58.350 196.600 ;
        RECT 58.520 196.325 58.770 196.785 ;
        RECT 58.940 196.285 59.190 196.615 ;
        RECT 59.405 196.285 60.085 196.615 ;
        RECT 58.940 196.155 59.110 196.285 ;
        RECT 58.715 195.985 59.110 196.155 ;
        RECT 58.085 194.765 58.545 195.815 ;
        RECT 58.715 194.625 58.885 195.985 ;
        RECT 59.280 195.725 59.745 196.115 ;
        RECT 59.055 194.915 59.405 195.535 ;
        RECT 59.575 195.135 59.745 195.725 ;
        RECT 59.915 195.505 60.085 196.285 ;
        RECT 60.255 196.185 60.425 196.525 ;
        RECT 60.660 196.355 60.990 196.785 ;
        RECT 61.160 196.185 61.330 196.525 ;
        RECT 61.625 196.325 61.995 196.785 ;
        RECT 60.255 196.015 61.330 196.185 ;
        RECT 62.165 196.155 62.335 196.615 ;
        RECT 62.570 196.275 63.440 196.615 ;
        RECT 63.610 196.325 63.860 196.785 ;
        RECT 61.775 195.985 62.335 196.155 ;
        RECT 61.775 195.845 61.945 195.985 ;
        RECT 60.445 195.675 61.945 195.845 ;
        RECT 62.640 195.815 63.100 196.105 ;
        RECT 59.915 195.335 61.605 195.505 ;
        RECT 59.575 194.915 59.930 195.135 ;
        RECT 60.100 194.625 60.270 195.335 ;
        RECT 60.475 194.915 61.265 195.165 ;
        RECT 61.435 195.155 61.605 195.335 ;
        RECT 61.775 194.985 61.945 195.675 ;
        RECT 58.215 194.235 58.545 194.595 ;
        RECT 58.715 194.455 59.210 194.625 ;
        RECT 59.415 194.455 60.270 194.625 ;
        RECT 61.145 194.235 61.475 194.695 ;
        RECT 61.685 194.595 61.945 194.985 ;
        RECT 62.135 195.805 63.100 195.815 ;
        RECT 63.270 195.895 63.440 196.275 ;
        RECT 64.030 196.235 64.200 196.525 ;
        RECT 64.380 196.405 64.710 196.785 ;
        RECT 64.030 196.065 64.830 196.235 ;
        RECT 62.135 195.645 62.810 195.805 ;
        RECT 63.270 195.725 64.490 195.895 ;
        RECT 62.135 194.855 62.345 195.645 ;
        RECT 63.270 195.635 63.440 195.725 ;
        RECT 62.515 194.855 62.865 195.475 ;
        RECT 63.035 195.465 63.440 195.635 ;
        RECT 63.035 194.685 63.205 195.465 ;
        RECT 63.375 195.015 63.595 195.295 ;
        RECT 63.775 195.185 64.315 195.555 ;
        RECT 64.660 195.445 64.830 196.065 ;
        RECT 65.005 195.725 65.175 196.785 ;
        RECT 65.385 195.775 65.675 196.615 ;
        RECT 65.845 195.945 66.015 196.785 ;
        RECT 66.225 195.775 66.475 196.615 ;
        RECT 66.685 195.945 66.855 196.785 ;
        RECT 65.385 195.605 67.110 195.775 ;
        RECT 63.375 194.845 63.905 195.015 ;
        RECT 61.685 194.425 62.035 194.595 ;
        RECT 62.255 194.405 63.205 194.685 ;
        RECT 63.375 194.235 63.565 194.675 ;
        RECT 63.735 194.615 63.905 194.845 ;
        RECT 64.075 194.785 64.315 195.185 ;
        RECT 64.485 195.435 64.830 195.445 ;
        RECT 64.485 195.225 66.515 195.435 ;
        RECT 64.485 194.970 64.810 195.225 ;
        RECT 66.700 195.055 67.110 195.605 ;
        RECT 64.485 194.615 64.805 194.970 ;
        RECT 63.735 194.445 64.805 194.615 ;
        RECT 65.005 194.235 65.175 195.045 ;
        RECT 65.345 194.885 67.110 195.055 ;
        RECT 67.335 195.710 67.605 196.615 ;
        RECT 67.775 196.025 68.105 196.785 ;
        RECT 68.285 195.855 68.455 196.615 ;
        RECT 67.335 194.910 67.505 195.710 ;
        RECT 67.790 195.685 68.455 195.855 ;
        RECT 69.175 195.695 72.685 196.785 ;
        RECT 67.790 195.540 67.960 195.685 ;
        RECT 67.675 195.210 67.960 195.540 ;
        RECT 67.790 194.955 67.960 195.210 ;
        RECT 68.195 195.135 68.525 195.505 ;
        RECT 69.175 195.175 70.865 195.695 ;
        RECT 72.895 195.645 73.125 196.785 ;
        RECT 73.295 195.635 73.625 196.615 ;
        RECT 73.795 195.645 74.005 196.785 ;
        RECT 74.235 196.275 74.535 196.785 ;
        RECT 74.705 196.105 75.035 196.615 ;
        RECT 75.205 196.275 75.835 196.785 ;
        RECT 76.415 196.275 76.795 196.445 ;
        RECT 76.965 196.275 77.265 196.785 ;
        RECT 76.625 196.105 76.795 196.275 ;
        RECT 74.235 195.935 76.455 196.105 ;
        RECT 71.035 195.005 72.685 195.525 ;
        RECT 72.875 195.225 73.205 195.475 ;
        RECT 65.345 194.405 65.675 194.885 ;
        RECT 65.845 194.235 66.015 194.705 ;
        RECT 66.185 194.405 66.515 194.885 ;
        RECT 66.685 194.235 66.855 194.705 ;
        RECT 67.335 194.405 67.595 194.910 ;
        RECT 67.790 194.785 68.455 194.955 ;
        RECT 67.775 194.235 68.105 194.615 ;
        RECT 68.285 194.405 68.455 194.785 ;
        RECT 69.175 194.235 72.685 195.005 ;
        RECT 72.895 194.235 73.125 195.055 ;
        RECT 73.375 195.035 73.625 195.635 ;
        RECT 73.295 194.405 73.625 195.035 ;
        RECT 73.795 194.235 74.005 195.055 ;
        RECT 74.235 194.975 74.405 195.935 ;
        RECT 74.575 195.595 76.115 195.765 ;
        RECT 74.575 195.145 74.820 195.595 ;
        RECT 75.080 195.225 75.775 195.425 ;
        RECT 75.945 195.395 76.115 195.595 ;
        RECT 76.285 195.735 76.455 195.935 ;
        RECT 76.625 195.905 77.285 196.105 ;
        RECT 76.285 195.565 76.945 195.735 ;
        RECT 75.945 195.225 76.545 195.395 ;
        RECT 76.775 195.145 76.945 195.565 ;
        RECT 74.235 194.430 74.700 194.975 ;
        RECT 75.205 194.235 75.375 195.055 ;
        RECT 75.545 194.975 76.455 195.055 ;
        RECT 77.115 194.975 77.285 195.905 ;
        RECT 77.455 195.620 77.745 196.785 ;
        RECT 78.380 196.350 83.725 196.785 ;
        RECT 84.270 196.445 84.525 196.475 ;
        RECT 79.970 195.100 80.320 196.350 ;
        RECT 84.185 196.275 84.525 196.445 ;
        RECT 84.270 195.805 84.525 196.275 ;
        RECT 84.705 195.985 84.990 196.785 ;
        RECT 85.170 196.065 85.500 196.575 ;
        RECT 75.545 194.885 76.795 194.975 ;
        RECT 75.545 194.405 75.875 194.885 ;
        RECT 76.285 194.805 76.795 194.885 ;
        RECT 76.045 194.235 76.395 194.625 ;
        RECT 76.565 194.405 76.795 194.805 ;
        RECT 76.965 194.495 77.285 194.975 ;
        RECT 77.455 194.235 77.745 194.960 ;
        RECT 81.800 194.780 82.140 195.610 ;
        RECT 84.270 194.945 84.450 195.805 ;
        RECT 85.170 195.475 85.420 196.065 ;
        RECT 85.770 195.915 85.940 196.525 ;
        RECT 86.110 196.095 86.440 196.785 ;
        RECT 86.670 196.235 86.910 196.525 ;
        RECT 87.110 196.405 87.530 196.785 ;
        RECT 87.710 196.315 88.340 196.565 ;
        RECT 88.810 196.405 89.140 196.785 ;
        RECT 87.710 196.235 87.880 196.315 ;
        RECT 89.310 196.235 89.480 196.525 ;
        RECT 89.660 196.405 90.040 196.785 ;
        RECT 90.280 196.400 91.110 196.570 ;
        RECT 86.670 196.065 87.880 196.235 ;
        RECT 84.620 195.145 85.420 195.475 ;
        RECT 78.380 194.235 83.725 194.780 ;
        RECT 84.270 194.415 84.525 194.945 ;
        RECT 84.705 194.235 84.990 194.695 ;
        RECT 85.170 194.495 85.420 195.145 ;
        RECT 85.620 195.895 85.940 195.915 ;
        RECT 85.620 195.725 87.540 195.895 ;
        RECT 85.620 194.830 85.810 195.725 ;
        RECT 87.710 195.555 87.880 196.065 ;
        RECT 88.050 195.805 88.570 196.115 ;
        RECT 85.980 195.385 87.880 195.555 ;
        RECT 85.980 195.325 86.310 195.385 ;
        RECT 86.460 195.155 86.790 195.215 ;
        RECT 86.130 194.885 86.790 195.155 ;
        RECT 85.620 194.500 85.940 194.830 ;
        RECT 86.120 194.235 86.780 194.715 ;
        RECT 86.980 194.625 87.150 195.385 ;
        RECT 88.050 195.215 88.230 195.625 ;
        RECT 87.320 195.045 87.650 195.165 ;
        RECT 88.400 195.045 88.570 195.805 ;
        RECT 87.320 194.875 88.570 195.045 ;
        RECT 88.740 195.985 90.110 196.235 ;
        RECT 88.740 195.215 88.930 195.985 ;
        RECT 89.860 195.725 90.110 195.985 ;
        RECT 89.100 195.555 89.350 195.715 ;
        RECT 90.280 195.555 90.450 196.400 ;
        RECT 91.345 196.115 91.515 196.615 ;
        RECT 91.685 196.285 92.015 196.785 ;
        RECT 90.620 195.725 91.120 196.105 ;
        RECT 91.345 195.945 92.040 196.115 ;
        RECT 89.100 195.385 90.450 195.555 ;
        RECT 90.030 195.345 90.450 195.385 ;
        RECT 88.740 194.875 89.160 195.215 ;
        RECT 89.450 194.885 89.860 195.215 ;
        RECT 86.980 194.455 87.830 194.625 ;
        RECT 88.390 194.235 88.710 194.695 ;
        RECT 88.910 194.445 89.160 194.875 ;
        RECT 89.450 194.235 89.860 194.675 ;
        RECT 90.030 194.615 90.200 195.345 ;
        RECT 90.370 194.795 90.720 195.165 ;
        RECT 90.900 194.855 91.120 195.725 ;
        RECT 91.290 195.155 91.700 195.775 ;
        RECT 91.870 194.975 92.040 195.945 ;
        RECT 91.345 194.785 92.040 194.975 ;
        RECT 90.030 194.415 91.045 194.615 ;
        RECT 91.345 194.455 91.515 194.785 ;
        RECT 91.685 194.235 92.015 194.615 ;
        RECT 92.230 194.495 92.455 196.615 ;
        RECT 92.625 196.285 92.955 196.785 ;
        RECT 93.125 196.115 93.295 196.615 ;
        RECT 92.630 195.945 93.295 196.115 ;
        RECT 92.630 194.955 92.860 195.945 ;
        RECT 93.030 195.125 93.380 195.775 ;
        RECT 94.020 195.595 94.275 196.475 ;
        RECT 94.445 195.645 94.750 196.785 ;
        RECT 95.090 196.405 95.420 196.785 ;
        RECT 95.600 196.235 95.770 196.525 ;
        RECT 95.940 196.325 96.190 196.785 ;
        RECT 94.970 196.065 95.770 196.235 ;
        RECT 96.360 196.275 97.230 196.615 ;
        RECT 92.630 194.785 93.295 194.955 ;
        RECT 92.625 194.235 92.955 194.615 ;
        RECT 93.125 194.495 93.295 194.785 ;
        RECT 94.020 194.945 94.230 195.595 ;
        RECT 94.970 195.475 95.140 196.065 ;
        RECT 96.360 195.895 96.530 196.275 ;
        RECT 97.465 196.155 97.635 196.615 ;
        RECT 97.805 196.325 98.175 196.785 ;
        RECT 98.470 196.185 98.640 196.525 ;
        RECT 98.810 196.355 99.140 196.785 ;
        RECT 99.375 196.185 99.545 196.525 ;
        RECT 95.310 195.725 96.530 195.895 ;
        RECT 96.700 195.815 97.160 196.105 ;
        RECT 97.465 195.985 98.025 196.155 ;
        RECT 98.470 196.015 99.545 196.185 ;
        RECT 99.715 196.285 100.395 196.615 ;
        RECT 100.610 196.285 100.860 196.615 ;
        RECT 101.030 196.325 101.280 196.785 ;
        RECT 97.855 195.845 98.025 195.985 ;
        RECT 96.700 195.805 97.665 195.815 ;
        RECT 96.360 195.635 96.530 195.725 ;
        RECT 96.990 195.645 97.665 195.805 ;
        RECT 94.400 195.445 95.140 195.475 ;
        RECT 94.400 195.145 95.315 195.445 ;
        RECT 94.990 194.970 95.315 195.145 ;
        RECT 94.020 194.415 94.275 194.945 ;
        RECT 94.445 194.235 94.750 194.695 ;
        RECT 94.995 194.615 95.315 194.970 ;
        RECT 95.485 195.185 96.025 195.555 ;
        RECT 96.360 195.465 96.765 195.635 ;
        RECT 95.485 194.785 95.725 195.185 ;
        RECT 96.205 195.015 96.425 195.295 ;
        RECT 95.895 194.845 96.425 195.015 ;
        RECT 95.895 194.615 96.065 194.845 ;
        RECT 96.595 194.685 96.765 195.465 ;
        RECT 96.935 194.855 97.285 195.475 ;
        RECT 97.455 194.855 97.665 195.645 ;
        RECT 97.855 195.675 99.355 195.845 ;
        RECT 97.855 194.985 98.025 195.675 ;
        RECT 99.715 195.505 99.885 196.285 ;
        RECT 100.690 196.155 100.860 196.285 ;
        RECT 98.195 195.335 99.885 195.505 ;
        RECT 100.055 195.725 100.520 196.115 ;
        RECT 100.690 195.985 101.085 196.155 ;
        RECT 98.195 195.155 98.365 195.335 ;
        RECT 94.995 194.445 96.065 194.615 ;
        RECT 96.235 194.235 96.425 194.675 ;
        RECT 96.595 194.405 97.545 194.685 ;
        RECT 97.855 194.595 98.115 194.985 ;
        RECT 98.535 194.915 99.325 195.165 ;
        RECT 97.765 194.425 98.115 194.595 ;
        RECT 98.325 194.235 98.655 194.695 ;
        RECT 99.530 194.625 99.700 195.335 ;
        RECT 100.055 195.135 100.225 195.725 ;
        RECT 99.870 194.915 100.225 195.135 ;
        RECT 100.395 194.915 100.745 195.535 ;
        RECT 100.915 194.625 101.085 195.985 ;
        RECT 101.450 195.815 101.775 196.600 ;
        RECT 101.255 194.765 101.715 195.815 ;
        RECT 99.530 194.455 100.385 194.625 ;
        RECT 100.590 194.455 101.085 194.625 ;
        RECT 101.255 194.235 101.585 194.595 ;
        RECT 101.945 194.495 102.115 196.615 ;
        RECT 102.285 196.285 102.615 196.785 ;
        RECT 102.785 196.115 103.040 196.615 ;
        RECT 102.290 195.945 103.040 196.115 ;
        RECT 102.290 194.955 102.520 195.945 ;
        RECT 102.690 195.125 103.040 195.775 ;
        RECT 103.215 195.620 103.505 196.785 ;
        RECT 104.600 196.350 109.945 196.785 ;
        RECT 106.190 195.100 106.540 196.350 ;
        RECT 110.175 195.645 110.385 196.785 ;
        RECT 110.555 195.635 110.885 196.615 ;
        RECT 111.055 195.645 111.285 196.785 ;
        RECT 102.290 194.785 103.040 194.955 ;
        RECT 102.285 194.235 102.615 194.615 ;
        RECT 102.785 194.495 103.040 194.785 ;
        RECT 103.215 194.235 103.505 194.960 ;
        RECT 108.020 194.780 108.360 195.610 ;
        RECT 104.600 194.235 109.945 194.780 ;
        RECT 110.175 194.235 110.385 195.055 ;
        RECT 110.555 195.035 110.805 195.635 ;
        RECT 111.500 195.595 111.755 196.475 ;
        RECT 111.925 195.645 112.230 196.785 ;
        RECT 112.570 196.405 112.900 196.785 ;
        RECT 113.080 196.235 113.250 196.525 ;
        RECT 113.420 196.325 113.670 196.785 ;
        RECT 112.450 196.065 113.250 196.235 ;
        RECT 113.840 196.275 114.710 196.615 ;
        RECT 110.975 195.225 111.305 195.475 ;
        RECT 110.555 194.405 110.885 195.035 ;
        RECT 111.055 194.235 111.285 195.055 ;
        RECT 111.500 194.945 111.710 195.595 ;
        RECT 112.450 195.475 112.620 196.065 ;
        RECT 113.840 195.895 114.010 196.275 ;
        RECT 114.945 196.155 115.115 196.615 ;
        RECT 115.285 196.325 115.655 196.785 ;
        RECT 115.950 196.185 116.120 196.525 ;
        RECT 116.290 196.355 116.620 196.785 ;
        RECT 116.855 196.185 117.025 196.525 ;
        RECT 112.790 195.725 114.010 195.895 ;
        RECT 114.180 195.815 114.640 196.105 ;
        RECT 114.945 195.985 115.505 196.155 ;
        RECT 115.950 196.015 117.025 196.185 ;
        RECT 117.195 196.285 117.875 196.615 ;
        RECT 118.090 196.285 118.340 196.615 ;
        RECT 118.510 196.325 118.760 196.785 ;
        RECT 115.335 195.845 115.505 195.985 ;
        RECT 114.180 195.805 115.145 195.815 ;
        RECT 113.840 195.635 114.010 195.725 ;
        RECT 114.470 195.645 115.145 195.805 ;
        RECT 111.880 195.445 112.620 195.475 ;
        RECT 111.880 195.145 112.795 195.445 ;
        RECT 112.470 194.970 112.795 195.145 ;
        RECT 111.500 194.415 111.755 194.945 ;
        RECT 111.925 194.235 112.230 194.695 ;
        RECT 112.475 194.615 112.795 194.970 ;
        RECT 112.965 195.185 113.505 195.555 ;
        RECT 113.840 195.465 114.245 195.635 ;
        RECT 112.965 194.785 113.205 195.185 ;
        RECT 113.685 195.015 113.905 195.295 ;
        RECT 113.375 194.845 113.905 195.015 ;
        RECT 113.375 194.615 113.545 194.845 ;
        RECT 114.075 194.685 114.245 195.465 ;
        RECT 114.415 194.855 114.765 195.475 ;
        RECT 114.935 194.855 115.145 195.645 ;
        RECT 115.335 195.675 116.835 195.845 ;
        RECT 115.335 194.985 115.505 195.675 ;
        RECT 117.195 195.505 117.365 196.285 ;
        RECT 118.170 196.155 118.340 196.285 ;
        RECT 115.675 195.335 117.365 195.505 ;
        RECT 117.535 195.725 118.000 196.115 ;
        RECT 118.170 195.985 118.565 196.155 ;
        RECT 115.675 195.155 115.845 195.335 ;
        RECT 112.475 194.445 113.545 194.615 ;
        RECT 113.715 194.235 113.905 194.675 ;
        RECT 114.075 194.405 115.025 194.685 ;
        RECT 115.335 194.595 115.595 194.985 ;
        RECT 116.015 194.915 116.805 195.165 ;
        RECT 115.245 194.425 115.595 194.595 ;
        RECT 115.805 194.235 116.135 194.695 ;
        RECT 117.010 194.625 117.180 195.335 ;
        RECT 117.535 195.135 117.705 195.725 ;
        RECT 117.350 194.915 117.705 195.135 ;
        RECT 117.875 194.915 118.225 195.535 ;
        RECT 118.395 194.625 118.565 195.985 ;
        RECT 118.930 195.815 119.255 196.600 ;
        RECT 118.735 194.765 119.195 195.815 ;
        RECT 117.010 194.455 117.865 194.625 ;
        RECT 118.070 194.455 118.565 194.625 ;
        RECT 118.735 194.235 119.065 194.595 ;
        RECT 119.425 194.495 119.595 196.615 ;
        RECT 119.765 196.285 120.095 196.785 ;
        RECT 120.265 196.115 120.520 196.615 ;
        RECT 119.770 195.945 120.520 196.115 ;
        RECT 119.770 194.955 120.000 195.945 ;
        RECT 120.170 195.125 120.520 195.775 ;
        RECT 120.695 195.695 122.365 196.785 ;
        RECT 122.540 196.350 127.885 196.785 ;
        RECT 120.695 195.175 121.445 195.695 ;
        RECT 121.615 195.005 122.365 195.525 ;
        RECT 124.130 195.100 124.480 196.350 ;
        RECT 128.055 195.695 129.265 196.785 ;
        RECT 119.770 194.785 120.520 194.955 ;
        RECT 119.765 194.235 120.095 194.615 ;
        RECT 120.265 194.495 120.520 194.785 ;
        RECT 120.695 194.235 122.365 195.005 ;
        RECT 125.960 194.780 126.300 195.610 ;
        RECT 128.055 195.155 128.575 195.695 ;
        RECT 128.745 194.985 129.265 195.525 ;
        RECT 122.540 194.235 127.885 194.780 ;
        RECT 128.055 194.235 129.265 194.985 ;
        RECT 9.290 194.065 129.350 194.235 ;
        RECT 9.375 193.315 10.585 194.065 ;
        RECT 9.375 192.775 9.895 193.315 ;
        RECT 11.215 193.295 12.885 194.065 ;
        RECT 13.055 193.340 13.345 194.065 ;
        RECT 14.435 193.295 17.945 194.065 ;
        RECT 18.120 193.520 23.465 194.065 ;
        RECT 23.640 193.520 28.985 194.065 ;
        RECT 29.160 193.520 34.505 194.065 ;
        RECT 10.065 192.605 10.585 193.145 ;
        RECT 9.375 191.515 10.585 192.605 ;
        RECT 11.215 192.605 11.965 193.125 ;
        RECT 12.135 192.775 12.885 193.295 ;
        RECT 11.215 191.515 12.885 192.605 ;
        RECT 13.055 191.515 13.345 192.680 ;
        RECT 14.435 192.605 16.125 193.125 ;
        RECT 16.295 192.775 17.945 193.295 ;
        RECT 14.435 191.515 17.945 192.605 ;
        RECT 19.710 191.950 20.060 193.200 ;
        RECT 21.540 192.690 21.880 193.520 ;
        RECT 25.230 191.950 25.580 193.200 ;
        RECT 27.060 192.690 27.400 193.520 ;
        RECT 30.750 191.950 31.100 193.200 ;
        RECT 32.580 192.690 32.920 193.520 ;
        RECT 34.950 193.255 35.195 193.860 ;
        RECT 35.415 193.530 35.925 194.065 ;
        RECT 34.675 193.085 35.905 193.255 ;
        RECT 34.675 192.275 35.015 193.085 ;
        RECT 35.185 192.520 35.935 192.710 ;
        RECT 18.120 191.515 23.465 191.950 ;
        RECT 23.640 191.515 28.985 191.950 ;
        RECT 29.160 191.515 34.505 191.950 ;
        RECT 34.675 191.865 35.190 192.275 ;
        RECT 35.425 191.515 35.595 192.275 ;
        RECT 35.765 191.855 35.935 192.520 ;
        RECT 36.105 192.535 36.295 193.895 ;
        RECT 36.465 193.045 36.740 193.895 ;
        RECT 36.930 193.530 37.460 193.895 ;
        RECT 37.885 193.665 38.215 194.065 ;
        RECT 37.285 193.495 37.460 193.530 ;
        RECT 36.465 192.875 36.745 193.045 ;
        RECT 36.465 192.735 36.740 192.875 ;
        RECT 36.945 192.535 37.115 193.335 ;
        RECT 36.105 192.365 37.115 192.535 ;
        RECT 37.285 193.325 38.215 193.495 ;
        RECT 38.385 193.325 38.640 193.895 ;
        RECT 38.815 193.340 39.105 194.065 ;
        RECT 39.280 193.515 39.535 193.805 ;
        RECT 39.705 193.685 40.035 194.065 ;
        RECT 39.280 193.345 40.030 193.515 ;
        RECT 37.285 192.195 37.455 193.325 ;
        RECT 38.045 193.155 38.215 193.325 ;
        RECT 36.330 192.025 37.455 192.195 ;
        RECT 37.625 192.825 37.820 193.155 ;
        RECT 38.045 192.825 38.300 193.155 ;
        RECT 37.625 191.855 37.795 192.825 ;
        RECT 38.470 192.655 38.640 193.325 ;
        RECT 35.765 191.685 37.795 191.855 ;
        RECT 37.965 191.515 38.135 192.655 ;
        RECT 38.305 191.685 38.640 192.655 ;
        RECT 38.815 191.515 39.105 192.680 ;
        RECT 39.280 192.525 39.630 193.175 ;
        RECT 39.800 192.355 40.030 193.345 ;
        RECT 39.280 192.185 40.030 192.355 ;
        RECT 39.280 191.685 39.535 192.185 ;
        RECT 39.705 191.515 40.035 192.015 ;
        RECT 40.205 191.685 40.375 193.805 ;
        RECT 40.735 193.705 41.065 194.065 ;
        RECT 41.235 193.675 41.730 193.845 ;
        RECT 41.935 193.675 42.790 193.845 ;
        RECT 40.605 192.485 41.065 193.535 ;
        RECT 40.545 191.700 40.870 192.485 ;
        RECT 41.235 192.315 41.405 193.675 ;
        RECT 41.575 192.765 41.925 193.385 ;
        RECT 42.095 193.165 42.450 193.385 ;
        RECT 42.095 192.575 42.265 193.165 ;
        RECT 42.620 192.965 42.790 193.675 ;
        RECT 43.665 193.605 43.995 194.065 ;
        RECT 44.205 193.705 44.555 193.875 ;
        RECT 42.995 193.135 43.785 193.385 ;
        RECT 44.205 193.315 44.465 193.705 ;
        RECT 44.775 193.615 45.725 193.895 ;
        RECT 45.895 193.625 46.085 194.065 ;
        RECT 46.255 193.685 47.325 193.855 ;
        RECT 43.955 192.965 44.125 193.145 ;
        RECT 41.235 192.145 41.630 192.315 ;
        RECT 41.800 192.185 42.265 192.575 ;
        RECT 42.435 192.795 44.125 192.965 ;
        RECT 41.460 192.015 41.630 192.145 ;
        RECT 42.435 192.015 42.605 192.795 ;
        RECT 44.295 192.625 44.465 193.315 ;
        RECT 42.965 192.455 44.465 192.625 ;
        RECT 44.655 192.655 44.865 193.445 ;
        RECT 45.035 192.825 45.385 193.445 ;
        RECT 45.555 192.835 45.725 193.615 ;
        RECT 46.255 193.455 46.425 193.685 ;
        RECT 45.895 193.285 46.425 193.455 ;
        RECT 45.895 193.005 46.115 193.285 ;
        RECT 46.595 193.115 46.835 193.515 ;
        RECT 45.555 192.665 45.960 192.835 ;
        RECT 46.295 192.745 46.835 193.115 ;
        RECT 47.005 193.330 47.325 193.685 ;
        RECT 47.570 193.605 47.875 194.065 ;
        RECT 48.045 193.355 48.300 193.885 ;
        RECT 47.005 193.155 47.330 193.330 ;
        RECT 47.005 192.855 47.920 193.155 ;
        RECT 47.180 192.825 47.920 192.855 ;
        RECT 44.655 192.495 45.330 192.655 ;
        RECT 45.790 192.575 45.960 192.665 ;
        RECT 44.655 192.485 45.620 192.495 ;
        RECT 44.295 192.315 44.465 192.455 ;
        RECT 41.040 191.515 41.290 191.975 ;
        RECT 41.460 191.685 41.710 192.015 ;
        RECT 41.925 191.685 42.605 192.015 ;
        RECT 42.775 192.115 43.850 192.285 ;
        RECT 44.295 192.145 44.855 192.315 ;
        RECT 45.160 192.195 45.620 192.485 ;
        RECT 45.790 192.405 47.010 192.575 ;
        RECT 42.775 191.775 42.945 192.115 ;
        RECT 43.180 191.515 43.510 191.945 ;
        RECT 43.680 191.775 43.850 192.115 ;
        RECT 44.145 191.515 44.515 191.975 ;
        RECT 44.685 191.685 44.855 192.145 ;
        RECT 45.790 192.025 45.960 192.405 ;
        RECT 47.180 192.235 47.350 192.825 ;
        RECT 48.090 192.705 48.300 193.355 ;
        RECT 45.090 191.685 45.960 192.025 ;
        RECT 46.550 192.065 47.350 192.235 ;
        RECT 46.130 191.515 46.380 191.975 ;
        RECT 46.550 191.775 46.720 192.065 ;
        RECT 46.900 191.515 47.230 191.895 ;
        RECT 47.570 191.515 47.875 192.655 ;
        RECT 48.045 191.825 48.300 192.705 ;
        RECT 48.940 193.355 49.195 193.885 ;
        RECT 49.365 193.605 49.670 194.065 ;
        RECT 49.915 193.685 50.985 193.855 ;
        RECT 48.940 192.705 49.150 193.355 ;
        RECT 49.915 193.330 50.235 193.685 ;
        RECT 49.910 193.155 50.235 193.330 ;
        RECT 49.320 192.855 50.235 193.155 ;
        RECT 50.405 193.115 50.645 193.515 ;
        RECT 50.815 193.455 50.985 193.685 ;
        RECT 51.155 193.625 51.345 194.065 ;
        RECT 51.515 193.615 52.465 193.895 ;
        RECT 52.685 193.705 53.035 193.875 ;
        RECT 50.815 193.285 51.345 193.455 ;
        RECT 49.320 192.825 50.060 192.855 ;
        RECT 48.940 191.825 49.195 192.705 ;
        RECT 49.365 191.515 49.670 192.655 ;
        RECT 49.890 192.235 50.060 192.825 ;
        RECT 50.405 192.745 50.945 193.115 ;
        RECT 51.125 193.005 51.345 193.285 ;
        RECT 51.515 192.835 51.685 193.615 ;
        RECT 51.280 192.665 51.685 192.835 ;
        RECT 51.855 192.825 52.205 193.445 ;
        RECT 51.280 192.575 51.450 192.665 ;
        RECT 52.375 192.655 52.585 193.445 ;
        RECT 50.230 192.405 51.450 192.575 ;
        RECT 51.910 192.495 52.585 192.655 ;
        RECT 49.890 192.065 50.690 192.235 ;
        RECT 50.010 191.515 50.340 191.895 ;
        RECT 50.520 191.775 50.690 192.065 ;
        RECT 51.280 192.025 51.450 192.405 ;
        RECT 51.620 192.485 52.585 192.495 ;
        RECT 52.775 193.315 53.035 193.705 ;
        RECT 53.245 193.605 53.575 194.065 ;
        RECT 54.450 193.675 55.305 193.845 ;
        RECT 55.510 193.675 56.005 193.845 ;
        RECT 56.175 193.705 56.505 194.065 ;
        RECT 52.775 192.625 52.945 193.315 ;
        RECT 53.115 192.965 53.285 193.145 ;
        RECT 53.455 193.135 54.245 193.385 ;
        RECT 54.450 192.965 54.620 193.675 ;
        RECT 54.790 193.165 55.145 193.385 ;
        RECT 53.115 192.795 54.805 192.965 ;
        RECT 51.620 192.195 52.080 192.485 ;
        RECT 52.775 192.455 54.275 192.625 ;
        RECT 52.775 192.315 52.945 192.455 ;
        RECT 52.385 192.145 52.945 192.315 ;
        RECT 50.860 191.515 51.110 191.975 ;
        RECT 51.280 191.685 52.150 192.025 ;
        RECT 52.385 191.685 52.555 192.145 ;
        RECT 53.390 192.115 54.465 192.285 ;
        RECT 52.725 191.515 53.095 191.975 ;
        RECT 53.390 191.775 53.560 192.115 ;
        RECT 53.730 191.515 54.060 191.945 ;
        RECT 54.295 191.775 54.465 192.115 ;
        RECT 54.635 192.015 54.805 192.795 ;
        RECT 54.975 192.575 55.145 193.165 ;
        RECT 55.315 192.765 55.665 193.385 ;
        RECT 54.975 192.185 55.440 192.575 ;
        RECT 55.835 192.315 56.005 193.675 ;
        RECT 56.175 192.485 56.635 193.535 ;
        RECT 55.610 192.145 56.005 192.315 ;
        RECT 55.610 192.015 55.780 192.145 ;
        RECT 54.635 191.685 55.315 192.015 ;
        RECT 55.530 191.685 55.780 192.015 ;
        RECT 55.950 191.515 56.200 191.975 ;
        RECT 56.370 191.700 56.695 192.485 ;
        RECT 56.865 191.685 57.035 193.805 ;
        RECT 57.205 193.685 57.535 194.065 ;
        RECT 57.705 193.515 57.960 193.805 ;
        RECT 57.210 193.345 57.960 193.515 ;
        RECT 57.210 192.355 57.440 193.345 ;
        RECT 58.595 193.295 62.105 194.065 ;
        RECT 57.610 192.525 57.960 193.175 ;
        RECT 58.595 192.605 60.285 193.125 ;
        RECT 60.455 192.775 62.105 193.295 ;
        RECT 62.335 193.245 62.545 194.065 ;
        RECT 62.715 193.265 63.045 193.895 ;
        RECT 62.715 192.665 62.965 193.265 ;
        RECT 63.215 193.245 63.445 194.065 ;
        RECT 64.575 193.340 64.865 194.065 ;
        RECT 65.495 193.415 65.755 193.895 ;
        RECT 65.925 193.525 66.175 194.065 ;
        RECT 63.135 192.825 63.465 193.075 ;
        RECT 57.210 192.185 57.960 192.355 ;
        RECT 57.205 191.515 57.535 192.015 ;
        RECT 57.705 191.685 57.960 192.185 ;
        RECT 58.595 191.515 62.105 192.605 ;
        RECT 62.335 191.515 62.545 192.655 ;
        RECT 62.715 191.685 63.045 192.665 ;
        RECT 63.215 191.515 63.445 192.655 ;
        RECT 64.575 191.515 64.865 192.680 ;
        RECT 65.495 192.385 65.665 193.415 ;
        RECT 66.345 193.385 66.565 193.845 ;
        RECT 66.315 193.360 66.565 193.385 ;
        RECT 65.835 192.765 66.065 193.160 ;
        RECT 66.235 192.935 66.565 193.360 ;
        RECT 66.735 193.685 67.625 193.855 ;
        RECT 66.735 192.960 66.905 193.685 ;
        RECT 67.075 193.130 67.625 193.515 ;
        RECT 67.795 193.325 68.490 193.895 ;
        RECT 68.660 193.325 69.010 193.850 ;
        RECT 66.735 192.890 67.625 192.960 ;
        RECT 66.730 192.865 67.625 192.890 ;
        RECT 66.720 192.850 67.625 192.865 ;
        RECT 66.715 192.835 67.625 192.850 ;
        RECT 66.705 192.830 67.625 192.835 ;
        RECT 66.700 192.820 67.625 192.830 ;
        RECT 66.695 192.810 67.625 192.820 ;
        RECT 66.685 192.805 67.625 192.810 ;
        RECT 66.675 192.795 67.625 192.805 ;
        RECT 66.665 192.790 67.625 192.795 ;
        RECT 66.665 192.785 67.000 192.790 ;
        RECT 66.650 192.780 67.000 192.785 ;
        RECT 66.635 192.770 67.000 192.780 ;
        RECT 66.610 192.765 67.000 192.770 ;
        RECT 65.835 192.760 67.000 192.765 ;
        RECT 65.835 192.725 66.970 192.760 ;
        RECT 65.835 192.700 66.935 192.725 ;
        RECT 65.835 192.670 66.905 192.700 ;
        RECT 65.835 192.640 66.885 192.670 ;
        RECT 65.835 192.610 66.865 192.640 ;
        RECT 65.835 192.600 66.795 192.610 ;
        RECT 65.835 192.590 66.770 192.600 ;
        RECT 65.835 192.575 66.750 192.590 ;
        RECT 65.835 192.560 66.730 192.575 ;
        RECT 65.940 192.550 66.725 192.560 ;
        RECT 65.940 192.515 66.710 192.550 ;
        RECT 65.495 191.685 65.770 192.385 ;
        RECT 65.940 192.265 66.695 192.515 ;
        RECT 66.865 192.195 67.195 192.440 ;
        RECT 67.365 192.340 67.625 192.790 ;
        RECT 67.795 192.485 68.035 193.155 ;
        RECT 68.215 192.655 68.385 193.325 ;
        RECT 68.660 193.155 68.865 193.325 ;
        RECT 69.200 193.155 69.415 193.850 ;
        RECT 69.585 193.325 69.920 194.065 ;
        RECT 70.095 193.265 70.405 194.065 ;
        RECT 70.610 193.265 71.305 193.895 ;
        RECT 71.480 193.355 71.735 193.885 ;
        RECT 71.905 193.605 72.210 194.065 ;
        RECT 72.455 193.685 73.525 193.855 ;
        RECT 68.555 192.825 68.865 193.155 ;
        RECT 69.035 192.825 69.415 193.155 ;
        RECT 69.615 192.825 69.900 193.155 ;
        RECT 70.105 192.825 70.440 193.095 ;
        RECT 70.610 192.665 70.780 193.265 ;
        RECT 70.950 192.825 71.285 193.075 ;
        RECT 71.480 192.705 71.690 193.355 ;
        RECT 72.455 193.330 72.775 193.685 ;
        RECT 72.450 193.155 72.775 193.330 ;
        RECT 71.860 192.855 72.775 193.155 ;
        RECT 72.945 193.115 73.185 193.515 ;
        RECT 73.355 193.455 73.525 193.685 ;
        RECT 73.695 193.625 73.885 194.065 ;
        RECT 74.055 193.615 75.005 193.895 ;
        RECT 75.225 193.705 75.575 193.875 ;
        RECT 73.355 193.285 73.885 193.455 ;
        RECT 71.860 192.825 72.600 192.855 ;
        RECT 68.215 192.485 69.495 192.655 ;
        RECT 67.010 192.170 67.195 192.195 ;
        RECT 67.010 192.070 67.625 192.170 ;
        RECT 65.940 191.515 66.195 192.060 ;
        RECT 66.365 191.685 66.845 192.025 ;
        RECT 67.020 191.515 67.625 192.070 ;
        RECT 67.815 191.515 68.095 192.315 ;
        RECT 68.295 191.685 68.625 192.485 ;
        RECT 68.825 191.515 68.995 192.315 ;
        RECT 69.165 191.685 69.495 192.485 ;
        RECT 69.665 191.515 69.925 192.655 ;
        RECT 70.095 191.515 70.375 192.655 ;
        RECT 70.545 191.685 70.875 192.665 ;
        RECT 71.045 191.515 71.305 192.655 ;
        RECT 71.480 191.825 71.735 192.705 ;
        RECT 71.905 191.515 72.210 192.655 ;
        RECT 72.430 192.235 72.600 192.825 ;
        RECT 72.945 192.745 73.485 193.115 ;
        RECT 73.665 193.005 73.885 193.285 ;
        RECT 74.055 192.835 74.225 193.615 ;
        RECT 73.820 192.665 74.225 192.835 ;
        RECT 74.395 192.825 74.745 193.445 ;
        RECT 73.820 192.575 73.990 192.665 ;
        RECT 74.915 192.655 75.125 193.445 ;
        RECT 72.770 192.405 73.990 192.575 ;
        RECT 74.450 192.495 75.125 192.655 ;
        RECT 72.430 192.065 73.230 192.235 ;
        RECT 72.550 191.515 72.880 191.895 ;
        RECT 73.060 191.775 73.230 192.065 ;
        RECT 73.820 192.025 73.990 192.405 ;
        RECT 74.160 192.485 75.125 192.495 ;
        RECT 75.315 193.315 75.575 193.705 ;
        RECT 75.785 193.605 76.115 194.065 ;
        RECT 76.990 193.675 77.845 193.845 ;
        RECT 78.050 193.675 78.545 193.845 ;
        RECT 78.715 193.705 79.045 194.065 ;
        RECT 75.315 192.625 75.485 193.315 ;
        RECT 75.655 192.965 75.825 193.145 ;
        RECT 75.995 193.135 76.785 193.385 ;
        RECT 76.990 192.965 77.160 193.675 ;
        RECT 77.330 193.165 77.685 193.385 ;
        RECT 75.655 192.795 77.345 192.965 ;
        RECT 74.160 192.195 74.620 192.485 ;
        RECT 75.315 192.455 76.815 192.625 ;
        RECT 75.315 192.315 75.485 192.455 ;
        RECT 74.925 192.145 75.485 192.315 ;
        RECT 73.400 191.515 73.650 191.975 ;
        RECT 73.820 191.685 74.690 192.025 ;
        RECT 74.925 191.685 75.095 192.145 ;
        RECT 75.930 192.115 77.005 192.285 ;
        RECT 75.265 191.515 75.635 191.975 ;
        RECT 75.930 191.775 76.100 192.115 ;
        RECT 76.270 191.515 76.600 191.945 ;
        RECT 76.835 191.775 77.005 192.115 ;
        RECT 77.175 192.015 77.345 192.795 ;
        RECT 77.515 192.575 77.685 193.165 ;
        RECT 77.855 192.765 78.205 193.385 ;
        RECT 77.515 192.185 77.980 192.575 ;
        RECT 78.375 192.315 78.545 193.675 ;
        RECT 78.715 192.485 79.175 193.535 ;
        RECT 78.150 192.145 78.545 192.315 ;
        RECT 78.150 192.015 78.320 192.145 ;
        RECT 77.175 191.685 77.855 192.015 ;
        RECT 78.070 191.685 78.320 192.015 ;
        RECT 78.490 191.515 78.740 191.975 ;
        RECT 78.910 191.700 79.235 192.485 ;
        RECT 79.405 191.685 79.575 193.805 ;
        RECT 79.745 193.685 80.075 194.065 ;
        RECT 80.245 193.515 80.500 193.805 ;
        RECT 79.750 193.345 80.500 193.515 ;
        RECT 81.050 193.355 81.305 193.885 ;
        RECT 81.485 193.605 81.770 194.065 ;
        RECT 79.750 192.355 79.980 193.345 ;
        RECT 80.150 192.525 80.500 193.175 ;
        RECT 81.050 192.495 81.230 193.355 ;
        RECT 81.950 193.155 82.200 193.805 ;
        RECT 81.400 192.825 82.200 193.155 ;
        RECT 79.750 192.185 80.500 192.355 ;
        RECT 79.745 191.515 80.075 192.015 ;
        RECT 80.245 191.685 80.500 192.185 ;
        RECT 81.050 192.025 81.305 192.495 ;
        RECT 80.965 191.855 81.305 192.025 ;
        RECT 81.050 191.825 81.305 191.855 ;
        RECT 81.485 191.515 81.770 192.315 ;
        RECT 81.950 192.235 82.200 192.825 ;
        RECT 82.400 193.470 82.720 193.800 ;
        RECT 82.900 193.585 83.560 194.065 ;
        RECT 83.760 193.675 84.610 193.845 ;
        RECT 82.400 192.575 82.590 193.470 ;
        RECT 82.910 193.145 83.570 193.415 ;
        RECT 83.240 193.085 83.570 193.145 ;
        RECT 82.760 192.915 83.090 192.975 ;
        RECT 83.760 192.915 83.930 193.675 ;
        RECT 85.170 193.605 85.490 194.065 ;
        RECT 85.690 193.425 85.940 193.855 ;
        RECT 86.230 193.625 86.640 194.065 ;
        RECT 86.810 193.685 87.825 193.885 ;
        RECT 84.100 193.255 85.350 193.425 ;
        RECT 84.100 193.135 84.430 193.255 ;
        RECT 82.760 192.745 84.660 192.915 ;
        RECT 82.400 192.405 84.320 192.575 ;
        RECT 82.400 192.385 82.720 192.405 ;
        RECT 81.950 191.725 82.280 192.235 ;
        RECT 82.550 191.775 82.720 192.385 ;
        RECT 84.490 192.235 84.660 192.745 ;
        RECT 84.830 192.675 85.010 193.085 ;
        RECT 85.180 192.495 85.350 193.255 ;
        RECT 82.890 191.515 83.220 192.205 ;
        RECT 83.450 192.065 84.660 192.235 ;
        RECT 84.830 192.185 85.350 192.495 ;
        RECT 85.520 193.085 85.940 193.425 ;
        RECT 86.230 193.085 86.640 193.415 ;
        RECT 85.520 192.315 85.710 193.085 ;
        RECT 86.810 192.955 86.980 193.685 ;
        RECT 88.125 193.515 88.295 193.845 ;
        RECT 88.465 193.685 88.795 194.065 ;
        RECT 87.150 193.135 87.500 193.505 ;
        RECT 86.810 192.915 87.230 192.955 ;
        RECT 85.880 192.745 87.230 192.915 ;
        RECT 85.880 192.585 86.130 192.745 ;
        RECT 86.640 192.315 86.890 192.575 ;
        RECT 85.520 192.065 86.890 192.315 ;
        RECT 83.450 191.775 83.690 192.065 ;
        RECT 84.490 191.985 84.660 192.065 ;
        RECT 83.890 191.515 84.310 191.895 ;
        RECT 84.490 191.735 85.120 191.985 ;
        RECT 85.590 191.515 85.920 191.895 ;
        RECT 86.090 191.775 86.260 192.065 ;
        RECT 87.060 191.900 87.230 192.745 ;
        RECT 87.680 192.575 87.900 193.445 ;
        RECT 88.125 193.325 88.820 193.515 ;
        RECT 87.400 192.195 87.900 192.575 ;
        RECT 88.070 192.525 88.480 193.145 ;
        RECT 88.650 192.355 88.820 193.325 ;
        RECT 88.125 192.185 88.820 192.355 ;
        RECT 86.440 191.515 86.820 191.895 ;
        RECT 87.060 191.730 87.890 191.900 ;
        RECT 88.125 191.685 88.295 192.185 ;
        RECT 88.465 191.515 88.795 192.015 ;
        RECT 89.010 191.685 89.235 193.805 ;
        RECT 89.405 193.685 89.735 194.065 ;
        RECT 89.905 193.515 90.075 193.805 ;
        RECT 89.410 193.345 90.075 193.515 ;
        RECT 89.410 192.355 89.640 193.345 ;
        RECT 90.335 193.340 90.625 194.065 ;
        RECT 90.855 193.245 91.065 194.065 ;
        RECT 91.235 193.265 91.565 193.895 ;
        RECT 89.810 192.525 90.160 193.175 ;
        RECT 89.410 192.185 90.075 192.355 ;
        RECT 89.405 191.515 89.735 192.015 ;
        RECT 89.905 191.685 90.075 192.185 ;
        RECT 90.335 191.515 90.625 192.680 ;
        RECT 91.235 192.665 91.485 193.265 ;
        RECT 91.735 193.245 91.965 194.065 ;
        RECT 92.235 193.245 92.445 194.065 ;
        RECT 92.615 193.265 92.945 193.895 ;
        RECT 91.655 192.825 91.985 193.075 ;
        RECT 92.615 192.665 92.865 193.265 ;
        RECT 93.115 193.245 93.345 194.065 ;
        RECT 93.555 193.390 93.815 193.895 ;
        RECT 93.995 193.685 94.325 194.065 ;
        RECT 94.505 193.515 94.675 193.895 ;
        RECT 93.035 192.825 93.365 193.075 ;
        RECT 90.855 191.515 91.065 192.655 ;
        RECT 91.235 191.685 91.565 192.665 ;
        RECT 91.735 191.515 91.965 192.655 ;
        RECT 92.235 191.515 92.445 192.655 ;
        RECT 92.615 191.685 92.945 192.665 ;
        RECT 93.115 191.515 93.345 192.655 ;
        RECT 93.555 192.590 93.725 193.390 ;
        RECT 94.010 193.345 94.675 193.515 ;
        RECT 94.010 193.090 94.180 193.345 ;
        RECT 95.670 193.255 95.915 193.860 ;
        RECT 96.135 193.530 96.645 194.065 ;
        RECT 93.895 192.760 94.180 193.090 ;
        RECT 94.415 192.795 94.745 193.165 ;
        RECT 95.395 193.085 96.625 193.255 ;
        RECT 94.010 192.615 94.180 192.760 ;
        RECT 93.555 191.685 93.825 192.590 ;
        RECT 94.010 192.445 94.675 192.615 ;
        RECT 93.995 191.515 94.325 192.275 ;
        RECT 94.505 191.685 94.675 192.445 ;
        RECT 95.395 192.275 95.735 193.085 ;
        RECT 95.905 192.520 96.655 192.710 ;
        RECT 95.395 191.865 95.910 192.275 ;
        RECT 96.145 191.515 96.315 192.275 ;
        RECT 96.485 191.855 96.655 192.520 ;
        RECT 96.825 192.535 97.015 193.895 ;
        RECT 97.185 193.045 97.460 193.895 ;
        RECT 97.650 193.530 98.180 193.895 ;
        RECT 98.605 193.665 98.935 194.065 ;
        RECT 98.005 193.495 98.180 193.530 ;
        RECT 97.185 192.875 97.465 193.045 ;
        RECT 97.185 192.735 97.460 192.875 ;
        RECT 97.665 192.535 97.835 193.335 ;
        RECT 96.825 192.365 97.835 192.535 ;
        RECT 98.005 193.325 98.935 193.495 ;
        RECT 99.105 193.325 99.360 193.895 ;
        RECT 98.005 192.195 98.175 193.325 ;
        RECT 98.765 193.155 98.935 193.325 ;
        RECT 97.050 192.025 98.175 192.195 ;
        RECT 98.345 192.825 98.540 193.155 ;
        RECT 98.765 192.825 99.020 193.155 ;
        RECT 98.345 191.855 98.515 192.825 ;
        RECT 99.190 192.655 99.360 193.325 ;
        RECT 99.535 193.315 100.745 194.065 ;
        RECT 96.485 191.685 98.515 191.855 ;
        RECT 98.685 191.515 98.855 192.655 ;
        RECT 99.025 191.685 99.360 192.655 ;
        RECT 99.535 192.605 100.055 193.145 ;
        RECT 100.225 192.775 100.745 193.315 ;
        RECT 100.975 193.245 101.185 194.065 ;
        RECT 101.355 193.265 101.685 193.895 ;
        RECT 101.355 192.665 101.605 193.265 ;
        RECT 101.855 193.245 102.085 194.065 ;
        RECT 103.215 193.295 106.725 194.065 ;
        RECT 101.775 192.825 102.105 193.075 ;
        RECT 99.535 191.515 100.745 192.605 ;
        RECT 100.975 191.515 101.185 192.655 ;
        RECT 101.355 191.685 101.685 192.665 ;
        RECT 101.855 191.515 102.085 192.655 ;
        RECT 103.215 192.605 104.905 193.125 ;
        RECT 105.075 192.775 106.725 193.295 ;
        RECT 106.900 193.355 107.155 193.885 ;
        RECT 107.325 193.605 107.630 194.065 ;
        RECT 107.875 193.685 108.945 193.855 ;
        RECT 106.900 192.705 107.110 193.355 ;
        RECT 107.875 193.330 108.195 193.685 ;
        RECT 107.870 193.155 108.195 193.330 ;
        RECT 107.280 192.855 108.195 193.155 ;
        RECT 108.365 193.115 108.605 193.515 ;
        RECT 108.775 193.455 108.945 193.685 ;
        RECT 109.115 193.625 109.305 194.065 ;
        RECT 109.475 193.615 110.425 193.895 ;
        RECT 110.645 193.705 110.995 193.875 ;
        RECT 108.775 193.285 109.305 193.455 ;
        RECT 107.280 192.825 108.020 192.855 ;
        RECT 103.215 191.515 106.725 192.605 ;
        RECT 106.900 191.825 107.155 192.705 ;
        RECT 107.325 191.515 107.630 192.655 ;
        RECT 107.850 192.235 108.020 192.825 ;
        RECT 108.365 192.745 108.905 193.115 ;
        RECT 109.085 193.005 109.305 193.285 ;
        RECT 109.475 192.835 109.645 193.615 ;
        RECT 109.240 192.665 109.645 192.835 ;
        RECT 109.815 192.825 110.165 193.445 ;
        RECT 109.240 192.575 109.410 192.665 ;
        RECT 110.335 192.655 110.545 193.445 ;
        RECT 108.190 192.405 109.410 192.575 ;
        RECT 109.870 192.495 110.545 192.655 ;
        RECT 107.850 192.065 108.650 192.235 ;
        RECT 107.970 191.515 108.300 191.895 ;
        RECT 108.480 191.775 108.650 192.065 ;
        RECT 109.240 192.025 109.410 192.405 ;
        RECT 109.580 192.485 110.545 192.495 ;
        RECT 110.735 193.315 110.995 193.705 ;
        RECT 111.205 193.605 111.535 194.065 ;
        RECT 112.410 193.675 113.265 193.845 ;
        RECT 113.470 193.675 113.965 193.845 ;
        RECT 114.135 193.705 114.465 194.065 ;
        RECT 110.735 192.625 110.905 193.315 ;
        RECT 111.075 192.965 111.245 193.145 ;
        RECT 111.415 193.135 112.205 193.385 ;
        RECT 112.410 192.965 112.580 193.675 ;
        RECT 112.750 193.165 113.105 193.385 ;
        RECT 111.075 192.795 112.765 192.965 ;
        RECT 109.580 192.195 110.040 192.485 ;
        RECT 110.735 192.455 112.235 192.625 ;
        RECT 110.735 192.315 110.905 192.455 ;
        RECT 110.345 192.145 110.905 192.315 ;
        RECT 108.820 191.515 109.070 191.975 ;
        RECT 109.240 191.685 110.110 192.025 ;
        RECT 110.345 191.685 110.515 192.145 ;
        RECT 111.350 192.115 112.425 192.285 ;
        RECT 110.685 191.515 111.055 191.975 ;
        RECT 111.350 191.775 111.520 192.115 ;
        RECT 111.690 191.515 112.020 191.945 ;
        RECT 112.255 191.775 112.425 192.115 ;
        RECT 112.595 192.015 112.765 192.795 ;
        RECT 112.935 192.575 113.105 193.165 ;
        RECT 113.275 192.765 113.625 193.385 ;
        RECT 112.935 192.185 113.400 192.575 ;
        RECT 113.795 192.315 113.965 193.675 ;
        RECT 114.135 192.485 114.595 193.535 ;
        RECT 113.570 192.145 113.965 192.315 ;
        RECT 113.570 192.015 113.740 192.145 ;
        RECT 112.595 191.685 113.275 192.015 ;
        RECT 113.490 191.685 113.740 192.015 ;
        RECT 113.910 191.515 114.160 191.975 ;
        RECT 114.330 191.700 114.655 192.485 ;
        RECT 114.825 191.685 114.995 193.805 ;
        RECT 115.165 193.685 115.495 194.065 ;
        RECT 115.665 193.515 115.920 193.805 ;
        RECT 115.170 193.345 115.920 193.515 ;
        RECT 115.170 192.355 115.400 193.345 ;
        RECT 116.095 193.340 116.385 194.065 ;
        RECT 116.645 193.515 116.815 193.895 ;
        RECT 116.995 193.685 117.325 194.065 ;
        RECT 116.645 193.345 117.310 193.515 ;
        RECT 117.505 193.390 117.765 193.895 ;
        RECT 115.570 192.525 115.920 193.175 ;
        RECT 116.575 192.795 116.905 193.165 ;
        RECT 117.140 193.090 117.310 193.345 ;
        RECT 117.140 192.760 117.425 193.090 ;
        RECT 115.170 192.185 115.920 192.355 ;
        RECT 115.165 191.515 115.495 192.015 ;
        RECT 115.665 191.685 115.920 192.185 ;
        RECT 116.095 191.515 116.385 192.680 ;
        RECT 117.140 192.615 117.310 192.760 ;
        RECT 116.645 192.445 117.310 192.615 ;
        RECT 117.595 192.590 117.765 193.390 ;
        RECT 118.855 193.295 122.365 194.065 ;
        RECT 122.540 193.520 127.885 194.065 ;
        RECT 116.645 191.685 116.815 192.445 ;
        RECT 116.995 191.515 117.325 192.275 ;
        RECT 117.495 191.685 117.765 192.590 ;
        RECT 118.855 192.605 120.545 193.125 ;
        RECT 120.715 192.775 122.365 193.295 ;
        RECT 118.855 191.515 122.365 192.605 ;
        RECT 124.130 191.950 124.480 193.200 ;
        RECT 125.960 192.690 126.300 193.520 ;
        RECT 128.055 193.315 129.265 194.065 ;
        RECT 128.055 192.605 128.575 193.145 ;
        RECT 128.745 192.775 129.265 193.315 ;
        RECT 122.540 191.515 127.885 191.950 ;
        RECT 128.055 191.515 129.265 192.605 ;
        RECT 9.290 191.345 129.350 191.515 ;
        RECT 9.375 190.255 10.585 191.345 ;
        RECT 9.375 189.545 9.895 190.085 ;
        RECT 10.065 189.715 10.585 190.255 ;
        RECT 11.215 190.255 14.725 191.345 ;
        RECT 14.900 190.910 20.245 191.345 ;
        RECT 20.420 190.910 25.765 191.345 ;
        RECT 11.215 189.735 12.905 190.255 ;
        RECT 13.075 189.565 14.725 190.085 ;
        RECT 16.490 189.660 16.840 190.910 ;
        RECT 9.375 188.795 10.585 189.545 ;
        RECT 11.215 188.795 14.725 189.565 ;
        RECT 18.320 189.340 18.660 190.170 ;
        RECT 22.010 189.660 22.360 190.910 ;
        RECT 25.935 190.180 26.225 191.345 ;
        RECT 26.855 190.255 29.445 191.345 ;
        RECT 23.840 189.340 24.180 190.170 ;
        RECT 26.855 189.735 28.065 190.255 ;
        RECT 29.655 190.205 29.885 191.345 ;
        RECT 30.055 190.195 30.385 191.175 ;
        RECT 30.555 190.205 30.765 191.345 ;
        RECT 31.370 190.365 31.625 191.035 ;
        RECT 31.805 190.545 32.090 191.345 ;
        RECT 32.270 190.625 32.600 191.135 ;
        RECT 28.235 189.565 29.445 190.085 ;
        RECT 29.635 189.785 29.965 190.035 ;
        RECT 14.900 188.795 20.245 189.340 ;
        RECT 20.420 188.795 25.765 189.340 ;
        RECT 25.935 188.795 26.225 189.520 ;
        RECT 26.855 188.795 29.445 189.565 ;
        RECT 29.655 188.795 29.885 189.615 ;
        RECT 30.135 189.595 30.385 190.195 ;
        RECT 30.055 188.965 30.385 189.595 ;
        RECT 30.555 188.795 30.765 189.615 ;
        RECT 31.370 189.505 31.550 190.365 ;
        RECT 32.270 190.035 32.520 190.625 ;
        RECT 32.870 190.475 33.040 191.085 ;
        RECT 33.210 190.655 33.540 191.345 ;
        RECT 33.770 190.795 34.010 191.085 ;
        RECT 34.210 190.965 34.630 191.345 ;
        RECT 34.810 190.875 35.440 191.125 ;
        RECT 35.910 190.965 36.240 191.345 ;
        RECT 34.810 190.795 34.980 190.875 ;
        RECT 36.410 190.795 36.580 191.085 ;
        RECT 36.760 190.965 37.140 191.345 ;
        RECT 37.380 190.960 38.210 191.130 ;
        RECT 33.770 190.625 34.980 190.795 ;
        RECT 31.720 189.705 32.520 190.035 ;
        RECT 31.370 189.305 31.625 189.505 ;
        RECT 31.285 189.135 31.625 189.305 ;
        RECT 31.370 188.975 31.625 189.135 ;
        RECT 31.805 188.795 32.090 189.255 ;
        RECT 32.270 189.055 32.520 189.705 ;
        RECT 32.720 190.455 33.040 190.475 ;
        RECT 32.720 190.285 34.640 190.455 ;
        RECT 32.720 189.390 32.910 190.285 ;
        RECT 34.810 190.115 34.980 190.625 ;
        RECT 35.150 190.365 35.670 190.675 ;
        RECT 33.080 189.945 34.980 190.115 ;
        RECT 33.080 189.885 33.410 189.945 ;
        RECT 33.560 189.715 33.890 189.775 ;
        RECT 33.230 189.445 33.890 189.715 ;
        RECT 32.720 189.060 33.040 189.390 ;
        RECT 33.220 188.795 33.880 189.275 ;
        RECT 34.080 189.185 34.250 189.945 ;
        RECT 35.150 189.775 35.330 190.185 ;
        RECT 34.420 189.605 34.750 189.725 ;
        RECT 35.500 189.605 35.670 190.365 ;
        RECT 34.420 189.435 35.670 189.605 ;
        RECT 35.840 190.545 37.210 190.795 ;
        RECT 35.840 189.775 36.030 190.545 ;
        RECT 36.960 190.285 37.210 190.545 ;
        RECT 36.200 190.115 36.450 190.275 ;
        RECT 37.380 190.115 37.550 190.960 ;
        RECT 38.445 190.675 38.615 191.175 ;
        RECT 38.785 190.845 39.115 191.345 ;
        RECT 37.720 190.285 38.220 190.665 ;
        RECT 38.445 190.505 39.140 190.675 ;
        RECT 36.200 189.945 37.550 190.115 ;
        RECT 37.130 189.905 37.550 189.945 ;
        RECT 35.840 189.435 36.260 189.775 ;
        RECT 36.550 189.445 36.960 189.775 ;
        RECT 34.080 189.015 34.930 189.185 ;
        RECT 35.490 188.795 35.810 189.255 ;
        RECT 36.010 189.005 36.260 189.435 ;
        RECT 36.550 188.795 36.960 189.235 ;
        RECT 37.130 189.175 37.300 189.905 ;
        RECT 37.470 189.355 37.820 189.725 ;
        RECT 38.000 189.415 38.220 190.285 ;
        RECT 38.390 189.715 38.800 190.335 ;
        RECT 38.970 189.535 39.140 190.505 ;
        RECT 38.445 189.345 39.140 189.535 ;
        RECT 37.130 188.975 38.145 189.175 ;
        RECT 38.445 189.015 38.615 189.345 ;
        RECT 38.785 188.795 39.115 189.175 ;
        RECT 39.330 189.055 39.555 191.175 ;
        RECT 39.725 190.845 40.055 191.345 ;
        RECT 40.225 190.675 40.395 191.175 ;
        RECT 39.730 190.505 40.395 190.675 ;
        RECT 39.730 189.515 39.960 190.505 ;
        RECT 40.130 189.685 40.480 190.335 ;
        RECT 40.655 190.270 40.925 191.175 ;
        RECT 41.095 190.585 41.425 191.345 ;
        RECT 41.605 190.415 41.775 191.175 ;
        RECT 39.730 189.345 40.395 189.515 ;
        RECT 39.725 188.795 40.055 189.175 ;
        RECT 40.225 189.055 40.395 189.345 ;
        RECT 40.655 189.470 40.825 190.270 ;
        RECT 41.110 190.245 41.775 190.415 ;
        RECT 41.110 190.100 41.280 190.245 ;
        RECT 40.995 189.770 41.280 190.100 ;
        RECT 42.500 190.155 42.755 191.035 ;
        RECT 42.925 190.205 43.230 191.345 ;
        RECT 43.570 190.965 43.900 191.345 ;
        RECT 44.080 190.795 44.250 191.085 ;
        RECT 44.420 190.885 44.670 191.345 ;
        RECT 43.450 190.625 44.250 190.795 ;
        RECT 44.840 190.835 45.710 191.175 ;
        RECT 41.110 189.515 41.280 189.770 ;
        RECT 41.515 189.695 41.845 190.065 ;
        RECT 40.655 188.965 40.915 189.470 ;
        RECT 41.110 189.345 41.775 189.515 ;
        RECT 41.095 188.795 41.425 189.175 ;
        RECT 41.605 188.965 41.775 189.345 ;
        RECT 42.500 189.505 42.710 190.155 ;
        RECT 43.450 190.035 43.620 190.625 ;
        RECT 44.840 190.455 45.010 190.835 ;
        RECT 45.945 190.715 46.115 191.175 ;
        RECT 46.285 190.885 46.655 191.345 ;
        RECT 46.950 190.745 47.120 191.085 ;
        RECT 47.290 190.915 47.620 191.345 ;
        RECT 47.855 190.745 48.025 191.085 ;
        RECT 43.790 190.285 45.010 190.455 ;
        RECT 45.180 190.375 45.640 190.665 ;
        RECT 45.945 190.545 46.505 190.715 ;
        RECT 46.950 190.575 48.025 190.745 ;
        RECT 48.195 190.845 48.875 191.175 ;
        RECT 49.090 190.845 49.340 191.175 ;
        RECT 49.510 190.885 49.760 191.345 ;
        RECT 46.335 190.405 46.505 190.545 ;
        RECT 45.180 190.365 46.145 190.375 ;
        RECT 44.840 190.195 45.010 190.285 ;
        RECT 45.470 190.205 46.145 190.365 ;
        RECT 42.880 190.005 43.620 190.035 ;
        RECT 42.880 189.705 43.795 190.005 ;
        RECT 43.470 189.530 43.795 189.705 ;
        RECT 42.500 188.975 42.755 189.505 ;
        RECT 42.925 188.795 43.230 189.255 ;
        RECT 43.475 189.175 43.795 189.530 ;
        RECT 43.965 189.745 44.505 190.115 ;
        RECT 44.840 190.025 45.245 190.195 ;
        RECT 43.965 189.345 44.205 189.745 ;
        RECT 44.685 189.575 44.905 189.855 ;
        RECT 44.375 189.405 44.905 189.575 ;
        RECT 44.375 189.175 44.545 189.405 ;
        RECT 45.075 189.245 45.245 190.025 ;
        RECT 45.415 189.415 45.765 190.035 ;
        RECT 45.935 189.415 46.145 190.205 ;
        RECT 46.335 190.235 47.835 190.405 ;
        RECT 46.335 189.545 46.505 190.235 ;
        RECT 48.195 190.065 48.365 190.845 ;
        RECT 49.170 190.715 49.340 190.845 ;
        RECT 46.675 189.895 48.365 190.065 ;
        RECT 48.535 190.285 49.000 190.675 ;
        RECT 49.170 190.545 49.565 190.715 ;
        RECT 46.675 189.715 46.845 189.895 ;
        RECT 43.475 189.005 44.545 189.175 ;
        RECT 44.715 188.795 44.905 189.235 ;
        RECT 45.075 188.965 46.025 189.245 ;
        RECT 46.335 189.155 46.595 189.545 ;
        RECT 47.015 189.475 47.805 189.725 ;
        RECT 46.245 188.985 46.595 189.155 ;
        RECT 46.805 188.795 47.135 189.255 ;
        RECT 48.010 189.185 48.180 189.895 ;
        RECT 48.535 189.695 48.705 190.285 ;
        RECT 48.350 189.475 48.705 189.695 ;
        RECT 48.875 189.475 49.225 190.095 ;
        RECT 49.395 189.185 49.565 190.545 ;
        RECT 49.930 190.375 50.255 191.160 ;
        RECT 49.735 189.325 50.195 190.375 ;
        RECT 48.010 189.015 48.865 189.185 ;
        RECT 49.070 189.015 49.565 189.185 ;
        RECT 49.735 188.795 50.065 189.155 ;
        RECT 50.425 189.055 50.595 191.175 ;
        RECT 50.765 190.845 51.095 191.345 ;
        RECT 51.265 190.675 51.520 191.175 ;
        RECT 50.770 190.505 51.520 190.675 ;
        RECT 50.770 189.515 51.000 190.505 ;
        RECT 51.170 189.685 51.520 190.335 ;
        RECT 51.695 190.180 51.985 191.345 ;
        RECT 52.215 190.205 52.425 191.345 ;
        RECT 52.595 190.195 52.925 191.175 ;
        RECT 53.095 190.205 53.325 191.345 ;
        RECT 53.535 190.255 56.125 191.345 ;
        RECT 56.300 190.910 61.645 191.345 ;
        RECT 50.770 189.345 51.520 189.515 ;
        RECT 50.765 188.795 51.095 189.175 ;
        RECT 51.265 189.055 51.520 189.345 ;
        RECT 51.695 188.795 51.985 189.520 ;
        RECT 52.215 188.795 52.425 189.615 ;
        RECT 52.595 189.595 52.845 190.195 ;
        RECT 53.015 189.785 53.345 190.035 ;
        RECT 53.535 189.735 54.745 190.255 ;
        RECT 52.595 188.965 52.925 189.595 ;
        RECT 53.095 188.795 53.325 189.615 ;
        RECT 54.915 189.565 56.125 190.085 ;
        RECT 57.890 189.660 58.240 190.910 ;
        RECT 62.115 190.705 62.445 191.135 ;
        RECT 61.990 190.535 62.445 190.705 ;
        RECT 62.625 190.705 62.875 191.125 ;
        RECT 63.105 190.875 63.435 191.345 ;
        RECT 63.665 190.705 63.915 191.125 ;
        RECT 62.625 190.535 63.915 190.705 ;
        RECT 53.535 188.795 56.125 189.565 ;
        RECT 59.720 189.340 60.060 190.170 ;
        RECT 61.990 189.535 62.160 190.535 ;
        RECT 62.330 189.705 62.575 190.365 ;
        RECT 62.790 189.705 63.055 190.365 ;
        RECT 63.250 189.705 63.535 190.365 ;
        RECT 63.710 190.035 63.925 190.365 ;
        RECT 64.105 190.205 64.355 191.345 ;
        RECT 64.525 190.285 64.855 191.135 ;
        RECT 63.710 189.705 64.015 190.035 ;
        RECT 64.185 189.705 64.495 190.035 ;
        RECT 64.185 189.535 64.355 189.705 ;
        RECT 61.990 189.365 64.355 189.535 ;
        RECT 64.665 189.520 64.855 190.285 ;
        RECT 65.035 190.205 65.295 191.345 ;
        RECT 65.535 190.835 67.150 191.165 ;
        RECT 65.545 190.035 65.715 190.595 ;
        RECT 65.975 190.495 67.150 190.665 ;
        RECT 67.320 190.545 67.600 191.345 ;
        RECT 65.975 190.205 66.305 190.495 ;
        RECT 66.980 190.375 67.150 190.495 ;
        RECT 66.475 190.035 66.720 190.325 ;
        RECT 66.980 190.205 67.640 190.375 ;
        RECT 67.810 190.205 68.085 191.175 ;
        RECT 67.470 190.035 67.640 190.205 ;
        RECT 65.040 189.785 65.375 190.035 ;
        RECT 65.545 189.705 66.260 190.035 ;
        RECT 66.475 189.705 67.300 190.035 ;
        RECT 67.470 189.705 67.745 190.035 ;
        RECT 65.545 189.615 65.795 189.705 ;
        RECT 56.300 188.795 61.645 189.340 ;
        RECT 62.145 188.795 62.475 189.195 ;
        RECT 62.645 189.025 62.975 189.365 ;
        RECT 64.025 188.795 64.355 189.195 ;
        RECT 64.525 189.010 64.855 189.520 ;
        RECT 65.035 188.795 65.295 189.615 ;
        RECT 65.465 189.195 65.795 189.615 ;
        RECT 67.470 189.535 67.640 189.705 ;
        RECT 65.975 189.365 67.640 189.535 ;
        RECT 67.915 189.470 68.085 190.205 ;
        RECT 65.975 188.965 66.235 189.365 ;
        RECT 66.405 188.795 66.735 189.195 ;
        RECT 66.905 189.015 67.075 189.365 ;
        RECT 67.245 188.795 67.620 189.195 ;
        RECT 67.810 189.125 68.085 189.470 ;
        RECT 68.255 190.205 68.530 191.175 ;
        RECT 68.740 190.545 69.020 191.345 ;
        RECT 69.190 190.835 70.805 191.165 ;
        RECT 69.190 190.495 70.365 190.665 ;
        RECT 69.190 190.375 69.360 190.495 ;
        RECT 68.700 190.205 69.360 190.375 ;
        RECT 68.255 189.470 68.425 190.205 ;
        RECT 68.700 190.035 68.870 190.205 ;
        RECT 69.620 190.035 69.865 190.325 ;
        RECT 70.035 190.205 70.365 190.495 ;
        RECT 70.625 190.035 70.795 190.595 ;
        RECT 71.045 190.205 71.305 191.345 ;
        RECT 71.660 190.375 72.050 190.550 ;
        RECT 72.535 190.545 72.865 191.345 ;
        RECT 73.035 190.555 73.570 191.175 ;
        RECT 71.660 190.205 73.085 190.375 ;
        RECT 68.595 189.705 68.870 190.035 ;
        RECT 69.040 189.705 69.865 190.035 ;
        RECT 70.080 189.705 70.795 190.035 ;
        RECT 70.965 189.785 71.300 190.035 ;
        RECT 68.700 189.535 68.870 189.705 ;
        RECT 70.545 189.615 70.795 189.705 ;
        RECT 68.255 189.125 68.530 189.470 ;
        RECT 68.700 189.365 70.365 189.535 ;
        RECT 68.720 188.795 69.095 189.195 ;
        RECT 69.265 189.015 69.435 189.365 ;
        RECT 69.605 188.795 69.935 189.195 ;
        RECT 70.105 188.965 70.365 189.365 ;
        RECT 70.545 189.195 70.875 189.615 ;
        RECT 71.045 188.795 71.305 189.615 ;
        RECT 71.535 189.475 71.890 190.035 ;
        RECT 72.060 189.305 72.230 190.205 ;
        RECT 72.400 189.475 72.665 190.035 ;
        RECT 72.915 189.705 73.085 190.205 ;
        RECT 73.255 189.535 73.570 190.555 ;
        RECT 71.640 188.795 71.880 189.305 ;
        RECT 72.060 188.975 72.340 189.305 ;
        RECT 72.570 188.795 72.785 189.305 ;
        RECT 72.955 188.965 73.570 189.535 ;
        RECT 73.775 190.475 74.050 191.175 ;
        RECT 74.220 190.800 74.475 191.345 ;
        RECT 74.645 190.835 75.125 191.175 ;
        RECT 75.300 190.790 75.905 191.345 ;
        RECT 75.290 190.690 75.905 190.790 ;
        RECT 75.290 190.665 75.475 190.690 ;
        RECT 73.775 189.445 73.945 190.475 ;
        RECT 74.220 190.345 74.975 190.595 ;
        RECT 75.145 190.420 75.475 190.665 ;
        RECT 74.220 190.310 74.990 190.345 ;
        RECT 74.220 190.300 75.005 190.310 ;
        RECT 74.115 190.285 75.010 190.300 ;
        RECT 74.115 190.270 75.030 190.285 ;
        RECT 74.115 190.260 75.050 190.270 ;
        RECT 74.115 190.250 75.075 190.260 ;
        RECT 74.115 190.220 75.145 190.250 ;
        RECT 74.115 190.190 75.165 190.220 ;
        RECT 74.115 190.160 75.185 190.190 ;
        RECT 74.115 190.135 75.215 190.160 ;
        RECT 74.115 190.100 75.250 190.135 ;
        RECT 74.115 190.095 75.280 190.100 ;
        RECT 74.115 189.700 74.345 190.095 ;
        RECT 74.890 190.090 75.280 190.095 ;
        RECT 74.915 190.080 75.280 190.090 ;
        RECT 74.930 190.075 75.280 190.080 ;
        RECT 74.945 190.070 75.280 190.075 ;
        RECT 75.645 190.070 75.905 190.520 ;
        RECT 74.945 190.065 75.905 190.070 ;
        RECT 74.955 190.055 75.905 190.065 ;
        RECT 74.965 190.050 75.905 190.055 ;
        RECT 74.975 190.040 75.905 190.050 ;
        RECT 74.980 190.030 75.905 190.040 ;
        RECT 74.985 190.025 75.905 190.030 ;
        RECT 74.995 190.010 75.905 190.025 ;
        RECT 75.000 189.995 75.905 190.010 ;
        RECT 75.010 189.970 75.905 189.995 ;
        RECT 74.515 189.500 74.845 189.925 ;
        RECT 74.595 189.475 74.845 189.500 ;
        RECT 73.775 188.965 74.035 189.445 ;
        RECT 74.205 188.795 74.455 189.335 ;
        RECT 74.625 189.015 74.845 189.475 ;
        RECT 75.015 189.900 75.905 189.970 ;
        RECT 76.075 190.255 77.285 191.345 ;
        RECT 75.015 189.175 75.185 189.900 ;
        RECT 75.355 189.345 75.905 189.730 ;
        RECT 76.075 189.715 76.595 190.255 ;
        RECT 77.455 190.180 77.745 191.345 ;
        RECT 77.915 190.255 80.505 191.345 ;
        RECT 80.680 190.910 86.025 191.345 ;
        RECT 76.765 189.545 77.285 190.085 ;
        RECT 77.915 189.735 79.125 190.255 ;
        RECT 79.295 189.565 80.505 190.085 ;
        RECT 82.270 189.660 82.620 190.910 ;
        RECT 86.195 190.585 86.710 190.995 ;
        RECT 86.945 190.585 87.115 191.345 ;
        RECT 87.285 191.005 89.315 191.175 ;
        RECT 75.015 189.005 75.905 189.175 ;
        RECT 76.075 188.795 77.285 189.545 ;
        RECT 77.455 188.795 77.745 189.520 ;
        RECT 77.915 188.795 80.505 189.565 ;
        RECT 84.100 189.340 84.440 190.170 ;
        RECT 86.195 189.775 86.535 190.585 ;
        RECT 87.285 190.340 87.455 191.005 ;
        RECT 87.850 190.665 88.975 190.835 ;
        RECT 86.705 190.150 87.455 190.340 ;
        RECT 87.625 190.325 88.635 190.495 ;
        RECT 86.195 189.605 87.425 189.775 ;
        RECT 80.680 188.795 86.025 189.340 ;
        RECT 86.470 189.000 86.715 189.605 ;
        RECT 86.935 188.795 87.445 189.330 ;
        RECT 87.625 188.965 87.815 190.325 ;
        RECT 87.985 189.305 88.260 190.125 ;
        RECT 88.465 189.525 88.635 190.325 ;
        RECT 88.805 189.535 88.975 190.665 ;
        RECT 89.145 190.035 89.315 191.005 ;
        RECT 89.485 190.205 89.655 191.345 ;
        RECT 89.825 190.205 90.160 191.175 ;
        RECT 89.145 189.705 89.340 190.035 ;
        RECT 89.565 189.705 89.820 190.035 ;
        RECT 89.565 189.535 89.735 189.705 ;
        RECT 89.990 189.535 90.160 190.205 ;
        RECT 88.805 189.365 89.735 189.535 ;
        RECT 88.805 189.330 88.980 189.365 ;
        RECT 87.985 189.135 88.265 189.305 ;
        RECT 87.985 188.965 88.260 189.135 ;
        RECT 88.450 188.965 88.980 189.330 ;
        RECT 89.405 188.795 89.735 189.195 ;
        RECT 89.905 188.965 90.160 189.535 ;
        RECT 90.335 190.270 90.605 191.175 ;
        RECT 90.775 190.585 91.105 191.345 ;
        RECT 91.285 190.415 91.455 191.175 ;
        RECT 90.335 189.470 90.505 190.270 ;
        RECT 90.790 190.245 91.455 190.415 ;
        RECT 92.175 190.255 93.845 191.345 ;
        RECT 94.020 190.675 94.275 191.175 ;
        RECT 94.445 190.845 94.775 191.345 ;
        RECT 94.020 190.505 94.770 190.675 ;
        RECT 90.790 190.100 90.960 190.245 ;
        RECT 90.675 189.770 90.960 190.100 ;
        RECT 90.790 189.515 90.960 189.770 ;
        RECT 91.195 189.695 91.525 190.065 ;
        RECT 92.175 189.735 92.925 190.255 ;
        RECT 93.095 189.565 93.845 190.085 ;
        RECT 94.020 189.685 94.370 190.335 ;
        RECT 90.335 188.965 90.595 189.470 ;
        RECT 90.790 189.345 91.455 189.515 ;
        RECT 90.775 188.795 91.105 189.175 ;
        RECT 91.285 188.965 91.455 189.345 ;
        RECT 92.175 188.795 93.845 189.565 ;
        RECT 94.540 189.515 94.770 190.505 ;
        RECT 94.020 189.345 94.770 189.515 ;
        RECT 94.020 189.055 94.275 189.345 ;
        RECT 94.445 188.795 94.775 189.175 ;
        RECT 94.945 189.055 95.115 191.175 ;
        RECT 95.285 190.375 95.610 191.160 ;
        RECT 95.780 190.885 96.030 191.345 ;
        RECT 96.200 190.845 96.450 191.175 ;
        RECT 96.665 190.845 97.345 191.175 ;
        RECT 96.200 190.715 96.370 190.845 ;
        RECT 95.975 190.545 96.370 190.715 ;
        RECT 95.345 189.325 95.805 190.375 ;
        RECT 95.975 189.185 96.145 190.545 ;
        RECT 96.540 190.285 97.005 190.675 ;
        RECT 96.315 189.475 96.665 190.095 ;
        RECT 96.835 189.695 97.005 190.285 ;
        RECT 97.175 190.065 97.345 190.845 ;
        RECT 97.515 190.745 97.685 191.085 ;
        RECT 97.920 190.915 98.250 191.345 ;
        RECT 98.420 190.745 98.590 191.085 ;
        RECT 98.885 190.885 99.255 191.345 ;
        RECT 97.515 190.575 98.590 190.745 ;
        RECT 99.425 190.715 99.595 191.175 ;
        RECT 99.830 190.835 100.700 191.175 ;
        RECT 100.870 190.885 101.120 191.345 ;
        RECT 99.035 190.545 99.595 190.715 ;
        RECT 99.035 190.405 99.205 190.545 ;
        RECT 97.705 190.235 99.205 190.405 ;
        RECT 99.900 190.375 100.360 190.665 ;
        RECT 97.175 189.895 98.865 190.065 ;
        RECT 96.835 189.475 97.190 189.695 ;
        RECT 97.360 189.185 97.530 189.895 ;
        RECT 97.735 189.475 98.525 189.725 ;
        RECT 98.695 189.715 98.865 189.895 ;
        RECT 99.035 189.545 99.205 190.235 ;
        RECT 95.475 188.795 95.805 189.155 ;
        RECT 95.975 189.015 96.470 189.185 ;
        RECT 96.675 189.015 97.530 189.185 ;
        RECT 98.405 188.795 98.735 189.255 ;
        RECT 98.945 189.155 99.205 189.545 ;
        RECT 99.395 190.365 100.360 190.375 ;
        RECT 100.530 190.455 100.700 190.835 ;
        RECT 101.290 190.795 101.460 191.085 ;
        RECT 101.640 190.965 101.970 191.345 ;
        RECT 101.290 190.625 102.090 190.795 ;
        RECT 99.395 190.205 100.070 190.365 ;
        RECT 100.530 190.285 101.750 190.455 ;
        RECT 99.395 189.415 99.605 190.205 ;
        RECT 100.530 190.195 100.700 190.285 ;
        RECT 99.775 189.415 100.125 190.035 ;
        RECT 100.295 190.025 100.700 190.195 ;
        RECT 100.295 189.245 100.465 190.025 ;
        RECT 100.635 189.575 100.855 189.855 ;
        RECT 101.035 189.745 101.575 190.115 ;
        RECT 101.920 190.035 102.090 190.625 ;
        RECT 102.310 190.205 102.615 191.345 ;
        RECT 102.785 190.155 103.040 191.035 ;
        RECT 103.215 190.180 103.505 191.345 ;
        RECT 103.675 190.255 104.885 191.345 ;
        RECT 105.060 190.910 110.405 191.345 ;
        RECT 101.920 190.005 102.660 190.035 ;
        RECT 100.635 189.405 101.165 189.575 ;
        RECT 98.945 188.985 99.295 189.155 ;
        RECT 99.515 188.965 100.465 189.245 ;
        RECT 100.635 188.795 100.825 189.235 ;
        RECT 100.995 189.175 101.165 189.405 ;
        RECT 101.335 189.345 101.575 189.745 ;
        RECT 101.745 189.705 102.660 190.005 ;
        RECT 101.745 189.530 102.070 189.705 ;
        RECT 101.745 189.175 102.065 189.530 ;
        RECT 102.830 189.505 103.040 190.155 ;
        RECT 103.675 189.715 104.195 190.255 ;
        RECT 104.365 189.545 104.885 190.085 ;
        RECT 106.650 189.660 107.000 190.910 ;
        RECT 110.575 190.585 111.090 190.995 ;
        RECT 111.325 190.585 111.495 191.345 ;
        RECT 111.665 191.005 113.695 191.175 ;
        RECT 100.995 189.005 102.065 189.175 ;
        RECT 102.310 188.795 102.615 189.255 ;
        RECT 102.785 188.975 103.040 189.505 ;
        RECT 103.215 188.795 103.505 189.520 ;
        RECT 103.675 188.795 104.885 189.545 ;
        RECT 108.480 189.340 108.820 190.170 ;
        RECT 110.575 189.775 110.915 190.585 ;
        RECT 111.665 190.340 111.835 191.005 ;
        RECT 112.230 190.665 113.355 190.835 ;
        RECT 111.085 190.150 111.835 190.340 ;
        RECT 112.005 190.325 113.015 190.495 ;
        RECT 110.575 189.605 111.805 189.775 ;
        RECT 105.060 188.795 110.405 189.340 ;
        RECT 110.850 189.000 111.095 189.605 ;
        RECT 111.315 188.795 111.825 189.330 ;
        RECT 112.005 188.965 112.195 190.325 ;
        RECT 112.365 189.305 112.640 190.125 ;
        RECT 112.845 189.525 113.015 190.325 ;
        RECT 113.185 189.535 113.355 190.665 ;
        RECT 113.525 190.035 113.695 191.005 ;
        RECT 113.865 190.205 114.035 191.345 ;
        RECT 114.205 190.205 114.540 191.175 ;
        RECT 113.525 189.705 113.720 190.035 ;
        RECT 113.945 189.705 114.200 190.035 ;
        RECT 113.945 189.535 114.115 189.705 ;
        RECT 114.370 189.535 114.540 190.205 ;
        RECT 113.185 189.365 114.115 189.535 ;
        RECT 113.185 189.330 113.360 189.365 ;
        RECT 112.365 189.135 112.645 189.305 ;
        RECT 112.365 188.965 112.640 189.135 ;
        RECT 112.830 188.965 113.360 189.330 ;
        RECT 113.785 188.795 114.115 189.195 ;
        RECT 114.285 188.965 114.540 189.535 ;
        RECT 114.715 190.270 114.985 191.175 ;
        RECT 115.155 190.585 115.485 191.345 ;
        RECT 115.665 190.415 115.835 191.175 ;
        RECT 117.020 190.910 122.365 191.345 ;
        RECT 122.540 190.910 127.885 191.345 ;
        RECT 114.715 189.470 114.885 190.270 ;
        RECT 115.170 190.245 115.835 190.415 ;
        RECT 115.170 190.100 115.340 190.245 ;
        RECT 115.055 189.770 115.340 190.100 ;
        RECT 115.170 189.515 115.340 189.770 ;
        RECT 115.575 189.695 115.905 190.065 ;
        RECT 118.610 189.660 118.960 190.910 ;
        RECT 114.715 188.965 114.975 189.470 ;
        RECT 115.170 189.345 115.835 189.515 ;
        RECT 115.155 188.795 115.485 189.175 ;
        RECT 115.665 188.965 115.835 189.345 ;
        RECT 120.440 189.340 120.780 190.170 ;
        RECT 124.130 189.660 124.480 190.910 ;
        RECT 128.055 190.255 129.265 191.345 ;
        RECT 125.960 189.340 126.300 190.170 ;
        RECT 128.055 189.715 128.575 190.255 ;
        RECT 128.745 189.545 129.265 190.085 ;
        RECT 117.020 188.795 122.365 189.340 ;
        RECT 122.540 188.795 127.885 189.340 ;
        RECT 128.055 188.795 129.265 189.545 ;
        RECT 9.290 188.625 129.350 188.795 ;
        RECT 9.375 187.875 10.585 188.625 ;
        RECT 9.375 187.335 9.895 187.875 ;
        RECT 11.215 187.855 12.885 188.625 ;
        RECT 13.055 187.900 13.345 188.625 ;
        RECT 13.515 187.875 14.725 188.625 ;
        RECT 14.900 188.080 20.245 188.625 ;
        RECT 10.065 187.165 10.585 187.705 ;
        RECT 9.375 186.075 10.585 187.165 ;
        RECT 11.215 187.165 11.965 187.685 ;
        RECT 12.135 187.335 12.885 187.855 ;
        RECT 11.215 186.075 12.885 187.165 ;
        RECT 13.055 186.075 13.345 187.240 ;
        RECT 13.515 187.165 14.035 187.705 ;
        RECT 14.205 187.335 14.725 187.875 ;
        RECT 13.515 186.075 14.725 187.165 ;
        RECT 16.490 186.510 16.840 187.760 ;
        RECT 18.320 187.250 18.660 188.080 ;
        RECT 20.455 187.805 20.685 188.625 ;
        RECT 20.855 187.825 21.185 188.455 ;
        RECT 20.435 187.385 20.765 187.635 ;
        RECT 20.935 187.225 21.185 187.825 ;
        RECT 21.355 187.805 21.565 188.625 ;
        RECT 21.800 187.915 22.055 188.445 ;
        RECT 22.225 188.165 22.530 188.625 ;
        RECT 22.775 188.245 23.845 188.415 ;
        RECT 14.900 186.075 20.245 186.510 ;
        RECT 20.455 186.075 20.685 187.215 ;
        RECT 20.855 186.245 21.185 187.225 ;
        RECT 21.800 187.265 22.010 187.915 ;
        RECT 22.775 187.890 23.095 188.245 ;
        RECT 22.770 187.715 23.095 187.890 ;
        RECT 22.180 187.415 23.095 187.715 ;
        RECT 23.265 187.675 23.505 188.075 ;
        RECT 23.675 188.015 23.845 188.245 ;
        RECT 24.015 188.185 24.205 188.625 ;
        RECT 24.375 188.175 25.325 188.455 ;
        RECT 25.545 188.265 25.895 188.435 ;
        RECT 23.675 187.845 24.205 188.015 ;
        RECT 22.180 187.385 22.920 187.415 ;
        RECT 21.355 186.075 21.565 187.215 ;
        RECT 21.800 186.385 22.055 187.265 ;
        RECT 22.225 186.075 22.530 187.215 ;
        RECT 22.750 186.795 22.920 187.385 ;
        RECT 23.265 187.305 23.805 187.675 ;
        RECT 23.985 187.565 24.205 187.845 ;
        RECT 24.375 187.395 24.545 188.175 ;
        RECT 24.140 187.225 24.545 187.395 ;
        RECT 24.715 187.385 25.065 188.005 ;
        RECT 24.140 187.135 24.310 187.225 ;
        RECT 25.235 187.215 25.445 188.005 ;
        RECT 23.090 186.965 24.310 187.135 ;
        RECT 24.770 187.055 25.445 187.215 ;
        RECT 22.750 186.625 23.550 186.795 ;
        RECT 22.870 186.075 23.200 186.455 ;
        RECT 23.380 186.335 23.550 186.625 ;
        RECT 24.140 186.585 24.310 186.965 ;
        RECT 24.480 187.045 25.445 187.055 ;
        RECT 25.635 187.875 25.895 188.265 ;
        RECT 26.105 188.165 26.435 188.625 ;
        RECT 27.310 188.235 28.165 188.405 ;
        RECT 28.370 188.235 28.865 188.405 ;
        RECT 29.035 188.265 29.365 188.625 ;
        RECT 25.635 187.185 25.805 187.875 ;
        RECT 25.975 187.525 26.145 187.705 ;
        RECT 26.315 187.695 27.105 187.945 ;
        RECT 27.310 187.525 27.480 188.235 ;
        RECT 27.650 187.725 28.005 187.945 ;
        RECT 25.975 187.355 27.665 187.525 ;
        RECT 24.480 186.755 24.940 187.045 ;
        RECT 25.635 187.015 27.135 187.185 ;
        RECT 25.635 186.875 25.805 187.015 ;
        RECT 25.245 186.705 25.805 186.875 ;
        RECT 23.720 186.075 23.970 186.535 ;
        RECT 24.140 186.245 25.010 186.585 ;
        RECT 25.245 186.245 25.415 186.705 ;
        RECT 26.250 186.675 27.325 186.845 ;
        RECT 25.585 186.075 25.955 186.535 ;
        RECT 26.250 186.335 26.420 186.675 ;
        RECT 26.590 186.075 26.920 186.505 ;
        RECT 27.155 186.335 27.325 186.675 ;
        RECT 27.495 186.575 27.665 187.355 ;
        RECT 27.835 187.135 28.005 187.725 ;
        RECT 28.175 187.325 28.525 187.945 ;
        RECT 27.835 186.745 28.300 187.135 ;
        RECT 28.695 186.875 28.865 188.235 ;
        RECT 29.035 187.045 29.495 188.095 ;
        RECT 28.470 186.705 28.865 186.875 ;
        RECT 28.470 186.575 28.640 186.705 ;
        RECT 27.495 186.245 28.175 186.575 ;
        RECT 28.390 186.245 28.640 186.575 ;
        RECT 28.810 186.075 29.060 186.535 ;
        RECT 29.230 186.260 29.555 187.045 ;
        RECT 29.725 186.245 29.895 188.365 ;
        RECT 30.065 188.245 30.395 188.625 ;
        RECT 30.565 188.075 30.820 188.365 ;
        RECT 30.070 187.905 30.820 188.075 ;
        RECT 30.995 187.950 31.255 188.455 ;
        RECT 31.435 188.245 31.765 188.625 ;
        RECT 31.945 188.075 32.115 188.455 ;
        RECT 30.070 186.915 30.300 187.905 ;
        RECT 30.470 187.085 30.820 187.735 ;
        RECT 30.995 187.150 31.165 187.950 ;
        RECT 31.450 187.905 32.115 188.075 ;
        RECT 31.450 187.650 31.620 187.905 ;
        RECT 32.375 187.855 34.045 188.625 ;
        RECT 31.335 187.320 31.620 187.650 ;
        RECT 31.855 187.355 32.185 187.725 ;
        RECT 31.450 187.175 31.620 187.320 ;
        RECT 30.070 186.745 30.820 186.915 ;
        RECT 30.065 186.075 30.395 186.575 ;
        RECT 30.565 186.245 30.820 186.745 ;
        RECT 30.995 186.245 31.265 187.150 ;
        RECT 31.450 187.005 32.115 187.175 ;
        RECT 31.435 186.075 31.765 186.835 ;
        RECT 31.945 186.245 32.115 187.005 ;
        RECT 32.375 187.165 33.125 187.685 ;
        RECT 33.295 187.335 34.045 187.855 ;
        RECT 34.490 187.815 34.735 188.420 ;
        RECT 34.955 188.090 35.465 188.625 ;
        RECT 34.215 187.645 35.445 187.815 ;
        RECT 32.375 186.075 34.045 187.165 ;
        RECT 34.215 186.835 34.555 187.645 ;
        RECT 34.725 187.080 35.475 187.270 ;
        RECT 34.215 186.425 34.730 186.835 ;
        RECT 34.965 186.075 35.135 186.835 ;
        RECT 35.305 186.415 35.475 187.080 ;
        RECT 35.645 187.095 35.835 188.455 ;
        RECT 36.005 188.285 36.280 188.455 ;
        RECT 36.005 188.115 36.285 188.285 ;
        RECT 36.005 187.295 36.280 188.115 ;
        RECT 36.470 188.090 37.000 188.455 ;
        RECT 37.425 188.225 37.755 188.625 ;
        RECT 36.825 188.055 37.000 188.090 ;
        RECT 36.485 187.095 36.655 187.895 ;
        RECT 35.645 186.925 36.655 187.095 ;
        RECT 36.825 187.885 37.755 188.055 ;
        RECT 37.925 187.885 38.180 188.455 ;
        RECT 38.815 187.900 39.105 188.625 ;
        RECT 36.825 186.755 36.995 187.885 ;
        RECT 37.585 187.715 37.755 187.885 ;
        RECT 35.870 186.585 36.995 186.755 ;
        RECT 37.165 187.385 37.360 187.715 ;
        RECT 37.585 187.385 37.840 187.715 ;
        RECT 37.165 186.415 37.335 187.385 ;
        RECT 38.010 187.215 38.180 187.885 ;
        RECT 39.735 187.855 42.325 188.625 ;
        RECT 42.500 188.080 47.845 188.625 ;
        RECT 35.305 186.245 37.335 186.415 ;
        RECT 37.505 186.075 37.675 187.215 ;
        RECT 37.845 186.245 38.180 187.215 ;
        RECT 38.815 186.075 39.105 187.240 ;
        RECT 39.735 187.165 40.945 187.685 ;
        RECT 41.115 187.335 42.325 187.855 ;
        RECT 39.735 186.075 42.325 187.165 ;
        RECT 44.090 186.510 44.440 187.760 ;
        RECT 45.920 187.250 46.260 188.080 ;
        RECT 48.105 188.075 48.275 188.455 ;
        RECT 48.455 188.245 48.785 188.625 ;
        RECT 48.105 187.905 48.770 188.075 ;
        RECT 48.965 187.950 49.225 188.455 ;
        RECT 48.035 187.355 48.365 187.725 ;
        RECT 48.600 187.650 48.770 187.905 ;
        RECT 48.600 187.320 48.885 187.650 ;
        RECT 48.600 187.175 48.770 187.320 ;
        RECT 48.105 187.005 48.770 187.175 ;
        RECT 49.055 187.150 49.225 187.950 ;
        RECT 49.670 187.815 49.915 188.420 ;
        RECT 50.135 188.090 50.645 188.625 ;
        RECT 42.500 186.075 47.845 186.510 ;
        RECT 48.105 186.245 48.275 187.005 ;
        RECT 48.455 186.075 48.785 186.835 ;
        RECT 48.955 186.245 49.225 187.150 ;
        RECT 49.395 187.645 50.625 187.815 ;
        RECT 49.395 186.835 49.735 187.645 ;
        RECT 49.905 187.080 50.655 187.270 ;
        RECT 49.395 186.425 49.910 186.835 ;
        RECT 50.145 186.075 50.315 186.835 ;
        RECT 50.485 186.415 50.655 187.080 ;
        RECT 50.825 187.095 51.015 188.455 ;
        RECT 51.185 187.945 51.460 188.455 ;
        RECT 51.650 188.090 52.180 188.455 ;
        RECT 52.605 188.225 52.935 188.625 ;
        RECT 52.005 188.055 52.180 188.090 ;
        RECT 51.185 187.775 51.465 187.945 ;
        RECT 51.185 187.295 51.460 187.775 ;
        RECT 51.665 187.095 51.835 187.895 ;
        RECT 50.825 186.925 51.835 187.095 ;
        RECT 52.005 187.885 52.935 188.055 ;
        RECT 53.105 187.885 53.360 188.455 ;
        RECT 53.540 188.080 58.885 188.625 ;
        RECT 59.060 188.080 64.405 188.625 ;
        RECT 52.005 186.755 52.175 187.885 ;
        RECT 52.765 187.715 52.935 187.885 ;
        RECT 51.050 186.585 52.175 186.755 ;
        RECT 52.345 187.385 52.540 187.715 ;
        RECT 52.765 187.385 53.020 187.715 ;
        RECT 52.345 186.415 52.515 187.385 ;
        RECT 53.190 187.215 53.360 187.885 ;
        RECT 50.485 186.245 52.515 186.415 ;
        RECT 52.685 186.075 52.855 187.215 ;
        RECT 53.025 186.245 53.360 187.215 ;
        RECT 55.130 186.510 55.480 187.760 ;
        RECT 56.960 187.250 57.300 188.080 ;
        RECT 60.650 186.510 61.000 187.760 ;
        RECT 62.480 187.250 62.820 188.080 ;
        RECT 64.575 187.900 64.865 188.625 ;
        RECT 65.955 187.855 69.465 188.625 ;
        RECT 53.540 186.075 58.885 186.510 ;
        RECT 59.060 186.075 64.405 186.510 ;
        RECT 64.575 186.075 64.865 187.240 ;
        RECT 65.955 187.165 67.645 187.685 ;
        RECT 67.815 187.335 69.465 187.855 ;
        RECT 69.640 187.785 69.900 188.625 ;
        RECT 70.075 187.880 70.330 188.455 ;
        RECT 70.500 188.245 70.830 188.625 ;
        RECT 71.045 188.075 71.215 188.455 ;
        RECT 70.500 187.905 71.215 188.075 ;
        RECT 71.480 187.915 71.735 188.445 ;
        RECT 71.905 188.165 72.210 188.625 ;
        RECT 72.455 188.245 73.525 188.415 ;
        RECT 65.955 186.075 69.465 187.165 ;
        RECT 69.640 186.075 69.900 187.225 ;
        RECT 70.075 187.150 70.245 187.880 ;
        RECT 70.500 187.715 70.670 187.905 ;
        RECT 70.415 187.385 70.670 187.715 ;
        RECT 70.500 187.175 70.670 187.385 ;
        RECT 70.950 187.355 71.305 187.725 ;
        RECT 71.480 187.265 71.690 187.915 ;
        RECT 72.455 187.890 72.775 188.245 ;
        RECT 72.450 187.715 72.775 187.890 ;
        RECT 71.860 187.415 72.775 187.715 ;
        RECT 72.945 187.675 73.185 188.075 ;
        RECT 73.355 188.015 73.525 188.245 ;
        RECT 73.695 188.185 73.885 188.625 ;
        RECT 74.055 188.175 75.005 188.455 ;
        RECT 75.225 188.265 75.575 188.435 ;
        RECT 73.355 187.845 73.885 188.015 ;
        RECT 71.860 187.385 72.600 187.415 ;
        RECT 70.075 186.245 70.330 187.150 ;
        RECT 70.500 187.005 71.215 187.175 ;
        RECT 70.500 186.075 70.830 186.835 ;
        RECT 71.045 186.245 71.215 187.005 ;
        RECT 71.480 186.385 71.735 187.265 ;
        RECT 71.905 186.075 72.210 187.215 ;
        RECT 72.430 186.795 72.600 187.385 ;
        RECT 72.945 187.305 73.485 187.675 ;
        RECT 73.665 187.565 73.885 187.845 ;
        RECT 74.055 187.395 74.225 188.175 ;
        RECT 73.820 187.225 74.225 187.395 ;
        RECT 74.395 187.385 74.745 188.005 ;
        RECT 73.820 187.135 73.990 187.225 ;
        RECT 74.915 187.215 75.125 188.005 ;
        RECT 72.770 186.965 73.990 187.135 ;
        RECT 74.450 187.055 75.125 187.215 ;
        RECT 72.430 186.625 73.230 186.795 ;
        RECT 72.550 186.075 72.880 186.455 ;
        RECT 73.060 186.335 73.230 186.625 ;
        RECT 73.820 186.585 73.990 186.965 ;
        RECT 74.160 187.045 75.125 187.055 ;
        RECT 75.315 187.875 75.575 188.265 ;
        RECT 75.785 188.165 76.115 188.625 ;
        RECT 76.990 188.235 77.845 188.405 ;
        RECT 78.050 188.235 78.545 188.405 ;
        RECT 78.715 188.265 79.045 188.625 ;
        RECT 75.315 187.185 75.485 187.875 ;
        RECT 75.655 187.525 75.825 187.705 ;
        RECT 75.995 187.695 76.785 187.945 ;
        RECT 76.990 187.525 77.160 188.235 ;
        RECT 77.330 187.725 77.685 187.945 ;
        RECT 75.655 187.355 77.345 187.525 ;
        RECT 74.160 186.755 74.620 187.045 ;
        RECT 75.315 187.015 76.815 187.185 ;
        RECT 75.315 186.875 75.485 187.015 ;
        RECT 74.925 186.705 75.485 186.875 ;
        RECT 73.400 186.075 73.650 186.535 ;
        RECT 73.820 186.245 74.690 186.585 ;
        RECT 74.925 186.245 75.095 186.705 ;
        RECT 75.930 186.675 77.005 186.845 ;
        RECT 75.265 186.075 75.635 186.535 ;
        RECT 75.930 186.335 76.100 186.675 ;
        RECT 76.270 186.075 76.600 186.505 ;
        RECT 76.835 186.335 77.005 186.675 ;
        RECT 77.175 186.575 77.345 187.355 ;
        RECT 77.515 187.135 77.685 187.725 ;
        RECT 77.855 187.325 78.205 187.945 ;
        RECT 77.515 186.745 77.980 187.135 ;
        RECT 78.375 186.875 78.545 188.235 ;
        RECT 78.715 187.045 79.175 188.095 ;
        RECT 78.150 186.705 78.545 186.875 ;
        RECT 78.150 186.575 78.320 186.705 ;
        RECT 77.175 186.245 77.855 186.575 ;
        RECT 78.070 186.245 78.320 186.575 ;
        RECT 78.490 186.075 78.740 186.535 ;
        RECT 78.910 186.260 79.235 187.045 ;
        RECT 79.405 186.245 79.575 188.365 ;
        RECT 79.745 188.245 80.075 188.625 ;
        RECT 80.245 188.075 80.500 188.365 ;
        RECT 79.750 187.905 80.500 188.075 ;
        RECT 79.750 186.915 79.980 187.905 ;
        RECT 80.675 187.875 81.885 188.625 ;
        RECT 80.150 187.085 80.500 187.735 ;
        RECT 80.675 187.165 81.195 187.705 ;
        RECT 81.365 187.335 81.885 187.875 ;
        RECT 82.055 187.855 85.565 188.625 ;
        RECT 82.055 187.165 83.745 187.685 ;
        RECT 83.915 187.335 85.565 187.855 ;
        RECT 86.010 187.815 86.255 188.420 ;
        RECT 86.475 188.090 86.985 188.625 ;
        RECT 85.735 187.645 86.965 187.815 ;
        RECT 79.750 186.745 80.500 186.915 ;
        RECT 79.745 186.075 80.075 186.575 ;
        RECT 80.245 186.245 80.500 186.745 ;
        RECT 80.675 186.075 81.885 187.165 ;
        RECT 82.055 186.075 85.565 187.165 ;
        RECT 85.735 186.835 86.075 187.645 ;
        RECT 86.245 187.080 86.995 187.270 ;
        RECT 85.735 186.425 86.250 186.835 ;
        RECT 86.485 186.075 86.655 186.835 ;
        RECT 86.825 186.415 86.995 187.080 ;
        RECT 87.165 187.095 87.355 188.455 ;
        RECT 87.525 187.605 87.800 188.455 ;
        RECT 87.990 188.090 88.520 188.455 ;
        RECT 88.945 188.225 89.275 188.625 ;
        RECT 88.345 188.055 88.520 188.090 ;
        RECT 87.525 187.435 87.805 187.605 ;
        RECT 87.525 187.295 87.800 187.435 ;
        RECT 88.005 187.095 88.175 187.895 ;
        RECT 87.165 186.925 88.175 187.095 ;
        RECT 88.345 187.885 89.275 188.055 ;
        RECT 89.445 187.885 89.700 188.455 ;
        RECT 90.335 187.900 90.625 188.625 ;
        RECT 88.345 186.755 88.515 187.885 ;
        RECT 89.105 187.715 89.275 187.885 ;
        RECT 87.390 186.585 88.515 186.755 ;
        RECT 88.685 187.385 88.880 187.715 ;
        RECT 89.105 187.385 89.360 187.715 ;
        RECT 88.685 186.415 88.855 187.385 ;
        RECT 89.530 187.215 89.700 187.885 ;
        RECT 90.795 187.875 92.005 188.625 ;
        RECT 86.825 186.245 88.855 186.415 ;
        RECT 89.025 186.075 89.195 187.215 ;
        RECT 89.365 186.245 89.700 187.215 ;
        RECT 90.335 186.075 90.625 187.240 ;
        RECT 90.795 187.165 91.315 187.705 ;
        RECT 91.485 187.335 92.005 187.875 ;
        RECT 92.175 187.855 95.685 188.625 ;
        RECT 95.860 188.080 101.205 188.625 ;
        RECT 92.175 187.165 93.865 187.685 ;
        RECT 94.035 187.335 95.685 187.855 ;
        RECT 90.795 186.075 92.005 187.165 ;
        RECT 92.175 186.075 95.685 187.165 ;
        RECT 97.450 186.510 97.800 187.760 ;
        RECT 99.280 187.250 99.620 188.080 ;
        RECT 101.375 187.950 101.635 188.455 ;
        RECT 101.815 188.245 102.145 188.625 ;
        RECT 102.325 188.075 102.495 188.455 ;
        RECT 101.375 187.150 101.545 187.950 ;
        RECT 101.830 187.905 102.495 188.075 ;
        RECT 101.830 187.650 102.000 187.905 ;
        RECT 102.760 187.885 103.015 188.455 ;
        RECT 103.185 188.225 103.515 188.625 ;
        RECT 103.940 188.090 104.470 188.455 ;
        RECT 103.940 188.055 104.115 188.090 ;
        RECT 103.185 187.885 104.115 188.055 ;
        RECT 101.715 187.320 102.000 187.650 ;
        RECT 102.235 187.355 102.565 187.725 ;
        RECT 101.830 187.175 102.000 187.320 ;
        RECT 102.760 187.215 102.930 187.885 ;
        RECT 103.185 187.715 103.355 187.885 ;
        RECT 103.100 187.385 103.355 187.715 ;
        RECT 103.580 187.385 103.775 187.715 ;
        RECT 95.860 186.075 101.205 186.510 ;
        RECT 101.375 186.245 101.645 187.150 ;
        RECT 101.830 187.005 102.495 187.175 ;
        RECT 101.815 186.075 102.145 186.835 ;
        RECT 102.325 186.245 102.495 187.005 ;
        RECT 102.760 186.245 103.095 187.215 ;
        RECT 103.265 186.075 103.435 187.215 ;
        RECT 103.605 186.415 103.775 187.385 ;
        RECT 103.945 186.755 104.115 187.885 ;
        RECT 104.285 187.095 104.455 187.895 ;
        RECT 104.660 187.605 104.935 188.455 ;
        RECT 104.655 187.435 104.935 187.605 ;
        RECT 104.660 187.295 104.935 187.435 ;
        RECT 105.105 187.095 105.295 188.455 ;
        RECT 105.475 188.090 105.985 188.625 ;
        RECT 106.205 187.815 106.450 188.420 ;
        RECT 106.895 187.855 109.485 188.625 ;
        RECT 105.495 187.645 106.725 187.815 ;
        RECT 104.285 186.925 105.295 187.095 ;
        RECT 105.465 187.080 106.215 187.270 ;
        RECT 103.945 186.585 105.070 186.755 ;
        RECT 105.465 186.415 105.635 187.080 ;
        RECT 106.385 186.835 106.725 187.645 ;
        RECT 103.605 186.245 105.635 186.415 ;
        RECT 105.805 186.075 105.975 186.835 ;
        RECT 106.210 186.425 106.725 186.835 ;
        RECT 106.895 187.165 108.105 187.685 ;
        RECT 108.275 187.335 109.485 187.855 ;
        RECT 109.930 187.815 110.175 188.420 ;
        RECT 110.395 188.090 110.905 188.625 ;
        RECT 109.655 187.645 110.885 187.815 ;
        RECT 106.895 186.075 109.485 187.165 ;
        RECT 109.655 186.835 109.995 187.645 ;
        RECT 110.165 187.080 110.915 187.270 ;
        RECT 109.655 186.425 110.170 186.835 ;
        RECT 110.405 186.075 110.575 186.835 ;
        RECT 110.745 186.415 110.915 187.080 ;
        RECT 111.085 187.095 111.275 188.455 ;
        RECT 111.445 188.285 111.720 188.455 ;
        RECT 111.445 188.115 111.725 188.285 ;
        RECT 111.445 187.295 111.720 188.115 ;
        RECT 111.910 188.090 112.440 188.455 ;
        RECT 112.865 188.225 113.195 188.625 ;
        RECT 112.265 188.055 112.440 188.090 ;
        RECT 111.925 187.095 112.095 187.895 ;
        RECT 111.085 186.925 112.095 187.095 ;
        RECT 112.265 187.885 113.195 188.055 ;
        RECT 113.365 187.885 113.620 188.455 ;
        RECT 112.265 186.755 112.435 187.885 ;
        RECT 113.025 187.715 113.195 187.885 ;
        RECT 111.310 186.585 112.435 186.755 ;
        RECT 112.605 187.385 112.800 187.715 ;
        RECT 113.025 187.385 113.280 187.715 ;
        RECT 112.605 186.415 112.775 187.385 ;
        RECT 113.450 187.215 113.620 187.885 ;
        RECT 114.255 187.855 115.925 188.625 ;
        RECT 116.095 187.900 116.385 188.625 ;
        RECT 117.020 188.080 122.365 188.625 ;
        RECT 122.540 188.080 127.885 188.625 ;
        RECT 110.745 186.245 112.775 186.415 ;
        RECT 112.945 186.075 113.115 187.215 ;
        RECT 113.285 186.245 113.620 187.215 ;
        RECT 114.255 187.165 115.005 187.685 ;
        RECT 115.175 187.335 115.925 187.855 ;
        RECT 114.255 186.075 115.925 187.165 ;
        RECT 116.095 186.075 116.385 187.240 ;
        RECT 118.610 186.510 118.960 187.760 ;
        RECT 120.440 187.250 120.780 188.080 ;
        RECT 124.130 186.510 124.480 187.760 ;
        RECT 125.960 187.250 126.300 188.080 ;
        RECT 128.055 187.875 129.265 188.625 ;
        RECT 128.055 187.165 128.575 187.705 ;
        RECT 128.745 187.335 129.265 187.875 ;
        RECT 117.020 186.075 122.365 186.510 ;
        RECT 122.540 186.075 127.885 186.510 ;
        RECT 128.055 186.075 129.265 187.165 ;
        RECT 9.290 185.905 129.350 186.075 ;
        RECT 9.375 184.815 10.585 185.905 ;
        RECT 9.375 184.105 9.895 184.645 ;
        RECT 10.065 184.275 10.585 184.815 ;
        RECT 11.215 184.815 14.725 185.905 ;
        RECT 14.900 185.470 20.245 185.905 ;
        RECT 20.420 185.470 25.765 185.905 ;
        RECT 11.215 184.295 12.905 184.815 ;
        RECT 13.075 184.125 14.725 184.645 ;
        RECT 16.490 184.220 16.840 185.470 ;
        RECT 9.375 183.355 10.585 184.105 ;
        RECT 11.215 183.355 14.725 184.125 ;
        RECT 18.320 183.900 18.660 184.730 ;
        RECT 22.010 184.220 22.360 185.470 ;
        RECT 25.935 184.740 26.225 185.905 ;
        RECT 26.395 185.145 26.910 185.555 ;
        RECT 27.145 185.145 27.315 185.905 ;
        RECT 27.485 185.565 29.515 185.735 ;
        RECT 23.840 183.900 24.180 184.730 ;
        RECT 26.395 184.335 26.735 185.145 ;
        RECT 27.485 184.900 27.655 185.565 ;
        RECT 28.050 185.225 29.175 185.395 ;
        RECT 26.905 184.710 27.655 184.900 ;
        RECT 27.825 184.885 28.835 185.055 ;
        RECT 26.395 184.165 27.625 184.335 ;
        RECT 14.900 183.355 20.245 183.900 ;
        RECT 20.420 183.355 25.765 183.900 ;
        RECT 25.935 183.355 26.225 184.080 ;
        RECT 26.670 183.560 26.915 184.165 ;
        RECT 27.135 183.355 27.645 183.890 ;
        RECT 27.825 183.525 28.015 184.885 ;
        RECT 28.185 183.865 28.460 184.685 ;
        RECT 28.665 184.085 28.835 184.885 ;
        RECT 29.005 184.095 29.175 185.225 ;
        RECT 29.345 184.595 29.515 185.565 ;
        RECT 29.685 184.765 29.855 185.905 ;
        RECT 30.025 184.765 30.360 185.735 ;
        RECT 29.345 184.265 29.540 184.595 ;
        RECT 29.765 184.265 30.020 184.595 ;
        RECT 29.765 184.095 29.935 184.265 ;
        RECT 30.190 184.095 30.360 184.765 ;
        RECT 30.535 184.815 34.045 185.905 ;
        RECT 30.535 184.295 32.225 184.815 ;
        RECT 34.220 184.715 34.475 185.595 ;
        RECT 34.645 184.765 34.950 185.905 ;
        RECT 35.290 185.525 35.620 185.905 ;
        RECT 35.800 185.355 35.970 185.645 ;
        RECT 36.140 185.445 36.390 185.905 ;
        RECT 35.170 185.185 35.970 185.355 ;
        RECT 36.560 185.395 37.430 185.735 ;
        RECT 32.395 184.125 34.045 184.645 ;
        RECT 29.005 183.925 29.935 184.095 ;
        RECT 29.005 183.890 29.180 183.925 ;
        RECT 28.185 183.695 28.465 183.865 ;
        RECT 28.185 183.525 28.460 183.695 ;
        RECT 28.650 183.525 29.180 183.890 ;
        RECT 29.605 183.355 29.935 183.755 ;
        RECT 30.105 183.525 30.360 184.095 ;
        RECT 30.535 183.355 34.045 184.125 ;
        RECT 34.220 184.065 34.430 184.715 ;
        RECT 35.170 184.595 35.340 185.185 ;
        RECT 36.560 185.015 36.730 185.395 ;
        RECT 37.665 185.275 37.835 185.735 ;
        RECT 38.005 185.445 38.375 185.905 ;
        RECT 38.670 185.305 38.840 185.645 ;
        RECT 39.010 185.475 39.340 185.905 ;
        RECT 39.575 185.305 39.745 185.645 ;
        RECT 35.510 184.845 36.730 185.015 ;
        RECT 36.900 184.935 37.360 185.225 ;
        RECT 37.665 185.105 38.225 185.275 ;
        RECT 38.670 185.135 39.745 185.305 ;
        RECT 39.915 185.405 40.595 185.735 ;
        RECT 40.810 185.405 41.060 185.735 ;
        RECT 41.230 185.445 41.480 185.905 ;
        RECT 38.055 184.965 38.225 185.105 ;
        RECT 36.900 184.925 37.865 184.935 ;
        RECT 36.560 184.755 36.730 184.845 ;
        RECT 37.190 184.765 37.865 184.925 ;
        RECT 34.600 184.565 35.340 184.595 ;
        RECT 34.600 184.265 35.515 184.565 ;
        RECT 35.190 184.090 35.515 184.265 ;
        RECT 34.220 183.535 34.475 184.065 ;
        RECT 34.645 183.355 34.950 183.815 ;
        RECT 35.195 183.735 35.515 184.090 ;
        RECT 35.685 184.305 36.225 184.675 ;
        RECT 36.560 184.585 36.965 184.755 ;
        RECT 35.685 183.905 35.925 184.305 ;
        RECT 36.405 184.135 36.625 184.415 ;
        RECT 36.095 183.965 36.625 184.135 ;
        RECT 36.095 183.735 36.265 183.965 ;
        RECT 36.795 183.805 36.965 184.585 ;
        RECT 37.135 183.975 37.485 184.595 ;
        RECT 37.655 183.975 37.865 184.765 ;
        RECT 38.055 184.795 39.555 184.965 ;
        RECT 38.055 184.105 38.225 184.795 ;
        RECT 39.915 184.625 40.085 185.405 ;
        RECT 40.890 185.275 41.060 185.405 ;
        RECT 38.395 184.455 40.085 184.625 ;
        RECT 40.255 184.845 40.720 185.235 ;
        RECT 40.890 185.105 41.285 185.275 ;
        RECT 38.395 184.275 38.565 184.455 ;
        RECT 35.195 183.565 36.265 183.735 ;
        RECT 36.435 183.355 36.625 183.795 ;
        RECT 36.795 183.525 37.745 183.805 ;
        RECT 38.055 183.715 38.315 184.105 ;
        RECT 38.735 184.035 39.525 184.285 ;
        RECT 37.965 183.545 38.315 183.715 ;
        RECT 38.525 183.355 38.855 183.815 ;
        RECT 39.730 183.745 39.900 184.455 ;
        RECT 40.255 184.255 40.425 184.845 ;
        RECT 40.070 184.035 40.425 184.255 ;
        RECT 40.595 184.035 40.945 184.655 ;
        RECT 41.115 183.745 41.285 185.105 ;
        RECT 41.650 184.935 41.975 185.720 ;
        RECT 41.455 183.885 41.915 184.935 ;
        RECT 39.730 183.575 40.585 183.745 ;
        RECT 40.790 183.575 41.285 183.745 ;
        RECT 41.455 183.355 41.785 183.715 ;
        RECT 42.145 183.615 42.315 185.735 ;
        RECT 42.485 185.405 42.815 185.905 ;
        RECT 42.985 185.235 43.240 185.735 ;
        RECT 42.490 185.065 43.240 185.235 ;
        RECT 42.490 184.075 42.720 185.065 ;
        RECT 42.890 184.245 43.240 184.895 ;
        RECT 43.875 184.815 46.465 185.905 ;
        RECT 43.875 184.295 45.085 184.815 ;
        RECT 46.640 184.765 46.975 185.735 ;
        RECT 47.145 184.765 47.315 185.905 ;
        RECT 47.485 185.565 49.515 185.735 ;
        RECT 45.255 184.125 46.465 184.645 ;
        RECT 42.490 183.905 43.240 184.075 ;
        RECT 42.485 183.355 42.815 183.735 ;
        RECT 42.985 183.615 43.240 183.905 ;
        RECT 43.875 183.355 46.465 184.125 ;
        RECT 46.640 184.095 46.810 184.765 ;
        RECT 47.485 184.595 47.655 185.565 ;
        RECT 46.980 184.265 47.235 184.595 ;
        RECT 47.460 184.265 47.655 184.595 ;
        RECT 47.825 185.225 48.950 185.395 ;
        RECT 47.065 184.095 47.235 184.265 ;
        RECT 47.825 184.095 47.995 185.225 ;
        RECT 46.640 183.525 46.895 184.095 ;
        RECT 47.065 183.925 47.995 184.095 ;
        RECT 48.165 184.885 49.175 185.055 ;
        RECT 48.165 184.085 48.335 184.885 ;
        RECT 47.820 183.890 47.995 183.925 ;
        RECT 47.065 183.355 47.395 183.755 ;
        RECT 47.820 183.525 48.350 183.890 ;
        RECT 48.540 183.865 48.815 184.685 ;
        RECT 48.535 183.695 48.815 183.865 ;
        RECT 48.540 183.525 48.815 183.695 ;
        RECT 48.985 183.525 49.175 184.885 ;
        RECT 49.345 184.900 49.515 185.565 ;
        RECT 49.685 185.145 49.855 185.905 ;
        RECT 50.090 185.145 50.605 185.555 ;
        RECT 49.345 184.710 50.095 184.900 ;
        RECT 50.265 184.335 50.605 185.145 ;
        RECT 51.695 184.740 51.985 185.905 ;
        RECT 52.675 184.765 52.885 185.905 ;
        RECT 53.055 184.755 53.385 185.735 ;
        RECT 53.555 184.765 53.785 185.905 ;
        RECT 53.995 184.815 55.205 185.905 ;
        RECT 55.380 185.470 60.725 185.905 ;
        RECT 60.900 185.470 66.245 185.905 ;
        RECT 66.420 185.480 66.755 185.905 ;
        RECT 49.375 184.165 50.605 184.335 ;
        RECT 49.355 183.355 49.865 183.890 ;
        RECT 50.085 183.560 50.330 184.165 ;
        RECT 51.695 183.355 51.985 184.080 ;
        RECT 52.675 183.355 52.885 184.175 ;
        RECT 53.055 184.155 53.305 184.755 ;
        RECT 53.475 184.345 53.805 184.595 ;
        RECT 53.995 184.275 54.515 184.815 ;
        RECT 53.055 183.525 53.385 184.155 ;
        RECT 53.555 183.355 53.785 184.175 ;
        RECT 54.685 184.105 55.205 184.645 ;
        RECT 56.970 184.220 57.320 185.470 ;
        RECT 53.995 183.355 55.205 184.105 ;
        RECT 58.800 183.900 59.140 184.730 ;
        RECT 62.490 184.220 62.840 185.470 ;
        RECT 66.925 185.300 67.110 185.705 ;
        RECT 66.445 185.125 67.110 185.300 ;
        RECT 67.315 185.125 67.645 185.905 ;
        RECT 64.320 183.900 64.660 184.730 ;
        RECT 66.445 184.095 66.785 185.125 ;
        RECT 67.815 184.935 68.085 185.705 ;
        RECT 66.955 184.765 68.085 184.935 ;
        RECT 66.955 184.265 67.205 184.765 ;
        RECT 66.445 183.925 67.130 184.095 ;
        RECT 67.385 184.015 67.745 184.595 ;
        RECT 55.380 183.355 60.725 183.900 ;
        RECT 60.900 183.355 66.245 183.900 ;
        RECT 66.420 183.355 66.755 183.755 ;
        RECT 66.925 183.525 67.130 183.925 ;
        RECT 67.915 183.855 68.085 184.765 ;
        RECT 67.340 183.355 67.615 183.835 ;
        RECT 67.825 183.525 68.085 183.855 ;
        RECT 68.255 184.765 68.515 185.735 ;
        RECT 68.710 185.495 69.040 185.905 ;
        RECT 69.240 185.315 69.410 185.735 ;
        RECT 69.625 185.495 70.295 185.905 ;
        RECT 70.530 185.315 70.700 185.735 ;
        RECT 71.005 185.465 71.335 185.905 ;
        RECT 68.685 185.145 70.700 185.315 ;
        RECT 71.505 185.285 71.680 185.735 ;
        RECT 68.255 184.075 68.425 184.765 ;
        RECT 68.685 184.595 68.855 185.145 ;
        RECT 68.595 184.265 68.855 184.595 ;
        RECT 68.255 183.610 68.595 184.075 ;
        RECT 69.025 183.935 69.365 184.965 ;
        RECT 69.555 183.865 69.825 184.965 ;
        RECT 68.260 183.565 68.595 183.610 ;
        RECT 68.765 183.355 69.095 183.735 ;
        RECT 69.555 183.695 69.865 183.865 ;
        RECT 69.555 183.690 69.825 183.695 ;
        RECT 70.050 183.690 70.330 184.965 ;
        RECT 70.530 183.855 70.700 185.145 ;
        RECT 71.050 185.115 71.680 185.285 ;
        RECT 71.050 184.595 71.220 185.115 ;
        RECT 70.870 184.265 71.220 184.595 ;
        RECT 71.400 184.265 71.765 184.945 ;
        RECT 71.935 184.815 73.605 185.905 ;
        RECT 73.865 184.975 74.035 185.735 ;
        RECT 74.215 185.145 74.545 185.905 ;
        RECT 71.935 184.295 72.685 184.815 ;
        RECT 73.865 184.805 74.530 184.975 ;
        RECT 74.715 184.830 74.985 185.735 ;
        RECT 74.360 184.660 74.530 184.805 ;
        RECT 71.050 184.095 71.220 184.265 ;
        RECT 72.855 184.125 73.605 184.645 ;
        RECT 73.795 184.255 74.125 184.625 ;
        RECT 74.360 184.330 74.645 184.660 ;
        RECT 71.050 183.925 71.680 184.095 ;
        RECT 70.530 183.525 70.760 183.855 ;
        RECT 71.005 183.355 71.335 183.735 ;
        RECT 71.505 183.525 71.680 183.925 ;
        RECT 71.935 183.355 73.605 184.125 ;
        RECT 74.360 184.075 74.530 184.330 ;
        RECT 73.865 183.905 74.530 184.075 ;
        RECT 74.815 184.030 74.985 184.830 ;
        RECT 75.215 184.765 75.425 185.905 ;
        RECT 75.595 184.755 75.925 185.735 ;
        RECT 76.095 184.765 76.325 185.905 ;
        RECT 73.865 183.525 74.035 183.905 ;
        RECT 74.215 183.355 74.545 183.735 ;
        RECT 74.725 183.525 74.985 184.030 ;
        RECT 75.215 183.355 75.425 184.175 ;
        RECT 75.595 184.155 75.845 184.755 ;
        RECT 77.455 184.740 77.745 185.905 ;
        RECT 78.375 184.815 80.965 185.905 ;
        RECT 81.140 185.470 86.485 185.905 ;
        RECT 76.015 184.345 76.345 184.595 ;
        RECT 78.375 184.295 79.585 184.815 ;
        RECT 75.595 183.525 75.925 184.155 ;
        RECT 76.095 183.355 76.325 184.175 ;
        RECT 79.755 184.125 80.965 184.645 ;
        RECT 82.730 184.220 83.080 185.470 ;
        RECT 86.655 185.145 87.170 185.555 ;
        RECT 87.405 185.145 87.575 185.905 ;
        RECT 87.745 185.565 89.775 185.735 ;
        RECT 77.455 183.355 77.745 184.080 ;
        RECT 78.375 183.355 80.965 184.125 ;
        RECT 84.560 183.900 84.900 184.730 ;
        RECT 86.655 184.335 86.995 185.145 ;
        RECT 87.745 184.900 87.915 185.565 ;
        RECT 88.310 185.225 89.435 185.395 ;
        RECT 87.165 184.710 87.915 184.900 ;
        RECT 88.085 184.885 89.095 185.055 ;
        RECT 86.655 184.165 87.885 184.335 ;
        RECT 81.140 183.355 86.485 183.900 ;
        RECT 86.930 183.560 87.175 184.165 ;
        RECT 87.395 183.355 87.905 183.890 ;
        RECT 88.085 183.525 88.275 184.885 ;
        RECT 88.445 183.865 88.720 184.685 ;
        RECT 88.925 184.085 89.095 184.885 ;
        RECT 89.265 184.095 89.435 185.225 ;
        RECT 89.605 184.595 89.775 185.565 ;
        RECT 89.945 184.765 90.115 185.905 ;
        RECT 90.285 184.765 90.620 185.735 ;
        RECT 89.605 184.265 89.800 184.595 ;
        RECT 90.025 184.265 90.280 184.595 ;
        RECT 90.025 184.095 90.195 184.265 ;
        RECT 90.450 184.095 90.620 184.765 ;
        RECT 90.795 184.815 92.005 185.905 ;
        RECT 92.175 184.815 95.685 185.905 ;
        RECT 95.855 185.145 96.370 185.555 ;
        RECT 96.605 185.145 96.775 185.905 ;
        RECT 96.945 185.565 98.975 185.735 ;
        RECT 90.795 184.275 91.315 184.815 ;
        RECT 91.485 184.105 92.005 184.645 ;
        RECT 92.175 184.295 93.865 184.815 ;
        RECT 94.035 184.125 95.685 184.645 ;
        RECT 95.855 184.335 96.195 185.145 ;
        RECT 96.945 184.900 97.115 185.565 ;
        RECT 97.510 185.225 98.635 185.395 ;
        RECT 96.365 184.710 97.115 184.900 ;
        RECT 97.285 184.885 98.295 185.055 ;
        RECT 95.855 184.165 97.085 184.335 ;
        RECT 89.265 183.925 90.195 184.095 ;
        RECT 89.265 183.890 89.440 183.925 ;
        RECT 88.445 183.695 88.725 183.865 ;
        RECT 88.445 183.525 88.720 183.695 ;
        RECT 88.910 183.525 89.440 183.890 ;
        RECT 89.865 183.355 90.195 183.755 ;
        RECT 90.365 183.525 90.620 184.095 ;
        RECT 90.795 183.355 92.005 184.105 ;
        RECT 92.175 183.355 95.685 184.125 ;
        RECT 96.130 183.560 96.375 184.165 ;
        RECT 96.595 183.355 97.105 183.890 ;
        RECT 97.285 183.525 97.475 184.885 ;
        RECT 97.645 184.205 97.920 184.685 ;
        RECT 97.645 184.035 97.925 184.205 ;
        RECT 98.125 184.085 98.295 184.885 ;
        RECT 98.465 184.095 98.635 185.225 ;
        RECT 98.805 184.595 98.975 185.565 ;
        RECT 99.145 184.765 99.315 185.905 ;
        RECT 99.485 184.765 99.820 185.735 ;
        RECT 98.805 184.265 99.000 184.595 ;
        RECT 99.225 184.265 99.480 184.595 ;
        RECT 99.225 184.095 99.395 184.265 ;
        RECT 99.650 184.095 99.820 184.765 ;
        RECT 100.455 184.815 103.045 185.905 ;
        RECT 100.455 184.295 101.665 184.815 ;
        RECT 103.215 184.740 103.505 185.905 ;
        RECT 103.675 184.815 105.345 185.905 ;
        RECT 105.520 185.470 110.865 185.905 ;
        RECT 111.040 185.470 116.385 185.905 ;
        RECT 101.835 184.125 103.045 184.645 ;
        RECT 103.675 184.295 104.425 184.815 ;
        RECT 104.595 184.125 105.345 184.645 ;
        RECT 107.110 184.220 107.460 185.470 ;
        RECT 97.645 183.525 97.920 184.035 ;
        RECT 98.465 183.925 99.395 184.095 ;
        RECT 98.465 183.890 98.640 183.925 ;
        RECT 98.110 183.525 98.640 183.890 ;
        RECT 99.065 183.355 99.395 183.755 ;
        RECT 99.565 183.525 99.820 184.095 ;
        RECT 100.455 183.355 103.045 184.125 ;
        RECT 103.215 183.355 103.505 184.080 ;
        RECT 103.675 183.355 105.345 184.125 ;
        RECT 108.940 183.900 109.280 184.730 ;
        RECT 112.630 184.220 112.980 185.470 ;
        RECT 116.595 184.765 116.825 185.905 ;
        RECT 116.995 184.755 117.325 185.735 ;
        RECT 117.495 184.765 117.705 185.905 ;
        RECT 117.975 184.765 118.205 185.905 ;
        RECT 118.375 184.755 118.705 185.735 ;
        RECT 118.875 184.765 119.085 185.905 ;
        RECT 120.325 184.975 120.495 185.735 ;
        RECT 120.675 185.145 121.005 185.905 ;
        RECT 120.325 184.805 120.990 184.975 ;
        RECT 121.175 184.830 121.445 185.735 ;
        RECT 122.540 185.470 127.885 185.905 ;
        RECT 114.460 183.900 114.800 184.730 ;
        RECT 116.575 184.345 116.905 184.595 ;
        RECT 105.520 183.355 110.865 183.900 ;
        RECT 111.040 183.355 116.385 183.900 ;
        RECT 116.595 183.355 116.825 184.175 ;
        RECT 117.075 184.155 117.325 184.755 ;
        RECT 117.955 184.345 118.285 184.595 ;
        RECT 116.995 183.525 117.325 184.155 ;
        RECT 117.495 183.355 117.705 184.175 ;
        RECT 117.975 183.355 118.205 184.175 ;
        RECT 118.455 184.155 118.705 184.755 ;
        RECT 120.820 184.660 120.990 184.805 ;
        RECT 120.255 184.255 120.585 184.625 ;
        RECT 120.820 184.330 121.105 184.660 ;
        RECT 118.375 183.525 118.705 184.155 ;
        RECT 118.875 183.355 119.085 184.175 ;
        RECT 120.820 184.075 120.990 184.330 ;
        RECT 120.325 183.905 120.990 184.075 ;
        RECT 121.275 184.030 121.445 184.830 ;
        RECT 124.130 184.220 124.480 185.470 ;
        RECT 128.055 184.815 129.265 185.905 ;
        RECT 120.325 183.525 120.495 183.905 ;
        RECT 120.675 183.355 121.005 183.735 ;
        RECT 121.185 183.525 121.445 184.030 ;
        RECT 125.960 183.900 126.300 184.730 ;
        RECT 128.055 184.275 128.575 184.815 ;
        RECT 128.745 184.105 129.265 184.645 ;
        RECT 122.540 183.355 127.885 183.900 ;
        RECT 128.055 183.355 129.265 184.105 ;
        RECT 9.290 183.185 129.350 183.355 ;
        RECT 9.375 182.435 10.585 183.185 ;
        RECT 9.375 181.895 9.895 182.435 ;
        RECT 11.215 182.415 12.885 183.185 ;
        RECT 13.055 182.460 13.345 183.185 ;
        RECT 13.975 182.415 15.645 183.185 ;
        RECT 15.820 182.640 21.165 183.185 ;
        RECT 10.065 181.725 10.585 182.265 ;
        RECT 9.375 180.635 10.585 181.725 ;
        RECT 11.215 181.725 11.965 182.245 ;
        RECT 12.135 181.895 12.885 182.415 ;
        RECT 11.215 180.635 12.885 181.725 ;
        RECT 13.055 180.635 13.345 181.800 ;
        RECT 13.975 181.725 14.725 182.245 ;
        RECT 14.895 181.895 15.645 182.415 ;
        RECT 13.975 180.635 15.645 181.725 ;
        RECT 17.410 181.070 17.760 182.320 ;
        RECT 19.240 181.810 19.580 182.640 ;
        RECT 21.375 182.365 21.605 183.185 ;
        RECT 21.775 182.385 22.105 183.015 ;
        RECT 21.355 181.945 21.685 182.195 ;
        RECT 21.855 181.785 22.105 182.385 ;
        RECT 22.275 182.365 22.485 183.185 ;
        RECT 22.715 182.415 26.225 183.185 ;
        RECT 15.820 180.635 21.165 181.070 ;
        RECT 21.375 180.635 21.605 181.775 ;
        RECT 21.775 180.805 22.105 181.785 ;
        RECT 22.275 180.635 22.485 181.775 ;
        RECT 22.715 181.725 24.405 182.245 ;
        RECT 24.575 181.895 26.225 182.415 ;
        RECT 26.395 182.510 26.655 183.015 ;
        RECT 26.835 182.805 27.165 183.185 ;
        RECT 27.345 182.635 27.515 183.015 ;
        RECT 22.715 180.635 26.225 181.725 ;
        RECT 26.395 181.710 26.565 182.510 ;
        RECT 26.850 182.465 27.515 182.635 ;
        RECT 26.850 182.210 27.020 182.465 ;
        RECT 27.775 182.415 30.365 183.185 ;
        RECT 30.540 182.640 35.885 183.185 ;
        RECT 26.735 181.880 27.020 182.210 ;
        RECT 27.255 181.915 27.585 182.285 ;
        RECT 26.850 181.735 27.020 181.880 ;
        RECT 26.395 180.805 26.665 181.710 ;
        RECT 26.850 181.565 27.515 181.735 ;
        RECT 26.835 180.635 27.165 181.395 ;
        RECT 27.345 180.805 27.515 181.565 ;
        RECT 27.775 181.725 28.985 182.245 ;
        RECT 29.155 181.895 30.365 182.415 ;
        RECT 27.775 180.635 30.365 181.725 ;
        RECT 32.130 181.070 32.480 182.320 ;
        RECT 33.960 181.810 34.300 182.640 ;
        RECT 36.095 182.365 36.325 183.185 ;
        RECT 36.495 182.385 36.825 183.015 ;
        RECT 36.075 181.945 36.405 182.195 ;
        RECT 36.575 181.785 36.825 182.385 ;
        RECT 36.995 182.365 37.205 183.185 ;
        RECT 37.525 182.635 37.695 183.015 ;
        RECT 37.875 182.805 38.205 183.185 ;
        RECT 37.525 182.465 38.190 182.635 ;
        RECT 38.385 182.510 38.645 183.015 ;
        RECT 37.455 181.915 37.785 182.285 ;
        RECT 38.020 182.210 38.190 182.465 ;
        RECT 30.540 180.635 35.885 181.070 ;
        RECT 36.095 180.635 36.325 181.775 ;
        RECT 36.495 180.805 36.825 181.785 ;
        RECT 38.020 181.880 38.305 182.210 ;
        RECT 36.995 180.635 37.205 181.775 ;
        RECT 38.020 181.735 38.190 181.880 ;
        RECT 37.525 181.565 38.190 181.735 ;
        RECT 38.475 181.710 38.645 182.510 ;
        RECT 38.815 182.460 39.105 183.185 ;
        RECT 39.280 182.445 39.535 183.015 ;
        RECT 39.705 182.785 40.035 183.185 ;
        RECT 40.460 182.650 40.990 183.015 ;
        RECT 41.180 182.845 41.455 183.015 ;
        RECT 41.175 182.675 41.455 182.845 ;
        RECT 40.460 182.615 40.635 182.650 ;
        RECT 39.705 182.445 40.635 182.615 ;
        RECT 37.525 180.805 37.695 181.565 ;
        RECT 37.875 180.635 38.205 181.395 ;
        RECT 38.375 180.805 38.645 181.710 ;
        RECT 38.815 180.635 39.105 181.800 ;
        RECT 39.280 181.775 39.450 182.445 ;
        RECT 39.705 182.275 39.875 182.445 ;
        RECT 39.620 181.945 39.875 182.275 ;
        RECT 40.100 181.945 40.295 182.275 ;
        RECT 39.280 180.805 39.615 181.775 ;
        RECT 39.785 180.635 39.955 181.775 ;
        RECT 40.125 180.975 40.295 181.945 ;
        RECT 40.465 181.315 40.635 182.445 ;
        RECT 40.805 181.655 40.975 182.455 ;
        RECT 41.180 181.855 41.455 182.675 ;
        RECT 41.625 181.655 41.815 183.015 ;
        RECT 41.995 182.650 42.505 183.185 ;
        RECT 42.725 182.375 42.970 182.980 ;
        RECT 43.880 182.640 49.225 183.185 ;
        RECT 42.015 182.205 43.245 182.375 ;
        RECT 40.805 181.485 41.815 181.655 ;
        RECT 41.985 181.640 42.735 181.830 ;
        RECT 40.465 181.145 41.590 181.315 ;
        RECT 41.985 180.975 42.155 181.640 ;
        RECT 42.905 181.395 43.245 182.205 ;
        RECT 40.125 180.805 42.155 180.975 ;
        RECT 42.325 180.635 42.495 181.395 ;
        RECT 42.730 180.985 43.245 181.395 ;
        RECT 45.470 181.070 45.820 182.320 ;
        RECT 47.300 181.810 47.640 182.640 ;
        RECT 49.400 182.475 49.655 183.005 ;
        RECT 49.825 182.725 50.130 183.185 ;
        RECT 50.375 182.805 51.445 182.975 ;
        RECT 49.400 181.825 49.610 182.475 ;
        RECT 50.375 182.450 50.695 182.805 ;
        RECT 50.370 182.275 50.695 182.450 ;
        RECT 49.780 181.975 50.695 182.275 ;
        RECT 50.865 182.235 51.105 182.635 ;
        RECT 51.275 182.575 51.445 182.805 ;
        RECT 51.615 182.745 51.805 183.185 ;
        RECT 51.975 182.735 52.925 183.015 ;
        RECT 53.145 182.825 53.495 182.995 ;
        RECT 51.275 182.405 51.805 182.575 ;
        RECT 49.780 181.945 50.520 181.975 ;
        RECT 43.880 180.635 49.225 181.070 ;
        RECT 49.400 180.945 49.655 181.825 ;
        RECT 49.825 180.635 50.130 181.775 ;
        RECT 50.350 181.355 50.520 181.945 ;
        RECT 50.865 181.865 51.405 182.235 ;
        RECT 51.585 182.125 51.805 182.405 ;
        RECT 51.975 181.955 52.145 182.735 ;
        RECT 51.740 181.785 52.145 181.955 ;
        RECT 52.315 181.945 52.665 182.565 ;
        RECT 51.740 181.695 51.910 181.785 ;
        RECT 52.835 181.775 53.045 182.565 ;
        RECT 50.690 181.525 51.910 181.695 ;
        RECT 52.370 181.615 53.045 181.775 ;
        RECT 50.350 181.185 51.150 181.355 ;
        RECT 50.470 180.635 50.800 181.015 ;
        RECT 50.980 180.895 51.150 181.185 ;
        RECT 51.740 181.145 51.910 181.525 ;
        RECT 52.080 181.605 53.045 181.615 ;
        RECT 53.235 182.435 53.495 182.825 ;
        RECT 53.705 182.725 54.035 183.185 ;
        RECT 54.910 182.795 55.765 182.965 ;
        RECT 55.970 182.795 56.465 182.965 ;
        RECT 56.635 182.825 56.965 183.185 ;
        RECT 53.235 181.745 53.405 182.435 ;
        RECT 53.575 182.085 53.745 182.265 ;
        RECT 53.915 182.255 54.705 182.505 ;
        RECT 54.910 182.085 55.080 182.795 ;
        RECT 55.250 182.285 55.605 182.505 ;
        RECT 53.575 181.915 55.265 182.085 ;
        RECT 52.080 181.315 52.540 181.605 ;
        RECT 53.235 181.575 54.735 181.745 ;
        RECT 53.235 181.435 53.405 181.575 ;
        RECT 52.845 181.265 53.405 181.435 ;
        RECT 51.320 180.635 51.570 181.095 ;
        RECT 51.740 180.805 52.610 181.145 ;
        RECT 52.845 180.805 53.015 181.265 ;
        RECT 53.850 181.235 54.925 181.405 ;
        RECT 53.185 180.635 53.555 181.095 ;
        RECT 53.850 180.895 54.020 181.235 ;
        RECT 54.190 180.635 54.520 181.065 ;
        RECT 54.755 180.895 54.925 181.235 ;
        RECT 55.095 181.135 55.265 181.915 ;
        RECT 55.435 181.695 55.605 182.285 ;
        RECT 55.775 181.885 56.125 182.505 ;
        RECT 55.435 181.305 55.900 181.695 ;
        RECT 56.295 181.435 56.465 182.795 ;
        RECT 56.635 181.605 57.095 182.655 ;
        RECT 56.070 181.265 56.465 181.435 ;
        RECT 56.070 181.135 56.240 181.265 ;
        RECT 55.095 180.805 55.775 181.135 ;
        RECT 55.990 180.805 56.240 181.135 ;
        RECT 56.410 180.635 56.660 181.095 ;
        RECT 56.830 180.820 57.155 181.605 ;
        RECT 57.325 180.805 57.495 182.925 ;
        RECT 57.665 182.805 57.995 183.185 ;
        RECT 58.165 182.635 58.420 182.925 ;
        RECT 59.060 182.640 64.405 183.185 ;
        RECT 57.670 182.465 58.420 182.635 ;
        RECT 57.670 181.475 57.900 182.465 ;
        RECT 58.070 181.645 58.420 182.295 ;
        RECT 57.670 181.305 58.420 181.475 ;
        RECT 57.665 180.635 57.995 181.135 ;
        RECT 58.165 180.805 58.420 181.305 ;
        RECT 60.650 181.070 61.000 182.320 ;
        RECT 62.480 181.810 62.820 182.640 ;
        RECT 64.575 182.460 64.865 183.185 ;
        RECT 65.960 182.785 66.295 183.185 ;
        RECT 66.465 182.615 66.670 183.015 ;
        RECT 66.880 182.705 67.155 183.185 ;
        RECT 67.365 182.685 67.625 183.015 ;
        RECT 65.985 182.445 66.670 182.615 ;
        RECT 59.060 180.635 64.405 181.070 ;
        RECT 64.575 180.635 64.865 181.800 ;
        RECT 65.985 181.415 66.325 182.445 ;
        RECT 66.495 181.775 66.745 182.275 ;
        RECT 66.925 181.945 67.285 182.525 ;
        RECT 67.455 181.775 67.625 182.685 ;
        RECT 66.495 181.605 67.625 181.775 ;
        RECT 65.985 181.240 66.650 181.415 ;
        RECT 65.960 180.635 66.295 181.060 ;
        RECT 66.465 180.835 66.650 181.240 ;
        RECT 66.855 180.635 67.185 181.415 ;
        RECT 67.355 180.835 67.625 181.605 ;
        RECT 67.795 180.805 68.055 183.015 ;
        RECT 68.225 182.805 68.555 183.185 ;
        RECT 68.765 182.275 68.960 182.850 ;
        RECT 69.230 182.275 69.415 182.855 ;
        RECT 68.225 181.355 68.395 182.275 ;
        RECT 68.705 181.945 68.960 182.275 ;
        RECT 69.185 181.945 69.415 182.275 ;
        RECT 69.665 182.845 71.145 183.015 ;
        RECT 69.665 181.945 69.835 182.845 ;
        RECT 70.005 182.345 70.555 182.675 ;
        RECT 70.745 182.515 71.145 182.845 ;
        RECT 71.325 182.805 71.655 183.185 ;
        RECT 71.965 182.685 72.225 183.015 ;
        RECT 68.765 181.635 68.960 181.945 ;
        RECT 69.230 181.635 69.415 181.945 ;
        RECT 70.005 181.355 70.175 182.345 ;
        RECT 70.745 182.035 70.915 182.515 ;
        RECT 71.495 182.325 71.705 182.505 ;
        RECT 71.085 182.155 71.705 182.325 ;
        RECT 68.225 181.185 70.175 181.355 ;
        RECT 70.345 181.865 70.915 182.035 ;
        RECT 72.055 181.985 72.225 182.685 ;
        RECT 73.355 182.365 73.585 183.185 ;
        RECT 73.755 182.385 74.085 183.015 ;
        RECT 70.345 181.355 70.515 181.865 ;
        RECT 71.095 181.815 72.225 181.985 ;
        RECT 73.335 181.945 73.665 182.195 ;
        RECT 71.095 181.695 71.265 181.815 ;
        RECT 70.685 181.525 71.265 181.695 ;
        RECT 70.345 181.185 71.085 181.355 ;
        RECT 71.535 181.315 71.885 181.645 ;
        RECT 68.225 180.635 68.555 181.015 ;
        RECT 68.980 180.805 69.150 181.185 ;
        RECT 69.410 180.635 69.740 181.015 ;
        RECT 69.935 180.805 70.105 181.185 ;
        RECT 70.315 180.635 70.645 181.015 ;
        RECT 70.895 180.805 71.085 181.185 ;
        RECT 72.055 181.135 72.225 181.815 ;
        RECT 73.835 181.785 74.085 182.385 ;
        RECT 74.255 182.365 74.465 183.185 ;
        RECT 74.755 182.365 74.965 183.185 ;
        RECT 75.135 182.385 75.465 183.015 ;
        RECT 71.325 180.635 71.655 181.015 ;
        RECT 71.965 180.805 72.225 181.135 ;
        RECT 73.355 180.635 73.585 181.775 ;
        RECT 73.755 180.805 74.085 181.785 ;
        RECT 75.135 181.785 75.385 182.385 ;
        RECT 75.635 182.365 75.865 183.185 ;
        RECT 76.075 182.435 77.285 183.185 ;
        RECT 75.555 181.945 75.885 182.195 ;
        RECT 74.255 180.635 74.465 181.775 ;
        RECT 74.755 180.635 74.965 181.775 ;
        RECT 75.135 180.805 75.465 181.785 ;
        RECT 75.635 180.635 75.865 181.775 ;
        RECT 76.075 181.725 76.595 182.265 ;
        RECT 76.765 181.895 77.285 182.435 ;
        RECT 77.455 182.415 80.965 183.185 ;
        RECT 77.455 181.725 79.145 182.245 ;
        RECT 79.315 181.895 80.965 182.415 ;
        RECT 81.140 182.475 81.395 183.005 ;
        RECT 81.565 182.725 81.870 183.185 ;
        RECT 82.115 182.805 83.185 182.975 ;
        RECT 81.140 181.825 81.350 182.475 ;
        RECT 82.115 182.450 82.435 182.805 ;
        RECT 82.110 182.275 82.435 182.450 ;
        RECT 81.520 181.975 82.435 182.275 ;
        RECT 82.605 182.235 82.845 182.635 ;
        RECT 83.015 182.575 83.185 182.805 ;
        RECT 83.355 182.745 83.545 183.185 ;
        RECT 83.715 182.735 84.665 183.015 ;
        RECT 84.885 182.825 85.235 182.995 ;
        RECT 83.015 182.405 83.545 182.575 ;
        RECT 81.520 181.945 82.260 181.975 ;
        RECT 76.075 180.635 77.285 181.725 ;
        RECT 77.455 180.635 80.965 181.725 ;
        RECT 81.140 180.945 81.395 181.825 ;
        RECT 81.565 180.635 81.870 181.775 ;
        RECT 82.090 181.355 82.260 181.945 ;
        RECT 82.605 181.865 83.145 182.235 ;
        RECT 83.325 182.125 83.545 182.405 ;
        RECT 83.715 181.955 83.885 182.735 ;
        RECT 83.480 181.785 83.885 181.955 ;
        RECT 84.055 181.945 84.405 182.565 ;
        RECT 83.480 181.695 83.650 181.785 ;
        RECT 84.575 181.775 84.785 182.565 ;
        RECT 82.430 181.525 83.650 181.695 ;
        RECT 84.110 181.615 84.785 181.775 ;
        RECT 82.090 181.185 82.890 181.355 ;
        RECT 82.210 180.635 82.540 181.015 ;
        RECT 82.720 180.895 82.890 181.185 ;
        RECT 83.480 181.145 83.650 181.525 ;
        RECT 83.820 181.605 84.785 181.615 ;
        RECT 84.975 182.435 85.235 182.825 ;
        RECT 85.445 182.725 85.775 183.185 ;
        RECT 86.650 182.795 87.505 182.965 ;
        RECT 87.710 182.795 88.205 182.965 ;
        RECT 88.375 182.825 88.705 183.185 ;
        RECT 84.975 181.745 85.145 182.435 ;
        RECT 85.315 182.085 85.485 182.265 ;
        RECT 85.655 182.255 86.445 182.505 ;
        RECT 86.650 182.085 86.820 182.795 ;
        RECT 86.990 182.285 87.345 182.505 ;
        RECT 85.315 181.915 87.005 182.085 ;
        RECT 83.820 181.315 84.280 181.605 ;
        RECT 84.975 181.575 86.475 181.745 ;
        RECT 84.975 181.435 85.145 181.575 ;
        RECT 84.585 181.265 85.145 181.435 ;
        RECT 83.060 180.635 83.310 181.095 ;
        RECT 83.480 180.805 84.350 181.145 ;
        RECT 84.585 180.805 84.755 181.265 ;
        RECT 85.590 181.235 86.665 181.405 ;
        RECT 84.925 180.635 85.295 181.095 ;
        RECT 85.590 180.895 85.760 181.235 ;
        RECT 85.930 180.635 86.260 181.065 ;
        RECT 86.495 180.895 86.665 181.235 ;
        RECT 86.835 181.135 87.005 181.915 ;
        RECT 87.175 181.695 87.345 182.285 ;
        RECT 87.515 181.885 87.865 182.505 ;
        RECT 87.175 181.305 87.640 181.695 ;
        RECT 88.035 181.435 88.205 182.795 ;
        RECT 88.375 181.605 88.835 182.655 ;
        RECT 87.810 181.265 88.205 181.435 ;
        RECT 87.810 181.135 87.980 181.265 ;
        RECT 86.835 180.805 87.515 181.135 ;
        RECT 87.730 180.805 87.980 181.135 ;
        RECT 88.150 180.635 88.400 181.095 ;
        RECT 88.570 180.820 88.895 181.605 ;
        RECT 89.065 180.805 89.235 182.925 ;
        RECT 89.405 182.805 89.735 183.185 ;
        RECT 89.905 182.635 90.160 182.925 ;
        RECT 89.410 182.465 90.160 182.635 ;
        RECT 89.410 181.475 89.640 182.465 ;
        RECT 90.335 182.460 90.625 183.185 ;
        RECT 90.795 182.510 91.055 183.015 ;
        RECT 91.235 182.805 91.565 183.185 ;
        RECT 91.745 182.635 91.915 183.015 ;
        RECT 89.810 181.645 90.160 182.295 ;
        RECT 89.410 181.305 90.160 181.475 ;
        RECT 89.405 180.635 89.735 181.135 ;
        RECT 89.905 180.805 90.160 181.305 ;
        RECT 90.335 180.635 90.625 181.800 ;
        RECT 90.795 181.710 90.965 182.510 ;
        RECT 91.250 182.465 91.915 182.635 ;
        RECT 92.640 182.475 92.895 183.005 ;
        RECT 93.065 182.725 93.370 183.185 ;
        RECT 93.615 182.805 94.685 182.975 ;
        RECT 91.250 182.210 91.420 182.465 ;
        RECT 91.135 181.880 91.420 182.210 ;
        RECT 91.655 181.915 91.985 182.285 ;
        RECT 91.250 181.735 91.420 181.880 ;
        RECT 92.640 181.825 92.850 182.475 ;
        RECT 93.615 182.450 93.935 182.805 ;
        RECT 93.610 182.275 93.935 182.450 ;
        RECT 93.020 181.975 93.935 182.275 ;
        RECT 94.105 182.235 94.345 182.635 ;
        RECT 94.515 182.575 94.685 182.805 ;
        RECT 94.855 182.745 95.045 183.185 ;
        RECT 95.215 182.735 96.165 183.015 ;
        RECT 96.385 182.825 96.735 182.995 ;
        RECT 94.515 182.405 95.045 182.575 ;
        RECT 93.020 181.945 93.760 181.975 ;
        RECT 90.795 180.805 91.065 181.710 ;
        RECT 91.250 181.565 91.915 181.735 ;
        RECT 91.235 180.635 91.565 181.395 ;
        RECT 91.745 180.805 91.915 181.565 ;
        RECT 92.640 180.945 92.895 181.825 ;
        RECT 93.065 180.635 93.370 181.775 ;
        RECT 93.590 181.355 93.760 181.945 ;
        RECT 94.105 181.865 94.645 182.235 ;
        RECT 94.825 182.125 95.045 182.405 ;
        RECT 95.215 181.955 95.385 182.735 ;
        RECT 94.980 181.785 95.385 181.955 ;
        RECT 95.555 181.945 95.905 182.565 ;
        RECT 94.980 181.695 95.150 181.785 ;
        RECT 96.075 181.775 96.285 182.565 ;
        RECT 93.930 181.525 95.150 181.695 ;
        RECT 95.610 181.615 96.285 181.775 ;
        RECT 93.590 181.185 94.390 181.355 ;
        RECT 93.710 180.635 94.040 181.015 ;
        RECT 94.220 180.895 94.390 181.185 ;
        RECT 94.980 181.145 95.150 181.525 ;
        RECT 95.320 181.605 96.285 181.615 ;
        RECT 96.475 182.435 96.735 182.825 ;
        RECT 96.945 182.725 97.275 183.185 ;
        RECT 98.150 182.795 99.005 182.965 ;
        RECT 99.210 182.795 99.705 182.965 ;
        RECT 99.875 182.825 100.205 183.185 ;
        RECT 96.475 181.745 96.645 182.435 ;
        RECT 96.815 182.085 96.985 182.265 ;
        RECT 97.155 182.255 97.945 182.505 ;
        RECT 98.150 182.085 98.320 182.795 ;
        RECT 98.490 182.285 98.845 182.505 ;
        RECT 96.815 181.915 98.505 182.085 ;
        RECT 95.320 181.315 95.780 181.605 ;
        RECT 96.475 181.575 97.975 181.745 ;
        RECT 96.475 181.435 96.645 181.575 ;
        RECT 96.085 181.265 96.645 181.435 ;
        RECT 94.560 180.635 94.810 181.095 ;
        RECT 94.980 180.805 95.850 181.145 ;
        RECT 96.085 180.805 96.255 181.265 ;
        RECT 97.090 181.235 98.165 181.405 ;
        RECT 96.425 180.635 96.795 181.095 ;
        RECT 97.090 180.895 97.260 181.235 ;
        RECT 97.430 180.635 97.760 181.065 ;
        RECT 97.995 180.895 98.165 181.235 ;
        RECT 98.335 181.135 98.505 181.915 ;
        RECT 98.675 181.695 98.845 182.285 ;
        RECT 99.015 181.885 99.365 182.505 ;
        RECT 98.675 181.305 99.140 181.695 ;
        RECT 99.535 181.435 99.705 182.795 ;
        RECT 99.875 181.605 100.335 182.655 ;
        RECT 99.310 181.265 99.705 181.435 ;
        RECT 99.310 181.135 99.480 181.265 ;
        RECT 98.335 180.805 99.015 181.135 ;
        RECT 99.230 180.805 99.480 181.135 ;
        RECT 99.650 180.635 99.900 181.095 ;
        RECT 100.070 180.820 100.395 181.605 ;
        RECT 100.565 180.805 100.735 182.925 ;
        RECT 100.905 182.805 101.235 183.185 ;
        RECT 101.405 182.635 101.660 182.925 ;
        RECT 100.910 182.465 101.660 182.635 ;
        RECT 100.910 181.475 101.140 182.465 ;
        RECT 102.755 182.415 106.265 183.185 ;
        RECT 106.440 182.640 111.785 183.185 ;
        RECT 101.310 181.645 101.660 182.295 ;
        RECT 102.755 181.725 104.445 182.245 ;
        RECT 104.615 181.895 106.265 182.415 ;
        RECT 100.910 181.305 101.660 181.475 ;
        RECT 100.905 180.635 101.235 181.135 ;
        RECT 101.405 180.805 101.660 181.305 ;
        RECT 102.755 180.635 106.265 181.725 ;
        RECT 108.030 181.070 108.380 182.320 ;
        RECT 109.860 181.810 110.200 182.640 ;
        RECT 112.230 182.375 112.475 182.980 ;
        RECT 112.695 182.650 113.205 183.185 ;
        RECT 111.955 182.205 113.185 182.375 ;
        RECT 111.955 181.395 112.295 182.205 ;
        RECT 112.465 181.640 113.215 181.830 ;
        RECT 106.440 180.635 111.785 181.070 ;
        RECT 111.955 180.985 112.470 181.395 ;
        RECT 112.705 180.635 112.875 181.395 ;
        RECT 113.045 180.975 113.215 181.640 ;
        RECT 113.385 181.655 113.575 183.015 ;
        RECT 113.745 182.505 114.020 183.015 ;
        RECT 114.210 182.650 114.740 183.015 ;
        RECT 115.165 182.785 115.495 183.185 ;
        RECT 114.565 182.615 114.740 182.650 ;
        RECT 113.745 182.335 114.025 182.505 ;
        RECT 113.745 181.855 114.020 182.335 ;
        RECT 114.225 181.655 114.395 182.455 ;
        RECT 113.385 181.485 114.395 181.655 ;
        RECT 114.565 182.445 115.495 182.615 ;
        RECT 115.665 182.445 115.920 183.015 ;
        RECT 116.095 182.460 116.385 183.185 ;
        RECT 116.560 182.475 116.815 183.005 ;
        RECT 116.985 182.725 117.290 183.185 ;
        RECT 117.535 182.805 118.605 182.975 ;
        RECT 114.565 181.315 114.735 182.445 ;
        RECT 115.325 182.275 115.495 182.445 ;
        RECT 113.610 181.145 114.735 181.315 ;
        RECT 114.905 181.945 115.100 182.275 ;
        RECT 115.325 181.945 115.580 182.275 ;
        RECT 114.905 180.975 115.075 181.945 ;
        RECT 115.750 181.775 115.920 182.445 ;
        RECT 116.560 181.825 116.770 182.475 ;
        RECT 117.535 182.450 117.855 182.805 ;
        RECT 117.530 182.275 117.855 182.450 ;
        RECT 116.940 181.975 117.855 182.275 ;
        RECT 118.025 182.235 118.265 182.635 ;
        RECT 118.435 182.575 118.605 182.805 ;
        RECT 118.775 182.745 118.965 183.185 ;
        RECT 119.135 182.735 120.085 183.015 ;
        RECT 120.305 182.825 120.655 182.995 ;
        RECT 118.435 182.405 118.965 182.575 ;
        RECT 116.940 181.945 117.680 181.975 ;
        RECT 113.045 180.805 115.075 180.975 ;
        RECT 115.245 180.635 115.415 181.775 ;
        RECT 115.585 180.805 115.920 181.775 ;
        RECT 116.095 180.635 116.385 181.800 ;
        RECT 116.560 180.945 116.815 181.825 ;
        RECT 116.985 180.635 117.290 181.775 ;
        RECT 117.510 181.355 117.680 181.945 ;
        RECT 118.025 181.865 118.565 182.235 ;
        RECT 118.745 182.125 118.965 182.405 ;
        RECT 119.135 181.955 119.305 182.735 ;
        RECT 118.900 181.785 119.305 181.955 ;
        RECT 119.475 181.945 119.825 182.565 ;
        RECT 118.900 181.695 119.070 181.785 ;
        RECT 119.995 181.775 120.205 182.565 ;
        RECT 117.850 181.525 119.070 181.695 ;
        RECT 119.530 181.615 120.205 181.775 ;
        RECT 117.510 181.185 118.310 181.355 ;
        RECT 117.630 180.635 117.960 181.015 ;
        RECT 118.140 180.895 118.310 181.185 ;
        RECT 118.900 181.145 119.070 181.525 ;
        RECT 119.240 181.605 120.205 181.615 ;
        RECT 120.395 182.435 120.655 182.825 ;
        RECT 120.865 182.725 121.195 183.185 ;
        RECT 122.070 182.795 122.925 182.965 ;
        RECT 123.130 182.795 123.625 182.965 ;
        RECT 123.795 182.825 124.125 183.185 ;
        RECT 120.395 181.745 120.565 182.435 ;
        RECT 120.735 182.085 120.905 182.265 ;
        RECT 121.075 182.255 121.865 182.505 ;
        RECT 122.070 182.085 122.240 182.795 ;
        RECT 122.410 182.285 122.765 182.505 ;
        RECT 120.735 181.915 122.425 182.085 ;
        RECT 119.240 181.315 119.700 181.605 ;
        RECT 120.395 181.575 121.895 181.745 ;
        RECT 120.395 181.435 120.565 181.575 ;
        RECT 120.005 181.265 120.565 181.435 ;
        RECT 118.480 180.635 118.730 181.095 ;
        RECT 118.900 180.805 119.770 181.145 ;
        RECT 120.005 180.805 120.175 181.265 ;
        RECT 121.010 181.235 122.085 181.405 ;
        RECT 120.345 180.635 120.715 181.095 ;
        RECT 121.010 180.895 121.180 181.235 ;
        RECT 121.350 180.635 121.680 181.065 ;
        RECT 121.915 180.895 122.085 181.235 ;
        RECT 122.255 181.135 122.425 181.915 ;
        RECT 122.595 181.695 122.765 182.285 ;
        RECT 122.935 181.885 123.285 182.505 ;
        RECT 122.595 181.305 123.060 181.695 ;
        RECT 123.455 181.435 123.625 182.795 ;
        RECT 123.795 181.605 124.255 182.655 ;
        RECT 123.230 181.265 123.625 181.435 ;
        RECT 123.230 181.135 123.400 181.265 ;
        RECT 122.255 180.805 122.935 181.135 ;
        RECT 123.150 180.805 123.400 181.135 ;
        RECT 123.570 180.635 123.820 181.095 ;
        RECT 123.990 180.820 124.315 181.605 ;
        RECT 124.485 180.805 124.655 182.925 ;
        RECT 124.825 182.805 125.155 183.185 ;
        RECT 125.325 182.635 125.580 182.925 ;
        RECT 124.830 182.465 125.580 182.635 ;
        RECT 124.830 181.475 125.060 182.465 ;
        RECT 126.215 182.415 127.885 183.185 ;
        RECT 128.055 182.435 129.265 183.185 ;
        RECT 125.230 181.645 125.580 182.295 ;
        RECT 126.215 181.725 126.965 182.245 ;
        RECT 127.135 181.895 127.885 182.415 ;
        RECT 128.055 181.725 128.575 182.265 ;
        RECT 128.745 181.895 129.265 182.435 ;
        RECT 124.830 181.305 125.580 181.475 ;
        RECT 124.825 180.635 125.155 181.135 ;
        RECT 125.325 180.805 125.580 181.305 ;
        RECT 126.215 180.635 127.885 181.725 ;
        RECT 128.055 180.635 129.265 181.725 ;
        RECT 9.290 180.465 129.350 180.635 ;
        RECT 9.375 179.375 10.585 180.465 ;
        RECT 11.220 180.030 16.565 180.465 ;
        RECT 9.375 178.665 9.895 179.205 ;
        RECT 10.065 178.835 10.585 179.375 ;
        RECT 12.810 178.780 13.160 180.030 ;
        RECT 16.740 179.795 16.995 180.295 ;
        RECT 17.165 179.965 17.495 180.465 ;
        RECT 16.740 179.625 17.490 179.795 ;
        RECT 9.375 177.915 10.585 178.665 ;
        RECT 14.640 178.460 14.980 179.290 ;
        RECT 16.740 178.805 17.090 179.455 ;
        RECT 17.260 178.635 17.490 179.625 ;
        RECT 16.740 178.465 17.490 178.635 ;
        RECT 11.220 177.915 16.565 178.460 ;
        RECT 16.740 178.175 16.995 178.465 ;
        RECT 17.165 177.915 17.495 178.295 ;
        RECT 17.665 178.175 17.835 180.295 ;
        RECT 18.005 179.495 18.330 180.280 ;
        RECT 18.500 180.005 18.750 180.465 ;
        RECT 18.920 179.965 19.170 180.295 ;
        RECT 19.385 179.965 20.065 180.295 ;
        RECT 18.920 179.835 19.090 179.965 ;
        RECT 18.695 179.665 19.090 179.835 ;
        RECT 18.065 178.445 18.525 179.495 ;
        RECT 18.695 178.305 18.865 179.665 ;
        RECT 19.260 179.405 19.725 179.795 ;
        RECT 19.035 178.595 19.385 179.215 ;
        RECT 19.555 178.815 19.725 179.405 ;
        RECT 19.895 179.185 20.065 179.965 ;
        RECT 20.235 179.865 20.405 180.205 ;
        RECT 20.640 180.035 20.970 180.465 ;
        RECT 21.140 179.865 21.310 180.205 ;
        RECT 21.605 180.005 21.975 180.465 ;
        RECT 20.235 179.695 21.310 179.865 ;
        RECT 22.145 179.835 22.315 180.295 ;
        RECT 22.550 179.955 23.420 180.295 ;
        RECT 23.590 180.005 23.840 180.465 ;
        RECT 21.755 179.665 22.315 179.835 ;
        RECT 21.755 179.525 21.925 179.665 ;
        RECT 20.425 179.355 21.925 179.525 ;
        RECT 22.620 179.495 23.080 179.785 ;
        RECT 19.895 179.015 21.585 179.185 ;
        RECT 19.555 178.595 19.910 178.815 ;
        RECT 20.080 178.305 20.250 179.015 ;
        RECT 20.455 178.595 21.245 178.845 ;
        RECT 21.415 178.835 21.585 179.015 ;
        RECT 21.755 178.665 21.925 179.355 ;
        RECT 18.195 177.915 18.525 178.275 ;
        RECT 18.695 178.135 19.190 178.305 ;
        RECT 19.395 178.135 20.250 178.305 ;
        RECT 21.125 177.915 21.455 178.375 ;
        RECT 21.665 178.275 21.925 178.665 ;
        RECT 22.115 179.485 23.080 179.495 ;
        RECT 23.250 179.575 23.420 179.955 ;
        RECT 24.010 179.915 24.180 180.205 ;
        RECT 24.360 180.085 24.690 180.465 ;
        RECT 24.010 179.745 24.810 179.915 ;
        RECT 22.115 179.325 22.790 179.485 ;
        RECT 23.250 179.405 24.470 179.575 ;
        RECT 22.115 178.535 22.325 179.325 ;
        RECT 23.250 179.315 23.420 179.405 ;
        RECT 22.495 178.535 22.845 179.155 ;
        RECT 23.015 179.145 23.420 179.315 ;
        RECT 23.015 178.365 23.185 179.145 ;
        RECT 23.355 178.695 23.575 178.975 ;
        RECT 23.755 178.865 24.295 179.235 ;
        RECT 24.640 179.155 24.810 179.745 ;
        RECT 25.030 179.325 25.335 180.465 ;
        RECT 25.505 179.275 25.760 180.155 ;
        RECT 25.935 179.300 26.225 180.465 ;
        RECT 26.400 179.325 26.735 180.295 ;
        RECT 26.905 179.325 27.075 180.465 ;
        RECT 27.245 180.125 29.275 180.295 ;
        RECT 24.640 179.125 25.380 179.155 ;
        RECT 23.355 178.525 23.885 178.695 ;
        RECT 21.665 178.105 22.015 178.275 ;
        RECT 22.235 178.085 23.185 178.365 ;
        RECT 23.355 177.915 23.545 178.355 ;
        RECT 23.715 178.295 23.885 178.525 ;
        RECT 24.055 178.465 24.295 178.865 ;
        RECT 24.465 178.825 25.380 179.125 ;
        RECT 24.465 178.650 24.790 178.825 ;
        RECT 24.465 178.295 24.785 178.650 ;
        RECT 25.550 178.625 25.760 179.275 ;
        RECT 26.400 178.655 26.570 179.325 ;
        RECT 27.245 179.155 27.415 180.125 ;
        RECT 26.740 178.825 26.995 179.155 ;
        RECT 27.220 178.825 27.415 179.155 ;
        RECT 27.585 179.785 28.710 179.955 ;
        RECT 26.825 178.655 26.995 178.825 ;
        RECT 27.585 178.655 27.755 179.785 ;
        RECT 23.715 178.125 24.785 178.295 ;
        RECT 25.030 177.915 25.335 178.375 ;
        RECT 25.505 178.095 25.760 178.625 ;
        RECT 25.935 177.915 26.225 178.640 ;
        RECT 26.400 178.085 26.655 178.655 ;
        RECT 26.825 178.485 27.755 178.655 ;
        RECT 27.925 179.445 28.935 179.615 ;
        RECT 27.925 178.645 28.095 179.445 ;
        RECT 28.300 178.765 28.575 179.245 ;
        RECT 28.295 178.595 28.575 178.765 ;
        RECT 27.580 178.450 27.755 178.485 ;
        RECT 26.825 177.915 27.155 178.315 ;
        RECT 27.580 178.085 28.110 178.450 ;
        RECT 28.300 178.085 28.575 178.595 ;
        RECT 28.745 178.085 28.935 179.445 ;
        RECT 29.105 179.460 29.275 180.125 ;
        RECT 29.445 179.705 29.615 180.465 ;
        RECT 29.850 179.705 30.365 180.115 ;
        RECT 29.105 179.270 29.855 179.460 ;
        RECT 30.025 178.895 30.365 179.705 ;
        RECT 29.135 178.725 30.365 178.895 ;
        RECT 30.535 179.325 30.875 180.295 ;
        RECT 31.045 179.325 31.215 180.465 ;
        RECT 31.485 179.665 31.735 180.465 ;
        RECT 32.380 179.495 32.710 180.295 ;
        RECT 33.010 179.665 33.340 180.465 ;
        RECT 33.510 179.495 33.840 180.295 ;
        RECT 31.405 179.325 33.840 179.495 ;
        RECT 34.215 179.325 34.555 180.295 ;
        RECT 34.725 179.325 34.895 180.465 ;
        RECT 35.165 179.665 35.415 180.465 ;
        RECT 36.060 179.495 36.390 180.295 ;
        RECT 36.690 179.665 37.020 180.465 ;
        RECT 37.190 179.495 37.520 180.295 ;
        RECT 35.085 179.325 37.520 179.495 ;
        RECT 38.355 179.375 41.865 180.465 ;
        RECT 42.040 180.030 47.385 180.465 ;
        RECT 30.535 178.765 30.710 179.325 ;
        RECT 31.405 179.075 31.575 179.325 ;
        RECT 30.880 178.905 31.575 179.075 ;
        RECT 31.750 178.905 32.170 179.105 ;
        RECT 32.340 178.905 32.670 179.105 ;
        RECT 32.840 178.905 33.170 179.105 ;
        RECT 29.115 177.915 29.625 178.450 ;
        RECT 29.845 178.120 30.090 178.725 ;
        RECT 30.535 178.715 30.765 178.765 ;
        RECT 30.535 178.085 30.875 178.715 ;
        RECT 31.045 177.915 31.295 178.715 ;
        RECT 31.485 178.565 32.710 178.735 ;
        RECT 31.485 178.085 31.815 178.565 ;
        RECT 31.985 177.915 32.210 178.375 ;
        RECT 32.380 178.085 32.710 178.565 ;
        RECT 33.340 178.695 33.510 179.325 ;
        RECT 33.695 178.905 34.045 179.155 ;
        RECT 34.215 178.765 34.390 179.325 ;
        RECT 35.085 179.075 35.255 179.325 ;
        RECT 34.560 178.905 35.255 179.075 ;
        RECT 35.430 178.905 35.850 179.105 ;
        RECT 36.020 178.905 36.350 179.105 ;
        RECT 36.520 178.905 36.850 179.105 ;
        RECT 34.215 178.715 34.445 178.765 ;
        RECT 33.340 178.085 33.840 178.695 ;
        RECT 34.215 178.085 34.555 178.715 ;
        RECT 34.725 177.915 34.975 178.715 ;
        RECT 35.165 178.565 36.390 178.735 ;
        RECT 35.165 178.085 35.495 178.565 ;
        RECT 35.665 177.915 35.890 178.375 ;
        RECT 36.060 178.085 36.390 178.565 ;
        RECT 37.020 178.695 37.190 179.325 ;
        RECT 37.375 178.905 37.725 179.155 ;
        RECT 38.355 178.855 40.045 179.375 ;
        RECT 37.020 178.085 37.520 178.695 ;
        RECT 40.215 178.685 41.865 179.205 ;
        RECT 43.630 178.780 43.980 180.030 ;
        RECT 47.555 179.705 48.070 180.115 ;
        RECT 48.305 179.705 48.475 180.465 ;
        RECT 48.645 180.125 50.675 180.295 ;
        RECT 38.355 177.915 41.865 178.685 ;
        RECT 45.460 178.460 45.800 179.290 ;
        RECT 47.555 178.895 47.895 179.705 ;
        RECT 48.645 179.460 48.815 180.125 ;
        RECT 49.210 179.785 50.335 179.955 ;
        RECT 48.065 179.270 48.815 179.460 ;
        RECT 48.985 179.445 49.995 179.615 ;
        RECT 47.555 178.725 48.785 178.895 ;
        RECT 42.040 177.915 47.385 178.460 ;
        RECT 47.830 178.120 48.075 178.725 ;
        RECT 48.295 177.915 48.805 178.450 ;
        RECT 48.985 178.085 49.175 179.445 ;
        RECT 49.345 178.425 49.620 179.245 ;
        RECT 49.825 178.645 49.995 179.445 ;
        RECT 50.165 178.655 50.335 179.785 ;
        RECT 50.505 179.155 50.675 180.125 ;
        RECT 50.845 179.325 51.015 180.465 ;
        RECT 51.185 179.325 51.520 180.295 ;
        RECT 50.505 178.825 50.700 179.155 ;
        RECT 50.925 178.825 51.180 179.155 ;
        RECT 50.925 178.655 51.095 178.825 ;
        RECT 51.350 178.655 51.520 179.325 ;
        RECT 51.695 179.300 51.985 180.465 ;
        RECT 53.165 179.535 53.335 180.295 ;
        RECT 53.515 179.705 53.845 180.465 ;
        RECT 53.165 179.365 53.830 179.535 ;
        RECT 54.015 179.390 54.285 180.295 ;
        RECT 54.510 179.595 54.795 180.465 ;
        RECT 54.965 179.835 55.225 180.295 ;
        RECT 55.400 180.005 55.655 180.465 ;
        RECT 55.825 179.835 56.085 180.295 ;
        RECT 54.965 179.665 56.085 179.835 ;
        RECT 56.255 179.665 56.565 180.465 ;
        RECT 54.965 179.415 55.225 179.665 ;
        RECT 56.735 179.495 57.045 180.295 ;
        RECT 57.220 180.030 62.565 180.465 ;
        RECT 62.740 180.030 68.085 180.465 ;
        RECT 53.660 179.220 53.830 179.365 ;
        RECT 53.095 178.815 53.425 179.185 ;
        RECT 53.660 178.890 53.945 179.220 ;
        RECT 50.165 178.485 51.095 178.655 ;
        RECT 50.165 178.450 50.340 178.485 ;
        RECT 49.345 178.255 49.625 178.425 ;
        RECT 49.345 178.085 49.620 178.255 ;
        RECT 49.810 178.085 50.340 178.450 ;
        RECT 50.765 177.915 51.095 178.315 ;
        RECT 51.265 178.085 51.520 178.655 ;
        RECT 51.695 177.915 51.985 178.640 ;
        RECT 53.660 178.635 53.830 178.890 ;
        RECT 53.165 178.465 53.830 178.635 ;
        RECT 54.115 178.590 54.285 179.390 ;
        RECT 53.165 178.085 53.335 178.465 ;
        RECT 53.515 177.915 53.845 178.295 ;
        RECT 54.025 178.085 54.285 178.590 ;
        RECT 54.470 179.245 55.225 179.415 ;
        RECT 56.015 179.325 57.045 179.495 ;
        RECT 54.470 178.735 54.875 179.245 ;
        RECT 56.015 179.075 56.185 179.325 ;
        RECT 55.045 178.905 56.185 179.075 ;
        RECT 54.470 178.565 56.120 178.735 ;
        RECT 56.355 178.585 56.705 179.155 ;
        RECT 54.515 177.915 54.795 178.395 ;
        RECT 54.965 178.175 55.225 178.565 ;
        RECT 55.400 177.915 55.655 178.395 ;
        RECT 55.825 178.175 56.120 178.565 ;
        RECT 56.875 178.415 57.045 179.325 ;
        RECT 58.810 178.780 59.160 180.030 ;
        RECT 60.640 178.460 60.980 179.290 ;
        RECT 64.330 178.780 64.680 180.030 ;
        RECT 66.160 178.460 66.500 179.290 ;
        RECT 68.260 179.275 68.515 180.155 ;
        RECT 68.685 179.325 68.990 180.465 ;
        RECT 69.330 180.085 69.660 180.465 ;
        RECT 69.840 179.915 70.010 180.205 ;
        RECT 70.180 180.005 70.430 180.465 ;
        RECT 69.210 179.745 70.010 179.915 ;
        RECT 70.600 179.955 71.470 180.295 ;
        RECT 68.260 178.625 68.470 179.275 ;
        RECT 69.210 179.155 69.380 179.745 ;
        RECT 70.600 179.575 70.770 179.955 ;
        RECT 71.705 179.835 71.875 180.295 ;
        RECT 72.045 180.005 72.415 180.465 ;
        RECT 72.710 179.865 72.880 180.205 ;
        RECT 73.050 180.035 73.380 180.465 ;
        RECT 73.615 179.865 73.785 180.205 ;
        RECT 69.550 179.405 70.770 179.575 ;
        RECT 70.940 179.495 71.400 179.785 ;
        RECT 71.705 179.665 72.265 179.835 ;
        RECT 72.710 179.695 73.785 179.865 ;
        RECT 73.955 179.965 74.635 180.295 ;
        RECT 74.850 179.965 75.100 180.295 ;
        RECT 75.270 180.005 75.520 180.465 ;
        RECT 72.095 179.525 72.265 179.665 ;
        RECT 70.940 179.485 71.905 179.495 ;
        RECT 70.600 179.315 70.770 179.405 ;
        RECT 71.230 179.325 71.905 179.485 ;
        RECT 68.640 179.125 69.380 179.155 ;
        RECT 68.640 178.825 69.555 179.125 ;
        RECT 69.230 178.650 69.555 178.825 ;
        RECT 56.300 177.915 56.575 178.395 ;
        RECT 56.745 178.085 57.045 178.415 ;
        RECT 57.220 177.915 62.565 178.460 ;
        RECT 62.740 177.915 68.085 178.460 ;
        RECT 68.260 178.095 68.515 178.625 ;
        RECT 68.685 177.915 68.990 178.375 ;
        RECT 69.235 178.295 69.555 178.650 ;
        RECT 69.725 178.865 70.265 179.235 ;
        RECT 70.600 179.145 71.005 179.315 ;
        RECT 69.725 178.465 69.965 178.865 ;
        RECT 70.445 178.695 70.665 178.975 ;
        RECT 70.135 178.525 70.665 178.695 ;
        RECT 70.135 178.295 70.305 178.525 ;
        RECT 70.835 178.365 71.005 179.145 ;
        RECT 71.175 178.535 71.525 179.155 ;
        RECT 71.695 178.535 71.905 179.325 ;
        RECT 72.095 179.355 73.595 179.525 ;
        RECT 72.095 178.665 72.265 179.355 ;
        RECT 73.955 179.185 74.125 179.965 ;
        RECT 74.930 179.835 75.100 179.965 ;
        RECT 72.435 179.015 74.125 179.185 ;
        RECT 74.295 179.405 74.760 179.795 ;
        RECT 74.930 179.665 75.325 179.835 ;
        RECT 72.435 178.835 72.605 179.015 ;
        RECT 69.235 178.125 70.305 178.295 ;
        RECT 70.475 177.915 70.665 178.355 ;
        RECT 70.835 178.085 71.785 178.365 ;
        RECT 72.095 178.275 72.355 178.665 ;
        RECT 72.775 178.595 73.565 178.845 ;
        RECT 72.005 178.105 72.355 178.275 ;
        RECT 72.565 177.915 72.895 178.375 ;
        RECT 73.770 178.305 73.940 179.015 ;
        RECT 74.295 178.815 74.465 179.405 ;
        RECT 74.110 178.595 74.465 178.815 ;
        RECT 74.635 178.595 74.985 179.215 ;
        RECT 75.155 178.305 75.325 179.665 ;
        RECT 75.690 179.495 76.015 180.280 ;
        RECT 75.495 178.445 75.955 179.495 ;
        RECT 73.770 178.135 74.625 178.305 ;
        RECT 74.830 178.135 75.325 178.305 ;
        RECT 75.495 177.915 75.825 178.275 ;
        RECT 76.185 178.175 76.355 180.295 ;
        RECT 76.525 179.965 76.855 180.465 ;
        RECT 77.025 179.795 77.280 180.295 ;
        RECT 76.530 179.625 77.280 179.795 ;
        RECT 76.530 178.635 76.760 179.625 ;
        RECT 76.930 178.805 77.280 179.455 ;
        RECT 77.455 179.300 77.745 180.465 ;
        RECT 78.375 179.375 80.965 180.465 ;
        RECT 81.135 179.495 81.445 180.295 ;
        RECT 81.615 179.665 81.925 180.465 ;
        RECT 82.095 179.835 82.355 180.295 ;
        RECT 82.525 180.005 82.780 180.465 ;
        RECT 82.955 179.835 83.215 180.295 ;
        RECT 82.095 179.665 83.215 179.835 ;
        RECT 78.375 178.855 79.585 179.375 ;
        RECT 81.135 179.325 82.165 179.495 ;
        RECT 79.755 178.685 80.965 179.205 ;
        RECT 76.530 178.465 77.280 178.635 ;
        RECT 76.525 177.915 76.855 178.295 ;
        RECT 77.025 178.175 77.280 178.465 ;
        RECT 77.455 177.915 77.745 178.640 ;
        RECT 78.375 177.915 80.965 178.685 ;
        RECT 81.135 178.415 81.305 179.325 ;
        RECT 81.475 178.585 81.825 179.155 ;
        RECT 81.995 179.075 82.165 179.325 ;
        RECT 82.955 179.415 83.215 179.665 ;
        RECT 83.385 179.595 83.670 180.465 ;
        RECT 82.955 179.245 83.710 179.415 ;
        RECT 81.995 178.905 83.135 179.075 ;
        RECT 83.305 178.735 83.710 179.245 ;
        RECT 83.895 179.375 87.405 180.465 ;
        RECT 83.895 178.855 85.585 179.375 ;
        RECT 87.635 179.325 87.845 180.465 ;
        RECT 88.015 179.315 88.345 180.295 ;
        RECT 88.515 179.325 88.745 180.465 ;
        RECT 89.880 180.030 95.225 180.465 ;
        RECT 82.060 178.565 83.710 178.735 ;
        RECT 85.755 178.685 87.405 179.205 ;
        RECT 81.135 178.085 81.435 178.415 ;
        RECT 81.605 177.915 81.880 178.395 ;
        RECT 82.060 178.175 82.355 178.565 ;
        RECT 82.525 177.915 82.780 178.395 ;
        RECT 82.955 178.175 83.215 178.565 ;
        RECT 83.385 177.915 83.665 178.395 ;
        RECT 83.895 177.915 87.405 178.685 ;
        RECT 87.635 177.915 87.845 178.735 ;
        RECT 88.015 178.715 88.265 179.315 ;
        RECT 88.435 178.905 88.765 179.155 ;
        RECT 91.470 178.780 91.820 180.030 ;
        RECT 95.455 179.325 95.665 180.465 ;
        RECT 95.835 179.315 96.165 180.295 ;
        RECT 96.335 179.325 96.565 180.465 ;
        RECT 97.235 179.375 98.905 180.465 ;
        RECT 99.165 179.535 99.335 180.295 ;
        RECT 99.515 179.705 99.845 180.465 ;
        RECT 88.015 178.085 88.345 178.715 ;
        RECT 88.515 177.915 88.745 178.735 ;
        RECT 93.300 178.460 93.640 179.290 ;
        RECT 89.880 177.915 95.225 178.460 ;
        RECT 95.455 177.915 95.665 178.735 ;
        RECT 95.835 178.715 96.085 179.315 ;
        RECT 96.255 178.905 96.585 179.155 ;
        RECT 97.235 178.855 97.985 179.375 ;
        RECT 99.165 179.365 99.830 179.535 ;
        RECT 100.015 179.390 100.285 180.295 ;
        RECT 99.660 179.220 99.830 179.365 ;
        RECT 95.835 178.085 96.165 178.715 ;
        RECT 96.335 177.915 96.565 178.735 ;
        RECT 98.155 178.685 98.905 179.205 ;
        RECT 99.095 178.815 99.425 179.185 ;
        RECT 99.660 178.890 99.945 179.220 ;
        RECT 97.235 177.915 98.905 178.685 ;
        RECT 99.660 178.635 99.830 178.890 ;
        RECT 99.165 178.465 99.830 178.635 ;
        RECT 100.115 178.590 100.285 179.390 ;
        RECT 100.455 179.375 103.045 180.465 ;
        RECT 100.455 178.855 101.665 179.375 ;
        RECT 103.215 179.300 103.505 180.465 ;
        RECT 103.675 179.375 105.345 180.465 ;
        RECT 101.835 178.685 103.045 179.205 ;
        RECT 103.675 178.855 104.425 179.375 ;
        RECT 105.515 179.325 105.855 180.295 ;
        RECT 106.025 179.325 106.195 180.465 ;
        RECT 106.465 179.665 106.715 180.465 ;
        RECT 107.360 179.495 107.690 180.295 ;
        RECT 107.990 179.665 108.320 180.465 ;
        RECT 108.490 179.495 108.820 180.295 ;
        RECT 106.385 179.325 108.820 179.495 ;
        RECT 109.195 179.375 111.785 180.465 ;
        RECT 111.955 179.705 112.470 180.115 ;
        RECT 112.705 179.705 112.875 180.465 ;
        RECT 113.045 180.125 115.075 180.295 ;
        RECT 104.595 178.685 105.345 179.205 ;
        RECT 99.165 178.085 99.335 178.465 ;
        RECT 99.515 177.915 99.845 178.295 ;
        RECT 100.025 178.085 100.285 178.590 ;
        RECT 100.455 177.915 103.045 178.685 ;
        RECT 103.215 177.915 103.505 178.640 ;
        RECT 103.675 177.915 105.345 178.685 ;
        RECT 105.515 178.765 105.690 179.325 ;
        RECT 106.385 179.075 106.555 179.325 ;
        RECT 105.860 178.905 106.555 179.075 ;
        RECT 106.730 178.905 107.150 179.105 ;
        RECT 107.320 178.905 107.650 179.105 ;
        RECT 107.820 178.905 108.150 179.105 ;
        RECT 105.515 178.715 105.745 178.765 ;
        RECT 105.515 178.085 105.855 178.715 ;
        RECT 106.025 177.915 106.275 178.715 ;
        RECT 106.465 178.565 107.690 178.735 ;
        RECT 106.465 178.085 106.795 178.565 ;
        RECT 106.965 177.915 107.190 178.375 ;
        RECT 107.360 178.085 107.690 178.565 ;
        RECT 108.320 178.695 108.490 179.325 ;
        RECT 108.675 178.905 109.025 179.155 ;
        RECT 109.195 178.855 110.405 179.375 ;
        RECT 108.320 178.085 108.820 178.695 ;
        RECT 110.575 178.685 111.785 179.205 ;
        RECT 111.955 178.895 112.295 179.705 ;
        RECT 113.045 179.460 113.215 180.125 ;
        RECT 113.610 179.785 114.735 179.955 ;
        RECT 112.465 179.270 113.215 179.460 ;
        RECT 113.385 179.445 114.395 179.615 ;
        RECT 111.955 178.725 113.185 178.895 ;
        RECT 109.195 177.915 111.785 178.685 ;
        RECT 112.230 178.120 112.475 178.725 ;
        RECT 112.695 177.915 113.205 178.450 ;
        RECT 113.385 178.085 113.575 179.445 ;
        RECT 113.745 178.425 114.020 179.245 ;
        RECT 114.225 178.645 114.395 179.445 ;
        RECT 114.565 178.655 114.735 179.785 ;
        RECT 114.905 179.155 115.075 180.125 ;
        RECT 115.245 179.325 115.415 180.465 ;
        RECT 115.585 179.325 115.920 180.295 ;
        RECT 114.905 178.825 115.100 179.155 ;
        RECT 115.325 178.825 115.580 179.155 ;
        RECT 115.325 178.655 115.495 178.825 ;
        RECT 115.750 178.655 115.920 179.325 ;
        RECT 114.565 178.485 115.495 178.655 ;
        RECT 114.565 178.450 114.740 178.485 ;
        RECT 113.745 178.255 114.025 178.425 ;
        RECT 113.745 178.085 114.020 178.255 ;
        RECT 114.210 178.085 114.740 178.450 ;
        RECT 115.165 177.915 115.495 178.315 ;
        RECT 115.665 178.085 115.920 178.655 ;
        RECT 116.100 179.275 116.355 180.155 ;
        RECT 116.525 179.325 116.830 180.465 ;
        RECT 117.170 180.085 117.500 180.465 ;
        RECT 117.680 179.915 117.850 180.205 ;
        RECT 118.020 180.005 118.270 180.465 ;
        RECT 117.050 179.745 117.850 179.915 ;
        RECT 118.440 179.955 119.310 180.295 ;
        RECT 116.100 178.625 116.310 179.275 ;
        RECT 117.050 179.155 117.220 179.745 ;
        RECT 118.440 179.575 118.610 179.955 ;
        RECT 119.545 179.835 119.715 180.295 ;
        RECT 119.885 180.005 120.255 180.465 ;
        RECT 120.550 179.865 120.720 180.205 ;
        RECT 120.890 180.035 121.220 180.465 ;
        RECT 121.455 179.865 121.625 180.205 ;
        RECT 117.390 179.405 118.610 179.575 ;
        RECT 118.780 179.495 119.240 179.785 ;
        RECT 119.545 179.665 120.105 179.835 ;
        RECT 120.550 179.695 121.625 179.865 ;
        RECT 121.795 179.965 122.475 180.295 ;
        RECT 122.690 179.965 122.940 180.295 ;
        RECT 123.110 180.005 123.360 180.465 ;
        RECT 119.935 179.525 120.105 179.665 ;
        RECT 118.780 179.485 119.745 179.495 ;
        RECT 118.440 179.315 118.610 179.405 ;
        RECT 119.070 179.325 119.745 179.485 ;
        RECT 116.480 179.125 117.220 179.155 ;
        RECT 116.480 178.825 117.395 179.125 ;
        RECT 117.070 178.650 117.395 178.825 ;
        RECT 116.100 178.095 116.355 178.625 ;
        RECT 116.525 177.915 116.830 178.375 ;
        RECT 117.075 178.295 117.395 178.650 ;
        RECT 117.565 178.865 118.105 179.235 ;
        RECT 118.440 179.145 118.845 179.315 ;
        RECT 117.565 178.465 117.805 178.865 ;
        RECT 118.285 178.695 118.505 178.975 ;
        RECT 117.975 178.525 118.505 178.695 ;
        RECT 117.975 178.295 118.145 178.525 ;
        RECT 118.675 178.365 118.845 179.145 ;
        RECT 119.015 178.535 119.365 179.155 ;
        RECT 119.535 178.535 119.745 179.325 ;
        RECT 119.935 179.355 121.435 179.525 ;
        RECT 119.935 178.665 120.105 179.355 ;
        RECT 121.795 179.185 121.965 179.965 ;
        RECT 122.770 179.835 122.940 179.965 ;
        RECT 120.275 179.015 121.965 179.185 ;
        RECT 122.135 179.405 122.600 179.795 ;
        RECT 122.770 179.665 123.165 179.835 ;
        RECT 120.275 178.835 120.445 179.015 ;
        RECT 117.075 178.125 118.145 178.295 ;
        RECT 118.315 177.915 118.505 178.355 ;
        RECT 118.675 178.085 119.625 178.365 ;
        RECT 119.935 178.275 120.195 178.665 ;
        RECT 120.615 178.595 121.405 178.845 ;
        RECT 119.845 178.105 120.195 178.275 ;
        RECT 120.405 177.915 120.735 178.375 ;
        RECT 121.610 178.305 121.780 179.015 ;
        RECT 122.135 178.815 122.305 179.405 ;
        RECT 121.950 178.595 122.305 178.815 ;
        RECT 122.475 178.595 122.825 179.215 ;
        RECT 122.995 178.305 123.165 179.665 ;
        RECT 123.530 179.495 123.855 180.280 ;
        RECT 123.335 178.445 123.795 179.495 ;
        RECT 121.610 178.135 122.465 178.305 ;
        RECT 122.670 178.135 123.165 178.305 ;
        RECT 123.335 177.915 123.665 178.275 ;
        RECT 124.025 178.175 124.195 180.295 ;
        RECT 124.365 179.965 124.695 180.465 ;
        RECT 124.865 179.795 125.120 180.295 ;
        RECT 124.370 179.625 125.120 179.795 ;
        RECT 124.370 178.635 124.600 179.625 ;
        RECT 124.770 178.805 125.120 179.455 ;
        RECT 125.295 179.375 127.885 180.465 ;
        RECT 128.055 179.375 129.265 180.465 ;
        RECT 125.295 178.855 126.505 179.375 ;
        RECT 126.675 178.685 127.885 179.205 ;
        RECT 128.055 178.835 128.575 179.375 ;
        RECT 124.370 178.465 125.120 178.635 ;
        RECT 124.365 177.915 124.695 178.295 ;
        RECT 124.865 178.175 125.120 178.465 ;
        RECT 125.295 177.915 127.885 178.685 ;
        RECT 128.745 178.665 129.265 179.205 ;
        RECT 128.055 177.915 129.265 178.665 ;
        RECT 9.290 177.745 129.350 177.915 ;
        RECT 9.375 176.995 10.585 177.745 ;
        RECT 9.375 176.455 9.895 176.995 ;
        RECT 11.215 176.975 12.885 177.745 ;
        RECT 13.055 177.020 13.345 177.745 ;
        RECT 13.975 176.975 15.645 177.745 ;
        RECT 15.820 177.200 21.165 177.745 ;
        RECT 10.065 176.285 10.585 176.825 ;
        RECT 9.375 175.195 10.585 176.285 ;
        RECT 11.215 176.285 11.965 176.805 ;
        RECT 12.135 176.455 12.885 176.975 ;
        RECT 11.215 175.195 12.885 176.285 ;
        RECT 13.055 175.195 13.345 176.360 ;
        RECT 13.975 176.285 14.725 176.805 ;
        RECT 14.895 176.455 15.645 176.975 ;
        RECT 13.975 175.195 15.645 176.285 ;
        RECT 17.410 175.630 17.760 176.880 ;
        RECT 19.240 176.370 19.580 177.200 ;
        RECT 21.375 176.925 21.605 177.745 ;
        RECT 21.775 176.945 22.105 177.575 ;
        RECT 21.355 176.505 21.685 176.755 ;
        RECT 21.855 176.345 22.105 176.945 ;
        RECT 22.275 176.925 22.485 177.745 ;
        RECT 22.720 177.035 22.975 177.565 ;
        RECT 23.145 177.285 23.450 177.745 ;
        RECT 23.695 177.365 24.765 177.535 ;
        RECT 15.820 175.195 21.165 175.630 ;
        RECT 21.375 175.195 21.605 176.335 ;
        RECT 21.775 175.365 22.105 176.345 ;
        RECT 22.720 176.385 22.930 177.035 ;
        RECT 23.695 177.010 24.015 177.365 ;
        RECT 23.690 176.835 24.015 177.010 ;
        RECT 23.100 176.535 24.015 176.835 ;
        RECT 24.185 176.795 24.425 177.195 ;
        RECT 24.595 177.135 24.765 177.365 ;
        RECT 24.935 177.305 25.125 177.745 ;
        RECT 25.295 177.295 26.245 177.575 ;
        RECT 26.465 177.385 26.815 177.555 ;
        RECT 24.595 176.965 25.125 177.135 ;
        RECT 23.100 176.505 23.840 176.535 ;
        RECT 22.275 175.195 22.485 176.335 ;
        RECT 22.720 175.505 22.975 176.385 ;
        RECT 23.145 175.195 23.450 176.335 ;
        RECT 23.670 175.915 23.840 176.505 ;
        RECT 24.185 176.425 24.725 176.795 ;
        RECT 24.905 176.685 25.125 176.965 ;
        RECT 25.295 176.515 25.465 177.295 ;
        RECT 25.060 176.345 25.465 176.515 ;
        RECT 25.635 176.505 25.985 177.125 ;
        RECT 25.060 176.255 25.230 176.345 ;
        RECT 26.155 176.335 26.365 177.125 ;
        RECT 24.010 176.085 25.230 176.255 ;
        RECT 25.690 176.175 26.365 176.335 ;
        RECT 23.670 175.745 24.470 175.915 ;
        RECT 23.790 175.195 24.120 175.575 ;
        RECT 24.300 175.455 24.470 175.745 ;
        RECT 25.060 175.705 25.230 176.085 ;
        RECT 25.400 176.165 26.365 176.175 ;
        RECT 26.555 176.995 26.815 177.385 ;
        RECT 27.025 177.285 27.355 177.745 ;
        RECT 28.230 177.355 29.085 177.525 ;
        RECT 29.290 177.355 29.785 177.525 ;
        RECT 29.955 177.385 30.285 177.745 ;
        RECT 26.555 176.305 26.725 176.995 ;
        RECT 26.895 176.645 27.065 176.825 ;
        RECT 27.235 176.815 28.025 177.065 ;
        RECT 28.230 176.645 28.400 177.355 ;
        RECT 28.570 176.845 28.925 177.065 ;
        RECT 26.895 176.475 28.585 176.645 ;
        RECT 25.400 175.875 25.860 176.165 ;
        RECT 26.555 176.135 28.055 176.305 ;
        RECT 26.555 175.995 26.725 176.135 ;
        RECT 26.165 175.825 26.725 175.995 ;
        RECT 24.640 175.195 24.890 175.655 ;
        RECT 25.060 175.365 25.930 175.705 ;
        RECT 26.165 175.365 26.335 175.825 ;
        RECT 27.170 175.795 28.245 175.965 ;
        RECT 26.505 175.195 26.875 175.655 ;
        RECT 27.170 175.455 27.340 175.795 ;
        RECT 27.510 175.195 27.840 175.625 ;
        RECT 28.075 175.455 28.245 175.795 ;
        RECT 28.415 175.695 28.585 176.475 ;
        RECT 28.755 176.255 28.925 176.845 ;
        RECT 29.095 176.445 29.445 177.065 ;
        RECT 28.755 175.865 29.220 176.255 ;
        RECT 29.615 175.995 29.785 177.355 ;
        RECT 29.955 176.165 30.415 177.215 ;
        RECT 29.390 175.825 29.785 175.995 ;
        RECT 29.390 175.695 29.560 175.825 ;
        RECT 28.415 175.365 29.095 175.695 ;
        RECT 29.310 175.365 29.560 175.695 ;
        RECT 29.730 175.195 29.980 175.655 ;
        RECT 30.150 175.380 30.475 176.165 ;
        RECT 30.645 175.365 30.815 177.485 ;
        RECT 30.985 177.365 31.315 177.745 ;
        RECT 31.485 177.195 31.740 177.485 ;
        RECT 30.990 177.025 31.740 177.195 ;
        RECT 30.990 176.035 31.220 177.025 ;
        RECT 31.920 177.005 32.175 177.575 ;
        RECT 32.345 177.345 32.675 177.745 ;
        RECT 33.100 177.210 33.630 177.575 ;
        RECT 33.820 177.405 34.095 177.575 ;
        RECT 33.815 177.235 34.095 177.405 ;
        RECT 33.100 177.175 33.275 177.210 ;
        RECT 32.345 177.005 33.275 177.175 ;
        RECT 31.390 176.205 31.740 176.855 ;
        RECT 31.920 176.335 32.090 177.005 ;
        RECT 32.345 176.835 32.515 177.005 ;
        RECT 32.260 176.505 32.515 176.835 ;
        RECT 32.740 176.505 32.935 176.835 ;
        RECT 30.990 175.865 31.740 176.035 ;
        RECT 30.985 175.195 31.315 175.695 ;
        RECT 31.485 175.365 31.740 175.865 ;
        RECT 31.920 175.365 32.255 176.335 ;
        RECT 32.425 175.195 32.595 176.335 ;
        RECT 32.765 175.535 32.935 176.505 ;
        RECT 33.105 175.875 33.275 177.005 ;
        RECT 33.445 176.215 33.615 177.015 ;
        RECT 33.820 176.415 34.095 177.235 ;
        RECT 34.265 176.215 34.455 177.575 ;
        RECT 34.635 177.210 35.145 177.745 ;
        RECT 35.365 176.935 35.610 177.540 ;
        RECT 36.055 176.975 38.645 177.745 ;
        RECT 38.815 177.020 39.105 177.745 ;
        RECT 39.735 176.975 41.405 177.745 ;
        RECT 34.655 176.765 35.885 176.935 ;
        RECT 33.445 176.045 34.455 176.215 ;
        RECT 34.625 176.200 35.375 176.390 ;
        RECT 33.105 175.705 34.230 175.875 ;
        RECT 34.625 175.535 34.795 176.200 ;
        RECT 35.545 175.955 35.885 176.765 ;
        RECT 32.765 175.365 34.795 175.535 ;
        RECT 34.965 175.195 35.135 175.955 ;
        RECT 35.370 175.545 35.885 175.955 ;
        RECT 36.055 176.285 37.265 176.805 ;
        RECT 37.435 176.455 38.645 176.975 ;
        RECT 36.055 175.195 38.645 176.285 ;
        RECT 38.815 175.195 39.105 176.360 ;
        RECT 39.735 176.285 40.485 176.805 ;
        RECT 40.655 176.455 41.405 176.975 ;
        RECT 41.575 176.945 41.915 177.575 ;
        RECT 42.085 176.945 42.335 177.745 ;
        RECT 42.525 177.095 42.855 177.575 ;
        RECT 43.025 177.285 43.250 177.745 ;
        RECT 43.420 177.095 43.750 177.575 ;
        RECT 41.575 176.335 41.750 176.945 ;
        RECT 42.525 176.925 43.750 177.095 ;
        RECT 44.380 176.965 44.880 177.575 ;
        RECT 41.920 176.585 42.615 176.755 ;
        RECT 42.445 176.335 42.615 176.585 ;
        RECT 42.790 176.555 43.210 176.755 ;
        RECT 43.380 176.555 43.710 176.755 ;
        RECT 43.880 176.555 44.210 176.755 ;
        RECT 44.380 176.335 44.550 176.965 ;
        RECT 45.530 176.935 45.775 177.540 ;
        RECT 45.995 177.210 46.505 177.745 ;
        RECT 45.255 176.765 46.485 176.935 ;
        RECT 44.735 176.505 45.085 176.755 ;
        RECT 39.735 175.195 41.405 176.285 ;
        RECT 41.575 175.365 41.915 176.335 ;
        RECT 42.085 175.195 42.255 176.335 ;
        RECT 42.445 176.165 44.880 176.335 ;
        RECT 42.525 175.195 42.775 175.995 ;
        RECT 43.420 175.365 43.750 176.165 ;
        RECT 44.050 175.195 44.380 175.995 ;
        RECT 44.550 175.365 44.880 176.165 ;
        RECT 45.255 175.955 45.595 176.765 ;
        RECT 45.765 176.200 46.515 176.390 ;
        RECT 45.255 175.545 45.770 175.955 ;
        RECT 46.005 175.195 46.175 175.955 ;
        RECT 46.345 175.535 46.515 176.200 ;
        RECT 46.685 176.215 46.875 177.575 ;
        RECT 47.045 176.725 47.320 177.575 ;
        RECT 47.510 177.210 48.040 177.575 ;
        RECT 48.465 177.345 48.795 177.745 ;
        RECT 47.865 177.175 48.040 177.210 ;
        RECT 47.045 176.555 47.325 176.725 ;
        RECT 47.045 176.415 47.320 176.555 ;
        RECT 47.525 176.215 47.695 177.015 ;
        RECT 46.685 176.045 47.695 176.215 ;
        RECT 47.865 177.005 48.795 177.175 ;
        RECT 48.965 177.005 49.220 177.575 ;
        RECT 47.865 175.875 48.035 177.005 ;
        RECT 48.625 176.835 48.795 177.005 ;
        RECT 46.910 175.705 48.035 175.875 ;
        RECT 48.205 176.505 48.400 176.835 ;
        RECT 48.625 176.505 48.880 176.835 ;
        RECT 48.205 175.535 48.375 176.505 ;
        RECT 49.050 176.335 49.220 177.005 ;
        RECT 46.345 175.365 48.375 175.535 ;
        RECT 48.545 175.195 48.715 176.335 ;
        RECT 48.885 175.365 49.220 176.335 ;
        RECT 49.400 177.035 49.655 177.565 ;
        RECT 49.825 177.285 50.130 177.745 ;
        RECT 50.375 177.365 51.445 177.535 ;
        RECT 49.400 176.385 49.610 177.035 ;
        RECT 50.375 177.010 50.695 177.365 ;
        RECT 50.370 176.835 50.695 177.010 ;
        RECT 49.780 176.535 50.695 176.835 ;
        RECT 50.865 176.795 51.105 177.195 ;
        RECT 51.275 177.135 51.445 177.365 ;
        RECT 51.615 177.305 51.805 177.745 ;
        RECT 51.975 177.295 52.925 177.575 ;
        RECT 53.145 177.385 53.495 177.555 ;
        RECT 51.275 176.965 51.805 177.135 ;
        RECT 49.780 176.505 50.520 176.535 ;
        RECT 49.400 175.505 49.655 176.385 ;
        RECT 49.825 175.195 50.130 176.335 ;
        RECT 50.350 175.915 50.520 176.505 ;
        RECT 50.865 176.425 51.405 176.795 ;
        RECT 51.585 176.685 51.805 176.965 ;
        RECT 51.975 176.515 52.145 177.295 ;
        RECT 51.740 176.345 52.145 176.515 ;
        RECT 52.315 176.505 52.665 177.125 ;
        RECT 51.740 176.255 51.910 176.345 ;
        RECT 52.835 176.335 53.045 177.125 ;
        RECT 50.690 176.085 51.910 176.255 ;
        RECT 52.370 176.175 53.045 176.335 ;
        RECT 50.350 175.745 51.150 175.915 ;
        RECT 50.470 175.195 50.800 175.575 ;
        RECT 50.980 175.455 51.150 175.745 ;
        RECT 51.740 175.705 51.910 176.085 ;
        RECT 52.080 176.165 53.045 176.175 ;
        RECT 53.235 176.995 53.495 177.385 ;
        RECT 53.705 177.285 54.035 177.745 ;
        RECT 54.910 177.355 55.765 177.525 ;
        RECT 55.970 177.355 56.465 177.525 ;
        RECT 56.635 177.385 56.965 177.745 ;
        RECT 53.235 176.305 53.405 176.995 ;
        RECT 53.575 176.645 53.745 176.825 ;
        RECT 53.915 176.815 54.705 177.065 ;
        RECT 54.910 176.645 55.080 177.355 ;
        RECT 55.250 176.845 55.605 177.065 ;
        RECT 53.575 176.475 55.265 176.645 ;
        RECT 52.080 175.875 52.540 176.165 ;
        RECT 53.235 176.135 54.735 176.305 ;
        RECT 53.235 175.995 53.405 176.135 ;
        RECT 52.845 175.825 53.405 175.995 ;
        RECT 51.320 175.195 51.570 175.655 ;
        RECT 51.740 175.365 52.610 175.705 ;
        RECT 52.845 175.365 53.015 175.825 ;
        RECT 53.850 175.795 54.925 175.965 ;
        RECT 53.185 175.195 53.555 175.655 ;
        RECT 53.850 175.455 54.020 175.795 ;
        RECT 54.190 175.195 54.520 175.625 ;
        RECT 54.755 175.455 54.925 175.795 ;
        RECT 55.095 175.695 55.265 176.475 ;
        RECT 55.435 176.255 55.605 176.845 ;
        RECT 55.775 176.445 56.125 177.065 ;
        RECT 55.435 175.865 55.900 176.255 ;
        RECT 56.295 175.995 56.465 177.355 ;
        RECT 56.635 176.165 57.095 177.215 ;
        RECT 56.070 175.825 56.465 175.995 ;
        RECT 56.070 175.695 56.240 175.825 ;
        RECT 55.095 175.365 55.775 175.695 ;
        RECT 55.990 175.365 56.240 175.695 ;
        RECT 56.410 175.195 56.660 175.655 ;
        RECT 56.830 175.380 57.155 176.165 ;
        RECT 57.325 175.365 57.495 177.485 ;
        RECT 57.665 177.365 57.995 177.745 ;
        RECT 58.165 177.195 58.420 177.485 ;
        RECT 57.670 177.025 58.420 177.195 ;
        RECT 57.670 176.035 57.900 177.025 ;
        RECT 59.055 176.975 62.565 177.745 ;
        RECT 58.070 176.205 58.420 176.855 ;
        RECT 59.055 176.285 60.745 176.805 ;
        RECT 60.915 176.455 62.565 176.975 ;
        RECT 62.740 176.905 63.000 177.745 ;
        RECT 63.175 177.000 63.430 177.575 ;
        RECT 63.600 177.365 63.930 177.745 ;
        RECT 64.145 177.195 64.315 177.575 ;
        RECT 63.600 177.025 64.315 177.195 ;
        RECT 57.670 175.865 58.420 176.035 ;
        RECT 57.665 175.195 57.995 175.695 ;
        RECT 58.165 175.365 58.420 175.865 ;
        RECT 59.055 175.195 62.565 176.285 ;
        RECT 62.740 175.195 63.000 176.345 ;
        RECT 63.175 176.270 63.345 177.000 ;
        RECT 63.600 176.835 63.770 177.025 ;
        RECT 64.575 177.020 64.865 177.745 ;
        RECT 65.035 176.995 66.245 177.745 ;
        RECT 66.685 177.350 67.015 177.745 ;
        RECT 67.185 177.175 67.385 177.530 ;
        RECT 67.555 177.345 67.885 177.745 ;
        RECT 68.055 177.175 68.255 177.520 ;
        RECT 63.515 176.505 63.770 176.835 ;
        RECT 63.600 176.295 63.770 176.505 ;
        RECT 64.050 176.475 64.405 176.845 ;
        RECT 63.175 175.365 63.430 176.270 ;
        RECT 63.600 176.125 64.315 176.295 ;
        RECT 63.600 175.195 63.930 175.955 ;
        RECT 64.145 175.365 64.315 176.125 ;
        RECT 64.575 175.195 64.865 176.360 ;
        RECT 65.035 176.285 65.555 176.825 ;
        RECT 65.725 176.455 66.245 176.995 ;
        RECT 66.415 177.005 68.255 177.175 ;
        RECT 68.425 177.005 68.755 177.745 ;
        RECT 68.990 177.175 69.160 177.425 ;
        RECT 68.990 177.005 69.465 177.175 ;
        RECT 65.035 175.195 66.245 176.285 ;
        RECT 66.415 175.380 66.675 177.005 ;
        RECT 66.855 176.035 67.075 176.835 ;
        RECT 67.315 176.215 67.615 176.835 ;
        RECT 67.785 176.215 68.115 176.835 ;
        RECT 68.285 176.215 68.605 176.835 ;
        RECT 68.775 176.215 69.125 176.835 ;
        RECT 69.295 176.035 69.465 177.005 ;
        RECT 70.095 176.975 71.765 177.745 ;
        RECT 71.940 177.200 77.285 177.745 ;
        RECT 66.855 175.825 69.465 176.035 ;
        RECT 70.095 176.285 70.845 176.805 ;
        RECT 71.015 176.455 71.765 176.975 ;
        RECT 68.425 175.195 68.755 175.645 ;
        RECT 70.095 175.195 71.765 176.285 ;
        RECT 73.530 175.630 73.880 176.880 ;
        RECT 75.360 176.370 75.700 177.200 ;
        RECT 77.545 177.095 77.715 177.575 ;
        RECT 77.895 177.265 78.135 177.745 ;
        RECT 78.385 177.095 78.555 177.575 ;
        RECT 78.725 177.265 79.055 177.745 ;
        RECT 79.225 177.095 79.395 177.575 ;
        RECT 77.545 176.925 78.180 177.095 ;
        RECT 78.385 176.925 79.395 177.095 ;
        RECT 79.565 176.945 79.895 177.745 ;
        RECT 80.215 176.945 80.555 177.575 ;
        RECT 80.725 176.945 80.975 177.745 ;
        RECT 81.165 177.095 81.495 177.575 ;
        RECT 81.665 177.285 81.890 177.745 ;
        RECT 82.060 177.095 82.390 177.575 ;
        RECT 78.010 176.755 78.180 176.925 ;
        RECT 78.895 176.895 79.395 176.925 ;
        RECT 77.460 176.515 77.840 176.755 ;
        RECT 78.010 176.585 78.510 176.755 ;
        RECT 78.010 176.345 78.180 176.585 ;
        RECT 78.900 176.385 79.395 176.895 ;
        RECT 77.465 176.175 78.180 176.345 ;
        RECT 78.385 176.215 79.395 176.385 ;
        RECT 71.940 175.195 77.285 175.630 ;
        RECT 77.465 175.365 77.795 176.175 ;
        RECT 77.965 175.195 78.205 175.995 ;
        RECT 78.385 175.365 78.555 176.215 ;
        RECT 78.725 175.195 79.055 175.995 ;
        RECT 79.225 175.365 79.395 176.215 ;
        RECT 79.565 175.195 79.895 176.345 ;
        RECT 80.215 176.335 80.390 176.945 ;
        RECT 81.165 176.925 82.390 177.095 ;
        RECT 83.020 176.965 83.520 177.575 ;
        RECT 83.985 177.095 84.155 177.575 ;
        RECT 84.335 177.265 84.575 177.745 ;
        RECT 84.825 177.095 84.995 177.575 ;
        RECT 85.165 177.265 85.495 177.745 ;
        RECT 85.665 177.095 85.835 177.575 ;
        RECT 80.560 176.585 81.255 176.755 ;
        RECT 81.085 176.335 81.255 176.585 ;
        RECT 81.430 176.555 81.850 176.755 ;
        RECT 82.020 176.555 82.350 176.755 ;
        RECT 82.520 176.555 82.850 176.755 ;
        RECT 83.020 176.335 83.190 176.965 ;
        RECT 83.985 176.925 84.620 177.095 ;
        RECT 84.825 176.925 85.835 177.095 ;
        RECT 86.005 176.945 86.335 177.745 ;
        RECT 86.655 176.975 90.165 177.745 ;
        RECT 90.335 177.020 90.625 177.745 ;
        RECT 91.255 176.975 92.925 177.745 ;
        RECT 93.100 177.200 98.445 177.745 ;
        RECT 84.450 176.755 84.620 176.925 ;
        RECT 85.335 176.895 85.835 176.925 ;
        RECT 83.375 176.505 83.725 176.755 ;
        RECT 83.900 176.515 84.280 176.755 ;
        RECT 84.450 176.585 84.950 176.755 ;
        RECT 84.450 176.345 84.620 176.585 ;
        RECT 85.340 176.385 85.835 176.895 ;
        RECT 80.215 175.365 80.555 176.335 ;
        RECT 80.725 175.195 80.895 176.335 ;
        RECT 81.085 176.165 83.520 176.335 ;
        RECT 81.165 175.195 81.415 175.995 ;
        RECT 82.060 175.365 82.390 176.165 ;
        RECT 82.690 175.195 83.020 175.995 ;
        RECT 83.190 175.365 83.520 176.165 ;
        RECT 83.905 176.175 84.620 176.345 ;
        RECT 84.825 176.215 85.835 176.385 ;
        RECT 83.905 175.365 84.235 176.175 ;
        RECT 84.405 175.195 84.645 175.995 ;
        RECT 84.825 175.365 84.995 176.215 ;
        RECT 85.165 175.195 85.495 175.995 ;
        RECT 85.665 175.365 85.835 176.215 ;
        RECT 86.005 175.195 86.335 176.345 ;
        RECT 86.655 176.285 88.345 176.805 ;
        RECT 88.515 176.455 90.165 176.975 ;
        RECT 86.655 175.195 90.165 176.285 ;
        RECT 90.335 175.195 90.625 176.360 ;
        RECT 91.255 176.285 92.005 176.805 ;
        RECT 92.175 176.455 92.925 176.975 ;
        RECT 91.255 175.195 92.925 176.285 ;
        RECT 94.690 175.630 95.040 176.880 ;
        RECT 96.520 176.370 96.860 177.200 ;
        RECT 98.615 176.945 98.955 177.575 ;
        RECT 99.125 176.945 99.375 177.745 ;
        RECT 99.565 177.095 99.895 177.575 ;
        RECT 100.065 177.285 100.290 177.745 ;
        RECT 100.460 177.095 100.790 177.575 ;
        RECT 98.615 176.335 98.790 176.945 ;
        RECT 99.565 176.925 100.790 177.095 ;
        RECT 101.420 176.965 101.920 177.575 ;
        RECT 102.755 176.975 104.425 177.745 ;
        RECT 98.960 176.585 99.655 176.755 ;
        RECT 99.485 176.335 99.655 176.585 ;
        RECT 99.830 176.555 100.250 176.755 ;
        RECT 100.420 176.555 100.750 176.755 ;
        RECT 100.920 176.555 101.250 176.755 ;
        RECT 101.420 176.335 101.590 176.965 ;
        RECT 101.775 176.505 102.125 176.755 ;
        RECT 93.100 175.195 98.445 175.630 ;
        RECT 98.615 175.365 98.955 176.335 ;
        RECT 99.125 175.195 99.295 176.335 ;
        RECT 99.485 176.165 101.920 176.335 ;
        RECT 99.565 175.195 99.815 175.995 ;
        RECT 100.460 175.365 100.790 176.165 ;
        RECT 101.090 175.195 101.420 175.995 ;
        RECT 101.590 175.365 101.920 176.165 ;
        RECT 102.755 176.285 103.505 176.805 ;
        RECT 103.675 176.455 104.425 176.975 ;
        RECT 104.595 176.945 104.935 177.575 ;
        RECT 105.105 176.945 105.355 177.745 ;
        RECT 105.545 177.095 105.875 177.575 ;
        RECT 106.045 177.285 106.270 177.745 ;
        RECT 106.440 177.095 106.770 177.575 ;
        RECT 104.595 176.335 104.770 176.945 ;
        RECT 105.545 176.925 106.770 177.095 ;
        RECT 107.400 176.965 107.900 177.575 ;
        RECT 104.940 176.585 105.635 176.755 ;
        RECT 105.465 176.335 105.635 176.585 ;
        RECT 105.810 176.555 106.230 176.755 ;
        RECT 106.400 176.555 106.730 176.755 ;
        RECT 106.900 176.555 107.230 176.755 ;
        RECT 107.400 176.335 107.570 176.965 ;
        RECT 108.275 176.945 108.615 177.575 ;
        RECT 108.785 176.945 109.035 177.745 ;
        RECT 109.225 177.095 109.555 177.575 ;
        RECT 109.725 177.285 109.950 177.745 ;
        RECT 110.120 177.095 110.450 177.575 ;
        RECT 107.755 176.505 108.105 176.755 ;
        RECT 108.275 176.335 108.450 176.945 ;
        RECT 109.225 176.925 110.450 177.095 ;
        RECT 111.080 176.965 111.580 177.575 ;
        RECT 112.160 176.965 112.660 177.575 ;
        RECT 108.620 176.585 109.315 176.755 ;
        RECT 109.145 176.335 109.315 176.585 ;
        RECT 109.490 176.555 109.910 176.755 ;
        RECT 110.080 176.555 110.410 176.755 ;
        RECT 110.580 176.555 110.910 176.755 ;
        RECT 111.080 176.335 111.250 176.965 ;
        RECT 111.435 176.505 111.785 176.755 ;
        RECT 111.955 176.505 112.305 176.755 ;
        RECT 112.490 176.335 112.660 176.965 ;
        RECT 113.290 177.095 113.620 177.575 ;
        RECT 113.790 177.285 114.015 177.745 ;
        RECT 114.185 177.095 114.515 177.575 ;
        RECT 113.290 176.925 114.515 177.095 ;
        RECT 114.705 176.945 114.955 177.745 ;
        RECT 115.125 176.945 115.465 177.575 ;
        RECT 116.095 177.020 116.385 177.745 ;
        RECT 117.015 176.975 120.525 177.745 ;
        RECT 120.785 177.195 120.955 177.575 ;
        RECT 121.135 177.365 121.465 177.745 ;
        RECT 120.785 177.025 121.450 177.195 ;
        RECT 121.645 177.070 121.905 177.575 ;
        RECT 122.540 177.200 127.885 177.745 ;
        RECT 112.830 176.555 113.160 176.755 ;
        RECT 113.330 176.555 113.660 176.755 ;
        RECT 113.830 176.555 114.250 176.755 ;
        RECT 114.425 176.585 115.120 176.755 ;
        RECT 114.425 176.335 114.595 176.585 ;
        RECT 115.290 176.335 115.465 176.945 ;
        RECT 102.755 175.195 104.425 176.285 ;
        RECT 104.595 175.365 104.935 176.335 ;
        RECT 105.105 175.195 105.275 176.335 ;
        RECT 105.465 176.165 107.900 176.335 ;
        RECT 105.545 175.195 105.795 175.995 ;
        RECT 106.440 175.365 106.770 176.165 ;
        RECT 107.070 175.195 107.400 175.995 ;
        RECT 107.570 175.365 107.900 176.165 ;
        RECT 108.275 175.365 108.615 176.335 ;
        RECT 108.785 175.195 108.955 176.335 ;
        RECT 109.145 176.165 111.580 176.335 ;
        RECT 109.225 175.195 109.475 175.995 ;
        RECT 110.120 175.365 110.450 176.165 ;
        RECT 110.750 175.195 111.080 175.995 ;
        RECT 111.250 175.365 111.580 176.165 ;
        RECT 112.160 176.165 114.595 176.335 ;
        RECT 112.160 175.365 112.490 176.165 ;
        RECT 112.660 175.195 112.990 175.995 ;
        RECT 113.290 175.365 113.620 176.165 ;
        RECT 114.265 175.195 114.515 175.995 ;
        RECT 114.785 175.195 114.955 176.335 ;
        RECT 115.125 175.365 115.465 176.335 ;
        RECT 116.095 175.195 116.385 176.360 ;
        RECT 117.015 176.285 118.705 176.805 ;
        RECT 118.875 176.455 120.525 176.975 ;
        RECT 120.715 176.475 121.045 176.845 ;
        RECT 121.280 176.770 121.450 177.025 ;
        RECT 121.280 176.440 121.565 176.770 ;
        RECT 121.280 176.295 121.450 176.440 ;
        RECT 117.015 175.195 120.525 176.285 ;
        RECT 120.785 176.125 121.450 176.295 ;
        RECT 121.735 176.270 121.905 177.070 ;
        RECT 120.785 175.365 120.955 176.125 ;
        RECT 121.135 175.195 121.465 175.955 ;
        RECT 121.635 175.365 121.905 176.270 ;
        RECT 124.130 175.630 124.480 176.880 ;
        RECT 125.960 176.370 126.300 177.200 ;
        RECT 128.055 176.995 129.265 177.745 ;
        RECT 128.055 176.285 128.575 176.825 ;
        RECT 128.745 176.455 129.265 176.995 ;
        RECT 122.540 175.195 127.885 175.630 ;
        RECT 128.055 175.195 129.265 176.285 ;
        RECT 9.290 175.025 129.350 175.195 ;
        RECT 9.375 173.935 10.585 175.025 ;
        RECT 9.375 173.225 9.895 173.765 ;
        RECT 10.065 173.395 10.585 173.935 ;
        RECT 11.215 173.935 14.725 175.025 ;
        RECT 14.900 174.590 20.245 175.025 ;
        RECT 20.420 174.590 25.765 175.025 ;
        RECT 11.215 173.415 12.905 173.935 ;
        RECT 13.075 173.245 14.725 173.765 ;
        RECT 16.490 173.340 16.840 174.590 ;
        RECT 9.375 172.475 10.585 173.225 ;
        RECT 11.215 172.475 14.725 173.245 ;
        RECT 18.320 173.020 18.660 173.850 ;
        RECT 22.010 173.340 22.360 174.590 ;
        RECT 25.935 173.860 26.225 175.025 ;
        RECT 26.395 173.935 27.605 175.025 ;
        RECT 27.775 173.935 31.285 175.025 ;
        RECT 31.455 173.950 31.725 174.855 ;
        RECT 31.895 174.265 32.225 175.025 ;
        RECT 32.405 174.095 32.575 174.855 ;
        RECT 23.840 173.020 24.180 173.850 ;
        RECT 26.395 173.395 26.915 173.935 ;
        RECT 27.085 173.225 27.605 173.765 ;
        RECT 27.775 173.415 29.465 173.935 ;
        RECT 29.635 173.245 31.285 173.765 ;
        RECT 14.900 172.475 20.245 173.020 ;
        RECT 20.420 172.475 25.765 173.020 ;
        RECT 25.935 172.475 26.225 173.200 ;
        RECT 26.395 172.475 27.605 173.225 ;
        RECT 27.775 172.475 31.285 173.245 ;
        RECT 31.455 173.150 31.625 173.950 ;
        RECT 31.910 173.925 32.575 174.095 ;
        RECT 31.910 173.780 32.080 173.925 ;
        RECT 31.795 173.450 32.080 173.780 ;
        RECT 32.835 173.885 33.175 174.855 ;
        RECT 33.345 173.885 33.515 175.025 ;
        RECT 33.785 174.225 34.035 175.025 ;
        RECT 34.680 174.055 35.010 174.855 ;
        RECT 35.310 174.225 35.640 175.025 ;
        RECT 35.810 174.055 36.140 174.855 ;
        RECT 33.705 173.885 36.140 174.055 ;
        RECT 36.975 173.885 37.315 174.855 ;
        RECT 37.485 173.885 37.655 175.025 ;
        RECT 37.925 174.225 38.175 175.025 ;
        RECT 38.820 174.055 39.150 174.855 ;
        RECT 39.450 174.225 39.780 175.025 ;
        RECT 39.950 174.055 40.280 174.855 ;
        RECT 37.845 173.885 40.280 174.055 ;
        RECT 40.655 173.885 40.995 174.855 ;
        RECT 41.165 173.885 41.335 175.025 ;
        RECT 41.605 174.225 41.855 175.025 ;
        RECT 42.500 174.055 42.830 174.855 ;
        RECT 43.130 174.225 43.460 175.025 ;
        RECT 43.630 174.055 43.960 174.855 ;
        RECT 41.525 173.885 43.960 174.055 ;
        RECT 44.335 173.885 44.675 174.855 ;
        RECT 44.845 173.885 45.015 175.025 ;
        RECT 45.285 174.225 45.535 175.025 ;
        RECT 46.180 174.055 46.510 174.855 ;
        RECT 46.810 174.225 47.140 175.025 ;
        RECT 47.310 174.055 47.640 174.855 ;
        RECT 45.205 173.885 47.640 174.055 ;
        RECT 48.015 173.885 48.355 174.855 ;
        RECT 48.525 173.885 48.695 175.025 ;
        RECT 48.965 174.225 49.215 175.025 ;
        RECT 49.860 174.055 50.190 174.855 ;
        RECT 50.490 174.225 50.820 175.025 ;
        RECT 50.990 174.055 51.320 174.855 ;
        RECT 48.885 173.885 51.320 174.055 ;
        RECT 31.910 173.195 32.080 173.450 ;
        RECT 32.315 173.375 32.645 173.745 ;
        RECT 32.835 173.275 33.010 173.885 ;
        RECT 33.705 173.635 33.875 173.885 ;
        RECT 33.180 173.465 33.875 173.635 ;
        RECT 34.050 173.465 34.470 173.665 ;
        RECT 34.640 173.465 34.970 173.665 ;
        RECT 35.140 173.465 35.470 173.665 ;
        RECT 31.455 172.645 31.715 173.150 ;
        RECT 31.910 173.025 32.575 173.195 ;
        RECT 31.895 172.475 32.225 172.855 ;
        RECT 32.405 172.645 32.575 173.025 ;
        RECT 32.835 172.645 33.175 173.275 ;
        RECT 33.345 172.475 33.595 173.275 ;
        RECT 33.785 173.125 35.010 173.295 ;
        RECT 33.785 172.645 34.115 173.125 ;
        RECT 34.285 172.475 34.510 172.935 ;
        RECT 34.680 172.645 35.010 173.125 ;
        RECT 35.640 173.255 35.810 173.885 ;
        RECT 35.995 173.465 36.345 173.715 ;
        RECT 36.975 173.275 37.150 173.885 ;
        RECT 37.845 173.635 38.015 173.885 ;
        RECT 37.320 173.465 38.015 173.635 ;
        RECT 38.190 173.465 38.610 173.665 ;
        RECT 38.780 173.465 39.110 173.665 ;
        RECT 39.280 173.465 39.610 173.665 ;
        RECT 35.640 172.645 36.140 173.255 ;
        RECT 36.975 172.645 37.315 173.275 ;
        RECT 37.485 172.475 37.735 173.275 ;
        RECT 37.925 173.125 39.150 173.295 ;
        RECT 37.925 172.645 38.255 173.125 ;
        RECT 38.425 172.475 38.650 172.935 ;
        RECT 38.820 172.645 39.150 173.125 ;
        RECT 39.780 173.255 39.950 173.885 ;
        RECT 40.135 173.465 40.485 173.715 ;
        RECT 40.655 173.275 40.830 173.885 ;
        RECT 41.525 173.635 41.695 173.885 ;
        RECT 41.000 173.465 41.695 173.635 ;
        RECT 41.870 173.465 42.290 173.665 ;
        RECT 42.460 173.465 42.790 173.665 ;
        RECT 42.960 173.465 43.290 173.665 ;
        RECT 39.780 172.645 40.280 173.255 ;
        RECT 40.655 172.645 40.995 173.275 ;
        RECT 41.165 172.475 41.415 173.275 ;
        RECT 41.605 173.125 42.830 173.295 ;
        RECT 41.605 172.645 41.935 173.125 ;
        RECT 42.105 172.475 42.330 172.935 ;
        RECT 42.500 172.645 42.830 173.125 ;
        RECT 43.460 173.255 43.630 173.885 ;
        RECT 43.815 173.465 44.165 173.715 ;
        RECT 44.335 173.275 44.510 173.885 ;
        RECT 45.205 173.635 45.375 173.885 ;
        RECT 44.680 173.465 45.375 173.635 ;
        RECT 45.550 173.465 45.970 173.665 ;
        RECT 46.140 173.465 46.470 173.665 ;
        RECT 46.640 173.465 46.970 173.665 ;
        RECT 43.460 172.645 43.960 173.255 ;
        RECT 44.335 172.645 44.675 173.275 ;
        RECT 44.845 172.475 45.095 173.275 ;
        RECT 45.285 173.125 46.510 173.295 ;
        RECT 45.285 172.645 45.615 173.125 ;
        RECT 45.785 172.475 46.010 172.935 ;
        RECT 46.180 172.645 46.510 173.125 ;
        RECT 47.140 173.255 47.310 173.885 ;
        RECT 47.495 173.465 47.845 173.715 ;
        RECT 48.015 173.275 48.190 173.885 ;
        RECT 48.885 173.635 49.055 173.885 ;
        RECT 48.360 173.465 49.055 173.635 ;
        RECT 49.230 173.465 49.650 173.665 ;
        RECT 49.820 173.465 50.150 173.665 ;
        RECT 50.320 173.465 50.650 173.665 ;
        RECT 47.140 172.645 47.640 173.255 ;
        RECT 48.015 172.645 48.355 173.275 ;
        RECT 48.525 172.475 48.775 173.275 ;
        RECT 48.965 173.125 50.190 173.295 ;
        RECT 48.965 172.645 49.295 173.125 ;
        RECT 49.465 172.475 49.690 172.935 ;
        RECT 49.860 172.645 50.190 173.125 ;
        RECT 50.820 173.255 50.990 173.885 ;
        RECT 51.695 173.860 51.985 175.025 ;
        RECT 52.675 173.885 52.885 175.025 ;
        RECT 53.055 173.875 53.385 174.855 ;
        RECT 53.555 173.885 53.785 175.025 ;
        RECT 55.005 174.095 55.175 174.855 ;
        RECT 55.355 174.265 55.685 175.025 ;
        RECT 55.005 173.925 55.670 174.095 ;
        RECT 55.855 173.950 56.125 174.855 ;
        RECT 51.175 173.465 51.525 173.715 ;
        RECT 50.820 172.645 51.320 173.255 ;
        RECT 51.695 172.475 51.985 173.200 ;
        RECT 52.675 172.475 52.885 173.295 ;
        RECT 53.055 173.275 53.305 173.875 ;
        RECT 55.500 173.780 55.670 173.925 ;
        RECT 53.475 173.465 53.805 173.715 ;
        RECT 54.935 173.375 55.265 173.745 ;
        RECT 55.500 173.450 55.785 173.780 ;
        RECT 53.055 172.645 53.385 173.275 ;
        RECT 53.555 172.475 53.785 173.295 ;
        RECT 55.500 173.195 55.670 173.450 ;
        RECT 55.005 173.025 55.670 173.195 ;
        RECT 55.955 173.150 56.125 173.950 ;
        RECT 56.295 173.935 59.805 175.025 ;
        RECT 56.295 173.415 57.985 173.935 ;
        RECT 59.980 173.875 60.240 175.025 ;
        RECT 60.415 173.950 60.670 174.855 ;
        RECT 60.840 174.265 61.170 175.025 ;
        RECT 61.385 174.095 61.555 174.855 ;
        RECT 58.155 173.245 59.805 173.765 ;
        RECT 55.005 172.645 55.175 173.025 ;
        RECT 55.355 172.475 55.685 172.855 ;
        RECT 55.865 172.645 56.125 173.150 ;
        RECT 56.295 172.475 59.805 173.245 ;
        RECT 59.980 172.475 60.240 173.315 ;
        RECT 60.415 173.220 60.585 173.950 ;
        RECT 60.840 173.925 61.555 174.095 ;
        RECT 60.840 173.715 61.010 173.925 ;
        RECT 61.820 173.875 62.080 175.025 ;
        RECT 62.255 173.950 62.510 174.855 ;
        RECT 62.680 174.265 63.010 175.025 ;
        RECT 63.225 174.095 63.395 174.855 ;
        RECT 64.365 174.575 64.695 175.025 ;
        RECT 60.755 173.385 61.010 173.715 ;
        RECT 60.415 172.645 60.670 173.220 ;
        RECT 60.840 173.195 61.010 173.385 ;
        RECT 61.290 173.375 61.645 173.745 ;
        RECT 60.840 173.025 61.555 173.195 ;
        RECT 60.840 172.475 61.170 172.855 ;
        RECT 61.385 172.645 61.555 173.025 ;
        RECT 61.820 172.475 62.080 173.315 ;
        RECT 62.255 173.220 62.425 173.950 ;
        RECT 62.680 173.925 63.395 174.095 ;
        RECT 63.655 174.185 66.265 174.395 ;
        RECT 62.680 173.715 62.850 173.925 ;
        RECT 62.595 173.385 62.850 173.715 ;
        RECT 62.255 172.645 62.510 173.220 ;
        RECT 62.680 173.195 62.850 173.385 ;
        RECT 63.130 173.375 63.485 173.745 ;
        RECT 63.655 173.215 63.825 174.185 ;
        RECT 63.995 173.385 64.345 174.005 ;
        RECT 64.515 173.385 64.835 174.005 ;
        RECT 65.005 173.385 65.335 174.005 ;
        RECT 65.505 173.385 65.805 174.005 ;
        RECT 66.045 173.385 66.265 174.185 ;
        RECT 66.445 173.215 66.705 174.840 ;
        RECT 62.680 173.025 63.395 173.195 ;
        RECT 63.655 173.045 64.130 173.215 ;
        RECT 62.680 172.475 63.010 172.855 ;
        RECT 63.225 172.645 63.395 173.025 ;
        RECT 63.960 172.795 64.130 173.045 ;
        RECT 64.365 172.475 64.695 173.215 ;
        RECT 64.865 173.045 66.705 173.215 ;
        RECT 66.875 173.215 67.135 174.840 ;
        RECT 68.885 174.575 69.215 175.025 ;
        RECT 67.315 174.185 69.925 174.395 ;
        RECT 67.315 173.385 67.535 174.185 ;
        RECT 67.775 173.385 68.075 174.005 ;
        RECT 68.245 173.385 68.575 174.005 ;
        RECT 68.745 173.385 69.065 174.005 ;
        RECT 69.235 173.385 69.585 174.005 ;
        RECT 69.755 173.215 69.925 174.185 ;
        RECT 70.095 173.935 71.765 175.025 ;
        RECT 71.940 174.590 77.285 175.025 ;
        RECT 70.095 173.415 70.845 173.935 ;
        RECT 71.015 173.245 71.765 173.765 ;
        RECT 73.530 173.340 73.880 174.590 ;
        RECT 77.455 173.860 77.745 175.025 ;
        RECT 78.375 173.935 80.045 175.025 ;
        RECT 66.875 173.045 68.715 173.215 ;
        RECT 64.865 172.700 65.065 173.045 ;
        RECT 65.235 172.475 65.565 172.875 ;
        RECT 65.735 172.690 65.935 173.045 ;
        RECT 66.105 172.475 66.435 172.870 ;
        RECT 67.145 172.475 67.475 172.870 ;
        RECT 67.645 172.690 67.845 173.045 ;
        RECT 68.015 172.475 68.345 172.875 ;
        RECT 68.515 172.700 68.715 173.045 ;
        RECT 68.885 172.475 69.215 173.215 ;
        RECT 69.450 173.045 69.925 173.215 ;
        RECT 69.450 172.795 69.620 173.045 ;
        RECT 70.095 172.475 71.765 173.245 ;
        RECT 75.360 173.020 75.700 173.850 ;
        RECT 78.375 173.415 79.125 173.935 ;
        RECT 80.215 173.885 80.555 174.855 ;
        RECT 80.725 173.885 80.895 175.025 ;
        RECT 81.165 174.225 81.415 175.025 ;
        RECT 82.060 174.055 82.390 174.855 ;
        RECT 82.690 174.225 83.020 175.025 ;
        RECT 83.190 174.055 83.520 174.855 ;
        RECT 81.085 173.885 83.520 174.055 ;
        RECT 83.895 173.885 84.235 174.855 ;
        RECT 84.405 173.885 84.575 175.025 ;
        RECT 84.845 174.225 85.095 175.025 ;
        RECT 85.740 174.055 86.070 174.855 ;
        RECT 86.370 174.225 86.700 175.025 ;
        RECT 86.870 174.055 87.200 174.855 ;
        RECT 84.765 173.885 87.200 174.055 ;
        RECT 87.575 173.935 88.785 175.025 ;
        RECT 88.960 174.590 94.305 175.025 ;
        RECT 79.295 173.245 80.045 173.765 ;
        RECT 71.940 172.475 77.285 173.020 ;
        RECT 77.455 172.475 77.745 173.200 ;
        RECT 78.375 172.475 80.045 173.245 ;
        RECT 80.215 173.275 80.390 173.885 ;
        RECT 81.085 173.635 81.255 173.885 ;
        RECT 80.560 173.465 81.255 173.635 ;
        RECT 81.430 173.465 81.850 173.665 ;
        RECT 82.020 173.465 82.350 173.665 ;
        RECT 82.520 173.465 82.850 173.665 ;
        RECT 80.215 172.645 80.555 173.275 ;
        RECT 80.725 172.475 80.975 173.275 ;
        RECT 81.165 173.125 82.390 173.295 ;
        RECT 81.165 172.645 81.495 173.125 ;
        RECT 81.665 172.475 81.890 172.935 ;
        RECT 82.060 172.645 82.390 173.125 ;
        RECT 83.020 173.255 83.190 173.885 ;
        RECT 83.375 173.465 83.725 173.715 ;
        RECT 83.895 173.275 84.070 173.885 ;
        RECT 84.765 173.635 84.935 173.885 ;
        RECT 84.240 173.465 84.935 173.635 ;
        RECT 85.110 173.465 85.530 173.665 ;
        RECT 85.700 173.465 86.030 173.665 ;
        RECT 86.200 173.465 86.530 173.665 ;
        RECT 83.020 172.645 83.520 173.255 ;
        RECT 83.895 172.645 84.235 173.275 ;
        RECT 84.405 172.475 84.655 173.275 ;
        RECT 84.845 173.125 86.070 173.295 ;
        RECT 84.845 172.645 85.175 173.125 ;
        RECT 85.345 172.475 85.570 172.935 ;
        RECT 85.740 172.645 86.070 173.125 ;
        RECT 86.700 173.255 86.870 173.885 ;
        RECT 87.055 173.465 87.405 173.715 ;
        RECT 87.575 173.395 88.095 173.935 ;
        RECT 86.700 172.645 87.200 173.255 ;
        RECT 88.265 173.225 88.785 173.765 ;
        RECT 90.550 173.340 90.900 174.590 ;
        RECT 94.515 173.885 94.745 175.025 ;
        RECT 94.915 173.875 95.245 174.855 ;
        RECT 95.415 173.885 95.625 175.025 ;
        RECT 95.855 173.935 97.525 175.025 ;
        RECT 97.700 174.590 103.045 175.025 ;
        RECT 87.575 172.475 88.785 173.225 ;
        RECT 92.380 173.020 92.720 173.850 ;
        RECT 94.495 173.465 94.825 173.715 ;
        RECT 88.960 172.475 94.305 173.020 ;
        RECT 94.515 172.475 94.745 173.295 ;
        RECT 94.995 173.275 95.245 173.875 ;
        RECT 95.855 173.415 96.605 173.935 ;
        RECT 94.915 172.645 95.245 173.275 ;
        RECT 95.415 172.475 95.625 173.295 ;
        RECT 96.775 173.245 97.525 173.765 ;
        RECT 99.290 173.340 99.640 174.590 ;
        RECT 103.215 173.860 103.505 175.025 ;
        RECT 104.595 173.935 108.105 175.025 ;
        RECT 95.855 172.475 97.525 173.245 ;
        RECT 101.120 173.020 101.460 173.850 ;
        RECT 104.595 173.415 106.285 173.935 ;
        RECT 108.275 173.885 108.615 174.855 ;
        RECT 108.785 173.885 108.955 175.025 ;
        RECT 109.225 174.225 109.475 175.025 ;
        RECT 110.120 174.055 110.450 174.855 ;
        RECT 110.750 174.225 111.080 175.025 ;
        RECT 111.250 174.055 111.580 174.855 ;
        RECT 109.145 173.885 111.580 174.055 ;
        RECT 111.955 173.935 113.165 175.025 ;
        RECT 113.335 173.935 116.845 175.025 ;
        RECT 117.020 174.590 122.365 175.025 ;
        RECT 122.540 174.590 127.885 175.025 ;
        RECT 106.455 173.245 108.105 173.765 ;
        RECT 97.700 172.475 103.045 173.020 ;
        RECT 103.215 172.475 103.505 173.200 ;
        RECT 104.595 172.475 108.105 173.245 ;
        RECT 108.275 173.275 108.450 173.885 ;
        RECT 109.145 173.635 109.315 173.885 ;
        RECT 108.620 173.465 109.315 173.635 ;
        RECT 109.490 173.465 109.910 173.665 ;
        RECT 110.080 173.465 110.410 173.665 ;
        RECT 110.580 173.465 110.910 173.665 ;
        RECT 108.275 172.645 108.615 173.275 ;
        RECT 108.785 172.475 109.035 173.275 ;
        RECT 109.225 173.125 110.450 173.295 ;
        RECT 109.225 172.645 109.555 173.125 ;
        RECT 109.725 172.475 109.950 172.935 ;
        RECT 110.120 172.645 110.450 173.125 ;
        RECT 111.080 173.255 111.250 173.885 ;
        RECT 111.435 173.465 111.785 173.715 ;
        RECT 111.955 173.395 112.475 173.935 ;
        RECT 111.080 172.645 111.580 173.255 ;
        RECT 112.645 173.225 113.165 173.765 ;
        RECT 113.335 173.415 115.025 173.935 ;
        RECT 115.195 173.245 116.845 173.765 ;
        RECT 118.610 173.340 118.960 174.590 ;
        RECT 111.955 172.475 113.165 173.225 ;
        RECT 113.335 172.475 116.845 173.245 ;
        RECT 120.440 173.020 120.780 173.850 ;
        RECT 124.130 173.340 124.480 174.590 ;
        RECT 128.055 173.935 129.265 175.025 ;
        RECT 125.960 173.020 126.300 173.850 ;
        RECT 128.055 173.395 128.575 173.935 ;
        RECT 128.745 173.225 129.265 173.765 ;
        RECT 117.020 172.475 122.365 173.020 ;
        RECT 122.540 172.475 127.885 173.020 ;
        RECT 128.055 172.475 129.265 173.225 ;
        RECT 9.290 172.305 129.350 172.475 ;
        RECT 9.375 171.555 10.585 172.305 ;
        RECT 9.375 171.015 9.895 171.555 ;
        RECT 11.215 171.535 12.885 172.305 ;
        RECT 13.055 171.580 13.345 172.305 ;
        RECT 13.975 171.535 16.565 172.305 ;
        RECT 16.740 171.760 22.085 172.305 ;
        RECT 22.260 171.760 27.605 172.305 ;
        RECT 27.780 171.760 33.125 172.305 ;
        RECT 33.300 171.760 38.645 172.305 ;
        RECT 10.065 170.845 10.585 171.385 ;
        RECT 9.375 169.755 10.585 170.845 ;
        RECT 11.215 170.845 11.965 171.365 ;
        RECT 12.135 171.015 12.885 171.535 ;
        RECT 11.215 169.755 12.885 170.845 ;
        RECT 13.055 169.755 13.345 170.920 ;
        RECT 13.975 170.845 15.185 171.365 ;
        RECT 15.355 171.015 16.565 171.535 ;
        RECT 13.975 169.755 16.565 170.845 ;
        RECT 18.330 170.190 18.680 171.440 ;
        RECT 20.160 170.930 20.500 171.760 ;
        RECT 23.850 170.190 24.200 171.440 ;
        RECT 25.680 170.930 26.020 171.760 ;
        RECT 29.370 170.190 29.720 171.440 ;
        RECT 31.200 170.930 31.540 171.760 ;
        RECT 34.890 170.190 35.240 171.440 ;
        RECT 36.720 170.930 37.060 171.760 ;
        RECT 38.815 171.580 39.105 172.305 ;
        RECT 39.275 171.505 39.615 172.135 ;
        RECT 39.785 171.505 40.035 172.305 ;
        RECT 40.225 171.655 40.555 172.135 ;
        RECT 40.725 171.845 40.950 172.305 ;
        RECT 41.120 171.655 41.450 172.135 ;
        RECT 16.740 169.755 22.085 170.190 ;
        RECT 22.260 169.755 27.605 170.190 ;
        RECT 27.780 169.755 33.125 170.190 ;
        RECT 33.300 169.755 38.645 170.190 ;
        RECT 38.815 169.755 39.105 170.920 ;
        RECT 39.275 170.895 39.450 171.505 ;
        RECT 40.225 171.485 41.450 171.655 ;
        RECT 42.080 171.525 42.580 172.135 ;
        RECT 43.415 171.535 46.005 172.305 ;
        RECT 39.620 171.145 40.315 171.315 ;
        RECT 40.145 170.895 40.315 171.145 ;
        RECT 40.490 171.115 40.910 171.315 ;
        RECT 41.080 171.115 41.410 171.315 ;
        RECT 41.580 171.115 41.910 171.315 ;
        RECT 42.080 170.895 42.250 171.525 ;
        RECT 42.435 171.065 42.785 171.315 ;
        RECT 39.275 169.925 39.615 170.895 ;
        RECT 39.785 169.755 39.955 170.895 ;
        RECT 40.145 170.725 42.580 170.895 ;
        RECT 40.225 169.755 40.475 170.555 ;
        RECT 41.120 169.925 41.450 170.725 ;
        RECT 41.750 169.755 42.080 170.555 ;
        RECT 42.250 169.925 42.580 170.725 ;
        RECT 43.415 170.845 44.625 171.365 ;
        RECT 44.795 171.015 46.005 171.535 ;
        RECT 46.175 171.505 46.515 172.135 ;
        RECT 46.685 171.505 46.935 172.305 ;
        RECT 47.125 171.655 47.455 172.135 ;
        RECT 47.625 171.845 47.850 172.305 ;
        RECT 48.020 171.655 48.350 172.135 ;
        RECT 46.175 170.895 46.350 171.505 ;
        RECT 47.125 171.485 48.350 171.655 ;
        RECT 48.980 171.525 49.480 172.135 ;
        RECT 49.855 171.535 51.525 172.305 ;
        RECT 51.700 171.760 57.045 172.305 ;
        RECT 57.220 171.760 62.565 172.305 ;
        RECT 46.520 171.145 47.215 171.315 ;
        RECT 47.045 170.895 47.215 171.145 ;
        RECT 47.390 171.115 47.810 171.315 ;
        RECT 47.980 171.115 48.310 171.315 ;
        RECT 48.480 171.115 48.810 171.315 ;
        RECT 48.980 170.895 49.150 171.525 ;
        RECT 49.335 171.065 49.685 171.315 ;
        RECT 43.415 169.755 46.005 170.845 ;
        RECT 46.175 169.925 46.515 170.895 ;
        RECT 46.685 169.755 46.855 170.895 ;
        RECT 47.045 170.725 49.480 170.895 ;
        RECT 47.125 169.755 47.375 170.555 ;
        RECT 48.020 169.925 48.350 170.725 ;
        RECT 48.650 169.755 48.980 170.555 ;
        RECT 49.150 169.925 49.480 170.725 ;
        RECT 49.855 170.845 50.605 171.365 ;
        RECT 50.775 171.015 51.525 171.535 ;
        RECT 49.855 169.755 51.525 170.845 ;
        RECT 53.290 170.190 53.640 171.440 ;
        RECT 55.120 170.930 55.460 171.760 ;
        RECT 58.810 170.190 59.160 171.440 ;
        RECT 60.640 170.930 60.980 171.760 ;
        RECT 62.825 171.755 62.995 172.135 ;
        RECT 63.210 171.925 63.540 172.305 ;
        RECT 62.825 171.585 63.540 171.755 ;
        RECT 62.735 171.035 63.090 171.405 ;
        RECT 63.370 171.395 63.540 171.585 ;
        RECT 63.710 171.560 63.965 172.135 ;
        RECT 63.370 171.065 63.625 171.395 ;
        RECT 63.370 170.855 63.540 171.065 ;
        RECT 62.825 170.685 63.540 170.855 ;
        RECT 63.795 170.830 63.965 171.560 ;
        RECT 64.140 171.465 64.400 172.305 ;
        RECT 64.575 171.580 64.865 172.305 ;
        RECT 65.105 171.945 65.435 172.305 ;
        RECT 65.965 171.945 66.295 172.305 ;
        RECT 66.825 171.945 67.155 172.305 ;
        RECT 67.385 171.945 69.455 172.135 ;
        RECT 67.385 171.925 68.505 171.945 ;
        RECT 65.605 171.755 65.795 171.875 ;
        RECT 65.095 171.315 65.435 171.625 ;
        RECT 65.605 171.545 68.145 171.755 ;
        RECT 68.315 171.500 68.505 171.925 ;
        RECT 69.635 171.805 69.895 172.135 ;
        RECT 70.205 171.925 70.535 172.305 ;
        RECT 70.715 171.965 72.195 172.135 ;
        RECT 65.095 171.145 66.045 171.315 ;
        RECT 65.095 171.095 65.990 171.145 ;
        RECT 66.215 171.035 67.185 171.315 ;
        RECT 67.645 171.025 68.505 171.315 ;
        RECT 51.700 169.755 57.045 170.190 ;
        RECT 57.220 169.755 62.565 170.190 ;
        RECT 62.825 169.925 62.995 170.685 ;
        RECT 63.210 169.755 63.540 170.515 ;
        RECT 63.710 169.925 63.965 170.830 ;
        RECT 64.140 169.755 64.400 170.905 ;
        RECT 64.575 169.755 64.865 170.920 ;
        RECT 65.105 170.695 66.225 170.865 ;
        RECT 68.675 170.850 69.005 171.720 ;
        RECT 65.105 169.925 65.365 170.695 ;
        RECT 65.535 169.755 65.865 170.525 ;
        RECT 66.035 170.095 66.225 170.695 ;
        RECT 66.395 170.680 69.005 170.850 ;
        RECT 66.395 170.265 66.725 170.680 ;
        RECT 66.895 170.095 67.155 170.290 ;
        RECT 66.035 169.925 67.155 170.095 ;
        RECT 67.385 169.755 67.715 170.475 ;
        RECT 67.885 169.925 68.075 170.680 ;
        RECT 68.245 169.755 68.575 170.475 ;
        RECT 68.745 169.925 69.005 170.680 ;
        RECT 69.175 170.420 69.465 171.395 ;
        RECT 69.635 171.105 69.805 171.805 ;
        RECT 70.715 171.635 71.115 171.965 ;
        RECT 70.155 171.445 70.365 171.625 ;
        RECT 70.155 171.275 70.775 171.445 ;
        RECT 70.945 171.155 71.115 171.635 ;
        RECT 71.305 171.465 71.855 171.795 ;
        RECT 69.635 170.935 70.765 171.105 ;
        RECT 70.945 170.985 71.515 171.155 ;
        RECT 69.635 170.255 69.805 170.935 ;
        RECT 70.595 170.815 70.765 170.935 ;
        RECT 69.975 170.435 70.325 170.765 ;
        RECT 70.595 170.645 71.175 170.815 ;
        RECT 71.345 170.475 71.515 170.985 ;
        RECT 70.775 170.305 71.515 170.475 ;
        RECT 71.685 170.475 71.855 171.465 ;
        RECT 72.025 171.065 72.195 171.965 ;
        RECT 72.445 171.395 72.630 171.975 ;
        RECT 72.900 171.395 73.095 171.970 ;
        RECT 73.305 171.925 73.635 172.305 ;
        RECT 72.445 171.065 72.675 171.395 ;
        RECT 72.900 171.065 73.155 171.395 ;
        RECT 72.445 170.755 72.630 171.065 ;
        RECT 72.900 170.755 73.095 171.065 ;
        RECT 73.465 170.475 73.635 171.395 ;
        RECT 71.685 170.305 73.635 170.475 ;
        RECT 69.175 169.755 69.435 170.215 ;
        RECT 69.635 169.925 69.895 170.255 ;
        RECT 70.205 169.755 70.535 170.135 ;
        RECT 70.775 169.925 70.965 170.305 ;
        RECT 71.215 169.755 71.545 170.135 ;
        RECT 71.755 169.925 71.925 170.305 ;
        RECT 72.120 169.755 72.450 170.135 ;
        RECT 72.710 169.925 72.880 170.305 ;
        RECT 73.305 169.755 73.635 170.135 ;
        RECT 73.805 169.925 74.065 172.135 ;
        RECT 74.700 171.760 80.045 172.305 ;
        RECT 76.290 170.190 76.640 171.440 ;
        RECT 78.120 170.930 78.460 171.760 ;
        RECT 80.215 171.505 80.555 172.135 ;
        RECT 80.725 171.505 80.975 172.305 ;
        RECT 81.165 171.655 81.495 172.135 ;
        RECT 81.665 171.845 81.890 172.305 ;
        RECT 82.060 171.655 82.390 172.135 ;
        RECT 80.215 170.895 80.390 171.505 ;
        RECT 81.165 171.485 82.390 171.655 ;
        RECT 83.020 171.525 83.520 172.135 ;
        RECT 84.820 171.760 90.165 172.305 ;
        RECT 80.560 171.145 81.255 171.315 ;
        RECT 81.085 170.895 81.255 171.145 ;
        RECT 81.430 171.115 81.850 171.315 ;
        RECT 82.020 171.115 82.350 171.315 ;
        RECT 82.520 171.115 82.850 171.315 ;
        RECT 83.020 170.895 83.190 171.525 ;
        RECT 83.375 171.065 83.725 171.315 ;
        RECT 74.700 169.755 80.045 170.190 ;
        RECT 80.215 169.925 80.555 170.895 ;
        RECT 80.725 169.755 80.895 170.895 ;
        RECT 81.085 170.725 83.520 170.895 ;
        RECT 81.165 169.755 81.415 170.555 ;
        RECT 82.060 169.925 82.390 170.725 ;
        RECT 82.690 169.755 83.020 170.555 ;
        RECT 83.190 169.925 83.520 170.725 ;
        RECT 86.410 170.190 86.760 171.440 ;
        RECT 88.240 170.930 88.580 171.760 ;
        RECT 90.335 171.580 90.625 172.305 ;
        RECT 91.260 171.755 91.515 172.045 ;
        RECT 91.685 171.925 92.015 172.305 ;
        RECT 91.260 171.585 92.010 171.755 ;
        RECT 84.820 169.755 90.165 170.190 ;
        RECT 90.335 169.755 90.625 170.920 ;
        RECT 91.260 170.765 91.610 171.415 ;
        RECT 91.780 170.595 92.010 171.585 ;
        RECT 91.260 170.425 92.010 170.595 ;
        RECT 91.260 169.925 91.515 170.425 ;
        RECT 91.685 169.755 92.015 170.255 ;
        RECT 92.185 169.925 92.355 172.045 ;
        RECT 92.715 171.945 93.045 172.305 ;
        RECT 93.215 171.915 93.710 172.085 ;
        RECT 93.915 171.915 94.770 172.085 ;
        RECT 92.585 170.725 93.045 171.775 ;
        RECT 92.525 169.940 92.850 170.725 ;
        RECT 93.215 170.555 93.385 171.915 ;
        RECT 93.555 171.005 93.905 171.625 ;
        RECT 94.075 171.405 94.430 171.625 ;
        RECT 94.075 170.815 94.245 171.405 ;
        RECT 94.600 171.205 94.770 171.915 ;
        RECT 95.645 171.845 95.975 172.305 ;
        RECT 96.185 171.945 96.535 172.115 ;
        RECT 94.975 171.375 95.765 171.625 ;
        RECT 96.185 171.555 96.445 171.945 ;
        RECT 96.755 171.855 97.705 172.135 ;
        RECT 97.875 171.865 98.065 172.305 ;
        RECT 98.235 171.925 99.305 172.095 ;
        RECT 95.935 171.205 96.105 171.385 ;
        RECT 93.215 170.385 93.610 170.555 ;
        RECT 93.780 170.425 94.245 170.815 ;
        RECT 94.415 171.035 96.105 171.205 ;
        RECT 93.440 170.255 93.610 170.385 ;
        RECT 94.415 170.255 94.585 171.035 ;
        RECT 96.275 170.865 96.445 171.555 ;
        RECT 94.945 170.695 96.445 170.865 ;
        RECT 96.635 170.895 96.845 171.685 ;
        RECT 97.015 171.065 97.365 171.685 ;
        RECT 97.535 171.075 97.705 171.855 ;
        RECT 98.235 171.695 98.405 171.925 ;
        RECT 97.875 171.525 98.405 171.695 ;
        RECT 97.875 171.245 98.095 171.525 ;
        RECT 98.575 171.355 98.815 171.755 ;
        RECT 97.535 170.905 97.940 171.075 ;
        RECT 98.275 170.985 98.815 171.355 ;
        RECT 98.985 171.570 99.305 171.925 ;
        RECT 99.550 171.845 99.855 172.305 ;
        RECT 100.025 171.595 100.280 172.125 ;
        RECT 98.985 171.395 99.310 171.570 ;
        RECT 98.985 171.095 99.900 171.395 ;
        RECT 99.160 171.065 99.900 171.095 ;
        RECT 96.635 170.735 97.310 170.895 ;
        RECT 97.770 170.815 97.940 170.905 ;
        RECT 96.635 170.725 97.600 170.735 ;
        RECT 96.275 170.555 96.445 170.695 ;
        RECT 93.020 169.755 93.270 170.215 ;
        RECT 93.440 169.925 93.690 170.255 ;
        RECT 93.905 169.925 94.585 170.255 ;
        RECT 94.755 170.355 95.830 170.525 ;
        RECT 96.275 170.385 96.835 170.555 ;
        RECT 97.140 170.435 97.600 170.725 ;
        RECT 97.770 170.645 98.990 170.815 ;
        RECT 94.755 170.015 94.925 170.355 ;
        RECT 95.160 169.755 95.490 170.185 ;
        RECT 95.660 170.015 95.830 170.355 ;
        RECT 96.125 169.755 96.495 170.215 ;
        RECT 96.665 169.925 96.835 170.385 ;
        RECT 97.770 170.265 97.940 170.645 ;
        RECT 99.160 170.475 99.330 171.065 ;
        RECT 100.070 170.945 100.280 171.595 ;
        RECT 100.455 171.555 101.665 172.305 ;
        RECT 97.070 169.925 97.940 170.265 ;
        RECT 98.530 170.305 99.330 170.475 ;
        RECT 98.110 169.755 98.360 170.215 ;
        RECT 98.530 170.015 98.700 170.305 ;
        RECT 98.880 169.755 99.210 170.135 ;
        RECT 99.550 169.755 99.855 170.895 ;
        RECT 100.025 170.065 100.280 170.945 ;
        RECT 100.455 170.845 100.975 171.385 ;
        RECT 101.145 171.015 101.665 171.555 ;
        RECT 101.875 171.485 102.105 172.305 ;
        RECT 102.275 171.505 102.605 172.135 ;
        RECT 101.855 171.065 102.185 171.315 ;
        RECT 102.355 170.905 102.605 171.505 ;
        RECT 102.775 171.485 102.985 172.305 ;
        RECT 103.680 171.760 109.025 172.305 ;
        RECT 100.455 169.755 101.665 170.845 ;
        RECT 101.875 169.755 102.105 170.895 ;
        RECT 102.275 169.925 102.605 170.905 ;
        RECT 102.775 169.755 102.985 170.895 ;
        RECT 105.270 170.190 105.620 171.440 ;
        RECT 107.100 170.930 107.440 171.760 ;
        RECT 109.255 171.485 109.465 172.305 ;
        RECT 109.635 171.505 109.965 172.135 ;
        RECT 109.635 170.905 109.885 171.505 ;
        RECT 110.135 171.485 110.365 172.305 ;
        RECT 110.580 171.760 115.925 172.305 ;
        RECT 110.055 171.065 110.385 171.315 ;
        RECT 103.680 169.755 109.025 170.190 ;
        RECT 109.255 169.755 109.465 170.895 ;
        RECT 109.635 169.925 109.965 170.905 ;
        RECT 110.135 169.755 110.365 170.895 ;
        RECT 112.170 170.190 112.520 171.440 ;
        RECT 114.000 170.930 114.340 171.760 ;
        RECT 116.095 171.580 116.385 172.305 ;
        RECT 117.055 171.485 117.285 172.305 ;
        RECT 117.455 171.505 117.785 172.135 ;
        RECT 117.035 171.065 117.365 171.315 ;
        RECT 110.580 169.755 115.925 170.190 ;
        RECT 116.095 169.755 116.385 170.920 ;
        RECT 117.535 170.905 117.785 171.505 ;
        RECT 117.955 171.485 118.165 172.305 ;
        RECT 118.435 171.485 118.665 172.305 ;
        RECT 118.835 171.505 119.165 172.135 ;
        RECT 118.415 171.065 118.745 171.315 ;
        RECT 118.915 170.905 119.165 171.505 ;
        RECT 119.335 171.485 119.545 172.305 ;
        RECT 120.235 171.535 122.825 172.305 ;
        RECT 123.000 171.905 123.335 172.305 ;
        RECT 123.505 171.735 123.710 172.135 ;
        RECT 123.920 171.825 124.195 172.305 ;
        RECT 124.405 171.805 124.665 172.135 ;
        RECT 117.055 169.755 117.285 170.895 ;
        RECT 117.455 169.925 117.785 170.905 ;
        RECT 117.955 169.755 118.165 170.895 ;
        RECT 118.435 169.755 118.665 170.895 ;
        RECT 118.835 169.925 119.165 170.905 ;
        RECT 119.335 169.755 119.545 170.895 ;
        RECT 120.235 170.845 121.445 171.365 ;
        RECT 121.615 171.015 122.825 171.535 ;
        RECT 123.025 171.565 123.710 171.735 ;
        RECT 120.235 169.755 122.825 170.845 ;
        RECT 123.025 170.535 123.365 171.565 ;
        RECT 123.535 170.895 123.785 171.395 ;
        RECT 123.965 171.065 124.325 171.645 ;
        RECT 124.495 170.895 124.665 171.805 ;
        RECT 125.295 171.535 127.885 172.305 ;
        RECT 128.055 171.555 129.265 172.305 ;
        RECT 123.535 170.725 124.665 170.895 ;
        RECT 123.025 170.360 123.690 170.535 ;
        RECT 123.000 169.755 123.335 170.180 ;
        RECT 123.505 169.955 123.690 170.360 ;
        RECT 123.895 169.755 124.225 170.535 ;
        RECT 124.395 169.955 124.665 170.725 ;
        RECT 125.295 170.845 126.505 171.365 ;
        RECT 126.675 171.015 127.885 171.535 ;
        RECT 128.055 170.845 128.575 171.385 ;
        RECT 128.745 171.015 129.265 171.555 ;
        RECT 125.295 169.755 127.885 170.845 ;
        RECT 128.055 169.755 129.265 170.845 ;
        RECT 9.290 169.585 129.350 169.755 ;
        RECT 9.375 168.495 10.585 169.585 ;
        RECT 9.375 167.785 9.895 168.325 ;
        RECT 10.065 167.955 10.585 168.495 ;
        RECT 11.215 168.495 14.725 169.585 ;
        RECT 14.900 169.150 20.245 169.585 ;
        RECT 20.420 169.150 25.765 169.585 ;
        RECT 11.215 167.975 12.905 168.495 ;
        RECT 13.075 167.805 14.725 168.325 ;
        RECT 16.490 167.900 16.840 169.150 ;
        RECT 9.375 167.035 10.585 167.785 ;
        RECT 11.215 167.035 14.725 167.805 ;
        RECT 18.320 167.580 18.660 168.410 ;
        RECT 22.010 167.900 22.360 169.150 ;
        RECT 25.935 168.420 26.225 169.585 ;
        RECT 26.855 168.495 28.525 169.585 ;
        RECT 28.700 169.150 34.045 169.585 ;
        RECT 34.220 169.150 39.565 169.585 ;
        RECT 23.840 167.580 24.180 168.410 ;
        RECT 26.855 167.975 27.605 168.495 ;
        RECT 27.775 167.805 28.525 168.325 ;
        RECT 30.290 167.900 30.640 169.150 ;
        RECT 14.900 167.035 20.245 167.580 ;
        RECT 20.420 167.035 25.765 167.580 ;
        RECT 25.935 167.035 26.225 167.760 ;
        RECT 26.855 167.035 28.525 167.805 ;
        RECT 32.120 167.580 32.460 168.410 ;
        RECT 35.810 167.900 36.160 169.150 ;
        RECT 39.795 168.445 40.005 169.585 ;
        RECT 40.175 168.435 40.505 169.415 ;
        RECT 40.675 168.445 40.905 169.585 ;
        RECT 42.035 168.495 45.545 169.585 ;
        RECT 45.815 169.125 45.985 169.585 ;
        RECT 46.155 168.635 46.485 169.415 ;
        RECT 46.655 168.785 46.825 169.585 ;
        RECT 45.715 168.615 46.485 168.635 ;
        RECT 46.995 168.615 47.325 169.415 ;
        RECT 47.495 168.785 47.665 169.585 ;
        RECT 47.835 168.615 48.165 169.415 ;
        RECT 37.640 167.580 37.980 168.410 ;
        RECT 28.700 167.035 34.045 167.580 ;
        RECT 34.220 167.035 39.565 167.580 ;
        RECT 39.795 167.035 40.005 167.855 ;
        RECT 40.175 167.835 40.425 168.435 ;
        RECT 40.595 168.025 40.925 168.275 ;
        RECT 42.035 167.975 43.725 168.495 ;
        RECT 45.715 168.445 48.165 168.615 ;
        RECT 48.425 168.445 48.720 169.585 ;
        RECT 48.935 168.495 51.525 169.585 ;
        RECT 40.175 167.205 40.505 167.835 ;
        RECT 40.675 167.035 40.905 167.855 ;
        RECT 43.895 167.805 45.545 168.325 ;
        RECT 42.035 167.035 45.545 167.805 ;
        RECT 45.715 167.855 46.065 168.445 ;
        RECT 46.235 168.025 48.745 168.275 ;
        RECT 48.935 167.975 50.145 168.495 ;
        RECT 51.695 168.420 51.985 169.585 ;
        RECT 52.155 168.495 53.365 169.585 ;
        RECT 53.540 169.150 58.885 169.585 ;
        RECT 59.060 169.150 64.405 169.585 ;
        RECT 45.715 167.675 48.085 167.855 ;
        RECT 50.315 167.805 51.525 168.325 ;
        RECT 52.155 167.955 52.675 168.495 ;
        RECT 45.815 167.035 46.065 167.500 ;
        RECT 46.235 167.205 46.405 167.675 ;
        RECT 46.655 167.035 46.825 167.495 ;
        RECT 47.075 167.205 47.245 167.675 ;
        RECT 47.495 167.035 47.665 167.495 ;
        RECT 47.915 167.205 48.085 167.675 ;
        RECT 48.455 167.035 48.720 167.495 ;
        RECT 48.935 167.035 51.525 167.805 ;
        RECT 52.845 167.785 53.365 168.325 ;
        RECT 55.130 167.900 55.480 169.150 ;
        RECT 51.695 167.035 51.985 167.760 ;
        RECT 52.155 167.035 53.365 167.785 ;
        RECT 56.960 167.580 57.300 168.410 ;
        RECT 60.650 167.900 61.000 169.150 ;
        RECT 64.615 168.445 64.845 169.585 ;
        RECT 65.015 168.435 65.345 169.415 ;
        RECT 65.515 168.445 65.725 169.585 ;
        RECT 66.045 168.655 66.215 169.415 ;
        RECT 66.430 168.825 66.760 169.585 ;
        RECT 66.045 168.485 66.760 168.655 ;
        RECT 66.930 168.510 67.185 169.415 ;
        RECT 62.480 167.580 62.820 168.410 ;
        RECT 64.595 168.025 64.925 168.275 ;
        RECT 53.540 167.035 58.885 167.580 ;
        RECT 59.060 167.035 64.405 167.580 ;
        RECT 64.615 167.035 64.845 167.855 ;
        RECT 65.095 167.835 65.345 168.435 ;
        RECT 65.955 167.935 66.310 168.305 ;
        RECT 66.590 168.275 66.760 168.485 ;
        RECT 66.590 167.945 66.845 168.275 ;
        RECT 65.015 167.205 65.345 167.835 ;
        RECT 65.515 167.035 65.725 167.855 ;
        RECT 66.590 167.755 66.760 167.945 ;
        RECT 67.015 167.780 67.185 168.510 ;
        RECT 67.360 168.435 67.620 169.585 ;
        RECT 66.045 167.585 66.760 167.755 ;
        RECT 66.045 167.205 66.215 167.585 ;
        RECT 66.430 167.035 66.760 167.415 ;
        RECT 66.930 167.205 67.185 167.780 ;
        RECT 67.360 167.035 67.620 167.875 ;
        RECT 67.795 167.775 68.055 169.400 ;
        RECT 69.805 169.135 70.135 169.585 ;
        RECT 71.940 169.150 77.285 169.585 ;
        RECT 68.235 168.745 70.845 168.955 ;
        RECT 68.235 167.945 68.455 168.745 ;
        RECT 68.695 167.945 68.995 168.565 ;
        RECT 69.165 167.945 69.495 168.565 ;
        RECT 69.665 167.945 69.985 168.565 ;
        RECT 70.155 167.945 70.505 168.565 ;
        RECT 70.675 167.775 70.845 168.745 ;
        RECT 73.530 167.900 73.880 169.150 ;
        RECT 77.455 168.420 77.745 169.585 ;
        RECT 78.375 168.495 80.965 169.585 ;
        RECT 81.135 168.825 81.650 169.235 ;
        RECT 81.885 168.825 82.055 169.585 ;
        RECT 82.225 169.245 84.255 169.415 ;
        RECT 67.795 167.605 69.635 167.775 ;
        RECT 68.065 167.035 68.395 167.430 ;
        RECT 68.565 167.250 68.765 167.605 ;
        RECT 68.935 167.035 69.265 167.435 ;
        RECT 69.435 167.260 69.635 167.605 ;
        RECT 69.805 167.035 70.135 167.775 ;
        RECT 70.370 167.605 70.845 167.775 ;
        RECT 70.370 167.355 70.540 167.605 ;
        RECT 75.360 167.580 75.700 168.410 ;
        RECT 78.375 167.975 79.585 168.495 ;
        RECT 79.755 167.805 80.965 168.325 ;
        RECT 81.135 168.015 81.475 168.825 ;
        RECT 82.225 168.580 82.395 169.245 ;
        RECT 82.790 168.905 83.915 169.075 ;
        RECT 81.645 168.390 82.395 168.580 ;
        RECT 82.565 168.565 83.575 168.735 ;
        RECT 81.135 167.845 82.365 168.015 ;
        RECT 71.940 167.035 77.285 167.580 ;
        RECT 77.455 167.035 77.745 167.760 ;
        RECT 78.375 167.035 80.965 167.805 ;
        RECT 81.410 167.240 81.655 167.845 ;
        RECT 81.875 167.035 82.385 167.570 ;
        RECT 82.565 167.205 82.755 168.565 ;
        RECT 82.925 167.545 83.200 168.365 ;
        RECT 83.405 167.765 83.575 168.565 ;
        RECT 83.745 167.775 83.915 168.905 ;
        RECT 84.085 168.275 84.255 169.245 ;
        RECT 84.425 168.445 84.595 169.585 ;
        RECT 84.765 168.445 85.100 169.415 ;
        RECT 86.255 168.445 86.465 169.585 ;
        RECT 84.085 167.945 84.280 168.275 ;
        RECT 84.505 167.945 84.760 168.275 ;
        RECT 84.505 167.775 84.675 167.945 ;
        RECT 84.930 167.775 85.100 168.445 ;
        RECT 86.635 168.435 86.965 169.415 ;
        RECT 87.135 168.445 87.365 169.585 ;
        RECT 88.495 168.495 92.005 169.585 ;
        RECT 92.175 168.825 92.690 169.235 ;
        RECT 92.925 168.825 93.095 169.585 ;
        RECT 93.265 169.245 95.295 169.415 ;
        RECT 83.745 167.605 84.675 167.775 ;
        RECT 83.745 167.570 83.920 167.605 ;
        RECT 82.925 167.375 83.205 167.545 ;
        RECT 82.925 167.205 83.200 167.375 ;
        RECT 83.390 167.205 83.920 167.570 ;
        RECT 84.345 167.035 84.675 167.435 ;
        RECT 84.845 167.205 85.100 167.775 ;
        RECT 86.255 167.035 86.465 167.855 ;
        RECT 86.635 167.835 86.885 168.435 ;
        RECT 87.055 168.025 87.385 168.275 ;
        RECT 88.495 167.975 90.185 168.495 ;
        RECT 86.635 167.205 86.965 167.835 ;
        RECT 87.135 167.035 87.365 167.855 ;
        RECT 90.355 167.805 92.005 168.325 ;
        RECT 92.175 168.015 92.515 168.825 ;
        RECT 93.265 168.580 93.435 169.245 ;
        RECT 93.830 168.905 94.955 169.075 ;
        RECT 92.685 168.390 93.435 168.580 ;
        RECT 93.605 168.565 94.615 168.735 ;
        RECT 92.175 167.845 93.405 168.015 ;
        RECT 88.495 167.035 92.005 167.805 ;
        RECT 92.450 167.240 92.695 167.845 ;
        RECT 92.915 167.035 93.425 167.570 ;
        RECT 93.605 167.205 93.795 168.565 ;
        RECT 93.965 167.885 94.240 168.365 ;
        RECT 93.965 167.715 94.245 167.885 ;
        RECT 94.445 167.765 94.615 168.565 ;
        RECT 94.785 167.775 94.955 168.905 ;
        RECT 95.125 168.275 95.295 169.245 ;
        RECT 95.465 168.445 95.635 169.585 ;
        RECT 95.805 168.445 96.140 169.415 ;
        RECT 95.125 167.945 95.320 168.275 ;
        RECT 95.545 167.945 95.800 168.275 ;
        RECT 95.545 167.775 95.715 167.945 ;
        RECT 95.970 167.775 96.140 168.445 ;
        RECT 93.965 167.205 94.240 167.715 ;
        RECT 94.785 167.605 95.715 167.775 ;
        RECT 94.785 167.570 94.960 167.605 ;
        RECT 94.430 167.205 94.960 167.570 ;
        RECT 95.385 167.035 95.715 167.435 ;
        RECT 95.885 167.205 96.140 167.775 ;
        RECT 96.775 168.510 97.045 169.415 ;
        RECT 97.215 168.825 97.545 169.585 ;
        RECT 97.725 168.655 97.895 169.415 ;
        RECT 96.775 167.710 96.945 168.510 ;
        RECT 97.230 168.485 97.895 168.655 ;
        RECT 99.075 168.825 99.590 169.235 ;
        RECT 99.825 168.825 99.995 169.585 ;
        RECT 100.165 169.245 102.195 169.415 ;
        RECT 97.230 168.340 97.400 168.485 ;
        RECT 97.115 168.010 97.400 168.340 ;
        RECT 97.230 167.755 97.400 168.010 ;
        RECT 97.635 167.935 97.965 168.305 ;
        RECT 99.075 168.015 99.415 168.825 ;
        RECT 100.165 168.580 100.335 169.245 ;
        RECT 100.730 168.905 101.855 169.075 ;
        RECT 99.585 168.390 100.335 168.580 ;
        RECT 100.505 168.565 101.515 168.735 ;
        RECT 99.075 167.845 100.305 168.015 ;
        RECT 96.775 167.205 97.035 167.710 ;
        RECT 97.230 167.585 97.895 167.755 ;
        RECT 97.215 167.035 97.545 167.415 ;
        RECT 97.725 167.205 97.895 167.585 ;
        RECT 99.350 167.240 99.595 167.845 ;
        RECT 99.815 167.035 100.325 167.570 ;
        RECT 100.505 167.205 100.695 168.565 ;
        RECT 100.865 168.225 101.140 168.365 ;
        RECT 100.865 168.055 101.145 168.225 ;
        RECT 100.865 167.205 101.140 168.055 ;
        RECT 101.345 167.765 101.515 168.565 ;
        RECT 101.685 167.775 101.855 168.905 ;
        RECT 102.025 168.275 102.195 169.245 ;
        RECT 102.365 168.445 102.535 169.585 ;
        RECT 102.705 168.445 103.040 169.415 ;
        RECT 102.025 167.945 102.220 168.275 ;
        RECT 102.445 167.945 102.700 168.275 ;
        RECT 102.445 167.775 102.615 167.945 ;
        RECT 102.870 167.775 103.040 168.445 ;
        RECT 103.215 168.420 103.505 169.585 ;
        RECT 101.685 167.605 102.615 167.775 ;
        RECT 101.685 167.570 101.860 167.605 ;
        RECT 101.330 167.205 101.860 167.570 ;
        RECT 102.285 167.035 102.615 167.435 ;
        RECT 102.785 167.205 103.040 167.775 ;
        RECT 103.680 168.395 103.935 169.275 ;
        RECT 104.105 168.445 104.410 169.585 ;
        RECT 104.750 169.205 105.080 169.585 ;
        RECT 105.260 169.035 105.430 169.325 ;
        RECT 105.600 169.125 105.850 169.585 ;
        RECT 104.630 168.865 105.430 169.035 ;
        RECT 106.020 169.075 106.890 169.415 ;
        RECT 103.215 167.035 103.505 167.760 ;
        RECT 103.680 167.745 103.890 168.395 ;
        RECT 104.630 168.275 104.800 168.865 ;
        RECT 106.020 168.695 106.190 169.075 ;
        RECT 107.125 168.955 107.295 169.415 ;
        RECT 107.465 169.125 107.835 169.585 ;
        RECT 108.130 168.985 108.300 169.325 ;
        RECT 108.470 169.155 108.800 169.585 ;
        RECT 109.035 168.985 109.205 169.325 ;
        RECT 104.970 168.525 106.190 168.695 ;
        RECT 106.360 168.615 106.820 168.905 ;
        RECT 107.125 168.785 107.685 168.955 ;
        RECT 108.130 168.815 109.205 168.985 ;
        RECT 109.375 169.085 110.055 169.415 ;
        RECT 110.270 169.085 110.520 169.415 ;
        RECT 110.690 169.125 110.940 169.585 ;
        RECT 107.515 168.645 107.685 168.785 ;
        RECT 106.360 168.605 107.325 168.615 ;
        RECT 106.020 168.435 106.190 168.525 ;
        RECT 106.650 168.445 107.325 168.605 ;
        RECT 104.060 168.245 104.800 168.275 ;
        RECT 104.060 167.945 104.975 168.245 ;
        RECT 104.650 167.770 104.975 167.945 ;
        RECT 103.680 167.215 103.935 167.745 ;
        RECT 104.105 167.035 104.410 167.495 ;
        RECT 104.655 167.415 104.975 167.770 ;
        RECT 105.145 167.985 105.685 168.355 ;
        RECT 106.020 168.265 106.425 168.435 ;
        RECT 105.145 167.585 105.385 167.985 ;
        RECT 105.865 167.815 106.085 168.095 ;
        RECT 105.555 167.645 106.085 167.815 ;
        RECT 105.555 167.415 105.725 167.645 ;
        RECT 106.255 167.485 106.425 168.265 ;
        RECT 106.595 167.655 106.945 168.275 ;
        RECT 107.115 167.655 107.325 168.445 ;
        RECT 107.515 168.475 109.015 168.645 ;
        RECT 107.515 167.785 107.685 168.475 ;
        RECT 109.375 168.305 109.545 169.085 ;
        RECT 110.350 168.955 110.520 169.085 ;
        RECT 107.855 168.135 109.545 168.305 ;
        RECT 109.715 168.525 110.180 168.915 ;
        RECT 110.350 168.785 110.745 168.955 ;
        RECT 107.855 167.955 108.025 168.135 ;
        RECT 104.655 167.245 105.725 167.415 ;
        RECT 105.895 167.035 106.085 167.475 ;
        RECT 106.255 167.205 107.205 167.485 ;
        RECT 107.515 167.395 107.775 167.785 ;
        RECT 108.195 167.715 108.985 167.965 ;
        RECT 107.425 167.225 107.775 167.395 ;
        RECT 107.985 167.035 108.315 167.495 ;
        RECT 109.190 167.425 109.360 168.135 ;
        RECT 109.715 167.935 109.885 168.525 ;
        RECT 109.530 167.715 109.885 167.935 ;
        RECT 110.055 167.715 110.405 168.335 ;
        RECT 110.575 167.425 110.745 168.785 ;
        RECT 111.110 168.615 111.435 169.400 ;
        RECT 110.915 167.565 111.375 168.615 ;
        RECT 109.190 167.255 110.045 167.425 ;
        RECT 110.250 167.255 110.745 167.425 ;
        RECT 110.915 167.035 111.245 167.395 ;
        RECT 111.605 167.295 111.775 169.415 ;
        RECT 111.945 169.085 112.275 169.585 ;
        RECT 112.445 168.915 112.700 169.415 ;
        RECT 111.950 168.745 112.700 168.915 ;
        RECT 112.875 168.825 113.390 169.235 ;
        RECT 113.625 168.825 113.795 169.585 ;
        RECT 113.965 169.245 115.995 169.415 ;
        RECT 111.950 167.755 112.180 168.745 ;
        RECT 112.350 167.925 112.700 168.575 ;
        RECT 112.875 168.015 113.215 168.825 ;
        RECT 113.965 168.580 114.135 169.245 ;
        RECT 114.530 168.905 115.655 169.075 ;
        RECT 113.385 168.390 114.135 168.580 ;
        RECT 114.305 168.565 115.315 168.735 ;
        RECT 112.875 167.845 114.105 168.015 ;
        RECT 111.950 167.585 112.700 167.755 ;
        RECT 111.945 167.035 112.275 167.415 ;
        RECT 112.445 167.295 112.700 167.585 ;
        RECT 113.150 167.240 113.395 167.845 ;
        RECT 113.615 167.035 114.125 167.570 ;
        RECT 114.305 167.205 114.495 168.565 ;
        RECT 114.665 167.545 114.940 168.365 ;
        RECT 115.145 167.765 115.315 168.565 ;
        RECT 115.485 167.775 115.655 168.905 ;
        RECT 115.825 168.275 115.995 169.245 ;
        RECT 116.165 168.445 116.335 169.585 ;
        RECT 116.505 168.445 116.840 169.415 ;
        RECT 115.825 167.945 116.020 168.275 ;
        RECT 116.245 167.945 116.500 168.275 ;
        RECT 116.245 167.775 116.415 167.945 ;
        RECT 116.670 167.775 116.840 168.445 ;
        RECT 115.485 167.605 116.415 167.775 ;
        RECT 115.485 167.570 115.660 167.605 ;
        RECT 114.665 167.375 114.945 167.545 ;
        RECT 114.665 167.205 114.940 167.375 ;
        RECT 115.130 167.205 115.660 167.570 ;
        RECT 116.085 167.035 116.415 167.435 ;
        RECT 116.585 167.205 116.840 167.775 ;
        RECT 117.020 168.395 117.275 169.275 ;
        RECT 117.445 168.445 117.750 169.585 ;
        RECT 118.090 169.205 118.420 169.585 ;
        RECT 118.600 169.035 118.770 169.325 ;
        RECT 118.940 169.125 119.190 169.585 ;
        RECT 117.970 168.865 118.770 169.035 ;
        RECT 119.360 169.075 120.230 169.415 ;
        RECT 117.020 167.745 117.230 168.395 ;
        RECT 117.970 168.275 118.140 168.865 ;
        RECT 119.360 168.695 119.530 169.075 ;
        RECT 120.465 168.955 120.635 169.415 ;
        RECT 120.805 169.125 121.175 169.585 ;
        RECT 121.470 168.985 121.640 169.325 ;
        RECT 121.810 169.155 122.140 169.585 ;
        RECT 122.375 168.985 122.545 169.325 ;
        RECT 118.310 168.525 119.530 168.695 ;
        RECT 119.700 168.615 120.160 168.905 ;
        RECT 120.465 168.785 121.025 168.955 ;
        RECT 121.470 168.815 122.545 168.985 ;
        RECT 122.715 169.085 123.395 169.415 ;
        RECT 123.610 169.085 123.860 169.415 ;
        RECT 124.030 169.125 124.280 169.585 ;
        RECT 120.855 168.645 121.025 168.785 ;
        RECT 119.700 168.605 120.665 168.615 ;
        RECT 119.360 168.435 119.530 168.525 ;
        RECT 119.990 168.445 120.665 168.605 ;
        RECT 117.400 168.245 118.140 168.275 ;
        RECT 117.400 167.945 118.315 168.245 ;
        RECT 117.990 167.770 118.315 167.945 ;
        RECT 117.020 167.215 117.275 167.745 ;
        RECT 117.445 167.035 117.750 167.495 ;
        RECT 117.995 167.415 118.315 167.770 ;
        RECT 118.485 167.985 119.025 168.355 ;
        RECT 119.360 168.265 119.765 168.435 ;
        RECT 118.485 167.585 118.725 167.985 ;
        RECT 119.205 167.815 119.425 168.095 ;
        RECT 118.895 167.645 119.425 167.815 ;
        RECT 118.895 167.415 119.065 167.645 ;
        RECT 119.595 167.485 119.765 168.265 ;
        RECT 119.935 167.655 120.285 168.275 ;
        RECT 120.455 167.655 120.665 168.445 ;
        RECT 120.855 168.475 122.355 168.645 ;
        RECT 120.855 167.785 121.025 168.475 ;
        RECT 122.715 168.305 122.885 169.085 ;
        RECT 123.690 168.955 123.860 169.085 ;
        RECT 121.195 168.135 122.885 168.305 ;
        RECT 123.055 168.525 123.520 168.915 ;
        RECT 123.690 168.785 124.085 168.955 ;
        RECT 121.195 167.955 121.365 168.135 ;
        RECT 117.995 167.245 119.065 167.415 ;
        RECT 119.235 167.035 119.425 167.475 ;
        RECT 119.595 167.205 120.545 167.485 ;
        RECT 120.855 167.395 121.115 167.785 ;
        RECT 121.535 167.715 122.325 167.965 ;
        RECT 120.765 167.225 121.115 167.395 ;
        RECT 121.325 167.035 121.655 167.495 ;
        RECT 122.530 167.425 122.700 168.135 ;
        RECT 123.055 167.935 123.225 168.525 ;
        RECT 122.870 167.715 123.225 167.935 ;
        RECT 123.395 167.715 123.745 168.335 ;
        RECT 123.915 167.425 124.085 168.785 ;
        RECT 124.450 168.615 124.775 169.400 ;
        RECT 124.255 167.565 124.715 168.615 ;
        RECT 122.530 167.255 123.385 167.425 ;
        RECT 123.590 167.255 124.085 167.425 ;
        RECT 124.255 167.035 124.585 167.395 ;
        RECT 124.945 167.295 125.115 169.415 ;
        RECT 125.285 169.085 125.615 169.585 ;
        RECT 125.785 168.915 126.040 169.415 ;
        RECT 125.290 168.745 126.040 168.915 ;
        RECT 125.290 167.755 125.520 168.745 ;
        RECT 125.690 167.925 126.040 168.575 ;
        RECT 126.215 168.495 127.885 169.585 ;
        RECT 128.055 168.495 129.265 169.585 ;
        RECT 126.215 167.975 126.965 168.495 ;
        RECT 127.135 167.805 127.885 168.325 ;
        RECT 128.055 167.955 128.575 168.495 ;
        RECT 125.290 167.585 126.040 167.755 ;
        RECT 125.285 167.035 125.615 167.415 ;
        RECT 125.785 167.295 126.040 167.585 ;
        RECT 126.215 167.035 127.885 167.805 ;
        RECT 128.745 167.785 129.265 168.325 ;
        RECT 128.055 167.035 129.265 167.785 ;
        RECT 9.290 166.865 129.350 167.035 ;
        RECT 9.375 166.115 10.585 166.865 ;
        RECT 9.375 165.575 9.895 166.115 ;
        RECT 11.215 166.095 12.885 166.865 ;
        RECT 13.055 166.140 13.345 166.865 ;
        RECT 13.515 166.115 14.725 166.865 ;
        RECT 14.900 166.315 15.155 166.605 ;
        RECT 15.325 166.485 15.655 166.865 ;
        RECT 14.900 166.145 15.650 166.315 ;
        RECT 10.065 165.405 10.585 165.945 ;
        RECT 9.375 164.315 10.585 165.405 ;
        RECT 11.215 165.405 11.965 165.925 ;
        RECT 12.135 165.575 12.885 166.095 ;
        RECT 11.215 164.315 12.885 165.405 ;
        RECT 13.055 164.315 13.345 165.480 ;
        RECT 13.515 165.405 14.035 165.945 ;
        RECT 14.205 165.575 14.725 166.115 ;
        RECT 13.515 164.315 14.725 165.405 ;
        RECT 14.900 165.325 15.250 165.975 ;
        RECT 15.420 165.155 15.650 166.145 ;
        RECT 14.900 164.985 15.650 165.155 ;
        RECT 14.900 164.485 15.155 164.985 ;
        RECT 15.325 164.315 15.655 164.815 ;
        RECT 15.825 164.485 15.995 166.605 ;
        RECT 16.355 166.505 16.685 166.865 ;
        RECT 16.855 166.475 17.350 166.645 ;
        RECT 17.555 166.475 18.410 166.645 ;
        RECT 16.225 165.285 16.685 166.335 ;
        RECT 16.165 164.500 16.490 165.285 ;
        RECT 16.855 165.115 17.025 166.475 ;
        RECT 17.195 165.565 17.545 166.185 ;
        RECT 17.715 165.965 18.070 166.185 ;
        RECT 17.715 165.375 17.885 165.965 ;
        RECT 18.240 165.765 18.410 166.475 ;
        RECT 19.285 166.405 19.615 166.865 ;
        RECT 19.825 166.505 20.175 166.675 ;
        RECT 18.615 165.935 19.405 166.185 ;
        RECT 19.825 166.115 20.085 166.505 ;
        RECT 20.395 166.415 21.345 166.695 ;
        RECT 21.515 166.425 21.705 166.865 ;
        RECT 21.875 166.485 22.945 166.655 ;
        RECT 19.575 165.765 19.745 165.945 ;
        RECT 16.855 164.945 17.250 165.115 ;
        RECT 17.420 164.985 17.885 165.375 ;
        RECT 18.055 165.595 19.745 165.765 ;
        RECT 17.080 164.815 17.250 164.945 ;
        RECT 18.055 164.815 18.225 165.595 ;
        RECT 19.915 165.425 20.085 166.115 ;
        RECT 18.585 165.255 20.085 165.425 ;
        RECT 20.275 165.455 20.485 166.245 ;
        RECT 20.655 165.625 21.005 166.245 ;
        RECT 21.175 165.635 21.345 166.415 ;
        RECT 21.875 166.255 22.045 166.485 ;
        RECT 21.515 166.085 22.045 166.255 ;
        RECT 21.515 165.805 21.735 166.085 ;
        RECT 22.215 165.915 22.455 166.315 ;
        RECT 21.175 165.465 21.580 165.635 ;
        RECT 21.915 165.545 22.455 165.915 ;
        RECT 22.625 166.130 22.945 166.485 ;
        RECT 23.190 166.405 23.495 166.865 ;
        RECT 23.665 166.155 23.920 166.685 ;
        RECT 22.625 165.955 22.950 166.130 ;
        RECT 22.625 165.655 23.540 165.955 ;
        RECT 22.800 165.625 23.540 165.655 ;
        RECT 20.275 165.295 20.950 165.455 ;
        RECT 21.410 165.375 21.580 165.465 ;
        RECT 20.275 165.285 21.240 165.295 ;
        RECT 19.915 165.115 20.085 165.255 ;
        RECT 16.660 164.315 16.910 164.775 ;
        RECT 17.080 164.485 17.330 164.815 ;
        RECT 17.545 164.485 18.225 164.815 ;
        RECT 18.395 164.915 19.470 165.085 ;
        RECT 19.915 164.945 20.475 165.115 ;
        RECT 20.780 164.995 21.240 165.285 ;
        RECT 21.410 165.205 22.630 165.375 ;
        RECT 18.395 164.575 18.565 164.915 ;
        RECT 18.800 164.315 19.130 164.745 ;
        RECT 19.300 164.575 19.470 164.915 ;
        RECT 19.765 164.315 20.135 164.775 ;
        RECT 20.305 164.485 20.475 164.945 ;
        RECT 21.410 164.825 21.580 165.205 ;
        RECT 22.800 165.035 22.970 165.625 ;
        RECT 23.710 165.505 23.920 166.155 ;
        RECT 24.155 166.045 24.365 166.865 ;
        RECT 24.535 166.065 24.865 166.695 ;
        RECT 20.710 164.485 21.580 164.825 ;
        RECT 22.170 164.865 22.970 165.035 ;
        RECT 21.750 164.315 22.000 164.775 ;
        RECT 22.170 164.575 22.340 164.865 ;
        RECT 22.520 164.315 22.850 164.695 ;
        RECT 23.190 164.315 23.495 165.455 ;
        RECT 23.665 164.625 23.920 165.505 ;
        RECT 24.535 165.465 24.785 166.065 ;
        RECT 25.035 166.045 25.265 166.865 ;
        RECT 25.935 166.095 27.605 166.865 ;
        RECT 24.955 165.625 25.285 165.875 ;
        RECT 24.155 164.315 24.365 165.455 ;
        RECT 24.535 164.485 24.865 165.465 ;
        RECT 25.035 164.315 25.265 165.455 ;
        RECT 25.935 165.405 26.685 165.925 ;
        RECT 26.855 165.575 27.605 166.095 ;
        RECT 27.815 166.045 28.045 166.865 ;
        RECT 28.215 166.065 28.545 166.695 ;
        RECT 27.795 165.625 28.125 165.875 ;
        RECT 28.295 165.465 28.545 166.065 ;
        RECT 28.715 166.045 28.925 166.865 ;
        RECT 29.160 166.155 29.415 166.685 ;
        RECT 29.585 166.405 29.890 166.865 ;
        RECT 30.135 166.485 31.205 166.655 ;
        RECT 25.935 164.315 27.605 165.405 ;
        RECT 27.815 164.315 28.045 165.455 ;
        RECT 28.215 164.485 28.545 165.465 ;
        RECT 29.160 165.505 29.370 166.155 ;
        RECT 30.135 166.130 30.455 166.485 ;
        RECT 30.130 165.955 30.455 166.130 ;
        RECT 29.540 165.655 30.455 165.955 ;
        RECT 30.625 165.915 30.865 166.315 ;
        RECT 31.035 166.255 31.205 166.485 ;
        RECT 31.375 166.425 31.565 166.865 ;
        RECT 31.735 166.415 32.685 166.695 ;
        RECT 32.905 166.505 33.255 166.675 ;
        RECT 31.035 166.085 31.565 166.255 ;
        RECT 29.540 165.625 30.280 165.655 ;
        RECT 28.715 164.315 28.925 165.455 ;
        RECT 29.160 164.625 29.415 165.505 ;
        RECT 29.585 164.315 29.890 165.455 ;
        RECT 30.110 165.035 30.280 165.625 ;
        RECT 30.625 165.545 31.165 165.915 ;
        RECT 31.345 165.805 31.565 166.085 ;
        RECT 31.735 165.635 31.905 166.415 ;
        RECT 31.500 165.465 31.905 165.635 ;
        RECT 32.075 165.625 32.425 166.245 ;
        RECT 31.500 165.375 31.670 165.465 ;
        RECT 32.595 165.455 32.805 166.245 ;
        RECT 30.450 165.205 31.670 165.375 ;
        RECT 32.130 165.295 32.805 165.455 ;
        RECT 30.110 164.865 30.910 165.035 ;
        RECT 30.230 164.315 30.560 164.695 ;
        RECT 30.740 164.575 30.910 164.865 ;
        RECT 31.500 164.825 31.670 165.205 ;
        RECT 31.840 165.285 32.805 165.295 ;
        RECT 32.995 166.115 33.255 166.505 ;
        RECT 33.465 166.405 33.795 166.865 ;
        RECT 34.670 166.475 35.525 166.645 ;
        RECT 35.730 166.475 36.225 166.645 ;
        RECT 36.395 166.505 36.725 166.865 ;
        RECT 32.995 165.425 33.165 166.115 ;
        RECT 33.335 165.765 33.505 165.945 ;
        RECT 33.675 165.935 34.465 166.185 ;
        RECT 34.670 165.765 34.840 166.475 ;
        RECT 35.010 165.965 35.365 166.185 ;
        RECT 33.335 165.595 35.025 165.765 ;
        RECT 31.840 164.995 32.300 165.285 ;
        RECT 32.995 165.255 34.495 165.425 ;
        RECT 32.995 165.115 33.165 165.255 ;
        RECT 32.605 164.945 33.165 165.115 ;
        RECT 31.080 164.315 31.330 164.775 ;
        RECT 31.500 164.485 32.370 164.825 ;
        RECT 32.605 164.485 32.775 164.945 ;
        RECT 33.610 164.915 34.685 165.085 ;
        RECT 32.945 164.315 33.315 164.775 ;
        RECT 33.610 164.575 33.780 164.915 ;
        RECT 33.950 164.315 34.280 164.745 ;
        RECT 34.515 164.575 34.685 164.915 ;
        RECT 34.855 164.815 35.025 165.595 ;
        RECT 35.195 165.375 35.365 165.965 ;
        RECT 35.535 165.565 35.885 166.185 ;
        RECT 35.195 164.985 35.660 165.375 ;
        RECT 36.055 165.115 36.225 166.475 ;
        RECT 36.395 165.285 36.855 166.335 ;
        RECT 35.830 164.945 36.225 165.115 ;
        RECT 35.830 164.815 36.000 164.945 ;
        RECT 34.855 164.485 35.535 164.815 ;
        RECT 35.750 164.485 36.000 164.815 ;
        RECT 36.170 164.315 36.420 164.775 ;
        RECT 36.590 164.500 36.915 165.285 ;
        RECT 37.085 164.485 37.255 166.605 ;
        RECT 37.425 166.485 37.755 166.865 ;
        RECT 37.925 166.315 38.180 166.605 ;
        RECT 37.430 166.145 38.180 166.315 ;
        RECT 37.430 165.155 37.660 166.145 ;
        RECT 38.815 166.140 39.105 166.865 ;
        RECT 39.735 166.355 40.040 166.865 ;
        RECT 37.830 165.325 38.180 165.975 ;
        RECT 39.735 165.625 40.050 166.185 ;
        RECT 40.220 165.875 40.470 166.685 ;
        RECT 40.640 166.340 40.900 166.865 ;
        RECT 41.080 165.875 41.330 166.685 ;
        RECT 41.500 166.305 41.760 166.865 ;
        RECT 41.930 166.215 42.190 166.670 ;
        RECT 42.360 166.385 42.620 166.865 ;
        RECT 42.790 166.215 43.050 166.670 ;
        RECT 43.220 166.385 43.480 166.865 ;
        RECT 43.650 166.215 43.910 166.670 ;
        RECT 44.080 166.385 44.325 166.865 ;
        RECT 44.495 166.215 44.770 166.670 ;
        RECT 44.940 166.385 45.185 166.865 ;
        RECT 45.355 166.215 45.615 166.670 ;
        RECT 45.795 166.385 46.045 166.865 ;
        RECT 46.215 166.215 46.475 166.670 ;
        RECT 46.655 166.385 46.905 166.865 ;
        RECT 47.075 166.215 47.335 166.670 ;
        RECT 47.515 166.385 47.775 166.865 ;
        RECT 47.945 166.215 48.205 166.670 ;
        RECT 48.375 166.385 48.675 166.865 ;
        RECT 41.930 166.045 48.675 166.215 ;
        RECT 49.455 166.045 49.665 166.865 ;
        RECT 49.835 166.065 50.165 166.695 ;
        RECT 40.220 165.625 47.340 165.875 ;
        RECT 37.430 164.985 38.180 165.155 ;
        RECT 37.425 164.315 37.755 164.815 ;
        RECT 37.925 164.485 38.180 164.985 ;
        RECT 38.815 164.315 39.105 165.480 ;
        RECT 39.745 164.315 40.040 165.125 ;
        RECT 40.220 164.485 40.465 165.625 ;
        RECT 40.640 164.315 40.900 165.125 ;
        RECT 41.080 164.490 41.330 165.625 ;
        RECT 47.510 165.505 48.675 166.045 ;
        RECT 47.510 165.455 48.705 165.505 ;
        RECT 49.835 165.465 50.085 166.065 ;
        RECT 50.335 166.045 50.565 166.865 ;
        RECT 50.775 166.095 52.445 166.865 ;
        RECT 50.255 165.625 50.585 165.875 ;
        RECT 41.930 165.335 48.705 165.455 ;
        RECT 41.930 165.230 48.675 165.335 ;
        RECT 41.930 165.215 47.335 165.230 ;
        RECT 41.500 164.320 41.760 165.115 ;
        RECT 41.930 164.490 42.190 165.215 ;
        RECT 42.360 164.320 42.620 165.045 ;
        RECT 42.790 164.490 43.050 165.215 ;
        RECT 43.220 164.320 43.480 165.045 ;
        RECT 43.650 164.490 43.910 165.215 ;
        RECT 44.080 164.320 44.340 165.045 ;
        RECT 44.510 164.490 44.770 165.215 ;
        RECT 44.940 164.320 45.185 165.045 ;
        RECT 45.355 164.490 45.615 165.215 ;
        RECT 45.800 164.320 46.045 165.045 ;
        RECT 46.215 164.490 46.475 165.215 ;
        RECT 46.660 164.320 46.905 165.045 ;
        RECT 47.075 164.490 47.335 165.215 ;
        RECT 47.520 164.320 47.775 165.045 ;
        RECT 47.945 164.490 48.235 165.230 ;
        RECT 41.500 164.315 47.775 164.320 ;
        RECT 48.405 164.315 48.675 165.060 ;
        RECT 49.455 164.315 49.665 165.455 ;
        RECT 49.835 164.485 50.165 165.465 ;
        RECT 50.335 164.315 50.565 165.455 ;
        RECT 50.775 165.405 51.525 165.925 ;
        RECT 51.695 165.575 52.445 166.095 ;
        RECT 52.765 166.065 53.095 166.865 ;
        RECT 53.265 166.215 53.435 166.695 ;
        RECT 53.605 166.385 53.935 166.865 ;
        RECT 54.105 166.215 54.275 166.695 ;
        RECT 54.525 166.385 54.765 166.865 ;
        RECT 54.945 166.215 55.115 166.695 ;
        RECT 53.265 166.045 54.275 166.215 ;
        RECT 54.480 166.045 55.115 166.215 ;
        RECT 55.375 166.115 56.585 166.865 ;
        RECT 53.265 165.845 53.760 166.045 ;
        RECT 54.480 165.875 54.650 166.045 ;
        RECT 53.265 165.675 53.765 165.845 ;
        RECT 54.150 165.705 54.650 165.875 ;
        RECT 53.265 165.505 53.760 165.675 ;
        RECT 50.775 164.315 52.445 165.405 ;
        RECT 52.765 164.315 53.095 165.465 ;
        RECT 53.265 165.335 54.275 165.505 ;
        RECT 53.265 164.485 53.435 165.335 ;
        RECT 53.605 164.315 53.935 165.115 ;
        RECT 54.105 164.485 54.275 165.335 ;
        RECT 54.480 165.465 54.650 165.705 ;
        RECT 54.820 165.635 55.200 165.875 ;
        RECT 54.480 165.295 55.195 165.465 ;
        RECT 54.455 164.315 54.695 165.115 ;
        RECT 54.865 164.485 55.195 165.295 ;
        RECT 55.375 165.405 55.895 165.945 ;
        RECT 56.065 165.575 56.585 166.115 ;
        RECT 56.905 166.065 57.235 166.865 ;
        RECT 57.405 166.215 57.575 166.695 ;
        RECT 57.745 166.385 58.075 166.865 ;
        RECT 58.245 166.215 58.415 166.695 ;
        RECT 58.665 166.385 58.905 166.865 ;
        RECT 59.085 166.215 59.255 166.695 ;
        RECT 57.405 166.045 58.415 166.215 ;
        RECT 58.620 166.045 59.255 166.215 ;
        RECT 59.515 166.115 60.725 166.865 ;
        RECT 57.405 165.505 57.900 166.045 ;
        RECT 58.620 165.875 58.790 166.045 ;
        RECT 58.290 165.705 58.790 165.875 ;
        RECT 55.375 164.315 56.585 165.405 ;
        RECT 56.905 164.315 57.235 165.465 ;
        RECT 57.405 165.335 58.415 165.505 ;
        RECT 57.405 164.485 57.575 165.335 ;
        RECT 57.745 164.315 58.075 165.115 ;
        RECT 58.245 164.485 58.415 165.335 ;
        RECT 58.620 165.465 58.790 165.705 ;
        RECT 58.960 165.635 59.340 165.875 ;
        RECT 58.620 165.295 59.335 165.465 ;
        RECT 58.595 164.315 58.835 165.115 ;
        RECT 59.005 164.485 59.335 165.295 ;
        RECT 59.515 165.405 60.035 165.945 ;
        RECT 60.205 165.575 60.725 166.115 ;
        RECT 60.895 166.095 64.405 166.865 ;
        RECT 64.575 166.140 64.865 166.865 ;
        RECT 65.495 166.095 68.085 166.865 ;
        RECT 60.895 165.405 62.585 165.925 ;
        RECT 62.755 165.575 64.405 166.095 ;
        RECT 59.515 164.315 60.725 165.405 ;
        RECT 60.895 164.315 64.405 165.405 ;
        RECT 64.575 164.315 64.865 165.480 ;
        RECT 65.495 165.405 66.705 165.925 ;
        RECT 66.875 165.575 68.085 166.095 ;
        RECT 68.260 166.025 68.520 166.865 ;
        RECT 68.695 166.120 68.950 166.695 ;
        RECT 69.120 166.485 69.450 166.865 ;
        RECT 69.665 166.315 69.835 166.695 ;
        RECT 69.120 166.145 69.835 166.315 ;
        RECT 65.495 164.315 68.085 165.405 ;
        RECT 68.260 164.315 68.520 165.465 ;
        RECT 68.695 165.390 68.865 166.120 ;
        RECT 69.120 165.955 69.290 166.145 ;
        RECT 70.095 166.095 73.605 166.865 ;
        RECT 73.780 166.320 79.125 166.865 ;
        RECT 69.035 165.625 69.290 165.955 ;
        RECT 69.120 165.415 69.290 165.625 ;
        RECT 69.570 165.595 69.925 165.965 ;
        RECT 68.695 164.485 68.950 165.390 ;
        RECT 69.120 165.245 69.835 165.415 ;
        RECT 69.120 164.315 69.450 165.075 ;
        RECT 69.665 164.485 69.835 165.245 ;
        RECT 70.095 165.405 71.785 165.925 ;
        RECT 71.955 165.575 73.605 166.095 ;
        RECT 70.095 164.315 73.605 165.405 ;
        RECT 75.370 164.750 75.720 166.000 ;
        RECT 77.200 165.490 77.540 166.320 ;
        RECT 79.385 166.315 79.555 166.695 ;
        RECT 79.735 166.485 80.065 166.865 ;
        RECT 79.385 166.145 80.050 166.315 ;
        RECT 80.245 166.190 80.505 166.695 ;
        RECT 79.315 165.595 79.645 165.965 ;
        RECT 79.880 165.890 80.050 166.145 ;
        RECT 79.880 165.560 80.165 165.890 ;
        RECT 79.880 165.415 80.050 165.560 ;
        RECT 79.385 165.245 80.050 165.415 ;
        RECT 80.335 165.390 80.505 166.190 ;
        RECT 73.780 164.315 79.125 164.750 ;
        RECT 79.385 164.485 79.555 165.245 ;
        RECT 79.735 164.315 80.065 165.075 ;
        RECT 80.235 164.485 80.505 165.390 ;
        RECT 81.050 166.155 81.305 166.685 ;
        RECT 81.485 166.405 81.770 166.865 ;
        RECT 81.050 165.295 81.230 166.155 ;
        RECT 81.950 165.955 82.200 166.605 ;
        RECT 81.400 165.625 82.200 165.955 ;
        RECT 81.050 165.165 81.305 165.295 ;
        RECT 80.965 164.995 81.305 165.165 ;
        RECT 81.050 164.625 81.305 164.995 ;
        RECT 81.485 164.315 81.770 165.115 ;
        RECT 81.950 165.035 82.200 165.625 ;
        RECT 82.400 166.270 82.720 166.600 ;
        RECT 82.900 166.385 83.560 166.865 ;
        RECT 83.760 166.475 84.610 166.645 ;
        RECT 82.400 165.375 82.590 166.270 ;
        RECT 82.910 165.945 83.570 166.215 ;
        RECT 83.240 165.885 83.570 165.945 ;
        RECT 82.760 165.715 83.090 165.775 ;
        RECT 83.760 165.715 83.930 166.475 ;
        RECT 85.170 166.405 85.490 166.865 ;
        RECT 85.690 166.225 85.940 166.655 ;
        RECT 86.230 166.425 86.640 166.865 ;
        RECT 86.810 166.485 87.825 166.685 ;
        RECT 84.100 166.055 85.350 166.225 ;
        RECT 84.100 165.935 84.430 166.055 ;
        RECT 82.760 165.545 84.660 165.715 ;
        RECT 82.400 165.205 84.320 165.375 ;
        RECT 82.400 165.185 82.720 165.205 ;
        RECT 81.950 164.525 82.280 165.035 ;
        RECT 82.550 164.575 82.720 165.185 ;
        RECT 84.490 165.035 84.660 165.545 ;
        RECT 84.830 165.475 85.010 165.885 ;
        RECT 85.180 165.295 85.350 166.055 ;
        RECT 82.890 164.315 83.220 165.005 ;
        RECT 83.450 164.865 84.660 165.035 ;
        RECT 84.830 164.985 85.350 165.295 ;
        RECT 85.520 165.885 85.940 166.225 ;
        RECT 86.230 165.885 86.640 166.215 ;
        RECT 85.520 165.115 85.710 165.885 ;
        RECT 86.810 165.755 86.980 166.485 ;
        RECT 88.125 166.315 88.295 166.645 ;
        RECT 88.465 166.485 88.795 166.865 ;
        RECT 87.150 165.935 87.500 166.305 ;
        RECT 86.810 165.715 87.230 165.755 ;
        RECT 85.880 165.545 87.230 165.715 ;
        RECT 85.880 165.385 86.130 165.545 ;
        RECT 86.640 165.115 86.890 165.375 ;
        RECT 85.520 164.865 86.890 165.115 ;
        RECT 83.450 164.575 83.690 164.865 ;
        RECT 84.490 164.785 84.660 164.865 ;
        RECT 83.890 164.315 84.310 164.695 ;
        RECT 84.490 164.535 85.120 164.785 ;
        RECT 85.590 164.315 85.920 164.695 ;
        RECT 86.090 164.575 86.260 164.865 ;
        RECT 87.060 164.700 87.230 165.545 ;
        RECT 87.680 165.375 87.900 166.245 ;
        RECT 88.125 166.125 88.820 166.315 ;
        RECT 87.400 164.995 87.900 165.375 ;
        RECT 88.070 165.325 88.480 165.945 ;
        RECT 88.650 165.155 88.820 166.125 ;
        RECT 88.125 164.985 88.820 165.155 ;
        RECT 86.440 164.315 86.820 164.695 ;
        RECT 87.060 164.530 87.890 164.700 ;
        RECT 88.125 164.485 88.295 164.985 ;
        RECT 88.465 164.315 88.795 164.815 ;
        RECT 89.010 164.485 89.235 166.605 ;
        RECT 89.405 166.485 89.735 166.865 ;
        RECT 89.905 166.315 90.075 166.605 ;
        RECT 89.410 166.145 90.075 166.315 ;
        RECT 89.410 165.155 89.640 166.145 ;
        RECT 90.335 166.140 90.625 166.865 ;
        RECT 90.795 166.190 91.055 166.695 ;
        RECT 91.235 166.485 91.565 166.865 ;
        RECT 91.745 166.315 91.915 166.695 ;
        RECT 89.810 165.325 90.160 165.975 ;
        RECT 89.410 164.985 90.075 165.155 ;
        RECT 89.405 164.315 89.735 164.815 ;
        RECT 89.905 164.485 90.075 164.985 ;
        RECT 90.335 164.315 90.625 165.480 ;
        RECT 90.795 165.390 90.965 166.190 ;
        RECT 91.250 166.145 91.915 166.315 ;
        RECT 91.250 165.890 91.420 166.145 ;
        RECT 92.635 166.095 95.225 166.865 ;
        RECT 95.395 166.355 95.700 166.865 ;
        RECT 91.135 165.560 91.420 165.890 ;
        RECT 91.655 165.595 91.985 165.965 ;
        RECT 91.250 165.415 91.420 165.560 ;
        RECT 90.795 164.485 91.065 165.390 ;
        RECT 91.250 165.245 91.915 165.415 ;
        RECT 91.235 164.315 91.565 165.075 ;
        RECT 91.745 164.485 91.915 165.245 ;
        RECT 92.635 165.405 93.845 165.925 ;
        RECT 94.015 165.575 95.225 166.095 ;
        RECT 95.395 165.625 95.710 166.185 ;
        RECT 95.880 165.875 96.130 166.685 ;
        RECT 96.300 166.340 96.560 166.865 ;
        RECT 96.740 165.875 96.990 166.685 ;
        RECT 97.160 166.305 97.420 166.865 ;
        RECT 97.590 166.215 97.850 166.670 ;
        RECT 98.020 166.385 98.280 166.865 ;
        RECT 98.450 166.215 98.710 166.670 ;
        RECT 98.880 166.385 99.140 166.865 ;
        RECT 99.310 166.215 99.570 166.670 ;
        RECT 99.740 166.385 99.985 166.865 ;
        RECT 100.155 166.215 100.430 166.670 ;
        RECT 100.600 166.385 100.845 166.865 ;
        RECT 101.015 166.215 101.275 166.670 ;
        RECT 101.455 166.385 101.705 166.865 ;
        RECT 101.875 166.215 102.135 166.670 ;
        RECT 102.315 166.385 102.565 166.865 ;
        RECT 102.735 166.215 102.995 166.670 ;
        RECT 103.175 166.385 103.435 166.865 ;
        RECT 103.605 166.215 103.865 166.670 ;
        RECT 104.035 166.385 104.335 166.865 ;
        RECT 97.590 166.045 104.335 166.215 ;
        RECT 104.595 166.095 106.265 166.865 ;
        RECT 95.880 165.625 103.000 165.875 ;
        RECT 92.635 164.315 95.225 165.405 ;
        RECT 95.405 164.315 95.700 165.125 ;
        RECT 95.880 164.485 96.125 165.625 ;
        RECT 96.300 164.315 96.560 165.125 ;
        RECT 96.740 164.490 96.990 165.625 ;
        RECT 103.170 165.455 104.335 166.045 ;
        RECT 97.590 165.230 104.335 165.455 ;
        RECT 104.595 165.405 105.345 165.925 ;
        RECT 105.515 165.575 106.265 166.095 ;
        RECT 106.440 166.155 106.695 166.685 ;
        RECT 106.865 166.405 107.170 166.865 ;
        RECT 107.415 166.485 108.485 166.655 ;
        RECT 106.440 165.505 106.650 166.155 ;
        RECT 107.415 166.130 107.735 166.485 ;
        RECT 107.410 165.955 107.735 166.130 ;
        RECT 106.820 165.655 107.735 165.955 ;
        RECT 107.905 165.915 108.145 166.315 ;
        RECT 108.315 166.255 108.485 166.485 ;
        RECT 108.655 166.425 108.845 166.865 ;
        RECT 109.015 166.415 109.965 166.695 ;
        RECT 110.185 166.505 110.535 166.675 ;
        RECT 108.315 166.085 108.845 166.255 ;
        RECT 106.820 165.625 107.560 165.655 ;
        RECT 97.590 165.215 102.995 165.230 ;
        RECT 97.160 164.320 97.420 165.115 ;
        RECT 97.590 164.490 97.850 165.215 ;
        RECT 98.020 164.320 98.280 165.045 ;
        RECT 98.450 164.490 98.710 165.215 ;
        RECT 98.880 164.320 99.140 165.045 ;
        RECT 99.310 164.490 99.570 165.215 ;
        RECT 99.740 164.320 100.000 165.045 ;
        RECT 100.170 164.490 100.430 165.215 ;
        RECT 100.600 164.320 100.845 165.045 ;
        RECT 101.015 164.490 101.275 165.215 ;
        RECT 101.460 164.320 101.705 165.045 ;
        RECT 101.875 164.490 102.135 165.215 ;
        RECT 102.320 164.320 102.565 165.045 ;
        RECT 102.735 164.490 102.995 165.215 ;
        RECT 103.180 164.320 103.435 165.045 ;
        RECT 103.605 164.490 103.895 165.230 ;
        RECT 97.160 164.315 103.435 164.320 ;
        RECT 104.065 164.315 104.335 165.060 ;
        RECT 104.595 164.315 106.265 165.405 ;
        RECT 106.440 164.625 106.695 165.505 ;
        RECT 106.865 164.315 107.170 165.455 ;
        RECT 107.390 165.035 107.560 165.625 ;
        RECT 107.905 165.545 108.445 165.915 ;
        RECT 108.625 165.805 108.845 166.085 ;
        RECT 109.015 165.635 109.185 166.415 ;
        RECT 108.780 165.465 109.185 165.635 ;
        RECT 109.355 165.625 109.705 166.245 ;
        RECT 108.780 165.375 108.950 165.465 ;
        RECT 109.875 165.455 110.085 166.245 ;
        RECT 107.730 165.205 108.950 165.375 ;
        RECT 109.410 165.295 110.085 165.455 ;
        RECT 107.390 164.865 108.190 165.035 ;
        RECT 107.510 164.315 107.840 164.695 ;
        RECT 108.020 164.575 108.190 164.865 ;
        RECT 108.780 164.825 108.950 165.205 ;
        RECT 109.120 165.285 110.085 165.295 ;
        RECT 110.275 166.115 110.535 166.505 ;
        RECT 110.745 166.405 111.075 166.865 ;
        RECT 111.950 166.475 112.805 166.645 ;
        RECT 113.010 166.475 113.505 166.645 ;
        RECT 113.675 166.505 114.005 166.865 ;
        RECT 110.275 165.425 110.445 166.115 ;
        RECT 110.615 165.765 110.785 165.945 ;
        RECT 110.955 165.935 111.745 166.185 ;
        RECT 111.950 165.765 112.120 166.475 ;
        RECT 112.290 165.965 112.645 166.185 ;
        RECT 110.615 165.595 112.305 165.765 ;
        RECT 109.120 164.995 109.580 165.285 ;
        RECT 110.275 165.255 111.775 165.425 ;
        RECT 110.275 165.115 110.445 165.255 ;
        RECT 109.885 164.945 110.445 165.115 ;
        RECT 108.360 164.315 108.610 164.775 ;
        RECT 108.780 164.485 109.650 164.825 ;
        RECT 109.885 164.485 110.055 164.945 ;
        RECT 110.890 164.915 111.965 165.085 ;
        RECT 110.225 164.315 110.595 164.775 ;
        RECT 110.890 164.575 111.060 164.915 ;
        RECT 111.230 164.315 111.560 164.745 ;
        RECT 111.795 164.575 111.965 164.915 ;
        RECT 112.135 164.815 112.305 165.595 ;
        RECT 112.475 165.375 112.645 165.965 ;
        RECT 112.815 165.565 113.165 166.185 ;
        RECT 112.475 164.985 112.940 165.375 ;
        RECT 113.335 165.115 113.505 166.475 ;
        RECT 113.675 165.285 114.135 166.335 ;
        RECT 113.110 164.945 113.505 165.115 ;
        RECT 113.110 164.815 113.280 164.945 ;
        RECT 112.135 164.485 112.815 164.815 ;
        RECT 113.030 164.485 113.280 164.815 ;
        RECT 113.450 164.315 113.700 164.775 ;
        RECT 113.870 164.500 114.195 165.285 ;
        RECT 114.365 164.485 114.535 166.605 ;
        RECT 114.705 166.485 115.035 166.865 ;
        RECT 115.205 166.315 115.460 166.605 ;
        RECT 114.710 166.145 115.460 166.315 ;
        RECT 114.710 165.155 114.940 166.145 ;
        RECT 116.095 166.140 116.385 166.865 ;
        RECT 116.560 166.155 116.815 166.685 ;
        RECT 116.985 166.405 117.290 166.865 ;
        RECT 117.535 166.485 118.605 166.655 ;
        RECT 115.110 165.325 115.460 165.975 ;
        RECT 116.560 165.505 116.770 166.155 ;
        RECT 117.535 166.130 117.855 166.485 ;
        RECT 117.530 165.955 117.855 166.130 ;
        RECT 116.940 165.655 117.855 165.955 ;
        RECT 118.025 165.915 118.265 166.315 ;
        RECT 118.435 166.255 118.605 166.485 ;
        RECT 118.775 166.425 118.965 166.865 ;
        RECT 119.135 166.415 120.085 166.695 ;
        RECT 120.305 166.505 120.655 166.675 ;
        RECT 118.435 166.085 118.965 166.255 ;
        RECT 116.940 165.625 117.680 165.655 ;
        RECT 114.710 164.985 115.460 165.155 ;
        RECT 114.705 164.315 115.035 164.815 ;
        RECT 115.205 164.485 115.460 164.985 ;
        RECT 116.095 164.315 116.385 165.480 ;
        RECT 116.560 164.625 116.815 165.505 ;
        RECT 116.985 164.315 117.290 165.455 ;
        RECT 117.510 165.035 117.680 165.625 ;
        RECT 118.025 165.545 118.565 165.915 ;
        RECT 118.745 165.805 118.965 166.085 ;
        RECT 119.135 165.635 119.305 166.415 ;
        RECT 118.900 165.465 119.305 165.635 ;
        RECT 119.475 165.625 119.825 166.245 ;
        RECT 118.900 165.375 119.070 165.465 ;
        RECT 119.995 165.455 120.205 166.245 ;
        RECT 117.850 165.205 119.070 165.375 ;
        RECT 119.530 165.295 120.205 165.455 ;
        RECT 117.510 164.865 118.310 165.035 ;
        RECT 117.630 164.315 117.960 164.695 ;
        RECT 118.140 164.575 118.310 164.865 ;
        RECT 118.900 164.825 119.070 165.205 ;
        RECT 119.240 165.285 120.205 165.295 ;
        RECT 120.395 166.115 120.655 166.505 ;
        RECT 120.865 166.405 121.195 166.865 ;
        RECT 122.070 166.475 122.925 166.645 ;
        RECT 123.130 166.475 123.625 166.645 ;
        RECT 123.795 166.505 124.125 166.865 ;
        RECT 120.395 165.425 120.565 166.115 ;
        RECT 120.735 165.765 120.905 165.945 ;
        RECT 121.075 165.935 121.865 166.185 ;
        RECT 122.070 165.765 122.240 166.475 ;
        RECT 122.410 165.965 122.765 166.185 ;
        RECT 120.735 165.595 122.425 165.765 ;
        RECT 119.240 164.995 119.700 165.285 ;
        RECT 120.395 165.255 121.895 165.425 ;
        RECT 120.395 165.115 120.565 165.255 ;
        RECT 120.005 164.945 120.565 165.115 ;
        RECT 118.480 164.315 118.730 164.775 ;
        RECT 118.900 164.485 119.770 164.825 ;
        RECT 120.005 164.485 120.175 164.945 ;
        RECT 121.010 164.915 122.085 165.085 ;
        RECT 120.345 164.315 120.715 164.775 ;
        RECT 121.010 164.575 121.180 164.915 ;
        RECT 121.350 164.315 121.680 164.745 ;
        RECT 121.915 164.575 122.085 164.915 ;
        RECT 122.255 164.815 122.425 165.595 ;
        RECT 122.595 165.375 122.765 165.965 ;
        RECT 122.935 165.565 123.285 166.185 ;
        RECT 122.595 164.985 123.060 165.375 ;
        RECT 123.455 165.115 123.625 166.475 ;
        RECT 123.795 165.285 124.255 166.335 ;
        RECT 123.230 164.945 123.625 165.115 ;
        RECT 123.230 164.815 123.400 164.945 ;
        RECT 122.255 164.485 122.935 164.815 ;
        RECT 123.150 164.485 123.400 164.815 ;
        RECT 123.570 164.315 123.820 164.775 ;
        RECT 123.990 164.500 124.315 165.285 ;
        RECT 124.485 164.485 124.655 166.605 ;
        RECT 124.825 166.485 125.155 166.865 ;
        RECT 125.325 166.315 125.580 166.605 ;
        RECT 124.830 166.145 125.580 166.315 ;
        RECT 125.755 166.190 126.015 166.695 ;
        RECT 126.195 166.485 126.525 166.865 ;
        RECT 126.705 166.315 126.875 166.695 ;
        RECT 124.830 165.155 125.060 166.145 ;
        RECT 125.230 165.325 125.580 165.975 ;
        RECT 125.755 165.390 125.925 166.190 ;
        RECT 126.210 166.145 126.875 166.315 ;
        RECT 126.210 165.890 126.380 166.145 ;
        RECT 128.055 166.115 129.265 166.865 ;
        RECT 126.095 165.560 126.380 165.890 ;
        RECT 126.615 165.595 126.945 165.965 ;
        RECT 126.210 165.415 126.380 165.560 ;
        RECT 124.830 164.985 125.580 165.155 ;
        RECT 124.825 164.315 125.155 164.815 ;
        RECT 125.325 164.485 125.580 164.985 ;
        RECT 125.755 164.485 126.025 165.390 ;
        RECT 126.210 165.245 126.875 165.415 ;
        RECT 126.195 164.315 126.525 165.075 ;
        RECT 126.705 164.485 126.875 165.245 ;
        RECT 128.055 165.405 128.575 165.945 ;
        RECT 128.745 165.575 129.265 166.115 ;
        RECT 128.055 164.315 129.265 165.405 ;
        RECT 9.290 164.145 129.350 164.315 ;
        RECT 9.375 163.055 10.585 164.145 ;
        RECT 9.375 162.345 9.895 162.885 ;
        RECT 10.065 162.515 10.585 163.055 ;
        RECT 11.675 163.055 15.185 164.145 ;
        RECT 15.445 163.215 15.615 163.975 ;
        RECT 15.795 163.385 16.125 164.145 ;
        RECT 11.675 162.535 13.365 163.055 ;
        RECT 15.445 163.045 16.110 163.215 ;
        RECT 16.295 163.070 16.565 163.975 ;
        RECT 16.740 163.475 16.995 163.975 ;
        RECT 17.165 163.645 17.495 164.145 ;
        RECT 16.740 163.305 17.490 163.475 ;
        RECT 15.940 162.900 16.110 163.045 ;
        RECT 13.535 162.365 15.185 162.885 ;
        RECT 15.375 162.495 15.705 162.865 ;
        RECT 15.940 162.570 16.225 162.900 ;
        RECT 9.375 161.595 10.585 162.345 ;
        RECT 11.675 161.595 15.185 162.365 ;
        RECT 15.940 162.315 16.110 162.570 ;
        RECT 15.445 162.145 16.110 162.315 ;
        RECT 16.395 162.270 16.565 163.070 ;
        RECT 16.740 162.485 17.090 163.135 ;
        RECT 17.260 162.315 17.490 163.305 ;
        RECT 15.445 161.765 15.615 162.145 ;
        RECT 15.795 161.595 16.125 161.975 ;
        RECT 16.305 161.765 16.565 162.270 ;
        RECT 16.740 162.145 17.490 162.315 ;
        RECT 16.740 161.855 16.995 162.145 ;
        RECT 17.165 161.595 17.495 161.975 ;
        RECT 17.665 161.855 17.835 163.975 ;
        RECT 18.005 163.175 18.330 163.960 ;
        RECT 18.500 163.685 18.750 164.145 ;
        RECT 18.920 163.645 19.170 163.975 ;
        RECT 19.385 163.645 20.065 163.975 ;
        RECT 18.920 163.515 19.090 163.645 ;
        RECT 18.695 163.345 19.090 163.515 ;
        RECT 18.065 162.125 18.525 163.175 ;
        RECT 18.695 161.985 18.865 163.345 ;
        RECT 19.260 163.085 19.725 163.475 ;
        RECT 19.035 162.275 19.385 162.895 ;
        RECT 19.555 162.495 19.725 163.085 ;
        RECT 19.895 162.865 20.065 163.645 ;
        RECT 20.235 163.545 20.405 163.885 ;
        RECT 20.640 163.715 20.970 164.145 ;
        RECT 21.140 163.545 21.310 163.885 ;
        RECT 21.605 163.685 21.975 164.145 ;
        RECT 20.235 163.375 21.310 163.545 ;
        RECT 22.145 163.515 22.315 163.975 ;
        RECT 22.550 163.635 23.420 163.975 ;
        RECT 23.590 163.685 23.840 164.145 ;
        RECT 21.755 163.345 22.315 163.515 ;
        RECT 21.755 163.205 21.925 163.345 ;
        RECT 20.425 163.035 21.925 163.205 ;
        RECT 22.620 163.175 23.080 163.465 ;
        RECT 19.895 162.695 21.585 162.865 ;
        RECT 19.555 162.275 19.910 162.495 ;
        RECT 20.080 161.985 20.250 162.695 ;
        RECT 20.455 162.275 21.245 162.525 ;
        RECT 21.415 162.515 21.585 162.695 ;
        RECT 21.755 162.345 21.925 163.035 ;
        RECT 18.195 161.595 18.525 161.955 ;
        RECT 18.695 161.815 19.190 161.985 ;
        RECT 19.395 161.815 20.250 161.985 ;
        RECT 21.125 161.595 21.455 162.055 ;
        RECT 21.665 161.955 21.925 162.345 ;
        RECT 22.115 163.165 23.080 163.175 ;
        RECT 23.250 163.255 23.420 163.635 ;
        RECT 24.010 163.595 24.180 163.885 ;
        RECT 24.360 163.765 24.690 164.145 ;
        RECT 24.010 163.425 24.810 163.595 ;
        RECT 22.115 163.005 22.790 163.165 ;
        RECT 23.250 163.085 24.470 163.255 ;
        RECT 22.115 162.215 22.325 163.005 ;
        RECT 23.250 162.995 23.420 163.085 ;
        RECT 22.495 162.215 22.845 162.835 ;
        RECT 23.015 162.825 23.420 162.995 ;
        RECT 23.015 162.045 23.185 162.825 ;
        RECT 23.355 162.375 23.575 162.655 ;
        RECT 23.755 162.545 24.295 162.915 ;
        RECT 24.640 162.835 24.810 163.425 ;
        RECT 25.030 163.005 25.335 164.145 ;
        RECT 25.505 162.955 25.760 163.835 ;
        RECT 25.935 162.980 26.225 164.145 ;
        RECT 26.860 163.005 27.195 163.975 ;
        RECT 27.365 163.005 27.535 164.145 ;
        RECT 27.705 163.805 29.735 163.975 ;
        RECT 24.640 162.805 25.380 162.835 ;
        RECT 23.355 162.205 23.885 162.375 ;
        RECT 21.665 161.785 22.015 161.955 ;
        RECT 22.235 161.765 23.185 162.045 ;
        RECT 23.355 161.595 23.545 162.035 ;
        RECT 23.715 161.975 23.885 162.205 ;
        RECT 24.055 162.145 24.295 162.545 ;
        RECT 24.465 162.505 25.380 162.805 ;
        RECT 24.465 162.330 24.790 162.505 ;
        RECT 24.465 161.975 24.785 162.330 ;
        RECT 25.550 162.305 25.760 162.955 ;
        RECT 26.860 162.335 27.030 163.005 ;
        RECT 27.705 162.835 27.875 163.805 ;
        RECT 27.200 162.505 27.455 162.835 ;
        RECT 27.680 162.505 27.875 162.835 ;
        RECT 28.045 163.465 29.170 163.635 ;
        RECT 27.285 162.335 27.455 162.505 ;
        RECT 28.045 162.335 28.215 163.465 ;
        RECT 23.715 161.805 24.785 161.975 ;
        RECT 25.030 161.595 25.335 162.055 ;
        RECT 25.505 161.775 25.760 162.305 ;
        RECT 25.935 161.595 26.225 162.320 ;
        RECT 26.860 161.765 27.115 162.335 ;
        RECT 27.285 162.165 28.215 162.335 ;
        RECT 28.385 163.125 29.395 163.295 ;
        RECT 28.385 162.325 28.555 163.125 ;
        RECT 28.040 162.130 28.215 162.165 ;
        RECT 27.285 161.595 27.615 161.995 ;
        RECT 28.040 161.765 28.570 162.130 ;
        RECT 28.760 162.105 29.035 162.925 ;
        RECT 28.755 161.935 29.035 162.105 ;
        RECT 28.760 161.765 29.035 161.935 ;
        RECT 29.205 161.765 29.395 163.125 ;
        RECT 29.565 163.140 29.735 163.805 ;
        RECT 29.905 163.385 30.075 164.145 ;
        RECT 30.310 163.385 30.825 163.795 ;
        RECT 29.565 162.950 30.315 163.140 ;
        RECT 30.485 162.575 30.825 163.385 ;
        RECT 32.005 163.215 32.175 163.975 ;
        RECT 32.355 163.385 32.685 164.145 ;
        RECT 32.005 163.045 32.670 163.215 ;
        RECT 32.855 163.070 33.125 163.975 ;
        RECT 33.300 163.475 33.555 163.975 ;
        RECT 33.725 163.645 34.055 164.145 ;
        RECT 33.300 163.305 34.050 163.475 ;
        RECT 32.500 162.900 32.670 163.045 ;
        RECT 29.595 162.405 30.825 162.575 ;
        RECT 31.935 162.495 32.265 162.865 ;
        RECT 32.500 162.570 32.785 162.900 ;
        RECT 29.575 161.595 30.085 162.130 ;
        RECT 30.305 161.800 30.550 162.405 ;
        RECT 32.500 162.315 32.670 162.570 ;
        RECT 32.005 162.145 32.670 162.315 ;
        RECT 32.955 162.270 33.125 163.070 ;
        RECT 33.300 162.485 33.650 163.135 ;
        RECT 33.820 162.315 34.050 163.305 ;
        RECT 32.005 161.765 32.175 162.145 ;
        RECT 32.355 161.595 32.685 161.975 ;
        RECT 32.865 161.765 33.125 162.270 ;
        RECT 33.300 162.145 34.050 162.315 ;
        RECT 33.300 161.855 33.555 162.145 ;
        RECT 33.725 161.595 34.055 161.975 ;
        RECT 34.225 161.855 34.395 163.975 ;
        RECT 34.565 163.175 34.890 163.960 ;
        RECT 35.060 163.685 35.310 164.145 ;
        RECT 35.480 163.645 35.730 163.975 ;
        RECT 35.945 163.645 36.625 163.975 ;
        RECT 35.480 163.515 35.650 163.645 ;
        RECT 35.255 163.345 35.650 163.515 ;
        RECT 34.625 162.125 35.085 163.175 ;
        RECT 35.255 161.985 35.425 163.345 ;
        RECT 35.820 163.085 36.285 163.475 ;
        RECT 35.595 162.275 35.945 162.895 ;
        RECT 36.115 162.495 36.285 163.085 ;
        RECT 36.455 162.865 36.625 163.645 ;
        RECT 36.795 163.545 36.965 163.885 ;
        RECT 37.200 163.715 37.530 164.145 ;
        RECT 37.700 163.545 37.870 163.885 ;
        RECT 38.165 163.685 38.535 164.145 ;
        RECT 36.795 163.375 37.870 163.545 ;
        RECT 38.705 163.515 38.875 163.975 ;
        RECT 39.110 163.635 39.980 163.975 ;
        RECT 40.150 163.685 40.400 164.145 ;
        RECT 38.315 163.345 38.875 163.515 ;
        RECT 38.315 163.205 38.485 163.345 ;
        RECT 36.985 163.035 38.485 163.205 ;
        RECT 39.180 163.175 39.640 163.465 ;
        RECT 36.455 162.695 38.145 162.865 ;
        RECT 36.115 162.275 36.470 162.495 ;
        RECT 36.640 161.985 36.810 162.695 ;
        RECT 37.015 162.275 37.805 162.525 ;
        RECT 37.975 162.515 38.145 162.695 ;
        RECT 38.315 162.345 38.485 163.035 ;
        RECT 34.755 161.595 35.085 161.955 ;
        RECT 35.255 161.815 35.750 161.985 ;
        RECT 35.955 161.815 36.810 161.985 ;
        RECT 37.685 161.595 38.015 162.055 ;
        RECT 38.225 161.955 38.485 162.345 ;
        RECT 38.675 163.165 39.640 163.175 ;
        RECT 39.810 163.255 39.980 163.635 ;
        RECT 40.570 163.595 40.740 163.885 ;
        RECT 40.920 163.765 41.250 164.145 ;
        RECT 40.570 163.425 41.370 163.595 ;
        RECT 38.675 163.005 39.350 163.165 ;
        RECT 39.810 163.085 41.030 163.255 ;
        RECT 38.675 162.215 38.885 163.005 ;
        RECT 39.810 162.995 39.980 163.085 ;
        RECT 39.055 162.215 39.405 162.835 ;
        RECT 39.575 162.825 39.980 162.995 ;
        RECT 39.575 162.045 39.745 162.825 ;
        RECT 39.915 162.375 40.135 162.655 ;
        RECT 40.315 162.545 40.855 162.915 ;
        RECT 41.200 162.835 41.370 163.425 ;
        RECT 41.590 163.005 41.895 164.145 ;
        RECT 42.065 162.955 42.320 163.835 ;
        RECT 41.200 162.805 41.940 162.835 ;
        RECT 39.915 162.205 40.445 162.375 ;
        RECT 38.225 161.785 38.575 161.955 ;
        RECT 38.795 161.765 39.745 162.045 ;
        RECT 39.915 161.595 40.105 162.035 ;
        RECT 40.275 161.975 40.445 162.205 ;
        RECT 40.615 162.145 40.855 162.545 ;
        RECT 41.025 162.505 41.940 162.805 ;
        RECT 41.025 162.330 41.350 162.505 ;
        RECT 41.025 161.975 41.345 162.330 ;
        RECT 42.110 162.305 42.320 162.955 ;
        RECT 40.275 161.805 41.345 161.975 ;
        RECT 41.590 161.595 41.895 162.055 ;
        RECT 42.065 161.775 42.320 162.305 ;
        RECT 42.500 162.955 42.755 163.835 ;
        RECT 42.925 163.005 43.230 164.145 ;
        RECT 43.570 163.765 43.900 164.145 ;
        RECT 44.080 163.595 44.250 163.885 ;
        RECT 44.420 163.685 44.670 164.145 ;
        RECT 43.450 163.425 44.250 163.595 ;
        RECT 44.840 163.635 45.710 163.975 ;
        RECT 42.500 162.305 42.710 162.955 ;
        RECT 43.450 162.835 43.620 163.425 ;
        RECT 44.840 163.255 45.010 163.635 ;
        RECT 45.945 163.515 46.115 163.975 ;
        RECT 46.285 163.685 46.655 164.145 ;
        RECT 46.950 163.545 47.120 163.885 ;
        RECT 47.290 163.715 47.620 164.145 ;
        RECT 47.855 163.545 48.025 163.885 ;
        RECT 43.790 163.085 45.010 163.255 ;
        RECT 45.180 163.175 45.640 163.465 ;
        RECT 45.945 163.345 46.505 163.515 ;
        RECT 46.950 163.375 48.025 163.545 ;
        RECT 48.195 163.645 48.875 163.975 ;
        RECT 49.090 163.645 49.340 163.975 ;
        RECT 49.510 163.685 49.760 164.145 ;
        RECT 46.335 163.205 46.505 163.345 ;
        RECT 45.180 163.165 46.145 163.175 ;
        RECT 44.840 162.995 45.010 163.085 ;
        RECT 45.470 163.005 46.145 163.165 ;
        RECT 42.880 162.805 43.620 162.835 ;
        RECT 42.880 162.505 43.795 162.805 ;
        RECT 43.470 162.330 43.795 162.505 ;
        RECT 42.500 161.775 42.755 162.305 ;
        RECT 42.925 161.595 43.230 162.055 ;
        RECT 43.475 161.975 43.795 162.330 ;
        RECT 43.965 162.545 44.505 162.915 ;
        RECT 44.840 162.825 45.245 162.995 ;
        RECT 43.965 162.145 44.205 162.545 ;
        RECT 44.685 162.375 44.905 162.655 ;
        RECT 44.375 162.205 44.905 162.375 ;
        RECT 44.375 161.975 44.545 162.205 ;
        RECT 45.075 162.045 45.245 162.825 ;
        RECT 45.415 162.215 45.765 162.835 ;
        RECT 45.935 162.215 46.145 163.005 ;
        RECT 46.335 163.035 47.835 163.205 ;
        RECT 46.335 162.345 46.505 163.035 ;
        RECT 48.195 162.865 48.365 163.645 ;
        RECT 49.170 163.515 49.340 163.645 ;
        RECT 46.675 162.695 48.365 162.865 ;
        RECT 48.535 163.085 49.000 163.475 ;
        RECT 49.170 163.345 49.565 163.515 ;
        RECT 46.675 162.515 46.845 162.695 ;
        RECT 43.475 161.805 44.545 161.975 ;
        RECT 44.715 161.595 44.905 162.035 ;
        RECT 45.075 161.765 46.025 162.045 ;
        RECT 46.335 161.955 46.595 162.345 ;
        RECT 47.015 162.275 47.805 162.525 ;
        RECT 46.245 161.785 46.595 161.955 ;
        RECT 46.805 161.595 47.135 162.055 ;
        RECT 48.010 161.985 48.180 162.695 ;
        RECT 48.535 162.495 48.705 163.085 ;
        RECT 48.350 162.275 48.705 162.495 ;
        RECT 48.875 162.275 49.225 162.895 ;
        RECT 49.395 161.985 49.565 163.345 ;
        RECT 49.930 163.175 50.255 163.960 ;
        RECT 49.735 162.125 50.195 163.175 ;
        RECT 48.010 161.815 48.865 161.985 ;
        RECT 49.070 161.815 49.565 161.985 ;
        RECT 49.735 161.595 50.065 161.955 ;
        RECT 50.425 161.855 50.595 163.975 ;
        RECT 50.765 163.645 51.095 164.145 ;
        RECT 51.265 163.475 51.520 163.975 ;
        RECT 50.770 163.305 51.520 163.475 ;
        RECT 50.770 162.315 51.000 163.305 ;
        RECT 51.170 162.485 51.520 163.135 ;
        RECT 51.695 162.980 51.985 164.145 ;
        RECT 52.155 163.055 54.745 164.145 ;
        RECT 54.920 163.710 60.265 164.145 ;
        RECT 52.155 162.535 53.365 163.055 ;
        RECT 53.535 162.365 54.745 162.885 ;
        RECT 56.510 162.460 56.860 163.710 ;
        RECT 60.585 162.995 60.915 164.145 ;
        RECT 61.085 163.125 61.255 163.975 ;
        RECT 61.425 163.345 61.755 164.145 ;
        RECT 61.925 163.125 62.095 163.975 ;
        RECT 62.275 163.345 62.515 164.145 ;
        RECT 62.685 163.165 63.015 163.975 ;
        RECT 63.660 163.710 69.005 164.145 ;
        RECT 50.770 162.145 51.520 162.315 ;
        RECT 50.765 161.595 51.095 161.975 ;
        RECT 51.265 161.855 51.520 162.145 ;
        RECT 51.695 161.595 51.985 162.320 ;
        RECT 52.155 161.595 54.745 162.365 ;
        RECT 58.340 162.140 58.680 162.970 ;
        RECT 61.085 162.955 62.095 163.125 ;
        RECT 62.300 162.995 63.015 163.165 ;
        RECT 61.085 162.415 61.580 162.955 ;
        RECT 62.300 162.755 62.470 162.995 ;
        RECT 61.970 162.585 62.470 162.755 ;
        RECT 62.640 162.585 63.020 162.825 ;
        RECT 62.300 162.415 62.470 162.585 ;
        RECT 65.250 162.460 65.600 163.710 ;
        RECT 69.185 163.085 69.515 164.145 ;
        RECT 54.920 161.595 60.265 162.140 ;
        RECT 60.585 161.595 60.915 162.395 ;
        RECT 61.085 162.245 62.095 162.415 ;
        RECT 62.300 162.245 62.935 162.415 ;
        RECT 61.085 161.765 61.255 162.245 ;
        RECT 61.425 161.595 61.755 162.075 ;
        RECT 61.925 161.765 62.095 162.245 ;
        RECT 62.345 161.595 62.585 162.075 ;
        RECT 62.765 161.765 62.935 162.245 ;
        RECT 67.080 162.140 67.420 162.970 ;
        RECT 69.695 162.835 69.865 163.805 ;
        RECT 70.035 163.555 70.365 163.955 ;
        RECT 70.535 163.785 70.865 164.145 ;
        RECT 71.065 163.555 71.765 163.975 ;
        RECT 70.035 163.325 71.765 163.555 ;
        RECT 70.035 163.105 70.365 163.325 ;
        RECT 70.560 162.835 70.885 163.125 ;
        RECT 69.175 162.505 69.485 162.835 ;
        RECT 69.695 162.505 70.070 162.835 ;
        RECT 70.390 162.505 70.885 162.835 ;
        RECT 71.060 162.585 71.390 163.125 ;
        RECT 71.560 162.355 71.765 163.325 ;
        RECT 63.660 161.595 69.005 162.140 ;
        RECT 69.185 162.125 70.545 162.335 ;
        RECT 69.185 161.765 69.515 162.125 ;
        RECT 69.685 161.595 70.015 161.955 ;
        RECT 70.215 161.765 70.545 162.125 ;
        RECT 71.055 161.765 71.765 162.355 ;
        RECT 71.935 163.175 72.245 163.975 ;
        RECT 72.415 163.345 72.725 164.145 ;
        RECT 72.895 163.515 73.155 163.975 ;
        RECT 73.325 163.685 73.580 164.145 ;
        RECT 73.755 163.515 74.015 163.975 ;
        RECT 72.895 163.345 74.015 163.515 ;
        RECT 71.935 163.005 72.965 163.175 ;
        RECT 71.935 162.095 72.105 163.005 ;
        RECT 72.275 162.265 72.625 162.835 ;
        RECT 72.795 162.755 72.965 163.005 ;
        RECT 73.755 163.095 74.015 163.345 ;
        RECT 74.185 163.275 74.470 164.145 ;
        RECT 73.755 162.925 74.510 163.095 ;
        RECT 72.795 162.585 73.935 162.755 ;
        RECT 74.105 162.415 74.510 162.925 ;
        RECT 74.695 163.055 75.905 164.145 ;
        RECT 74.695 162.515 75.215 163.055 ;
        RECT 76.135 163.005 76.345 164.145 ;
        RECT 76.515 162.995 76.845 163.975 ;
        RECT 77.015 163.005 77.245 164.145 ;
        RECT 72.860 162.245 74.510 162.415 ;
        RECT 75.385 162.345 75.905 162.885 ;
        RECT 71.935 161.765 72.235 162.095 ;
        RECT 72.405 161.595 72.680 162.075 ;
        RECT 72.860 161.855 73.155 162.245 ;
        RECT 73.325 161.595 73.580 162.075 ;
        RECT 73.755 161.855 74.015 162.245 ;
        RECT 74.185 161.595 74.465 162.075 ;
        RECT 74.695 161.595 75.905 162.345 ;
        RECT 76.135 161.595 76.345 162.415 ;
        RECT 76.515 162.395 76.765 162.995 ;
        RECT 77.455 162.980 77.745 164.145 ;
        RECT 78.290 163.165 78.545 163.835 ;
        RECT 78.725 163.345 79.010 164.145 ;
        RECT 79.190 163.425 79.520 163.935 ;
        RECT 76.935 162.585 77.265 162.835 ;
        RECT 76.515 161.765 76.845 162.395 ;
        RECT 77.015 161.595 77.245 162.415 ;
        RECT 77.455 161.595 77.745 162.320 ;
        RECT 78.290 162.305 78.470 163.165 ;
        RECT 79.190 162.835 79.440 163.425 ;
        RECT 79.790 163.275 79.960 163.885 ;
        RECT 80.130 163.455 80.460 164.145 ;
        RECT 80.690 163.595 80.930 163.885 ;
        RECT 81.130 163.765 81.550 164.145 ;
        RECT 81.730 163.675 82.360 163.925 ;
        RECT 82.830 163.765 83.160 164.145 ;
        RECT 81.730 163.595 81.900 163.675 ;
        RECT 83.330 163.595 83.500 163.885 ;
        RECT 83.680 163.765 84.060 164.145 ;
        RECT 84.300 163.760 85.130 163.930 ;
        RECT 80.690 163.425 81.900 163.595 ;
        RECT 78.640 162.505 79.440 162.835 ;
        RECT 78.290 162.105 78.545 162.305 ;
        RECT 78.205 161.935 78.545 162.105 ;
        RECT 78.290 161.775 78.545 161.935 ;
        RECT 78.725 161.595 79.010 162.055 ;
        RECT 79.190 161.855 79.440 162.505 ;
        RECT 79.640 163.255 79.960 163.275 ;
        RECT 79.640 163.085 81.560 163.255 ;
        RECT 79.640 162.190 79.830 163.085 ;
        RECT 81.730 162.915 81.900 163.425 ;
        RECT 82.070 163.165 82.590 163.475 ;
        RECT 80.000 162.745 81.900 162.915 ;
        RECT 80.000 162.685 80.330 162.745 ;
        RECT 80.480 162.515 80.810 162.575 ;
        RECT 80.150 162.245 80.810 162.515 ;
        RECT 79.640 161.860 79.960 162.190 ;
        RECT 80.140 161.595 80.800 162.075 ;
        RECT 81.000 161.985 81.170 162.745 ;
        RECT 82.070 162.575 82.250 162.985 ;
        RECT 81.340 162.405 81.670 162.525 ;
        RECT 82.420 162.405 82.590 163.165 ;
        RECT 81.340 162.235 82.590 162.405 ;
        RECT 82.760 163.345 84.130 163.595 ;
        RECT 82.760 162.575 82.950 163.345 ;
        RECT 83.880 163.085 84.130 163.345 ;
        RECT 83.120 162.915 83.370 163.075 ;
        RECT 84.300 162.915 84.470 163.760 ;
        RECT 85.365 163.475 85.535 163.975 ;
        RECT 85.705 163.645 86.035 164.145 ;
        RECT 84.640 163.085 85.140 163.465 ;
        RECT 85.365 163.305 86.060 163.475 ;
        RECT 83.120 162.745 84.470 162.915 ;
        RECT 84.050 162.705 84.470 162.745 ;
        RECT 82.760 162.235 83.180 162.575 ;
        RECT 83.470 162.245 83.880 162.575 ;
        RECT 81.000 161.815 81.850 161.985 ;
        RECT 82.410 161.595 82.730 162.055 ;
        RECT 82.930 161.805 83.180 162.235 ;
        RECT 83.470 161.595 83.880 162.035 ;
        RECT 84.050 161.975 84.220 162.705 ;
        RECT 84.390 162.155 84.740 162.525 ;
        RECT 84.920 162.215 85.140 163.085 ;
        RECT 85.310 162.515 85.720 163.135 ;
        RECT 85.890 162.335 86.060 163.305 ;
        RECT 85.365 162.145 86.060 162.335 ;
        RECT 84.050 161.775 85.065 161.975 ;
        RECT 85.365 161.815 85.535 162.145 ;
        RECT 85.705 161.595 86.035 161.975 ;
        RECT 86.250 161.855 86.475 163.975 ;
        RECT 86.645 163.645 86.975 164.145 ;
        RECT 87.145 163.475 87.315 163.975 ;
        RECT 86.650 163.305 87.315 163.475 ;
        RECT 87.665 163.400 87.935 164.145 ;
        RECT 88.565 164.140 94.840 164.145 ;
        RECT 86.650 162.315 86.880 163.305 ;
        RECT 88.105 163.230 88.395 163.970 ;
        RECT 88.565 163.415 88.820 164.140 ;
        RECT 89.005 163.245 89.265 163.970 ;
        RECT 89.435 163.415 89.680 164.140 ;
        RECT 89.865 163.245 90.125 163.970 ;
        RECT 90.295 163.415 90.540 164.140 ;
        RECT 90.725 163.245 90.985 163.970 ;
        RECT 91.155 163.415 91.400 164.140 ;
        RECT 91.570 163.245 91.830 163.970 ;
        RECT 92.000 163.415 92.260 164.140 ;
        RECT 92.430 163.245 92.690 163.970 ;
        RECT 92.860 163.415 93.120 164.140 ;
        RECT 93.290 163.245 93.550 163.970 ;
        RECT 93.720 163.415 93.980 164.140 ;
        RECT 94.150 163.245 94.410 163.970 ;
        RECT 94.580 163.345 94.840 164.140 ;
        RECT 89.005 163.230 94.410 163.245 ;
        RECT 87.050 162.485 87.400 163.135 ;
        RECT 87.665 163.005 94.410 163.230 ;
        RECT 87.665 162.415 88.830 163.005 ;
        RECT 95.010 162.835 95.260 163.970 ;
        RECT 95.440 163.335 95.700 164.145 ;
        RECT 95.875 162.835 96.120 163.975 ;
        RECT 96.300 163.335 96.595 164.145 ;
        RECT 97.235 163.055 98.905 164.145 ;
        RECT 99.075 163.385 99.590 163.795 ;
        RECT 99.825 163.385 99.995 164.145 ;
        RECT 100.165 163.805 102.195 163.975 ;
        RECT 89.000 162.585 96.120 162.835 ;
        RECT 86.650 162.145 87.315 162.315 ;
        RECT 87.665 162.245 94.410 162.415 ;
        RECT 86.645 161.595 86.975 161.975 ;
        RECT 87.145 161.855 87.315 162.145 ;
        RECT 87.665 161.595 87.965 162.075 ;
        RECT 88.135 161.790 88.395 162.245 ;
        RECT 88.565 161.595 88.825 162.075 ;
        RECT 89.005 161.790 89.265 162.245 ;
        RECT 89.435 161.595 89.685 162.075 ;
        RECT 89.865 161.790 90.125 162.245 ;
        RECT 90.295 161.595 90.545 162.075 ;
        RECT 90.725 161.790 90.985 162.245 ;
        RECT 91.155 161.595 91.400 162.075 ;
        RECT 91.570 161.790 91.845 162.245 ;
        RECT 92.015 161.595 92.260 162.075 ;
        RECT 92.430 161.790 92.690 162.245 ;
        RECT 92.860 161.595 93.120 162.075 ;
        RECT 93.290 161.790 93.550 162.245 ;
        RECT 93.720 161.595 93.980 162.075 ;
        RECT 94.150 161.790 94.410 162.245 ;
        RECT 94.580 161.595 94.840 162.155 ;
        RECT 95.010 161.775 95.260 162.585 ;
        RECT 95.440 161.595 95.700 162.120 ;
        RECT 95.870 161.775 96.120 162.585 ;
        RECT 96.290 162.275 96.605 162.835 ;
        RECT 97.235 162.535 97.985 163.055 ;
        RECT 98.155 162.365 98.905 162.885 ;
        RECT 99.075 162.575 99.415 163.385 ;
        RECT 100.165 163.140 100.335 163.805 ;
        RECT 100.730 163.465 101.855 163.635 ;
        RECT 99.585 162.950 100.335 163.140 ;
        RECT 100.505 163.125 101.515 163.295 ;
        RECT 99.075 162.405 100.305 162.575 ;
        RECT 96.300 161.595 96.605 162.105 ;
        RECT 97.235 161.595 98.905 162.365 ;
        RECT 99.350 161.800 99.595 162.405 ;
        RECT 99.815 161.595 100.325 162.130 ;
        RECT 100.505 161.765 100.695 163.125 ;
        RECT 100.865 162.105 101.140 162.925 ;
        RECT 101.345 162.325 101.515 163.125 ;
        RECT 101.685 162.335 101.855 163.465 ;
        RECT 102.025 162.835 102.195 163.805 ;
        RECT 102.365 163.005 102.535 164.145 ;
        RECT 102.705 163.005 103.040 163.975 ;
        RECT 102.025 162.505 102.220 162.835 ;
        RECT 102.445 162.505 102.700 162.835 ;
        RECT 102.445 162.335 102.615 162.505 ;
        RECT 102.870 162.335 103.040 163.005 ;
        RECT 103.215 162.980 103.505 164.145 ;
        RECT 104.685 163.215 104.855 163.975 ;
        RECT 105.035 163.385 105.365 164.145 ;
        RECT 104.685 163.045 105.350 163.215 ;
        RECT 105.535 163.070 105.805 163.975 ;
        RECT 105.180 162.900 105.350 163.045 ;
        RECT 104.615 162.495 104.945 162.865 ;
        RECT 105.180 162.570 105.465 162.900 ;
        RECT 101.685 162.165 102.615 162.335 ;
        RECT 101.685 162.130 101.860 162.165 ;
        RECT 100.865 161.935 101.145 162.105 ;
        RECT 100.865 161.765 101.140 161.935 ;
        RECT 101.330 161.765 101.860 162.130 ;
        RECT 102.285 161.595 102.615 161.995 ;
        RECT 102.785 161.765 103.040 162.335 ;
        RECT 103.215 161.595 103.505 162.320 ;
        RECT 105.180 162.315 105.350 162.570 ;
        RECT 104.685 162.145 105.350 162.315 ;
        RECT 105.635 162.270 105.805 163.070 ;
        RECT 106.065 163.215 106.235 163.975 ;
        RECT 106.415 163.385 106.745 164.145 ;
        RECT 106.065 163.045 106.730 163.215 ;
        RECT 106.915 163.070 107.185 163.975 ;
        RECT 106.560 162.900 106.730 163.045 ;
        RECT 105.995 162.495 106.325 162.865 ;
        RECT 106.560 162.570 106.845 162.900 ;
        RECT 106.560 162.315 106.730 162.570 ;
        RECT 104.685 161.765 104.855 162.145 ;
        RECT 105.035 161.595 105.365 161.975 ;
        RECT 105.545 161.765 105.805 162.270 ;
        RECT 106.065 162.145 106.730 162.315 ;
        RECT 107.015 162.270 107.185 163.070 ;
        RECT 107.815 163.055 109.485 164.145 ;
        RECT 109.655 163.385 110.170 163.795 ;
        RECT 110.405 163.385 110.575 164.145 ;
        RECT 110.745 163.805 112.775 163.975 ;
        RECT 107.815 162.535 108.565 163.055 ;
        RECT 108.735 162.365 109.485 162.885 ;
        RECT 109.655 162.575 109.995 163.385 ;
        RECT 110.745 163.140 110.915 163.805 ;
        RECT 111.310 163.465 112.435 163.635 ;
        RECT 110.165 162.950 110.915 163.140 ;
        RECT 111.085 163.125 112.095 163.295 ;
        RECT 109.655 162.405 110.885 162.575 ;
        RECT 106.065 161.765 106.235 162.145 ;
        RECT 106.415 161.595 106.745 161.975 ;
        RECT 106.925 161.765 107.185 162.270 ;
        RECT 107.815 161.595 109.485 162.365 ;
        RECT 109.930 161.800 110.175 162.405 ;
        RECT 110.395 161.595 110.905 162.130 ;
        RECT 111.085 161.765 111.275 163.125 ;
        RECT 111.445 162.105 111.720 162.925 ;
        RECT 111.925 162.325 112.095 163.125 ;
        RECT 112.265 162.335 112.435 163.465 ;
        RECT 112.605 162.835 112.775 163.805 ;
        RECT 112.945 163.005 113.115 164.145 ;
        RECT 113.285 163.005 113.620 163.975 ;
        RECT 112.605 162.505 112.800 162.835 ;
        RECT 113.025 162.505 113.280 162.835 ;
        RECT 113.025 162.335 113.195 162.505 ;
        RECT 113.450 162.335 113.620 163.005 ;
        RECT 112.265 162.165 113.195 162.335 ;
        RECT 112.265 162.130 112.440 162.165 ;
        RECT 111.445 161.935 111.725 162.105 ;
        RECT 111.445 161.765 111.720 161.935 ;
        RECT 111.910 161.765 112.440 162.130 ;
        RECT 112.865 161.595 113.195 161.995 ;
        RECT 113.365 161.765 113.620 162.335 ;
        RECT 113.795 163.070 114.065 163.975 ;
        RECT 114.235 163.385 114.565 164.145 ;
        RECT 114.745 163.215 114.915 163.975 ;
        RECT 113.795 162.270 113.965 163.070 ;
        RECT 114.250 163.045 114.915 163.215 ;
        RECT 115.175 163.385 115.690 163.795 ;
        RECT 115.925 163.385 116.095 164.145 ;
        RECT 116.265 163.805 118.295 163.975 ;
        RECT 114.250 162.900 114.420 163.045 ;
        RECT 114.135 162.570 114.420 162.900 ;
        RECT 114.250 162.315 114.420 162.570 ;
        RECT 114.655 162.495 114.985 162.865 ;
        RECT 115.175 162.575 115.515 163.385 ;
        RECT 116.265 163.140 116.435 163.805 ;
        RECT 116.830 163.465 117.955 163.635 ;
        RECT 115.685 162.950 116.435 163.140 ;
        RECT 116.605 163.125 117.615 163.295 ;
        RECT 115.175 162.405 116.405 162.575 ;
        RECT 113.795 161.765 114.055 162.270 ;
        RECT 114.250 162.145 114.915 162.315 ;
        RECT 114.235 161.595 114.565 161.975 ;
        RECT 114.745 161.765 114.915 162.145 ;
        RECT 115.450 161.800 115.695 162.405 ;
        RECT 115.915 161.595 116.425 162.130 ;
        RECT 116.605 161.765 116.795 163.125 ;
        RECT 116.965 162.105 117.240 162.925 ;
        RECT 117.445 162.325 117.615 163.125 ;
        RECT 117.785 162.335 117.955 163.465 ;
        RECT 118.125 162.835 118.295 163.805 ;
        RECT 118.465 163.005 118.635 164.145 ;
        RECT 118.805 163.005 119.140 163.975 ;
        RECT 118.125 162.505 118.320 162.835 ;
        RECT 118.545 162.505 118.800 162.835 ;
        RECT 118.545 162.335 118.715 162.505 ;
        RECT 118.970 162.335 119.140 163.005 ;
        RECT 119.315 163.055 120.985 164.145 ;
        RECT 121.245 163.215 121.415 163.975 ;
        RECT 121.595 163.385 121.925 164.145 ;
        RECT 119.315 162.535 120.065 163.055 ;
        RECT 121.245 163.045 121.910 163.215 ;
        RECT 122.095 163.070 122.365 163.975 ;
        RECT 122.540 163.710 127.885 164.145 ;
        RECT 121.740 162.900 121.910 163.045 ;
        RECT 120.235 162.365 120.985 162.885 ;
        RECT 121.175 162.495 121.505 162.865 ;
        RECT 121.740 162.570 122.025 162.900 ;
        RECT 117.785 162.165 118.715 162.335 ;
        RECT 117.785 162.130 117.960 162.165 ;
        RECT 116.965 161.935 117.245 162.105 ;
        RECT 116.965 161.765 117.240 161.935 ;
        RECT 117.430 161.765 117.960 162.130 ;
        RECT 118.385 161.595 118.715 161.995 ;
        RECT 118.885 161.765 119.140 162.335 ;
        RECT 119.315 161.595 120.985 162.365 ;
        RECT 121.740 162.315 121.910 162.570 ;
        RECT 121.245 162.145 121.910 162.315 ;
        RECT 122.195 162.270 122.365 163.070 ;
        RECT 124.130 162.460 124.480 163.710 ;
        RECT 128.055 163.055 129.265 164.145 ;
        RECT 121.245 161.765 121.415 162.145 ;
        RECT 121.595 161.595 121.925 161.975 ;
        RECT 122.105 161.765 122.365 162.270 ;
        RECT 125.960 162.140 126.300 162.970 ;
        RECT 128.055 162.515 128.575 163.055 ;
        RECT 128.745 162.345 129.265 162.885 ;
        RECT 122.540 161.595 127.885 162.140 ;
        RECT 128.055 161.595 129.265 162.345 ;
        RECT 9.290 161.425 129.350 161.595 ;
        RECT 9.375 160.675 10.585 161.425 ;
        RECT 9.375 160.135 9.895 160.675 ;
        RECT 11.215 160.655 12.885 161.425 ;
        RECT 13.055 160.700 13.345 161.425 ;
        RECT 13.975 160.655 17.485 161.425 ;
        RECT 10.065 159.965 10.585 160.505 ;
        RECT 9.375 158.875 10.585 159.965 ;
        RECT 11.215 159.965 11.965 160.485 ;
        RECT 12.135 160.135 12.885 160.655 ;
        RECT 11.215 158.875 12.885 159.965 ;
        RECT 13.055 158.875 13.345 160.040 ;
        RECT 13.975 159.965 15.665 160.485 ;
        RECT 15.835 160.135 17.485 160.655 ;
        RECT 17.715 160.605 17.925 161.425 ;
        RECT 18.095 160.625 18.425 161.255 ;
        RECT 18.095 160.025 18.345 160.625 ;
        RECT 18.595 160.605 18.825 161.425 ;
        RECT 19.040 160.685 19.295 161.255 ;
        RECT 19.465 161.025 19.795 161.425 ;
        RECT 20.220 160.890 20.750 161.255 ;
        RECT 20.220 160.855 20.395 160.890 ;
        RECT 19.465 160.685 20.395 160.855 ;
        RECT 20.940 160.745 21.215 161.255 ;
        RECT 18.515 160.185 18.845 160.435 ;
        RECT 13.975 158.875 17.485 159.965 ;
        RECT 17.715 158.875 17.925 160.015 ;
        RECT 18.095 159.045 18.425 160.025 ;
        RECT 19.040 160.015 19.210 160.685 ;
        RECT 19.465 160.515 19.635 160.685 ;
        RECT 19.380 160.185 19.635 160.515 ;
        RECT 19.860 160.185 20.055 160.515 ;
        RECT 18.595 158.875 18.825 160.015 ;
        RECT 19.040 159.045 19.375 160.015 ;
        RECT 19.545 158.875 19.715 160.015 ;
        RECT 19.885 159.215 20.055 160.185 ;
        RECT 20.225 159.555 20.395 160.685 ;
        RECT 20.565 159.895 20.735 160.695 ;
        RECT 20.935 160.575 21.215 160.745 ;
        RECT 20.940 160.095 21.215 160.575 ;
        RECT 21.385 159.895 21.575 161.255 ;
        RECT 21.755 160.890 22.265 161.425 ;
        RECT 22.485 160.615 22.730 161.220 ;
        RECT 23.635 160.655 26.225 161.425 ;
        RECT 21.775 160.445 23.005 160.615 ;
        RECT 20.565 159.725 21.575 159.895 ;
        RECT 21.745 159.880 22.495 160.070 ;
        RECT 20.225 159.385 21.350 159.555 ;
        RECT 21.745 159.215 21.915 159.880 ;
        RECT 22.665 159.635 23.005 160.445 ;
        RECT 19.885 159.045 21.915 159.215 ;
        RECT 22.085 158.875 22.255 159.635 ;
        RECT 22.490 159.225 23.005 159.635 ;
        RECT 23.635 159.965 24.845 160.485 ;
        RECT 25.015 160.135 26.225 160.655 ;
        RECT 26.395 160.750 26.655 161.255 ;
        RECT 26.835 161.045 27.165 161.425 ;
        RECT 27.345 160.875 27.515 161.255 ;
        RECT 27.865 160.945 28.165 161.425 ;
        RECT 23.635 158.875 26.225 159.965 ;
        RECT 26.395 159.950 26.565 160.750 ;
        RECT 26.850 160.705 27.515 160.875 ;
        RECT 28.335 160.775 28.595 161.230 ;
        RECT 28.765 160.945 29.025 161.425 ;
        RECT 29.205 160.775 29.465 161.230 ;
        RECT 29.635 160.945 29.885 161.425 ;
        RECT 30.065 160.775 30.325 161.230 ;
        RECT 30.495 160.945 30.745 161.425 ;
        RECT 30.925 160.775 31.185 161.230 ;
        RECT 31.355 160.945 31.600 161.425 ;
        RECT 31.770 160.775 32.045 161.230 ;
        RECT 32.215 160.945 32.460 161.425 ;
        RECT 32.630 160.775 32.890 161.230 ;
        RECT 33.060 160.945 33.320 161.425 ;
        RECT 33.490 160.775 33.750 161.230 ;
        RECT 33.920 160.945 34.180 161.425 ;
        RECT 34.350 160.775 34.610 161.230 ;
        RECT 34.780 160.865 35.040 161.425 ;
        RECT 26.850 160.450 27.020 160.705 ;
        RECT 27.865 160.605 34.610 160.775 ;
        RECT 26.735 160.120 27.020 160.450 ;
        RECT 27.255 160.155 27.585 160.525 ;
        RECT 26.850 159.975 27.020 160.120 ;
        RECT 27.865 160.015 29.030 160.605 ;
        RECT 35.210 160.435 35.460 161.245 ;
        RECT 35.640 160.900 35.900 161.425 ;
        RECT 36.070 160.435 36.320 161.245 ;
        RECT 36.500 160.915 36.805 161.425 ;
        RECT 29.200 160.185 36.320 160.435 ;
        RECT 36.490 160.185 36.805 160.745 ;
        RECT 36.975 160.655 38.645 161.425 ;
        RECT 38.815 160.700 39.105 161.425 ;
        RECT 39.735 160.750 39.995 161.255 ;
        RECT 40.175 161.045 40.505 161.425 ;
        RECT 40.685 160.875 40.855 161.255 ;
        RECT 26.395 159.045 26.665 159.950 ;
        RECT 26.850 159.805 27.515 159.975 ;
        RECT 26.835 158.875 27.165 159.635 ;
        RECT 27.345 159.045 27.515 159.805 ;
        RECT 27.865 159.790 34.610 160.015 ;
        RECT 27.865 158.875 28.135 159.620 ;
        RECT 28.305 159.050 28.595 159.790 ;
        RECT 29.205 159.775 34.610 159.790 ;
        RECT 28.765 158.880 29.020 159.605 ;
        RECT 29.205 159.050 29.465 159.775 ;
        RECT 29.635 158.880 29.880 159.605 ;
        RECT 30.065 159.050 30.325 159.775 ;
        RECT 30.495 158.880 30.740 159.605 ;
        RECT 30.925 159.050 31.185 159.775 ;
        RECT 31.355 158.880 31.600 159.605 ;
        RECT 31.770 159.050 32.030 159.775 ;
        RECT 32.200 158.880 32.460 159.605 ;
        RECT 32.630 159.050 32.890 159.775 ;
        RECT 33.060 158.880 33.320 159.605 ;
        RECT 33.490 159.050 33.750 159.775 ;
        RECT 33.920 158.880 34.180 159.605 ;
        RECT 34.350 159.050 34.610 159.775 ;
        RECT 34.780 158.880 35.040 159.675 ;
        RECT 35.210 159.050 35.460 160.185 ;
        RECT 28.765 158.875 35.040 158.880 ;
        RECT 35.640 158.875 35.900 159.685 ;
        RECT 36.075 159.045 36.320 160.185 ;
        RECT 36.975 159.965 37.725 160.485 ;
        RECT 37.895 160.135 38.645 160.655 ;
        RECT 36.500 158.875 36.795 159.685 ;
        RECT 36.975 158.875 38.645 159.965 ;
        RECT 38.815 158.875 39.105 160.040 ;
        RECT 39.735 159.950 39.905 160.750 ;
        RECT 40.190 160.705 40.855 160.875 ;
        RECT 40.190 160.450 40.360 160.705 ;
        RECT 41.120 160.685 41.375 161.255 ;
        RECT 41.545 161.025 41.875 161.425 ;
        RECT 42.300 160.890 42.830 161.255 ;
        RECT 42.300 160.855 42.475 160.890 ;
        RECT 41.545 160.685 42.475 160.855 ;
        RECT 40.075 160.120 40.360 160.450 ;
        RECT 40.595 160.155 40.925 160.525 ;
        RECT 40.190 159.975 40.360 160.120 ;
        RECT 41.120 160.015 41.290 160.685 ;
        RECT 41.545 160.515 41.715 160.685 ;
        RECT 41.460 160.185 41.715 160.515 ;
        RECT 41.940 160.185 42.135 160.515 ;
        RECT 39.735 159.045 40.005 159.950 ;
        RECT 40.190 159.805 40.855 159.975 ;
        RECT 40.175 158.875 40.505 159.635 ;
        RECT 40.685 159.045 40.855 159.805 ;
        RECT 41.120 159.045 41.455 160.015 ;
        RECT 41.625 158.875 41.795 160.015 ;
        RECT 41.965 159.215 42.135 160.185 ;
        RECT 42.305 159.555 42.475 160.685 ;
        RECT 42.645 159.895 42.815 160.695 ;
        RECT 43.020 160.405 43.295 161.255 ;
        RECT 43.015 160.235 43.295 160.405 ;
        RECT 43.020 160.095 43.295 160.235 ;
        RECT 43.465 159.895 43.655 161.255 ;
        RECT 43.835 160.890 44.345 161.425 ;
        RECT 44.565 160.615 44.810 161.220 ;
        RECT 45.530 160.615 45.775 161.220 ;
        RECT 45.995 160.890 46.505 161.425 ;
        RECT 43.855 160.445 45.085 160.615 ;
        RECT 42.645 159.725 43.655 159.895 ;
        RECT 43.825 159.880 44.575 160.070 ;
        RECT 42.305 159.385 43.430 159.555 ;
        RECT 43.825 159.215 43.995 159.880 ;
        RECT 44.745 159.635 45.085 160.445 ;
        RECT 41.965 159.045 43.995 159.215 ;
        RECT 44.165 158.875 44.335 159.635 ;
        RECT 44.570 159.225 45.085 159.635 ;
        RECT 45.255 160.445 46.485 160.615 ;
        RECT 45.255 159.635 45.595 160.445 ;
        RECT 45.765 159.880 46.515 160.070 ;
        RECT 45.255 159.225 45.770 159.635 ;
        RECT 46.005 158.875 46.175 159.635 ;
        RECT 46.345 159.215 46.515 159.880 ;
        RECT 46.685 159.895 46.875 161.255 ;
        RECT 47.045 160.745 47.320 161.255 ;
        RECT 47.510 160.890 48.040 161.255 ;
        RECT 48.465 161.025 48.795 161.425 ;
        RECT 47.865 160.855 48.040 160.890 ;
        RECT 47.045 160.575 47.325 160.745 ;
        RECT 47.045 160.095 47.320 160.575 ;
        RECT 47.525 159.895 47.695 160.695 ;
        RECT 46.685 159.725 47.695 159.895 ;
        RECT 47.865 160.685 48.795 160.855 ;
        RECT 48.965 160.685 49.220 161.255 ;
        RECT 47.865 159.555 48.035 160.685 ;
        RECT 48.625 160.515 48.795 160.685 ;
        RECT 46.910 159.385 48.035 159.555 ;
        RECT 48.205 160.185 48.400 160.515 ;
        RECT 48.625 160.185 48.880 160.515 ;
        RECT 48.205 159.215 48.375 160.185 ;
        RECT 49.050 160.015 49.220 160.685 ;
        RECT 49.395 160.675 50.605 161.425 ;
        RECT 46.345 159.045 48.375 159.215 ;
        RECT 48.545 158.875 48.715 160.015 ;
        RECT 48.885 159.045 49.220 160.015 ;
        RECT 49.395 159.965 49.915 160.505 ;
        RECT 50.085 160.135 50.605 160.675 ;
        RECT 50.775 160.750 51.035 161.255 ;
        RECT 51.215 161.045 51.545 161.425 ;
        RECT 51.725 160.875 51.895 161.255 ;
        RECT 49.395 158.875 50.605 159.965 ;
        RECT 50.775 159.950 50.945 160.750 ;
        RECT 51.230 160.705 51.895 160.875 ;
        RECT 51.230 160.450 51.400 160.705 ;
        RECT 52.155 160.675 53.365 161.425 ;
        RECT 53.540 160.880 58.885 161.425 ;
        RECT 59.060 160.880 64.405 161.425 ;
        RECT 51.115 160.120 51.400 160.450 ;
        RECT 51.635 160.155 51.965 160.525 ;
        RECT 51.230 159.975 51.400 160.120 ;
        RECT 50.775 159.045 51.045 159.950 ;
        RECT 51.230 159.805 51.895 159.975 ;
        RECT 51.215 158.875 51.545 159.635 ;
        RECT 51.725 159.045 51.895 159.805 ;
        RECT 52.155 159.965 52.675 160.505 ;
        RECT 52.845 160.135 53.365 160.675 ;
        RECT 52.155 158.875 53.365 159.965 ;
        RECT 55.130 159.310 55.480 160.560 ;
        RECT 56.960 160.050 57.300 160.880 ;
        RECT 60.650 159.310 61.000 160.560 ;
        RECT 62.480 160.050 62.820 160.880 ;
        RECT 64.575 160.700 64.865 161.425 ;
        RECT 65.040 160.585 65.300 161.425 ;
        RECT 65.475 160.680 65.730 161.255 ;
        RECT 65.900 161.045 66.230 161.425 ;
        RECT 66.445 160.875 66.615 161.255 ;
        RECT 66.935 160.945 67.215 161.425 ;
        RECT 65.900 160.705 66.615 160.875 ;
        RECT 67.385 160.775 67.645 161.165 ;
        RECT 67.820 160.945 68.075 161.425 ;
        RECT 68.245 160.775 68.540 161.165 ;
        RECT 68.720 160.945 68.995 161.425 ;
        RECT 69.165 160.925 69.465 161.255 ;
        RECT 53.540 158.875 58.885 159.310 ;
        RECT 59.060 158.875 64.405 159.310 ;
        RECT 64.575 158.875 64.865 160.040 ;
        RECT 65.040 158.875 65.300 160.025 ;
        RECT 65.475 159.950 65.645 160.680 ;
        RECT 65.900 160.515 66.070 160.705 ;
        RECT 66.890 160.605 68.540 160.775 ;
        RECT 65.815 160.185 66.070 160.515 ;
        RECT 65.900 159.975 66.070 160.185 ;
        RECT 66.350 160.155 66.705 160.525 ;
        RECT 66.890 160.095 67.295 160.605 ;
        RECT 67.465 160.265 68.605 160.435 ;
        RECT 65.475 159.045 65.730 159.950 ;
        RECT 65.900 159.805 66.615 159.975 ;
        RECT 66.890 159.925 67.645 160.095 ;
        RECT 65.900 158.875 66.230 159.635 ;
        RECT 66.445 159.045 66.615 159.805 ;
        RECT 66.930 158.875 67.215 159.745 ;
        RECT 67.385 159.675 67.645 159.925 ;
        RECT 68.435 160.015 68.605 160.265 ;
        RECT 68.775 160.185 69.125 160.755 ;
        RECT 69.295 160.015 69.465 160.925 ;
        RECT 69.635 160.655 73.145 161.425 ;
        RECT 73.320 160.880 78.665 161.425 ;
        RECT 68.435 159.845 69.465 160.015 ;
        RECT 67.385 159.505 68.505 159.675 ;
        RECT 67.385 159.045 67.645 159.505 ;
        RECT 67.820 158.875 68.075 159.335 ;
        RECT 68.245 159.045 68.505 159.505 ;
        RECT 68.675 158.875 68.985 159.675 ;
        RECT 69.155 159.045 69.465 159.845 ;
        RECT 69.635 159.965 71.325 160.485 ;
        RECT 71.495 160.135 73.145 160.655 ;
        RECT 69.635 158.875 73.145 159.965 ;
        RECT 74.910 159.310 75.260 160.560 ;
        RECT 76.740 160.050 77.080 160.880 ;
        RECT 78.840 160.685 79.095 161.255 ;
        RECT 79.265 161.025 79.595 161.425 ;
        RECT 80.020 160.890 80.550 161.255 ;
        RECT 80.020 160.855 80.195 160.890 ;
        RECT 79.265 160.685 80.195 160.855 ;
        RECT 78.840 160.015 79.010 160.685 ;
        RECT 79.265 160.515 79.435 160.685 ;
        RECT 79.180 160.185 79.435 160.515 ;
        RECT 79.660 160.185 79.855 160.515 ;
        RECT 73.320 158.875 78.665 159.310 ;
        RECT 78.840 159.045 79.175 160.015 ;
        RECT 79.345 158.875 79.515 160.015 ;
        RECT 79.685 159.215 79.855 160.185 ;
        RECT 80.025 159.555 80.195 160.685 ;
        RECT 80.365 159.895 80.535 160.695 ;
        RECT 80.740 160.405 81.015 161.255 ;
        RECT 80.735 160.235 81.015 160.405 ;
        RECT 80.740 160.095 81.015 160.235 ;
        RECT 81.185 159.895 81.375 161.255 ;
        RECT 81.555 160.890 82.065 161.425 ;
        RECT 82.285 160.615 82.530 161.220 ;
        RECT 82.975 160.675 84.185 161.425 ;
        RECT 81.575 160.445 82.805 160.615 ;
        RECT 80.365 159.725 81.375 159.895 ;
        RECT 81.545 159.880 82.295 160.070 ;
        RECT 80.025 159.385 81.150 159.555 ;
        RECT 81.545 159.215 81.715 159.880 ;
        RECT 82.465 159.635 82.805 160.445 ;
        RECT 79.685 159.045 81.715 159.215 ;
        RECT 81.885 158.875 82.055 159.635 ;
        RECT 82.290 159.225 82.805 159.635 ;
        RECT 82.975 159.965 83.495 160.505 ;
        RECT 83.665 160.135 84.185 160.675 ;
        RECT 84.415 160.605 84.625 161.425 ;
        RECT 84.795 160.625 85.125 161.255 ;
        RECT 84.795 160.025 85.045 160.625 ;
        RECT 85.295 160.605 85.525 161.425 ;
        RECT 85.825 160.875 85.995 161.255 ;
        RECT 86.175 161.045 86.505 161.425 ;
        RECT 85.825 160.705 86.490 160.875 ;
        RECT 86.685 160.750 86.945 161.255 ;
        RECT 87.215 160.960 87.465 161.425 ;
        RECT 87.635 160.785 87.805 161.255 ;
        RECT 88.055 160.965 88.225 161.425 ;
        RECT 88.475 160.785 88.645 161.255 ;
        RECT 88.895 160.965 89.065 161.425 ;
        RECT 89.315 160.785 89.485 161.255 ;
        RECT 89.855 160.965 90.120 161.425 ;
        RECT 85.215 160.185 85.545 160.435 ;
        RECT 85.755 160.155 86.085 160.525 ;
        RECT 86.320 160.450 86.490 160.705 ;
        RECT 86.320 160.120 86.605 160.450 ;
        RECT 82.975 158.875 84.185 159.965 ;
        RECT 84.415 158.875 84.625 160.015 ;
        RECT 84.795 159.045 85.125 160.025 ;
        RECT 85.295 158.875 85.525 160.015 ;
        RECT 86.320 159.975 86.490 160.120 ;
        RECT 85.825 159.805 86.490 159.975 ;
        RECT 86.775 159.950 86.945 160.750 ;
        RECT 85.825 159.045 85.995 159.805 ;
        RECT 86.175 158.875 86.505 159.635 ;
        RECT 86.675 159.045 86.945 159.950 ;
        RECT 87.115 160.605 89.485 160.785 ;
        RECT 90.335 160.700 90.625 161.425 ;
        RECT 91.255 160.655 93.845 161.425 ;
        RECT 87.115 160.015 87.465 160.605 ;
        RECT 87.635 160.185 90.145 160.435 ;
        RECT 87.115 159.845 89.565 160.015 ;
        RECT 87.115 159.825 87.885 159.845 ;
        RECT 87.215 158.875 87.385 159.335 ;
        RECT 87.555 159.045 87.885 159.825 ;
        RECT 88.055 158.875 88.225 159.675 ;
        RECT 88.395 159.045 88.725 159.845 ;
        RECT 88.895 158.875 89.065 159.675 ;
        RECT 89.235 159.045 89.565 159.845 ;
        RECT 89.825 158.875 90.120 160.015 ;
        RECT 90.335 158.875 90.625 160.040 ;
        RECT 91.255 159.965 92.465 160.485 ;
        RECT 92.635 160.135 93.845 160.655 ;
        RECT 94.075 160.605 94.285 161.425 ;
        RECT 94.455 160.625 94.785 161.255 ;
        RECT 94.455 160.025 94.705 160.625 ;
        RECT 94.955 160.605 95.185 161.425 ;
        RECT 95.855 160.655 97.525 161.425 ;
        RECT 94.875 160.185 95.205 160.435 ;
        RECT 91.255 158.875 93.845 159.965 ;
        RECT 94.075 158.875 94.285 160.015 ;
        RECT 94.455 159.045 94.785 160.025 ;
        RECT 94.955 158.875 95.185 160.015 ;
        RECT 95.855 159.965 96.605 160.485 ;
        RECT 96.775 160.135 97.525 160.655 ;
        RECT 98.070 160.715 98.325 161.245 ;
        RECT 98.505 160.965 98.790 161.425 ;
        RECT 95.855 158.875 97.525 159.965 ;
        RECT 98.070 159.855 98.250 160.715 ;
        RECT 98.970 160.515 99.220 161.165 ;
        RECT 98.420 160.185 99.220 160.515 ;
        RECT 98.070 159.385 98.325 159.855 ;
        RECT 97.985 159.215 98.325 159.385 ;
        RECT 98.070 159.185 98.325 159.215 ;
        RECT 98.505 158.875 98.790 159.675 ;
        RECT 98.970 159.595 99.220 160.185 ;
        RECT 99.420 160.830 99.740 161.160 ;
        RECT 99.920 160.945 100.580 161.425 ;
        RECT 100.780 161.035 101.630 161.205 ;
        RECT 99.420 159.935 99.610 160.830 ;
        RECT 99.930 160.505 100.590 160.775 ;
        RECT 100.260 160.445 100.590 160.505 ;
        RECT 99.780 160.275 100.110 160.335 ;
        RECT 100.780 160.275 100.950 161.035 ;
        RECT 102.190 160.965 102.510 161.425 ;
        RECT 102.710 160.785 102.960 161.215 ;
        RECT 103.250 160.985 103.660 161.425 ;
        RECT 103.830 161.045 104.845 161.245 ;
        RECT 101.120 160.615 102.370 160.785 ;
        RECT 101.120 160.495 101.450 160.615 ;
        RECT 99.780 160.105 101.680 160.275 ;
        RECT 99.420 159.765 101.340 159.935 ;
        RECT 99.420 159.745 99.740 159.765 ;
        RECT 98.970 159.085 99.300 159.595 ;
        RECT 99.570 159.135 99.740 159.745 ;
        RECT 101.510 159.595 101.680 160.105 ;
        RECT 101.850 160.035 102.030 160.445 ;
        RECT 102.200 159.855 102.370 160.615 ;
        RECT 99.910 158.875 100.240 159.565 ;
        RECT 100.470 159.425 101.680 159.595 ;
        RECT 101.850 159.545 102.370 159.855 ;
        RECT 102.540 160.445 102.960 160.785 ;
        RECT 103.250 160.445 103.660 160.775 ;
        RECT 102.540 159.675 102.730 160.445 ;
        RECT 103.830 160.315 104.000 161.045 ;
        RECT 105.145 160.875 105.315 161.205 ;
        RECT 105.485 161.045 105.815 161.425 ;
        RECT 104.170 160.495 104.520 160.865 ;
        RECT 103.830 160.275 104.250 160.315 ;
        RECT 102.900 160.105 104.250 160.275 ;
        RECT 102.900 159.945 103.150 160.105 ;
        RECT 103.660 159.675 103.910 159.935 ;
        RECT 102.540 159.425 103.910 159.675 ;
        RECT 100.470 159.135 100.710 159.425 ;
        RECT 101.510 159.345 101.680 159.425 ;
        RECT 100.910 158.875 101.330 159.255 ;
        RECT 101.510 159.095 102.140 159.345 ;
        RECT 102.610 158.875 102.940 159.255 ;
        RECT 103.110 159.135 103.280 159.425 ;
        RECT 104.080 159.260 104.250 160.105 ;
        RECT 104.700 159.935 104.920 160.805 ;
        RECT 105.145 160.685 105.840 160.875 ;
        RECT 104.420 159.555 104.920 159.935 ;
        RECT 105.090 159.885 105.500 160.505 ;
        RECT 105.670 159.715 105.840 160.685 ;
        RECT 105.145 159.545 105.840 159.715 ;
        RECT 103.460 158.875 103.840 159.255 ;
        RECT 104.080 159.090 104.910 159.260 ;
        RECT 105.145 159.045 105.315 159.545 ;
        RECT 105.485 158.875 105.815 159.375 ;
        RECT 106.030 159.045 106.255 161.165 ;
        RECT 106.425 161.045 106.755 161.425 ;
        RECT 106.925 160.875 107.095 161.165 ;
        RECT 106.430 160.705 107.095 160.875 ;
        RECT 106.430 159.715 106.660 160.705 ;
        RECT 107.815 160.655 110.405 161.425 ;
        RECT 110.580 160.880 115.925 161.425 ;
        RECT 106.830 159.885 107.180 160.535 ;
        RECT 107.815 159.965 109.025 160.485 ;
        RECT 109.195 160.135 110.405 160.655 ;
        RECT 106.430 159.545 107.095 159.715 ;
        RECT 106.425 158.875 106.755 159.375 ;
        RECT 106.925 159.045 107.095 159.545 ;
        RECT 107.815 158.875 110.405 159.965 ;
        RECT 112.170 159.310 112.520 160.560 ;
        RECT 114.000 160.050 114.340 160.880 ;
        RECT 116.095 160.700 116.385 161.425 ;
        RECT 116.555 160.655 118.225 161.425 ;
        RECT 110.580 158.875 115.925 159.310 ;
        RECT 116.095 158.875 116.385 160.040 ;
        RECT 116.555 159.965 117.305 160.485 ;
        RECT 117.475 160.135 118.225 160.655 ;
        RECT 118.545 160.625 118.875 161.425 ;
        RECT 119.045 160.775 119.215 161.255 ;
        RECT 119.385 160.945 119.715 161.425 ;
        RECT 119.885 160.775 120.055 161.255 ;
        RECT 120.305 160.945 120.545 161.425 ;
        RECT 120.725 160.775 120.895 161.255 ;
        RECT 119.045 160.605 120.055 160.775 ;
        RECT 120.260 160.605 120.895 160.775 ;
        RECT 121.155 160.675 122.365 161.425 ;
        RECT 122.540 160.880 127.885 161.425 ;
        RECT 119.045 160.065 119.540 160.605 ;
        RECT 120.260 160.435 120.430 160.605 ;
        RECT 119.930 160.265 120.430 160.435 ;
        RECT 116.555 158.875 118.225 159.965 ;
        RECT 118.545 158.875 118.875 160.025 ;
        RECT 119.045 159.895 120.055 160.065 ;
        RECT 119.045 159.045 119.215 159.895 ;
        RECT 119.385 158.875 119.715 159.675 ;
        RECT 119.885 159.045 120.055 159.895 ;
        RECT 120.260 160.025 120.430 160.265 ;
        RECT 120.600 160.195 120.980 160.435 ;
        RECT 120.260 159.855 120.975 160.025 ;
        RECT 120.235 158.875 120.475 159.675 ;
        RECT 120.645 159.045 120.975 159.855 ;
        RECT 121.155 159.965 121.675 160.505 ;
        RECT 121.845 160.135 122.365 160.675 ;
        RECT 121.155 158.875 122.365 159.965 ;
        RECT 124.130 159.310 124.480 160.560 ;
        RECT 125.960 160.050 126.300 160.880 ;
        RECT 128.055 160.675 129.265 161.425 ;
        RECT 128.055 159.965 128.575 160.505 ;
        RECT 128.745 160.135 129.265 160.675 ;
        RECT 122.540 158.875 127.885 159.310 ;
        RECT 128.055 158.875 129.265 159.965 ;
        RECT 9.290 158.705 129.350 158.875 ;
        RECT 9.375 157.615 10.585 158.705 ;
        RECT 9.375 156.905 9.895 157.445 ;
        RECT 10.065 157.075 10.585 157.615 ;
        RECT 11.590 157.725 11.845 158.395 ;
        RECT 12.025 157.905 12.310 158.705 ;
        RECT 12.490 157.985 12.820 158.495 ;
        RECT 9.375 156.155 10.585 156.905 ;
        RECT 11.590 156.865 11.770 157.725 ;
        RECT 12.490 157.395 12.740 157.985 ;
        RECT 13.090 157.835 13.260 158.445 ;
        RECT 13.430 158.015 13.760 158.705 ;
        RECT 13.990 158.155 14.230 158.445 ;
        RECT 14.430 158.325 14.850 158.705 ;
        RECT 15.030 158.235 15.660 158.485 ;
        RECT 16.130 158.325 16.460 158.705 ;
        RECT 15.030 158.155 15.200 158.235 ;
        RECT 16.630 158.155 16.800 158.445 ;
        RECT 16.980 158.325 17.360 158.705 ;
        RECT 17.600 158.320 18.430 158.490 ;
        RECT 13.990 157.985 15.200 158.155 ;
        RECT 11.940 157.065 12.740 157.395 ;
        RECT 11.590 156.665 11.845 156.865 ;
        RECT 11.505 156.495 11.845 156.665 ;
        RECT 11.590 156.335 11.845 156.495 ;
        RECT 12.025 156.155 12.310 156.615 ;
        RECT 12.490 156.415 12.740 157.065 ;
        RECT 12.940 157.815 13.260 157.835 ;
        RECT 12.940 157.645 14.860 157.815 ;
        RECT 12.940 156.750 13.130 157.645 ;
        RECT 15.030 157.475 15.200 157.985 ;
        RECT 15.370 157.725 15.890 158.035 ;
        RECT 13.300 157.305 15.200 157.475 ;
        RECT 13.300 157.245 13.630 157.305 ;
        RECT 13.780 157.075 14.110 157.135 ;
        RECT 13.450 156.805 14.110 157.075 ;
        RECT 12.940 156.420 13.260 156.750 ;
        RECT 13.440 156.155 14.100 156.635 ;
        RECT 14.300 156.545 14.470 157.305 ;
        RECT 15.370 157.135 15.550 157.545 ;
        RECT 14.640 156.965 14.970 157.085 ;
        RECT 15.720 156.965 15.890 157.725 ;
        RECT 14.640 156.795 15.890 156.965 ;
        RECT 16.060 157.905 17.430 158.155 ;
        RECT 16.060 157.135 16.250 157.905 ;
        RECT 17.180 157.645 17.430 157.905 ;
        RECT 16.420 157.475 16.670 157.635 ;
        RECT 17.600 157.475 17.770 158.320 ;
        RECT 18.665 158.035 18.835 158.535 ;
        RECT 19.005 158.205 19.335 158.705 ;
        RECT 17.940 157.645 18.440 158.025 ;
        RECT 18.665 157.865 19.360 158.035 ;
        RECT 16.420 157.305 17.770 157.475 ;
        RECT 17.350 157.265 17.770 157.305 ;
        RECT 16.060 156.795 16.480 157.135 ;
        RECT 16.770 156.805 17.180 157.135 ;
        RECT 14.300 156.375 15.150 156.545 ;
        RECT 15.710 156.155 16.030 156.615 ;
        RECT 16.230 156.365 16.480 156.795 ;
        RECT 16.770 156.155 17.180 156.595 ;
        RECT 17.350 156.535 17.520 157.265 ;
        RECT 17.690 156.715 18.040 157.085 ;
        RECT 18.220 156.775 18.440 157.645 ;
        RECT 18.610 157.075 19.020 157.695 ;
        RECT 19.190 156.895 19.360 157.865 ;
        RECT 18.665 156.705 19.360 156.895 ;
        RECT 17.350 156.335 18.365 156.535 ;
        RECT 18.665 156.375 18.835 156.705 ;
        RECT 19.005 156.155 19.335 156.535 ;
        RECT 19.550 156.415 19.775 158.535 ;
        RECT 19.945 158.205 20.275 158.705 ;
        RECT 20.445 158.035 20.615 158.535 ;
        RECT 19.950 157.865 20.615 158.035 ;
        RECT 19.950 156.875 20.180 157.865 ;
        RECT 20.350 157.045 20.700 157.695 ;
        RECT 20.875 157.615 24.385 158.705 ;
        RECT 20.875 157.095 22.565 157.615 ;
        RECT 24.595 157.565 24.825 158.705 ;
        RECT 24.995 157.555 25.325 158.535 ;
        RECT 25.495 157.565 25.705 158.705 ;
        RECT 22.735 156.925 24.385 157.445 ;
        RECT 24.575 157.145 24.905 157.395 ;
        RECT 19.950 156.705 20.615 156.875 ;
        RECT 19.945 156.155 20.275 156.535 ;
        RECT 20.445 156.415 20.615 156.705 ;
        RECT 20.875 156.155 24.385 156.925 ;
        RECT 24.595 156.155 24.825 156.975 ;
        RECT 25.075 156.955 25.325 157.555 ;
        RECT 25.935 157.540 26.225 158.705 ;
        RECT 26.395 157.945 26.910 158.355 ;
        RECT 27.145 157.945 27.315 158.705 ;
        RECT 27.485 158.365 29.515 158.535 ;
        RECT 26.395 157.135 26.735 157.945 ;
        RECT 27.485 157.700 27.655 158.365 ;
        RECT 28.050 158.025 29.175 158.195 ;
        RECT 26.905 157.510 27.655 157.700 ;
        RECT 27.825 157.685 28.835 157.855 ;
        RECT 24.995 156.325 25.325 156.955 ;
        RECT 25.495 156.155 25.705 156.975 ;
        RECT 26.395 156.965 27.625 157.135 ;
        RECT 25.935 156.155 26.225 156.880 ;
        RECT 26.670 156.360 26.915 156.965 ;
        RECT 27.135 156.155 27.645 156.690 ;
        RECT 27.825 156.325 28.015 157.685 ;
        RECT 28.185 157.005 28.460 157.485 ;
        RECT 28.185 156.835 28.465 157.005 ;
        RECT 28.665 156.885 28.835 157.685 ;
        RECT 29.005 156.895 29.175 158.025 ;
        RECT 29.345 157.395 29.515 158.365 ;
        RECT 29.685 157.565 29.855 158.705 ;
        RECT 30.025 157.565 30.360 158.535 ;
        RECT 31.455 157.870 31.840 158.705 ;
        RECT 32.010 157.700 32.270 158.505 ;
        RECT 32.440 157.870 32.700 158.705 ;
        RECT 32.870 157.700 33.125 158.505 ;
        RECT 33.300 157.870 33.560 158.705 ;
        RECT 33.730 157.700 33.985 158.505 ;
        RECT 34.160 157.870 34.505 158.705 ;
        RECT 29.345 157.065 29.540 157.395 ;
        RECT 29.765 157.065 30.020 157.395 ;
        RECT 29.765 156.895 29.935 157.065 ;
        RECT 30.190 156.895 30.360 157.565 ;
        RECT 28.185 156.325 28.460 156.835 ;
        RECT 29.005 156.725 29.935 156.895 ;
        RECT 29.005 156.690 29.180 156.725 ;
        RECT 28.650 156.325 29.180 156.690 ;
        RECT 29.605 156.155 29.935 156.555 ;
        RECT 30.105 156.325 30.360 156.895 ;
        RECT 31.455 157.530 34.485 157.700 ;
        RECT 31.455 156.965 31.755 157.530 ;
        RECT 31.930 157.135 34.145 157.360 ;
        RECT 34.315 156.965 34.485 157.530 ;
        RECT 31.455 156.795 34.485 156.965 ;
        RECT 34.680 157.565 35.015 158.535 ;
        RECT 35.185 157.565 35.355 158.705 ;
        RECT 35.525 158.365 37.555 158.535 ;
        RECT 34.680 156.895 34.850 157.565 ;
        RECT 35.525 157.395 35.695 158.365 ;
        RECT 35.020 157.065 35.275 157.395 ;
        RECT 35.500 157.065 35.695 157.395 ;
        RECT 35.865 158.025 36.990 158.195 ;
        RECT 35.105 156.895 35.275 157.065 ;
        RECT 35.865 156.895 36.035 158.025 ;
        RECT 31.975 156.155 32.275 156.625 ;
        RECT 32.445 156.350 32.700 156.795 ;
        RECT 32.870 156.155 33.130 156.625 ;
        RECT 33.300 156.350 33.560 156.795 ;
        RECT 33.730 156.155 34.025 156.625 ;
        RECT 34.680 156.325 34.935 156.895 ;
        RECT 35.105 156.725 36.035 156.895 ;
        RECT 36.205 157.685 37.215 157.855 ;
        RECT 36.205 156.885 36.375 157.685 ;
        RECT 36.580 157.345 36.855 157.485 ;
        RECT 36.575 157.175 36.855 157.345 ;
        RECT 35.860 156.690 36.035 156.725 ;
        RECT 35.105 156.155 35.435 156.555 ;
        RECT 35.860 156.325 36.390 156.690 ;
        RECT 36.580 156.325 36.855 157.175 ;
        RECT 37.025 156.325 37.215 157.685 ;
        RECT 37.385 157.700 37.555 158.365 ;
        RECT 37.725 157.945 37.895 158.705 ;
        RECT 38.130 157.945 38.645 158.355 ;
        RECT 37.385 157.510 38.135 157.700 ;
        RECT 38.305 157.135 38.645 157.945 ;
        RECT 37.415 156.965 38.645 157.135 ;
        RECT 38.815 157.615 40.485 158.705 ;
        RECT 40.660 158.270 46.005 158.705 ;
        RECT 46.180 158.270 51.525 158.705 ;
        RECT 38.815 157.095 39.565 157.615 ;
        RECT 37.395 156.155 37.905 156.690 ;
        RECT 38.125 156.360 38.370 156.965 ;
        RECT 39.735 156.925 40.485 157.445 ;
        RECT 42.250 157.020 42.600 158.270 ;
        RECT 38.815 156.155 40.485 156.925 ;
        RECT 44.080 156.700 44.420 157.530 ;
        RECT 47.770 157.020 48.120 158.270 ;
        RECT 51.695 157.540 51.985 158.705 ;
        RECT 52.195 157.565 52.425 158.705 ;
        RECT 52.595 157.555 52.925 158.535 ;
        RECT 53.095 157.565 53.305 158.705 ;
        RECT 53.685 157.555 54.015 158.705 ;
        RECT 54.185 157.685 54.355 158.535 ;
        RECT 54.525 157.905 54.855 158.705 ;
        RECT 55.025 157.685 55.195 158.535 ;
        RECT 55.375 157.905 55.615 158.705 ;
        RECT 55.785 157.725 56.115 158.535 ;
        RECT 49.600 156.700 49.940 157.530 ;
        RECT 52.175 157.145 52.505 157.395 ;
        RECT 40.660 156.155 46.005 156.700 ;
        RECT 46.180 156.155 51.525 156.700 ;
        RECT 51.695 156.155 51.985 156.880 ;
        RECT 52.195 156.155 52.425 156.975 ;
        RECT 52.675 156.955 52.925 157.555 ;
        RECT 54.185 157.515 55.195 157.685 ;
        RECT 55.400 157.555 56.115 157.725 ;
        RECT 54.185 157.345 54.680 157.515 ;
        RECT 54.185 157.175 54.685 157.345 ;
        RECT 55.400 157.315 55.570 157.555 ;
        RECT 56.300 157.515 56.555 158.395 ;
        RECT 56.725 157.565 57.030 158.705 ;
        RECT 57.370 158.325 57.700 158.705 ;
        RECT 57.880 158.155 58.050 158.445 ;
        RECT 58.220 158.245 58.470 158.705 ;
        RECT 57.250 157.985 58.050 158.155 ;
        RECT 58.640 158.195 59.510 158.535 ;
        RECT 54.185 156.975 54.680 157.175 ;
        RECT 55.070 157.145 55.570 157.315 ;
        RECT 55.740 157.145 56.120 157.385 ;
        RECT 55.400 156.975 55.570 157.145 ;
        RECT 52.595 156.325 52.925 156.955 ;
        RECT 53.095 156.155 53.305 156.975 ;
        RECT 53.685 156.155 54.015 156.955 ;
        RECT 54.185 156.805 55.195 156.975 ;
        RECT 55.400 156.805 56.035 156.975 ;
        RECT 54.185 156.325 54.355 156.805 ;
        RECT 54.525 156.155 54.855 156.635 ;
        RECT 55.025 156.325 55.195 156.805 ;
        RECT 55.445 156.155 55.685 156.635 ;
        RECT 55.865 156.325 56.035 156.805 ;
        RECT 56.300 156.865 56.510 157.515 ;
        RECT 57.250 157.395 57.420 157.985 ;
        RECT 58.640 157.815 58.810 158.195 ;
        RECT 59.745 158.075 59.915 158.535 ;
        RECT 60.085 158.245 60.455 158.705 ;
        RECT 60.750 158.105 60.920 158.445 ;
        RECT 61.090 158.275 61.420 158.705 ;
        RECT 61.655 158.105 61.825 158.445 ;
        RECT 57.590 157.645 58.810 157.815 ;
        RECT 58.980 157.735 59.440 158.025 ;
        RECT 59.745 157.905 60.305 158.075 ;
        RECT 60.750 157.935 61.825 158.105 ;
        RECT 61.995 158.205 62.675 158.535 ;
        RECT 62.890 158.205 63.140 158.535 ;
        RECT 63.310 158.245 63.560 158.705 ;
        RECT 60.135 157.765 60.305 157.905 ;
        RECT 58.980 157.725 59.945 157.735 ;
        RECT 58.640 157.555 58.810 157.645 ;
        RECT 59.270 157.565 59.945 157.725 ;
        RECT 56.680 157.365 57.420 157.395 ;
        RECT 56.680 157.065 57.595 157.365 ;
        RECT 57.270 156.890 57.595 157.065 ;
        RECT 56.300 156.335 56.555 156.865 ;
        RECT 56.725 156.155 57.030 156.615 ;
        RECT 57.275 156.535 57.595 156.890 ;
        RECT 57.765 157.105 58.305 157.475 ;
        RECT 58.640 157.385 59.045 157.555 ;
        RECT 57.765 156.705 58.005 157.105 ;
        RECT 58.485 156.935 58.705 157.215 ;
        RECT 58.175 156.765 58.705 156.935 ;
        RECT 58.175 156.535 58.345 156.765 ;
        RECT 58.875 156.605 59.045 157.385 ;
        RECT 59.215 156.775 59.565 157.395 ;
        RECT 59.735 156.775 59.945 157.565 ;
        RECT 60.135 157.595 61.635 157.765 ;
        RECT 60.135 156.905 60.305 157.595 ;
        RECT 61.995 157.425 62.165 158.205 ;
        RECT 62.970 158.075 63.140 158.205 ;
        RECT 60.475 157.255 62.165 157.425 ;
        RECT 62.335 157.645 62.800 158.035 ;
        RECT 62.970 157.905 63.365 158.075 ;
        RECT 60.475 157.075 60.645 157.255 ;
        RECT 57.275 156.365 58.345 156.535 ;
        RECT 58.515 156.155 58.705 156.595 ;
        RECT 58.875 156.325 59.825 156.605 ;
        RECT 60.135 156.515 60.395 156.905 ;
        RECT 60.815 156.835 61.605 157.085 ;
        RECT 60.045 156.345 60.395 156.515 ;
        RECT 60.605 156.155 60.935 156.615 ;
        RECT 61.810 156.545 61.980 157.255 ;
        RECT 62.335 157.055 62.505 157.645 ;
        RECT 62.150 156.835 62.505 157.055 ;
        RECT 62.675 156.835 63.025 157.455 ;
        RECT 63.195 156.545 63.365 157.905 ;
        RECT 63.730 157.735 64.055 158.520 ;
        RECT 63.535 156.685 63.995 157.735 ;
        RECT 61.810 156.375 62.665 156.545 ;
        RECT 62.870 156.375 63.365 156.545 ;
        RECT 63.535 156.155 63.865 156.515 ;
        RECT 64.225 156.415 64.395 158.535 ;
        RECT 64.565 158.205 64.895 158.705 ;
        RECT 65.065 158.035 65.320 158.535 ;
        RECT 64.570 157.865 65.320 158.035 ;
        RECT 64.570 156.875 64.800 157.865 ;
        RECT 64.970 157.045 65.320 157.695 ;
        RECT 65.495 157.615 66.705 158.705 ;
        RECT 65.495 157.075 66.015 157.615 ;
        RECT 66.880 157.555 67.140 158.705 ;
        RECT 67.315 157.630 67.570 158.535 ;
        RECT 67.740 157.945 68.070 158.705 ;
        RECT 68.285 157.775 68.455 158.535 ;
        RECT 66.185 156.905 66.705 157.445 ;
        RECT 64.570 156.705 65.320 156.875 ;
        RECT 64.565 156.155 64.895 156.535 ;
        RECT 65.065 156.415 65.320 156.705 ;
        RECT 65.495 156.155 66.705 156.905 ;
        RECT 66.880 156.155 67.140 156.995 ;
        RECT 67.315 156.900 67.485 157.630 ;
        RECT 67.740 157.605 68.455 157.775 ;
        RECT 68.805 157.775 68.975 158.535 ;
        RECT 69.190 157.945 69.520 158.705 ;
        RECT 68.805 157.605 69.520 157.775 ;
        RECT 69.690 157.630 69.945 158.535 ;
        RECT 67.740 157.395 67.910 157.605 ;
        RECT 67.655 157.065 67.910 157.395 ;
        RECT 67.315 156.325 67.570 156.900 ;
        RECT 67.740 156.875 67.910 157.065 ;
        RECT 68.190 157.055 68.545 157.425 ;
        RECT 68.715 157.055 69.070 157.425 ;
        RECT 69.350 157.395 69.520 157.605 ;
        RECT 69.350 157.065 69.605 157.395 ;
        RECT 69.350 156.875 69.520 157.065 ;
        RECT 69.775 156.900 69.945 157.630 ;
        RECT 70.120 157.555 70.380 158.705 ;
        RECT 70.645 157.775 70.815 158.535 ;
        RECT 71.030 157.945 71.360 158.705 ;
        RECT 70.645 157.605 71.360 157.775 ;
        RECT 71.530 157.630 71.785 158.535 ;
        RECT 70.555 157.055 70.910 157.425 ;
        RECT 71.190 157.395 71.360 157.605 ;
        RECT 71.190 157.065 71.445 157.395 ;
        RECT 67.740 156.705 68.455 156.875 ;
        RECT 67.740 156.155 68.070 156.535 ;
        RECT 68.285 156.325 68.455 156.705 ;
        RECT 68.805 156.705 69.520 156.875 ;
        RECT 68.805 156.325 68.975 156.705 ;
        RECT 69.190 156.155 69.520 156.535 ;
        RECT 69.690 156.325 69.945 156.900 ;
        RECT 70.120 156.155 70.380 156.995 ;
        RECT 71.190 156.875 71.360 157.065 ;
        RECT 71.615 156.900 71.785 157.630 ;
        RECT 71.960 157.555 72.220 158.705 ;
        RECT 72.395 157.615 73.605 158.705 ;
        RECT 73.775 157.615 77.285 158.705 ;
        RECT 72.395 157.075 72.915 157.615 ;
        RECT 70.645 156.705 71.360 156.875 ;
        RECT 70.645 156.325 70.815 156.705 ;
        RECT 71.030 156.155 71.360 156.535 ;
        RECT 71.530 156.325 71.785 156.900 ;
        RECT 71.960 156.155 72.220 156.995 ;
        RECT 73.085 156.905 73.605 157.445 ;
        RECT 73.775 157.095 75.465 157.615 ;
        RECT 77.455 157.540 77.745 158.705 ;
        RECT 78.375 157.615 80.045 158.705 ;
        RECT 80.590 157.725 80.845 158.395 ;
        RECT 81.025 157.905 81.310 158.705 ;
        RECT 81.490 157.985 81.820 158.495 ;
        RECT 75.635 156.925 77.285 157.445 ;
        RECT 78.375 157.095 79.125 157.615 ;
        RECT 79.295 156.925 80.045 157.445 ;
        RECT 80.590 157.345 80.770 157.725 ;
        RECT 81.490 157.395 81.740 157.985 ;
        RECT 82.090 157.835 82.260 158.445 ;
        RECT 82.430 158.015 82.760 158.705 ;
        RECT 82.990 158.155 83.230 158.445 ;
        RECT 83.430 158.325 83.850 158.705 ;
        RECT 84.030 158.235 84.660 158.485 ;
        RECT 85.130 158.325 85.460 158.705 ;
        RECT 84.030 158.155 84.200 158.235 ;
        RECT 85.630 158.155 85.800 158.445 ;
        RECT 85.980 158.325 86.360 158.705 ;
        RECT 86.600 158.320 87.430 158.490 ;
        RECT 82.990 157.985 84.200 158.155 ;
        RECT 80.505 157.175 80.770 157.345 ;
        RECT 72.395 156.155 73.605 156.905 ;
        RECT 73.775 156.155 77.285 156.925 ;
        RECT 77.455 156.155 77.745 156.880 ;
        RECT 78.375 156.155 80.045 156.925 ;
        RECT 80.590 156.865 80.770 157.175 ;
        RECT 80.940 157.065 81.740 157.395 ;
        RECT 80.590 156.335 80.845 156.865 ;
        RECT 81.025 156.155 81.310 156.615 ;
        RECT 81.490 156.415 81.740 157.065 ;
        RECT 81.940 157.815 82.260 157.835 ;
        RECT 81.940 157.645 83.860 157.815 ;
        RECT 81.940 156.750 82.130 157.645 ;
        RECT 84.030 157.475 84.200 157.985 ;
        RECT 84.370 157.725 84.890 158.035 ;
        RECT 82.300 157.305 84.200 157.475 ;
        RECT 82.300 157.245 82.630 157.305 ;
        RECT 82.780 157.075 83.110 157.135 ;
        RECT 82.450 156.805 83.110 157.075 ;
        RECT 81.940 156.420 82.260 156.750 ;
        RECT 82.440 156.155 83.100 156.635 ;
        RECT 83.300 156.545 83.470 157.305 ;
        RECT 84.370 157.135 84.550 157.545 ;
        RECT 83.640 156.965 83.970 157.085 ;
        RECT 84.720 156.965 84.890 157.725 ;
        RECT 83.640 156.795 84.890 156.965 ;
        RECT 85.060 157.905 86.430 158.155 ;
        RECT 85.060 157.135 85.250 157.905 ;
        RECT 86.180 157.645 86.430 157.905 ;
        RECT 85.420 157.475 85.670 157.635 ;
        RECT 86.600 157.475 86.770 158.320 ;
        RECT 87.665 158.035 87.835 158.535 ;
        RECT 88.005 158.205 88.335 158.705 ;
        RECT 86.940 157.645 87.440 158.025 ;
        RECT 87.665 157.865 88.360 158.035 ;
        RECT 85.420 157.305 86.770 157.475 ;
        RECT 86.350 157.265 86.770 157.305 ;
        RECT 85.060 156.795 85.480 157.135 ;
        RECT 85.770 156.805 86.180 157.135 ;
        RECT 83.300 156.375 84.150 156.545 ;
        RECT 84.710 156.155 85.030 156.615 ;
        RECT 85.230 156.365 85.480 156.795 ;
        RECT 85.770 156.155 86.180 156.595 ;
        RECT 86.350 156.535 86.520 157.265 ;
        RECT 86.690 156.715 87.040 157.085 ;
        RECT 87.220 156.775 87.440 157.645 ;
        RECT 87.610 157.075 88.020 157.695 ;
        RECT 88.190 156.895 88.360 157.865 ;
        RECT 87.665 156.705 88.360 156.895 ;
        RECT 86.350 156.335 87.365 156.535 ;
        RECT 87.665 156.375 87.835 156.705 ;
        RECT 88.005 156.155 88.335 156.535 ;
        RECT 88.550 156.415 88.775 158.535 ;
        RECT 88.945 158.205 89.275 158.705 ;
        RECT 89.445 158.035 89.615 158.535 ;
        RECT 88.950 157.865 89.615 158.035 ;
        RECT 88.950 156.875 89.180 157.865 ;
        RECT 90.710 157.725 90.965 158.395 ;
        RECT 91.145 157.905 91.430 158.705 ;
        RECT 91.610 157.985 91.940 158.495 ;
        RECT 89.350 157.045 89.700 157.695 ;
        RECT 88.950 156.705 89.615 156.875 ;
        RECT 88.945 156.155 89.275 156.535 ;
        RECT 89.445 156.415 89.615 156.705 ;
        RECT 90.710 156.865 90.890 157.725 ;
        RECT 91.610 157.395 91.860 157.985 ;
        RECT 92.210 157.835 92.380 158.445 ;
        RECT 92.550 158.015 92.880 158.705 ;
        RECT 93.110 158.155 93.350 158.445 ;
        RECT 93.550 158.325 93.970 158.705 ;
        RECT 94.150 158.235 94.780 158.485 ;
        RECT 95.250 158.325 95.580 158.705 ;
        RECT 94.150 158.155 94.320 158.235 ;
        RECT 95.750 158.155 95.920 158.445 ;
        RECT 96.100 158.325 96.480 158.705 ;
        RECT 96.720 158.320 97.550 158.490 ;
        RECT 93.110 157.985 94.320 158.155 ;
        RECT 91.060 157.065 91.860 157.395 ;
        RECT 90.710 156.665 90.965 156.865 ;
        RECT 90.625 156.495 90.965 156.665 ;
        RECT 90.710 156.335 90.965 156.495 ;
        RECT 91.145 156.155 91.430 156.615 ;
        RECT 91.610 156.415 91.860 157.065 ;
        RECT 92.060 157.815 92.380 157.835 ;
        RECT 92.060 157.645 93.980 157.815 ;
        RECT 92.060 156.750 92.250 157.645 ;
        RECT 94.150 157.475 94.320 157.985 ;
        RECT 94.490 157.725 95.010 158.035 ;
        RECT 92.420 157.305 94.320 157.475 ;
        RECT 92.420 157.245 92.750 157.305 ;
        RECT 92.900 157.075 93.230 157.135 ;
        RECT 92.570 156.805 93.230 157.075 ;
        RECT 92.060 156.420 92.380 156.750 ;
        RECT 92.560 156.155 93.220 156.635 ;
        RECT 93.420 156.545 93.590 157.305 ;
        RECT 94.490 157.135 94.670 157.545 ;
        RECT 93.760 156.965 94.090 157.085 ;
        RECT 94.840 156.965 95.010 157.725 ;
        RECT 93.760 156.795 95.010 156.965 ;
        RECT 95.180 157.905 96.550 158.155 ;
        RECT 95.180 157.135 95.370 157.905 ;
        RECT 96.300 157.645 96.550 157.905 ;
        RECT 95.540 157.475 95.790 157.635 ;
        RECT 96.720 157.475 96.890 158.320 ;
        RECT 97.785 158.035 97.955 158.535 ;
        RECT 98.125 158.205 98.455 158.705 ;
        RECT 97.060 157.645 97.560 158.025 ;
        RECT 97.785 157.865 98.480 158.035 ;
        RECT 95.540 157.305 96.890 157.475 ;
        RECT 96.470 157.265 96.890 157.305 ;
        RECT 95.180 156.795 95.600 157.135 ;
        RECT 95.890 156.805 96.300 157.135 ;
        RECT 93.420 156.375 94.270 156.545 ;
        RECT 94.830 156.155 95.150 156.615 ;
        RECT 95.350 156.365 95.600 156.795 ;
        RECT 95.890 156.155 96.300 156.595 ;
        RECT 96.470 156.535 96.640 157.265 ;
        RECT 96.810 156.715 97.160 157.085 ;
        RECT 97.340 156.775 97.560 157.645 ;
        RECT 97.730 157.075 98.140 157.695 ;
        RECT 98.310 156.895 98.480 157.865 ;
        RECT 97.785 156.705 98.480 156.895 ;
        RECT 96.470 156.335 97.485 156.535 ;
        RECT 97.785 156.375 97.955 156.705 ;
        RECT 98.125 156.155 98.455 156.535 ;
        RECT 98.670 156.415 98.895 158.535 ;
        RECT 99.065 158.205 99.395 158.705 ;
        RECT 99.565 158.035 99.735 158.535 ;
        RECT 99.070 157.865 99.735 158.035 ;
        RECT 99.070 156.875 99.300 157.865 ;
        RECT 99.470 157.045 99.820 157.695 ;
        RECT 99.995 157.630 100.265 158.535 ;
        RECT 100.435 157.945 100.765 158.705 ;
        RECT 100.945 157.775 101.115 158.535 ;
        RECT 101.435 157.870 101.690 158.705 ;
        RECT 99.070 156.705 99.735 156.875 ;
        RECT 99.065 156.155 99.395 156.535 ;
        RECT 99.565 156.415 99.735 156.705 ;
        RECT 99.995 156.830 100.165 157.630 ;
        RECT 100.450 157.605 101.115 157.775 ;
        RECT 101.860 157.700 102.120 158.505 ;
        RECT 102.290 157.870 102.550 158.705 ;
        RECT 102.720 157.700 102.975 158.505 ;
        RECT 100.450 157.460 100.620 157.605 ;
        RECT 100.335 157.130 100.620 157.460 ;
        RECT 101.375 157.530 102.975 157.700 ;
        RECT 103.215 157.540 103.505 158.705 ;
        RECT 103.735 157.565 103.945 158.705 ;
        RECT 104.115 157.555 104.445 158.535 ;
        RECT 104.615 157.565 104.845 158.705 ;
        RECT 105.515 157.615 107.185 158.705 ;
        RECT 107.360 158.270 112.705 158.705 ;
        RECT 112.880 158.270 118.225 158.705 ;
        RECT 100.450 156.875 100.620 157.130 ;
        RECT 100.855 157.055 101.185 157.425 ;
        RECT 101.375 156.965 101.655 157.530 ;
        RECT 101.825 157.135 103.045 157.360 ;
        RECT 99.995 156.325 100.255 156.830 ;
        RECT 100.450 156.705 101.115 156.875 ;
        RECT 101.375 156.795 102.105 156.965 ;
        RECT 100.435 156.155 100.765 156.535 ;
        RECT 100.945 156.325 101.115 156.705 ;
        RECT 101.380 156.155 101.710 156.625 ;
        RECT 101.880 156.350 102.105 156.795 ;
        RECT 102.275 156.155 102.570 156.680 ;
        RECT 103.215 156.155 103.505 156.880 ;
        RECT 103.735 156.155 103.945 156.975 ;
        RECT 104.115 156.955 104.365 157.555 ;
        RECT 104.535 157.145 104.865 157.395 ;
        RECT 105.515 157.095 106.265 157.615 ;
        RECT 104.115 156.325 104.445 156.955 ;
        RECT 104.615 156.155 104.845 156.975 ;
        RECT 106.435 156.925 107.185 157.445 ;
        RECT 108.950 157.020 109.300 158.270 ;
        RECT 105.515 156.155 107.185 156.925 ;
        RECT 110.780 156.700 111.120 157.530 ;
        RECT 114.470 157.020 114.820 158.270 ;
        RECT 118.435 157.565 118.665 158.705 ;
        RECT 118.835 157.555 119.165 158.535 ;
        RECT 119.335 157.565 119.545 158.705 ;
        RECT 119.815 157.565 120.045 158.705 ;
        RECT 120.215 157.555 120.545 158.535 ;
        RECT 120.715 157.565 120.925 158.705 ;
        RECT 121.155 157.615 122.365 158.705 ;
        RECT 122.540 158.270 127.885 158.705 ;
        RECT 116.300 156.700 116.640 157.530 ;
        RECT 118.415 157.145 118.745 157.395 ;
        RECT 107.360 156.155 112.705 156.700 ;
        RECT 112.880 156.155 118.225 156.700 ;
        RECT 118.435 156.155 118.665 156.975 ;
        RECT 118.915 156.955 119.165 157.555 ;
        RECT 119.795 157.145 120.125 157.395 ;
        RECT 118.835 156.325 119.165 156.955 ;
        RECT 119.335 156.155 119.545 156.975 ;
        RECT 119.815 156.155 120.045 156.975 ;
        RECT 120.295 156.955 120.545 157.555 ;
        RECT 121.155 157.075 121.675 157.615 ;
        RECT 120.215 156.325 120.545 156.955 ;
        RECT 120.715 156.155 120.925 156.975 ;
        RECT 121.845 156.905 122.365 157.445 ;
        RECT 124.130 157.020 124.480 158.270 ;
        RECT 128.055 157.615 129.265 158.705 ;
        RECT 121.155 156.155 122.365 156.905 ;
        RECT 125.960 156.700 126.300 157.530 ;
        RECT 128.055 157.075 128.575 157.615 ;
        RECT 128.745 156.905 129.265 157.445 ;
        RECT 122.540 156.155 127.885 156.700 ;
        RECT 128.055 156.155 129.265 156.905 ;
        RECT 9.290 155.985 129.350 156.155 ;
        RECT 9.375 155.235 10.585 155.985 ;
        RECT 9.375 154.695 9.895 155.235 ;
        RECT 11.215 155.215 12.885 155.985 ;
        RECT 13.055 155.260 13.345 155.985 ;
        RECT 13.515 155.215 15.185 155.985 ;
        RECT 10.065 154.525 10.585 155.065 ;
        RECT 9.375 153.435 10.585 154.525 ;
        RECT 11.215 154.525 11.965 155.045 ;
        RECT 12.135 154.695 12.885 155.215 ;
        RECT 11.215 153.435 12.885 154.525 ;
        RECT 13.055 153.435 13.345 154.600 ;
        RECT 13.515 154.525 14.265 155.045 ;
        RECT 14.435 154.695 15.185 155.215 ;
        RECT 15.415 155.165 15.625 155.985 ;
        RECT 15.795 155.185 16.125 155.815 ;
        RECT 15.795 154.585 16.045 155.185 ;
        RECT 16.295 155.165 16.525 155.985 ;
        RECT 16.735 155.215 18.405 155.985 ;
        RECT 16.215 154.745 16.545 154.995 ;
        RECT 13.515 153.435 15.185 154.525 ;
        RECT 15.415 153.435 15.625 154.575 ;
        RECT 15.795 153.605 16.125 154.585 ;
        RECT 16.295 153.435 16.525 154.575 ;
        RECT 16.735 154.525 17.485 155.045 ;
        RECT 17.655 154.695 18.405 155.215 ;
        RECT 18.575 155.310 18.835 155.815 ;
        RECT 19.015 155.605 19.345 155.985 ;
        RECT 19.525 155.435 19.695 155.815 ;
        RECT 16.735 153.435 18.405 154.525 ;
        RECT 18.575 154.510 18.745 155.310 ;
        RECT 19.030 155.265 19.695 155.435 ;
        RECT 19.030 155.010 19.200 155.265 ;
        RECT 19.955 155.215 22.545 155.985 ;
        RECT 23.090 155.645 23.345 155.805 ;
        RECT 23.005 155.475 23.345 155.645 ;
        RECT 23.525 155.525 23.810 155.985 ;
        RECT 18.915 154.680 19.200 155.010 ;
        RECT 19.435 154.715 19.765 155.085 ;
        RECT 19.030 154.535 19.200 154.680 ;
        RECT 18.575 153.605 18.845 154.510 ;
        RECT 19.030 154.365 19.695 154.535 ;
        RECT 19.015 153.435 19.345 154.195 ;
        RECT 19.525 153.605 19.695 154.365 ;
        RECT 19.955 154.525 21.165 155.045 ;
        RECT 21.335 154.695 22.545 155.215 ;
        RECT 23.090 155.275 23.345 155.475 ;
        RECT 19.955 153.435 22.545 154.525 ;
        RECT 23.090 154.415 23.270 155.275 ;
        RECT 23.990 155.075 24.240 155.725 ;
        RECT 23.440 154.745 24.240 155.075 ;
        RECT 23.090 153.745 23.345 154.415 ;
        RECT 23.525 153.435 23.810 154.235 ;
        RECT 23.990 154.155 24.240 154.745 ;
        RECT 24.440 155.390 24.760 155.720 ;
        RECT 24.940 155.505 25.600 155.985 ;
        RECT 25.800 155.595 26.650 155.765 ;
        RECT 24.440 154.495 24.630 155.390 ;
        RECT 24.950 155.065 25.610 155.335 ;
        RECT 25.280 155.005 25.610 155.065 ;
        RECT 24.800 154.835 25.130 154.895 ;
        RECT 25.800 154.835 25.970 155.595 ;
        RECT 27.210 155.525 27.530 155.985 ;
        RECT 27.730 155.345 27.980 155.775 ;
        RECT 28.270 155.545 28.680 155.985 ;
        RECT 28.850 155.605 29.865 155.805 ;
        RECT 26.140 155.175 27.390 155.345 ;
        RECT 26.140 155.055 26.470 155.175 ;
        RECT 24.800 154.665 26.700 154.835 ;
        RECT 24.440 154.325 26.360 154.495 ;
        RECT 24.440 154.305 24.760 154.325 ;
        RECT 23.990 153.645 24.320 154.155 ;
        RECT 24.590 153.695 24.760 154.305 ;
        RECT 26.530 154.155 26.700 154.665 ;
        RECT 26.870 154.595 27.050 155.005 ;
        RECT 27.220 154.415 27.390 155.175 ;
        RECT 24.930 153.435 25.260 154.125 ;
        RECT 25.490 153.985 26.700 154.155 ;
        RECT 26.870 154.105 27.390 154.415 ;
        RECT 27.560 155.005 27.980 155.345 ;
        RECT 28.270 155.005 28.680 155.335 ;
        RECT 27.560 154.235 27.750 155.005 ;
        RECT 28.850 154.875 29.020 155.605 ;
        RECT 30.165 155.435 30.335 155.765 ;
        RECT 30.505 155.605 30.835 155.985 ;
        RECT 29.190 155.055 29.540 155.425 ;
        RECT 28.850 154.835 29.270 154.875 ;
        RECT 27.920 154.665 29.270 154.835 ;
        RECT 27.920 154.505 28.170 154.665 ;
        RECT 28.680 154.235 28.930 154.495 ;
        RECT 27.560 153.985 28.930 154.235 ;
        RECT 25.490 153.695 25.730 153.985 ;
        RECT 26.530 153.905 26.700 153.985 ;
        RECT 25.930 153.435 26.350 153.815 ;
        RECT 26.530 153.655 27.160 153.905 ;
        RECT 27.630 153.435 27.960 153.815 ;
        RECT 28.130 153.695 28.300 153.985 ;
        RECT 29.100 153.820 29.270 154.665 ;
        RECT 29.720 154.495 29.940 155.365 ;
        RECT 30.165 155.245 30.860 155.435 ;
        RECT 29.440 154.115 29.940 154.495 ;
        RECT 30.110 154.445 30.520 155.065 ;
        RECT 30.690 154.275 30.860 155.245 ;
        RECT 30.165 154.105 30.860 154.275 ;
        RECT 28.480 153.435 28.860 153.815 ;
        RECT 29.100 153.650 29.930 153.820 ;
        RECT 30.165 153.605 30.335 154.105 ;
        RECT 30.505 153.435 30.835 153.935 ;
        RECT 31.050 153.605 31.275 155.725 ;
        RECT 31.445 155.605 31.775 155.985 ;
        RECT 31.945 155.435 32.115 155.725 ;
        RECT 31.450 155.265 32.115 155.435 ;
        RECT 31.450 154.275 31.680 155.265 ;
        RECT 32.835 155.215 34.505 155.985 ;
        RECT 31.850 154.445 32.200 155.095 ;
        RECT 32.835 154.525 33.585 155.045 ;
        RECT 33.755 154.695 34.505 155.215 ;
        RECT 34.675 155.185 35.015 155.815 ;
        RECT 35.185 155.185 35.435 155.985 ;
        RECT 35.625 155.335 35.955 155.815 ;
        RECT 36.125 155.525 36.350 155.985 ;
        RECT 36.520 155.335 36.850 155.815 ;
        RECT 34.675 154.575 34.850 155.185 ;
        RECT 35.625 155.165 36.850 155.335 ;
        RECT 37.480 155.205 37.980 155.815 ;
        RECT 38.815 155.260 39.105 155.985 ;
        RECT 39.740 155.440 45.085 155.985 ;
        RECT 35.020 154.825 35.715 154.995 ;
        RECT 35.545 154.575 35.715 154.825 ;
        RECT 35.890 154.795 36.310 154.995 ;
        RECT 36.480 154.795 36.810 154.995 ;
        RECT 36.980 154.795 37.310 154.995 ;
        RECT 37.480 154.575 37.650 155.205 ;
        RECT 37.835 154.745 38.185 154.995 ;
        RECT 31.450 154.105 32.115 154.275 ;
        RECT 31.445 153.435 31.775 153.935 ;
        RECT 31.945 153.605 32.115 154.105 ;
        RECT 32.835 153.435 34.505 154.525 ;
        RECT 34.675 153.605 35.015 154.575 ;
        RECT 35.185 153.435 35.355 154.575 ;
        RECT 35.545 154.405 37.980 154.575 ;
        RECT 35.625 153.435 35.875 154.235 ;
        RECT 36.520 153.605 36.850 154.405 ;
        RECT 37.150 153.435 37.480 154.235 ;
        RECT 37.650 153.605 37.980 154.405 ;
        RECT 38.815 153.435 39.105 154.600 ;
        RECT 41.330 153.870 41.680 155.120 ;
        RECT 43.160 154.610 43.500 155.440 ;
        RECT 45.255 155.185 45.595 155.815 ;
        RECT 45.765 155.185 46.015 155.985 ;
        RECT 46.205 155.335 46.535 155.815 ;
        RECT 46.705 155.525 46.930 155.985 ;
        RECT 47.100 155.335 47.430 155.815 ;
        RECT 45.255 154.575 45.430 155.185 ;
        RECT 46.205 155.165 47.430 155.335 ;
        RECT 48.060 155.205 48.560 155.815 ;
        RECT 49.395 155.215 51.985 155.985 ;
        RECT 45.600 154.825 46.295 154.995 ;
        RECT 46.125 154.575 46.295 154.825 ;
        RECT 46.470 154.795 46.890 154.995 ;
        RECT 47.060 154.795 47.390 154.995 ;
        RECT 47.560 154.795 47.890 154.995 ;
        RECT 48.060 154.575 48.230 155.205 ;
        RECT 48.415 154.745 48.765 154.995 ;
        RECT 39.740 153.435 45.085 153.870 ;
        RECT 45.255 153.605 45.595 154.575 ;
        RECT 45.765 153.435 45.935 154.575 ;
        RECT 46.125 154.405 48.560 154.575 ;
        RECT 46.205 153.435 46.455 154.235 ;
        RECT 47.100 153.605 47.430 154.405 ;
        RECT 47.730 153.435 48.060 154.235 ;
        RECT 48.230 153.605 48.560 154.405 ;
        RECT 49.395 154.525 50.605 155.045 ;
        RECT 50.775 154.695 51.985 155.215 ;
        RECT 52.530 155.275 52.785 155.805 ;
        RECT 52.965 155.525 53.250 155.985 ;
        RECT 49.395 153.435 51.985 154.525 ;
        RECT 52.530 154.415 52.710 155.275 ;
        RECT 53.430 155.075 53.680 155.725 ;
        RECT 52.880 154.745 53.680 155.075 ;
        RECT 52.530 153.945 52.785 154.415 ;
        RECT 52.445 153.775 52.785 153.945 ;
        RECT 52.530 153.745 52.785 153.775 ;
        RECT 52.965 153.435 53.250 154.235 ;
        RECT 53.430 154.155 53.680 154.745 ;
        RECT 53.880 155.390 54.200 155.720 ;
        RECT 54.380 155.505 55.040 155.985 ;
        RECT 55.240 155.595 56.090 155.765 ;
        RECT 53.880 154.495 54.070 155.390 ;
        RECT 54.390 155.065 55.050 155.335 ;
        RECT 54.720 155.005 55.050 155.065 ;
        RECT 54.240 154.835 54.570 154.895 ;
        RECT 55.240 154.835 55.410 155.595 ;
        RECT 56.650 155.525 56.970 155.985 ;
        RECT 57.170 155.345 57.420 155.775 ;
        RECT 57.710 155.545 58.120 155.985 ;
        RECT 58.290 155.605 59.305 155.805 ;
        RECT 55.580 155.175 56.830 155.345 ;
        RECT 55.580 155.055 55.910 155.175 ;
        RECT 54.240 154.665 56.140 154.835 ;
        RECT 53.880 154.325 55.800 154.495 ;
        RECT 53.880 154.305 54.200 154.325 ;
        RECT 53.430 153.645 53.760 154.155 ;
        RECT 54.030 153.695 54.200 154.305 ;
        RECT 55.970 154.155 56.140 154.665 ;
        RECT 56.310 154.595 56.490 155.005 ;
        RECT 56.660 154.415 56.830 155.175 ;
        RECT 54.370 153.435 54.700 154.125 ;
        RECT 54.930 153.985 56.140 154.155 ;
        RECT 56.310 154.105 56.830 154.415 ;
        RECT 57.000 155.005 57.420 155.345 ;
        RECT 57.710 155.005 58.120 155.335 ;
        RECT 57.000 154.235 57.190 155.005 ;
        RECT 58.290 154.875 58.460 155.605 ;
        RECT 59.605 155.435 59.775 155.765 ;
        RECT 59.945 155.605 60.275 155.985 ;
        RECT 58.630 155.055 58.980 155.425 ;
        RECT 58.290 154.835 58.710 154.875 ;
        RECT 57.360 154.665 58.710 154.835 ;
        RECT 57.360 154.505 57.610 154.665 ;
        RECT 58.120 154.235 58.370 154.495 ;
        RECT 57.000 153.985 58.370 154.235 ;
        RECT 54.930 153.695 55.170 153.985 ;
        RECT 55.970 153.905 56.140 153.985 ;
        RECT 55.370 153.435 55.790 153.815 ;
        RECT 55.970 153.655 56.600 153.905 ;
        RECT 57.070 153.435 57.400 153.815 ;
        RECT 57.570 153.695 57.740 153.985 ;
        RECT 58.540 153.820 58.710 154.665 ;
        RECT 59.160 154.495 59.380 155.365 ;
        RECT 59.605 155.245 60.300 155.435 ;
        RECT 58.880 154.115 59.380 154.495 ;
        RECT 59.550 154.445 59.960 155.065 ;
        RECT 60.130 154.275 60.300 155.245 ;
        RECT 59.605 154.105 60.300 154.275 ;
        RECT 57.920 153.435 58.300 153.815 ;
        RECT 58.540 153.650 59.370 153.820 ;
        RECT 59.605 153.605 59.775 154.105 ;
        RECT 59.945 153.435 60.275 153.935 ;
        RECT 60.490 153.605 60.715 155.725 ;
        RECT 60.885 155.605 61.215 155.985 ;
        RECT 61.385 155.435 61.555 155.725 ;
        RECT 60.890 155.265 61.555 155.435 ;
        RECT 60.890 154.275 61.120 155.265 ;
        RECT 61.855 155.165 62.085 155.985 ;
        RECT 62.255 155.185 62.585 155.815 ;
        RECT 61.290 154.445 61.640 155.095 ;
        RECT 61.835 154.745 62.165 154.995 ;
        RECT 62.335 154.585 62.585 155.185 ;
        RECT 62.755 155.165 62.965 155.985 ;
        RECT 63.195 155.235 64.405 155.985 ;
        RECT 64.575 155.260 64.865 155.985 ;
        RECT 60.890 154.105 61.555 154.275 ;
        RECT 60.885 153.435 61.215 153.935 ;
        RECT 61.385 153.605 61.555 154.105 ;
        RECT 61.855 153.435 62.085 154.575 ;
        RECT 62.255 153.605 62.585 154.585 ;
        RECT 62.755 153.435 62.965 154.575 ;
        RECT 63.195 154.525 63.715 155.065 ;
        RECT 63.885 154.695 64.405 155.235 ;
        RECT 65.035 155.215 66.705 155.985 ;
        RECT 63.195 153.435 64.405 154.525 ;
        RECT 64.575 153.435 64.865 154.600 ;
        RECT 65.035 154.525 65.785 155.045 ;
        RECT 65.955 154.695 66.705 155.215 ;
        RECT 66.880 155.145 67.140 155.985 ;
        RECT 67.315 155.240 67.570 155.815 ;
        RECT 67.740 155.605 68.070 155.985 ;
        RECT 68.285 155.435 68.455 155.815 ;
        RECT 67.740 155.265 68.455 155.435 ;
        RECT 65.035 153.435 66.705 154.525 ;
        RECT 66.880 153.435 67.140 154.585 ;
        RECT 67.315 154.510 67.485 155.240 ;
        RECT 67.740 155.075 67.910 155.265 ;
        RECT 68.720 155.145 68.980 155.985 ;
        RECT 69.155 155.240 69.410 155.815 ;
        RECT 69.580 155.605 69.910 155.985 ;
        RECT 70.125 155.435 70.295 155.815 ;
        RECT 71.480 155.440 76.825 155.985 ;
        RECT 69.580 155.265 70.295 155.435 ;
        RECT 67.655 154.745 67.910 155.075 ;
        RECT 67.740 154.535 67.910 154.745 ;
        RECT 68.190 154.715 68.545 155.085 ;
        RECT 67.315 153.605 67.570 154.510 ;
        RECT 67.740 154.365 68.455 154.535 ;
        RECT 67.740 153.435 68.070 154.195 ;
        RECT 68.285 153.605 68.455 154.365 ;
        RECT 68.720 153.435 68.980 154.585 ;
        RECT 69.155 154.510 69.325 155.240 ;
        RECT 69.580 155.075 69.750 155.265 ;
        RECT 69.495 154.745 69.750 155.075 ;
        RECT 69.580 154.535 69.750 154.745 ;
        RECT 70.030 154.715 70.385 155.085 ;
        RECT 69.155 153.605 69.410 154.510 ;
        RECT 69.580 154.365 70.295 154.535 ;
        RECT 69.580 153.435 69.910 154.195 ;
        RECT 70.125 153.605 70.295 154.365 ;
        RECT 73.070 153.870 73.420 155.120 ;
        RECT 74.900 154.610 75.240 155.440 ;
        RECT 76.995 155.185 77.335 155.815 ;
        RECT 77.505 155.185 77.755 155.985 ;
        RECT 77.945 155.335 78.275 155.815 ;
        RECT 78.445 155.525 78.670 155.985 ;
        RECT 78.840 155.335 79.170 155.815 ;
        RECT 76.995 154.575 77.170 155.185 ;
        RECT 77.945 155.165 79.170 155.335 ;
        RECT 79.800 155.205 80.300 155.815 ;
        RECT 77.340 154.825 78.035 154.995 ;
        RECT 77.865 154.575 78.035 154.825 ;
        RECT 78.210 154.795 78.630 154.995 ;
        RECT 78.800 154.795 79.130 154.995 ;
        RECT 79.300 154.795 79.630 154.995 ;
        RECT 79.800 154.575 79.970 155.205 ;
        RECT 81.870 155.175 82.115 155.780 ;
        RECT 82.335 155.450 82.845 155.985 ;
        RECT 81.595 155.005 82.825 155.175 ;
        RECT 80.155 154.745 80.505 154.995 ;
        RECT 71.480 153.435 76.825 153.870 ;
        RECT 76.995 153.605 77.335 154.575 ;
        RECT 77.505 153.435 77.675 154.575 ;
        RECT 77.865 154.405 80.300 154.575 ;
        RECT 77.945 153.435 78.195 154.235 ;
        RECT 78.840 153.605 79.170 154.405 ;
        RECT 79.470 153.435 79.800 154.235 ;
        RECT 79.970 153.605 80.300 154.405 ;
        RECT 81.595 154.195 81.935 155.005 ;
        RECT 82.105 154.440 82.855 154.630 ;
        RECT 81.595 153.785 82.110 154.195 ;
        RECT 82.345 153.435 82.515 154.195 ;
        RECT 82.685 153.775 82.855 154.440 ;
        RECT 83.025 154.455 83.215 155.815 ;
        RECT 83.385 154.965 83.660 155.815 ;
        RECT 83.850 155.450 84.380 155.815 ;
        RECT 84.805 155.585 85.135 155.985 ;
        RECT 84.205 155.415 84.380 155.450 ;
        RECT 83.385 154.795 83.665 154.965 ;
        RECT 83.385 154.655 83.660 154.795 ;
        RECT 83.865 154.455 84.035 155.255 ;
        RECT 83.025 154.285 84.035 154.455 ;
        RECT 84.205 155.245 85.135 155.415 ;
        RECT 85.305 155.245 85.560 155.815 ;
        RECT 84.205 154.115 84.375 155.245 ;
        RECT 84.965 155.075 85.135 155.245 ;
        RECT 83.250 153.945 84.375 154.115 ;
        RECT 84.545 154.745 84.740 155.075 ;
        RECT 84.965 154.745 85.220 155.075 ;
        RECT 84.545 153.775 84.715 154.745 ;
        RECT 85.390 154.575 85.560 155.245 ;
        RECT 86.655 155.215 90.165 155.985 ;
        RECT 90.335 155.260 90.625 155.985 ;
        RECT 91.255 155.215 93.845 155.985 ;
        RECT 82.685 153.605 84.715 153.775 ;
        RECT 84.885 153.435 85.055 154.575 ;
        RECT 85.225 153.605 85.560 154.575 ;
        RECT 86.655 154.525 88.345 155.045 ;
        RECT 88.515 154.695 90.165 155.215 ;
        RECT 86.655 153.435 90.165 154.525 ;
        RECT 90.335 153.435 90.625 154.600 ;
        RECT 91.255 154.525 92.465 155.045 ;
        RECT 92.635 154.695 93.845 155.215 ;
        RECT 94.290 155.175 94.535 155.780 ;
        RECT 94.755 155.450 95.265 155.985 ;
        RECT 94.015 155.005 95.245 155.175 ;
        RECT 91.255 153.435 93.845 154.525 ;
        RECT 94.015 154.195 94.355 155.005 ;
        RECT 94.525 154.440 95.275 154.630 ;
        RECT 94.015 153.785 94.530 154.195 ;
        RECT 94.765 153.435 94.935 154.195 ;
        RECT 95.105 153.775 95.275 154.440 ;
        RECT 95.445 154.455 95.635 155.815 ;
        RECT 95.805 154.965 96.080 155.815 ;
        RECT 96.270 155.450 96.800 155.815 ;
        RECT 97.225 155.585 97.555 155.985 ;
        RECT 96.625 155.415 96.800 155.450 ;
        RECT 95.805 154.795 96.085 154.965 ;
        RECT 95.805 154.655 96.080 154.795 ;
        RECT 96.285 154.455 96.455 155.255 ;
        RECT 95.445 154.285 96.455 154.455 ;
        RECT 96.625 155.245 97.555 155.415 ;
        RECT 97.725 155.245 97.980 155.815 ;
        RECT 96.625 154.115 96.795 155.245 ;
        RECT 97.385 155.075 97.555 155.245 ;
        RECT 95.670 153.945 96.795 154.115 ;
        RECT 96.965 154.745 97.160 155.075 ;
        RECT 97.385 154.745 97.640 155.075 ;
        RECT 96.965 153.775 97.135 154.745 ;
        RECT 97.810 154.575 97.980 155.245 ;
        RECT 99.075 155.215 102.585 155.985 ;
        RECT 102.760 155.440 108.105 155.985 ;
        RECT 95.105 153.605 97.135 153.775 ;
        RECT 97.305 153.435 97.475 154.575 ;
        RECT 97.645 153.605 97.980 154.575 ;
        RECT 99.075 154.525 100.765 155.045 ;
        RECT 100.935 154.695 102.585 155.215 ;
        RECT 99.075 153.435 102.585 154.525 ;
        RECT 104.350 153.870 104.700 155.120 ;
        RECT 106.180 154.610 106.520 155.440 ;
        RECT 108.275 155.185 108.615 155.815 ;
        RECT 108.785 155.185 109.035 155.985 ;
        RECT 109.225 155.335 109.555 155.815 ;
        RECT 109.725 155.525 109.950 155.985 ;
        RECT 110.120 155.335 110.450 155.815 ;
        RECT 108.275 154.575 108.450 155.185 ;
        RECT 109.225 155.165 110.450 155.335 ;
        RECT 111.080 155.205 111.580 155.815 ;
        RECT 111.955 155.235 113.165 155.985 ;
        RECT 108.620 154.825 109.315 154.995 ;
        RECT 109.145 154.575 109.315 154.825 ;
        RECT 109.490 154.795 109.910 154.995 ;
        RECT 110.080 154.795 110.410 154.995 ;
        RECT 110.580 154.795 110.910 154.995 ;
        RECT 111.080 154.575 111.250 155.205 ;
        RECT 111.435 154.745 111.785 154.995 ;
        RECT 102.760 153.435 108.105 153.870 ;
        RECT 108.275 153.605 108.615 154.575 ;
        RECT 108.785 153.435 108.955 154.575 ;
        RECT 109.145 154.405 111.580 154.575 ;
        RECT 109.225 153.435 109.475 154.235 ;
        RECT 110.120 153.605 110.450 154.405 ;
        RECT 110.750 153.435 111.080 154.235 ;
        RECT 111.250 153.605 111.580 154.405 ;
        RECT 111.955 154.525 112.475 155.065 ;
        RECT 112.645 154.695 113.165 155.235 ;
        RECT 113.425 155.335 113.595 155.815 ;
        RECT 113.775 155.505 114.015 155.985 ;
        RECT 114.265 155.335 114.435 155.815 ;
        RECT 114.605 155.505 114.935 155.985 ;
        RECT 115.105 155.335 115.275 155.815 ;
        RECT 113.425 155.165 114.060 155.335 ;
        RECT 114.265 155.165 115.275 155.335 ;
        RECT 115.445 155.185 115.775 155.985 ;
        RECT 116.095 155.260 116.385 155.985 ;
        RECT 117.020 155.275 117.275 155.805 ;
        RECT 117.445 155.525 117.750 155.985 ;
        RECT 117.995 155.605 119.065 155.775 ;
        RECT 113.890 154.995 114.060 155.165 ;
        RECT 114.775 155.135 115.275 155.165 ;
        RECT 113.340 154.755 113.720 154.995 ;
        RECT 113.890 154.825 114.390 154.995 ;
        RECT 113.890 154.585 114.060 154.825 ;
        RECT 114.780 154.625 115.275 155.135 ;
        RECT 111.955 153.435 113.165 154.525 ;
        RECT 113.345 154.415 114.060 154.585 ;
        RECT 114.265 154.455 115.275 154.625 ;
        RECT 117.020 154.625 117.230 155.275 ;
        RECT 117.995 155.250 118.315 155.605 ;
        RECT 117.990 155.075 118.315 155.250 ;
        RECT 117.400 154.775 118.315 155.075 ;
        RECT 118.485 155.035 118.725 155.435 ;
        RECT 118.895 155.375 119.065 155.605 ;
        RECT 119.235 155.545 119.425 155.985 ;
        RECT 119.595 155.535 120.545 155.815 ;
        RECT 120.765 155.625 121.115 155.795 ;
        RECT 118.895 155.205 119.425 155.375 ;
        RECT 117.400 154.745 118.140 154.775 ;
        RECT 113.345 153.605 113.675 154.415 ;
        RECT 113.845 153.435 114.085 154.235 ;
        RECT 114.265 153.605 114.435 154.455 ;
        RECT 114.605 153.435 114.935 154.235 ;
        RECT 115.105 153.605 115.275 154.455 ;
        RECT 115.445 153.435 115.775 154.585 ;
        RECT 116.095 153.435 116.385 154.600 ;
        RECT 117.020 153.745 117.275 154.625 ;
        RECT 117.445 153.435 117.750 154.575 ;
        RECT 117.970 154.155 118.140 154.745 ;
        RECT 118.485 154.665 119.025 155.035 ;
        RECT 119.205 154.925 119.425 155.205 ;
        RECT 119.595 154.755 119.765 155.535 ;
        RECT 119.360 154.585 119.765 154.755 ;
        RECT 119.935 154.745 120.285 155.365 ;
        RECT 119.360 154.495 119.530 154.585 ;
        RECT 120.455 154.575 120.665 155.365 ;
        RECT 118.310 154.325 119.530 154.495 ;
        RECT 119.990 154.415 120.665 154.575 ;
        RECT 117.970 153.985 118.770 154.155 ;
        RECT 118.090 153.435 118.420 153.815 ;
        RECT 118.600 153.695 118.770 153.985 ;
        RECT 119.360 153.945 119.530 154.325 ;
        RECT 119.700 154.405 120.665 154.415 ;
        RECT 120.855 155.235 121.115 155.625 ;
        RECT 121.325 155.525 121.655 155.985 ;
        RECT 122.530 155.595 123.385 155.765 ;
        RECT 123.590 155.595 124.085 155.765 ;
        RECT 124.255 155.625 124.585 155.985 ;
        RECT 120.855 154.545 121.025 155.235 ;
        RECT 121.195 154.885 121.365 155.065 ;
        RECT 121.535 155.055 122.325 155.305 ;
        RECT 122.530 154.885 122.700 155.595 ;
        RECT 122.870 155.085 123.225 155.305 ;
        RECT 121.195 154.715 122.885 154.885 ;
        RECT 119.700 154.115 120.160 154.405 ;
        RECT 120.855 154.375 122.355 154.545 ;
        RECT 120.855 154.235 121.025 154.375 ;
        RECT 120.465 154.065 121.025 154.235 ;
        RECT 118.940 153.435 119.190 153.895 ;
        RECT 119.360 153.605 120.230 153.945 ;
        RECT 120.465 153.605 120.635 154.065 ;
        RECT 121.470 154.035 122.545 154.205 ;
        RECT 120.805 153.435 121.175 153.895 ;
        RECT 121.470 153.695 121.640 154.035 ;
        RECT 121.810 153.435 122.140 153.865 ;
        RECT 122.375 153.695 122.545 154.035 ;
        RECT 122.715 153.935 122.885 154.715 ;
        RECT 123.055 154.495 123.225 155.085 ;
        RECT 123.395 154.685 123.745 155.305 ;
        RECT 123.055 154.105 123.520 154.495 ;
        RECT 123.915 154.235 124.085 155.595 ;
        RECT 124.255 154.405 124.715 155.455 ;
        RECT 123.690 154.065 124.085 154.235 ;
        RECT 123.690 153.935 123.860 154.065 ;
        RECT 122.715 153.605 123.395 153.935 ;
        RECT 123.610 153.605 123.860 153.935 ;
        RECT 124.030 153.435 124.280 153.895 ;
        RECT 124.450 153.620 124.775 154.405 ;
        RECT 124.945 153.605 125.115 155.725 ;
        RECT 125.285 155.605 125.615 155.985 ;
        RECT 125.785 155.435 126.040 155.725 ;
        RECT 125.290 155.265 126.040 155.435 ;
        RECT 125.290 154.275 125.520 155.265 ;
        RECT 126.215 155.215 127.885 155.985 ;
        RECT 128.055 155.235 129.265 155.985 ;
        RECT 125.690 154.445 126.040 155.095 ;
        RECT 126.215 154.525 126.965 155.045 ;
        RECT 127.135 154.695 127.885 155.215 ;
        RECT 128.055 154.525 128.575 155.065 ;
        RECT 128.745 154.695 129.265 155.235 ;
        RECT 125.290 154.105 126.040 154.275 ;
        RECT 125.285 153.435 125.615 153.935 ;
        RECT 125.785 153.605 126.040 154.105 ;
        RECT 126.215 153.435 127.885 154.525 ;
        RECT 128.055 153.435 129.265 154.525 ;
        RECT 9.290 153.265 129.350 153.435 ;
        RECT 9.375 152.175 10.585 153.265 ;
        RECT 10.760 152.830 16.105 153.265 ;
        RECT 9.375 151.465 9.895 152.005 ;
        RECT 10.065 151.635 10.585 152.175 ;
        RECT 12.350 151.580 12.700 152.830 ;
        RECT 16.275 152.505 16.790 152.915 ;
        RECT 17.025 152.505 17.195 153.265 ;
        RECT 17.365 152.925 19.395 153.095 ;
        RECT 9.375 150.715 10.585 151.465 ;
        RECT 14.180 151.260 14.520 152.090 ;
        RECT 16.275 151.695 16.615 152.505 ;
        RECT 17.365 152.260 17.535 152.925 ;
        RECT 17.930 152.585 19.055 152.755 ;
        RECT 16.785 152.070 17.535 152.260 ;
        RECT 17.705 152.245 18.715 152.415 ;
        RECT 16.275 151.525 17.505 151.695 ;
        RECT 10.760 150.715 16.105 151.260 ;
        RECT 16.550 150.920 16.795 151.525 ;
        RECT 17.015 150.715 17.525 151.250 ;
        RECT 17.705 150.885 17.895 152.245 ;
        RECT 18.065 151.225 18.340 152.045 ;
        RECT 18.545 151.445 18.715 152.245 ;
        RECT 18.885 151.455 19.055 152.585 ;
        RECT 19.225 151.955 19.395 152.925 ;
        RECT 19.565 152.125 19.735 153.265 ;
        RECT 19.905 152.125 20.240 153.095 ;
        RECT 20.420 152.830 25.765 153.265 ;
        RECT 19.225 151.625 19.420 151.955 ;
        RECT 19.645 151.625 19.900 151.955 ;
        RECT 19.645 151.455 19.815 151.625 ;
        RECT 20.070 151.455 20.240 152.125 ;
        RECT 22.010 151.580 22.360 152.830 ;
        RECT 25.935 152.100 26.225 153.265 ;
        RECT 26.855 152.175 29.445 153.265 ;
        RECT 29.705 152.335 29.875 153.095 ;
        RECT 30.055 152.505 30.385 153.265 ;
        RECT 18.885 151.285 19.815 151.455 ;
        RECT 18.885 151.250 19.060 151.285 ;
        RECT 18.065 151.055 18.345 151.225 ;
        RECT 18.065 150.885 18.340 151.055 ;
        RECT 18.530 150.885 19.060 151.250 ;
        RECT 19.485 150.715 19.815 151.115 ;
        RECT 19.985 150.885 20.240 151.455 ;
        RECT 23.840 151.260 24.180 152.090 ;
        RECT 26.855 151.655 28.065 152.175 ;
        RECT 29.705 152.165 30.370 152.335 ;
        RECT 30.555 152.190 30.825 153.095 ;
        RECT 30.200 152.020 30.370 152.165 ;
        RECT 28.235 151.485 29.445 152.005 ;
        RECT 29.635 151.615 29.965 151.985 ;
        RECT 30.200 151.690 30.485 152.020 ;
        RECT 20.420 150.715 25.765 151.260 ;
        RECT 25.935 150.715 26.225 151.440 ;
        RECT 26.855 150.715 29.445 151.485 ;
        RECT 30.200 151.435 30.370 151.690 ;
        RECT 29.705 151.265 30.370 151.435 ;
        RECT 30.655 151.390 30.825 152.190 ;
        RECT 31.455 152.175 34.045 153.265 ;
        RECT 34.420 152.295 34.750 153.095 ;
        RECT 34.920 152.465 35.250 153.265 ;
        RECT 35.550 152.295 35.880 153.095 ;
        RECT 36.525 152.465 36.775 153.265 ;
        RECT 31.455 151.655 32.665 152.175 ;
        RECT 34.420 152.125 36.855 152.295 ;
        RECT 37.045 152.125 37.215 153.265 ;
        RECT 37.385 152.125 37.725 153.095 ;
        RECT 38.100 152.295 38.430 153.095 ;
        RECT 38.600 152.465 38.930 153.265 ;
        RECT 39.230 152.295 39.560 153.095 ;
        RECT 40.205 152.465 40.455 153.265 ;
        RECT 38.100 152.125 40.535 152.295 ;
        RECT 40.725 152.125 40.895 153.265 ;
        RECT 41.065 152.125 41.405 153.095 ;
        RECT 42.700 152.295 43.030 153.095 ;
        RECT 43.200 152.465 43.530 153.265 ;
        RECT 43.830 152.295 44.160 153.095 ;
        RECT 44.805 152.465 45.055 153.265 ;
        RECT 42.700 152.125 45.135 152.295 ;
        RECT 45.325 152.125 45.495 153.265 ;
        RECT 45.665 152.125 46.005 153.095 ;
        RECT 46.180 152.830 51.525 153.265 ;
        RECT 32.835 151.485 34.045 152.005 ;
        RECT 34.215 151.705 34.565 151.955 ;
        RECT 34.750 151.495 34.920 152.125 ;
        RECT 35.090 151.705 35.420 151.905 ;
        RECT 35.590 151.705 35.920 151.905 ;
        RECT 36.090 151.705 36.510 151.905 ;
        RECT 36.685 151.875 36.855 152.125 ;
        RECT 36.685 151.705 37.380 151.875 ;
        RECT 29.705 150.885 29.875 151.265 ;
        RECT 30.055 150.715 30.385 151.095 ;
        RECT 30.565 150.885 30.825 151.390 ;
        RECT 31.455 150.715 34.045 151.485 ;
        RECT 34.420 150.885 34.920 151.495 ;
        RECT 35.550 151.365 36.775 151.535 ;
        RECT 37.550 151.515 37.725 152.125 ;
        RECT 37.895 151.705 38.245 151.955 ;
        RECT 35.550 150.885 35.880 151.365 ;
        RECT 36.050 150.715 36.275 151.175 ;
        RECT 36.445 150.885 36.775 151.365 ;
        RECT 36.965 150.715 37.215 151.515 ;
        RECT 37.385 150.885 37.725 151.515 ;
        RECT 38.430 151.495 38.600 152.125 ;
        RECT 38.770 151.705 39.100 151.905 ;
        RECT 39.270 151.705 39.600 151.905 ;
        RECT 39.770 151.705 40.190 151.905 ;
        RECT 40.365 151.875 40.535 152.125 ;
        RECT 40.365 151.705 41.060 151.875 ;
        RECT 38.100 150.885 38.600 151.495 ;
        RECT 39.230 151.365 40.455 151.535 ;
        RECT 41.230 151.515 41.405 152.125 ;
        RECT 42.495 151.705 42.845 151.955 ;
        RECT 39.230 150.885 39.560 151.365 ;
        RECT 39.730 150.715 39.955 151.175 ;
        RECT 40.125 150.885 40.455 151.365 ;
        RECT 40.645 150.715 40.895 151.515 ;
        RECT 41.065 150.885 41.405 151.515 ;
        RECT 43.030 151.495 43.200 152.125 ;
        RECT 43.370 151.705 43.700 151.905 ;
        RECT 43.870 151.705 44.200 151.905 ;
        RECT 44.370 151.705 44.790 151.905 ;
        RECT 44.965 151.875 45.135 152.125 ;
        RECT 44.965 151.705 45.660 151.875 ;
        RECT 42.700 150.885 43.200 151.495 ;
        RECT 43.830 151.365 45.055 151.535 ;
        RECT 45.830 151.515 46.005 152.125 ;
        RECT 47.770 151.580 48.120 152.830 ;
        RECT 51.695 152.100 51.985 153.265 ;
        RECT 52.155 152.175 53.825 153.265 ;
        RECT 53.995 152.505 54.510 152.915 ;
        RECT 54.745 152.505 54.915 153.265 ;
        RECT 55.085 152.925 57.115 153.095 ;
        RECT 43.830 150.885 44.160 151.365 ;
        RECT 44.330 150.715 44.555 151.175 ;
        RECT 44.725 150.885 45.055 151.365 ;
        RECT 45.245 150.715 45.495 151.515 ;
        RECT 45.665 150.885 46.005 151.515 ;
        RECT 49.600 151.260 49.940 152.090 ;
        RECT 52.155 151.655 52.905 152.175 ;
        RECT 53.075 151.485 53.825 152.005 ;
        RECT 53.995 151.695 54.335 152.505 ;
        RECT 55.085 152.260 55.255 152.925 ;
        RECT 55.650 152.585 56.775 152.755 ;
        RECT 54.505 152.070 55.255 152.260 ;
        RECT 55.425 152.245 56.435 152.415 ;
        RECT 53.995 151.525 55.225 151.695 ;
        RECT 46.180 150.715 51.525 151.260 ;
        RECT 51.695 150.715 51.985 151.440 ;
        RECT 52.155 150.715 53.825 151.485 ;
        RECT 54.270 150.920 54.515 151.525 ;
        RECT 54.735 150.715 55.245 151.250 ;
        RECT 55.425 150.885 55.615 152.245 ;
        RECT 55.785 151.225 56.060 152.045 ;
        RECT 56.265 151.445 56.435 152.245 ;
        RECT 56.605 151.455 56.775 152.585 ;
        RECT 56.945 151.955 57.115 152.925 ;
        RECT 57.285 152.125 57.455 153.265 ;
        RECT 57.625 152.125 57.960 153.095 ;
        RECT 58.225 152.335 58.395 153.095 ;
        RECT 58.575 152.505 58.905 153.265 ;
        RECT 58.225 152.165 58.890 152.335 ;
        RECT 59.075 152.190 59.345 153.095 ;
        RECT 56.945 151.625 57.140 151.955 ;
        RECT 57.365 151.625 57.620 151.955 ;
        RECT 57.365 151.455 57.535 151.625 ;
        RECT 57.790 151.455 57.960 152.125 ;
        RECT 58.720 152.020 58.890 152.165 ;
        RECT 58.155 151.615 58.485 151.985 ;
        RECT 58.720 151.690 59.005 152.020 ;
        RECT 56.605 151.285 57.535 151.455 ;
        RECT 56.605 151.250 56.780 151.285 ;
        RECT 55.785 151.055 56.065 151.225 ;
        RECT 55.785 150.885 56.060 151.055 ;
        RECT 56.250 150.885 56.780 151.250 ;
        RECT 57.205 150.715 57.535 151.115 ;
        RECT 57.705 150.885 57.960 151.455 ;
        RECT 58.720 151.435 58.890 151.690 ;
        RECT 58.225 151.265 58.890 151.435 ;
        RECT 59.175 151.390 59.345 152.190 ;
        RECT 59.975 152.175 62.565 153.265 ;
        RECT 62.825 152.335 62.995 153.095 ;
        RECT 63.175 152.505 63.505 153.265 ;
        RECT 59.975 151.655 61.185 152.175 ;
        RECT 62.825 152.165 63.490 152.335 ;
        RECT 63.675 152.190 63.945 153.095 ;
        RECT 63.320 152.020 63.490 152.165 ;
        RECT 61.355 151.485 62.565 152.005 ;
        RECT 62.755 151.615 63.085 151.985 ;
        RECT 63.320 151.690 63.605 152.020 ;
        RECT 58.225 150.885 58.395 151.265 ;
        RECT 58.575 150.715 58.905 151.095 ;
        RECT 59.085 150.885 59.345 151.390 ;
        RECT 59.975 150.715 62.565 151.485 ;
        RECT 63.320 151.435 63.490 151.690 ;
        RECT 62.825 151.265 63.490 151.435 ;
        RECT 63.775 151.390 63.945 152.190 ;
        RECT 64.575 152.175 67.165 153.265 ;
        RECT 67.425 152.335 67.595 153.095 ;
        RECT 67.810 152.505 68.140 153.265 ;
        RECT 64.575 151.655 65.785 152.175 ;
        RECT 67.425 152.165 68.140 152.335 ;
        RECT 68.310 152.190 68.565 153.095 ;
        RECT 65.955 151.485 67.165 152.005 ;
        RECT 67.335 151.615 67.690 151.985 ;
        RECT 67.970 151.955 68.140 152.165 ;
        RECT 67.970 151.625 68.225 151.955 ;
        RECT 62.825 150.885 62.995 151.265 ;
        RECT 63.175 150.715 63.505 151.095 ;
        RECT 63.685 150.885 63.945 151.390 ;
        RECT 64.575 150.715 67.165 151.485 ;
        RECT 67.970 151.435 68.140 151.625 ;
        RECT 68.395 151.460 68.565 152.190 ;
        RECT 68.740 152.115 69.000 153.265 ;
        RECT 69.265 152.335 69.435 153.095 ;
        RECT 69.650 152.505 69.980 153.265 ;
        RECT 69.265 152.165 69.980 152.335 ;
        RECT 70.150 152.190 70.405 153.095 ;
        RECT 69.175 151.615 69.530 151.985 ;
        RECT 69.810 151.955 69.980 152.165 ;
        RECT 69.810 151.625 70.065 151.955 ;
        RECT 67.425 151.265 68.140 151.435 ;
        RECT 67.425 150.885 67.595 151.265 ;
        RECT 67.810 150.715 68.140 151.095 ;
        RECT 68.310 150.885 68.565 151.460 ;
        RECT 68.740 150.715 69.000 151.555 ;
        RECT 69.810 151.435 69.980 151.625 ;
        RECT 70.235 151.460 70.405 152.190 ;
        RECT 70.580 152.115 70.840 153.265 ;
        RECT 71.025 152.205 71.355 153.265 ;
        RECT 71.535 151.955 71.705 152.925 ;
        RECT 71.875 152.675 72.205 153.075 ;
        RECT 72.375 152.905 72.705 153.265 ;
        RECT 72.905 152.675 73.605 153.095 ;
        RECT 71.875 152.445 73.605 152.675 ;
        RECT 71.875 152.225 72.205 152.445 ;
        RECT 72.400 151.955 72.725 152.245 ;
        RECT 71.015 151.625 71.325 151.955 ;
        RECT 71.535 151.625 71.910 151.955 ;
        RECT 72.230 151.625 72.725 151.955 ;
        RECT 72.900 151.705 73.230 152.245 ;
        RECT 73.400 151.565 73.605 152.445 ;
        RECT 73.980 152.295 74.310 153.095 ;
        RECT 74.480 152.465 74.810 153.265 ;
        RECT 75.110 152.295 75.440 153.095 ;
        RECT 76.085 152.465 76.335 153.265 ;
        RECT 73.980 152.125 76.415 152.295 ;
        RECT 76.605 152.125 76.775 153.265 ;
        RECT 76.945 152.125 77.285 153.095 ;
        RECT 73.775 151.705 74.125 151.955 ;
        RECT 69.265 151.265 69.980 151.435 ;
        RECT 69.265 150.885 69.435 151.265 ;
        RECT 69.650 150.715 69.980 151.095 ;
        RECT 70.150 150.885 70.405 151.460 ;
        RECT 70.580 150.715 70.840 151.555 ;
        RECT 73.375 151.475 73.605 151.565 ;
        RECT 74.310 151.495 74.480 152.125 ;
        RECT 74.650 151.705 74.980 151.905 ;
        RECT 75.150 151.705 75.480 151.905 ;
        RECT 75.650 151.705 76.070 151.905 ;
        RECT 76.245 151.875 76.415 152.125 ;
        RECT 76.245 151.705 76.940 151.875 ;
        RECT 71.025 151.245 72.385 151.455 ;
        RECT 71.025 150.885 71.355 151.245 ;
        RECT 71.525 150.715 71.855 151.075 ;
        RECT 72.055 150.885 72.385 151.245 ;
        RECT 72.895 150.885 73.605 151.475 ;
        RECT 73.980 150.885 74.480 151.495 ;
        RECT 75.110 151.365 76.335 151.535 ;
        RECT 77.110 151.515 77.285 152.125 ;
        RECT 77.455 152.100 77.745 153.265 ;
        RECT 77.915 152.125 78.255 153.095 ;
        RECT 78.425 152.125 78.595 153.265 ;
        RECT 78.865 152.465 79.115 153.265 ;
        RECT 79.760 152.295 80.090 153.095 ;
        RECT 80.390 152.465 80.720 153.265 ;
        RECT 80.890 152.295 81.220 153.095 ;
        RECT 78.785 152.125 81.220 152.295 ;
        RECT 82.515 152.175 86.025 153.265 ;
        RECT 86.200 152.830 91.545 153.265 ;
        RECT 91.720 152.830 97.065 153.265 ;
        RECT 75.110 150.885 75.440 151.365 ;
        RECT 75.610 150.715 75.835 151.175 ;
        RECT 76.005 150.885 76.335 151.365 ;
        RECT 76.525 150.715 76.775 151.515 ;
        RECT 76.945 150.885 77.285 151.515 ;
        RECT 77.915 151.515 78.090 152.125 ;
        RECT 78.785 151.875 78.955 152.125 ;
        RECT 78.260 151.705 78.955 151.875 ;
        RECT 79.130 151.705 79.550 151.905 ;
        RECT 79.720 151.705 80.050 151.905 ;
        RECT 80.220 151.705 80.550 151.905 ;
        RECT 77.455 150.715 77.745 151.440 ;
        RECT 77.915 150.885 78.255 151.515 ;
        RECT 78.425 150.715 78.675 151.515 ;
        RECT 78.865 151.365 80.090 151.535 ;
        RECT 78.865 150.885 79.195 151.365 ;
        RECT 79.365 150.715 79.590 151.175 ;
        RECT 79.760 150.885 80.090 151.365 ;
        RECT 80.720 151.495 80.890 152.125 ;
        RECT 81.075 151.705 81.425 151.955 ;
        RECT 82.515 151.655 84.205 152.175 ;
        RECT 80.720 150.885 81.220 151.495 ;
        RECT 84.375 151.485 86.025 152.005 ;
        RECT 87.790 151.580 88.140 152.830 ;
        RECT 82.515 150.715 86.025 151.485 ;
        RECT 89.620 151.260 89.960 152.090 ;
        RECT 93.310 151.580 93.660 152.830 ;
        RECT 97.235 152.125 97.575 153.095 ;
        RECT 97.745 152.125 97.915 153.265 ;
        RECT 98.185 152.465 98.435 153.265 ;
        RECT 99.080 152.295 99.410 153.095 ;
        RECT 99.710 152.465 100.040 153.265 ;
        RECT 100.210 152.295 100.540 153.095 ;
        RECT 98.105 152.125 100.540 152.295 ;
        RECT 101.375 152.175 103.045 153.265 ;
        RECT 95.140 151.260 95.480 152.090 ;
        RECT 97.235 151.515 97.410 152.125 ;
        RECT 98.105 151.875 98.275 152.125 ;
        RECT 97.580 151.705 98.275 151.875 ;
        RECT 98.450 151.705 98.870 151.905 ;
        RECT 99.040 151.705 99.370 151.905 ;
        RECT 99.540 151.705 99.870 151.905 ;
        RECT 86.200 150.715 91.545 151.260 ;
        RECT 91.720 150.715 97.065 151.260 ;
        RECT 97.235 150.885 97.575 151.515 ;
        RECT 97.745 150.715 97.995 151.515 ;
        RECT 98.185 151.365 99.410 151.535 ;
        RECT 98.185 150.885 98.515 151.365 ;
        RECT 98.685 150.715 98.910 151.175 ;
        RECT 99.080 150.885 99.410 151.365 ;
        RECT 100.040 151.495 100.210 152.125 ;
        RECT 100.395 151.705 100.745 151.955 ;
        RECT 101.375 151.655 102.125 152.175 ;
        RECT 103.215 152.100 103.505 153.265 ;
        RECT 104.135 152.175 105.805 153.265 ;
        RECT 106.180 152.295 106.510 153.095 ;
        RECT 106.680 152.465 107.010 153.265 ;
        RECT 107.310 152.295 107.640 153.095 ;
        RECT 108.285 152.465 108.535 153.265 ;
        RECT 100.040 150.885 100.540 151.495 ;
        RECT 102.295 151.485 103.045 152.005 ;
        RECT 104.135 151.655 104.885 152.175 ;
        RECT 106.180 152.125 108.615 152.295 ;
        RECT 108.805 152.125 108.975 153.265 ;
        RECT 109.145 152.125 109.485 153.095 ;
        RECT 109.860 152.295 110.190 153.095 ;
        RECT 110.360 152.465 110.690 153.265 ;
        RECT 110.990 152.295 111.320 153.095 ;
        RECT 111.965 152.465 112.215 153.265 ;
        RECT 109.860 152.125 112.295 152.295 ;
        RECT 112.485 152.125 112.655 153.265 ;
        RECT 112.825 152.125 113.165 153.095 ;
        RECT 105.055 151.485 105.805 152.005 ;
        RECT 105.975 151.705 106.325 151.955 ;
        RECT 106.510 151.495 106.680 152.125 ;
        RECT 106.850 151.705 107.180 151.905 ;
        RECT 107.350 151.705 107.680 151.905 ;
        RECT 107.850 151.705 108.270 151.905 ;
        RECT 108.445 151.875 108.615 152.125 ;
        RECT 108.445 151.705 109.140 151.875 ;
        RECT 101.375 150.715 103.045 151.485 ;
        RECT 103.215 150.715 103.505 151.440 ;
        RECT 104.135 150.715 105.805 151.485 ;
        RECT 106.180 150.885 106.680 151.495 ;
        RECT 107.310 151.365 108.535 151.535 ;
        RECT 109.310 151.515 109.485 152.125 ;
        RECT 109.655 151.705 110.005 151.955 ;
        RECT 107.310 150.885 107.640 151.365 ;
        RECT 107.810 150.715 108.035 151.175 ;
        RECT 108.205 150.885 108.535 151.365 ;
        RECT 108.725 150.715 108.975 151.515 ;
        RECT 109.145 150.885 109.485 151.515 ;
        RECT 110.190 151.495 110.360 152.125 ;
        RECT 110.530 151.705 110.860 151.905 ;
        RECT 111.030 151.705 111.360 151.905 ;
        RECT 111.530 151.705 111.950 151.905 ;
        RECT 112.125 151.875 112.295 152.125 ;
        RECT 112.125 151.705 112.820 151.875 ;
        RECT 109.860 150.885 110.360 151.495 ;
        RECT 110.990 151.365 112.215 151.535 ;
        RECT 112.990 151.515 113.165 152.125 ;
        RECT 113.335 152.175 115.925 153.265 ;
        RECT 116.185 152.335 116.355 153.095 ;
        RECT 116.535 152.505 116.865 153.265 ;
        RECT 113.335 151.655 114.545 152.175 ;
        RECT 116.185 152.165 116.850 152.335 ;
        RECT 117.035 152.190 117.305 153.095 ;
        RECT 116.680 152.020 116.850 152.165 ;
        RECT 110.990 150.885 111.320 151.365 ;
        RECT 111.490 150.715 111.715 151.175 ;
        RECT 111.885 150.885 112.215 151.365 ;
        RECT 112.405 150.715 112.655 151.515 ;
        RECT 112.825 150.885 113.165 151.515 ;
        RECT 114.715 151.485 115.925 152.005 ;
        RECT 116.115 151.615 116.445 151.985 ;
        RECT 116.680 151.690 116.965 152.020 ;
        RECT 113.335 150.715 115.925 151.485 ;
        RECT 116.680 151.435 116.850 151.690 ;
        RECT 116.185 151.265 116.850 151.435 ;
        RECT 117.135 151.390 117.305 152.190 ;
        RECT 116.185 150.885 116.355 151.265 ;
        RECT 116.535 150.715 116.865 151.095 ;
        RECT 117.045 150.885 117.305 151.390 ;
        RECT 117.850 152.285 118.105 152.955 ;
        RECT 118.285 152.465 118.570 153.265 ;
        RECT 118.750 152.545 119.080 153.055 ;
        RECT 117.850 151.425 118.030 152.285 ;
        RECT 118.750 151.955 119.000 152.545 ;
        RECT 119.350 152.395 119.520 153.005 ;
        RECT 119.690 152.575 120.020 153.265 ;
        RECT 120.250 152.715 120.490 153.005 ;
        RECT 120.690 152.885 121.110 153.265 ;
        RECT 121.290 152.795 121.920 153.045 ;
        RECT 122.390 152.885 122.720 153.265 ;
        RECT 121.290 152.715 121.460 152.795 ;
        RECT 122.890 152.715 123.060 153.005 ;
        RECT 123.240 152.885 123.620 153.265 ;
        RECT 123.860 152.880 124.690 153.050 ;
        RECT 120.250 152.545 121.460 152.715 ;
        RECT 118.200 151.625 119.000 151.955 ;
        RECT 117.850 151.225 118.105 151.425 ;
        RECT 117.765 151.055 118.105 151.225 ;
        RECT 117.850 150.895 118.105 151.055 ;
        RECT 118.285 150.715 118.570 151.175 ;
        RECT 118.750 150.975 119.000 151.625 ;
        RECT 119.200 152.375 119.520 152.395 ;
        RECT 119.200 152.205 121.120 152.375 ;
        RECT 119.200 151.310 119.390 152.205 ;
        RECT 121.290 152.035 121.460 152.545 ;
        RECT 121.630 152.285 122.150 152.595 ;
        RECT 119.560 151.865 121.460 152.035 ;
        RECT 119.560 151.805 119.890 151.865 ;
        RECT 120.040 151.635 120.370 151.695 ;
        RECT 119.710 151.365 120.370 151.635 ;
        RECT 119.200 150.980 119.520 151.310 ;
        RECT 119.700 150.715 120.360 151.195 ;
        RECT 120.560 151.105 120.730 151.865 ;
        RECT 121.630 151.695 121.810 152.105 ;
        RECT 120.900 151.525 121.230 151.645 ;
        RECT 121.980 151.525 122.150 152.285 ;
        RECT 120.900 151.355 122.150 151.525 ;
        RECT 122.320 152.465 123.690 152.715 ;
        RECT 122.320 151.695 122.510 152.465 ;
        RECT 123.440 152.205 123.690 152.465 ;
        RECT 122.680 152.035 122.930 152.195 ;
        RECT 123.860 152.035 124.030 152.880 ;
        RECT 124.925 152.595 125.095 153.095 ;
        RECT 125.265 152.765 125.595 153.265 ;
        RECT 124.200 152.205 124.700 152.585 ;
        RECT 124.925 152.425 125.620 152.595 ;
        RECT 122.680 151.865 124.030 152.035 ;
        RECT 123.610 151.825 124.030 151.865 ;
        RECT 122.320 151.355 122.740 151.695 ;
        RECT 123.030 151.365 123.440 151.695 ;
        RECT 120.560 150.935 121.410 151.105 ;
        RECT 121.970 150.715 122.290 151.175 ;
        RECT 122.490 150.925 122.740 151.355 ;
        RECT 123.030 150.715 123.440 151.155 ;
        RECT 123.610 151.095 123.780 151.825 ;
        RECT 123.950 151.275 124.300 151.645 ;
        RECT 124.480 151.335 124.700 152.205 ;
        RECT 124.870 151.635 125.280 152.255 ;
        RECT 125.450 151.455 125.620 152.425 ;
        RECT 124.925 151.265 125.620 151.455 ;
        RECT 123.610 150.895 124.625 151.095 ;
        RECT 124.925 150.935 125.095 151.265 ;
        RECT 125.265 150.715 125.595 151.095 ;
        RECT 125.810 150.975 126.035 153.095 ;
        RECT 126.205 152.765 126.535 153.265 ;
        RECT 126.705 152.595 126.875 153.095 ;
        RECT 126.210 152.425 126.875 152.595 ;
        RECT 126.210 151.435 126.440 152.425 ;
        RECT 126.610 151.605 126.960 152.255 ;
        RECT 128.055 152.175 129.265 153.265 ;
        RECT 128.055 151.635 128.575 152.175 ;
        RECT 128.745 151.465 129.265 152.005 ;
        RECT 126.210 151.265 126.875 151.435 ;
        RECT 126.205 150.715 126.535 151.095 ;
        RECT 126.705 150.975 126.875 151.265 ;
        RECT 128.055 150.715 129.265 151.465 ;
        RECT 9.290 150.545 129.350 150.715 ;
        RECT 9.375 149.795 10.585 150.545 ;
        RECT 9.375 149.255 9.895 149.795 ;
        RECT 11.215 149.775 12.885 150.545 ;
        RECT 13.055 149.820 13.345 150.545 ;
        RECT 10.065 149.085 10.585 149.625 ;
        RECT 9.375 147.995 10.585 149.085 ;
        RECT 11.215 149.085 11.965 149.605 ;
        RECT 12.135 149.255 12.885 149.775 ;
        RECT 13.575 149.725 13.785 150.545 ;
        RECT 13.955 149.745 14.285 150.375 ;
        RECT 11.215 147.995 12.885 149.085 ;
        RECT 13.055 147.995 13.345 149.160 ;
        RECT 13.955 149.145 14.205 149.745 ;
        RECT 14.455 149.725 14.685 150.545 ;
        RECT 14.985 149.995 15.155 150.375 ;
        RECT 15.335 150.165 15.665 150.545 ;
        RECT 14.985 149.825 15.650 149.995 ;
        RECT 15.845 149.870 16.105 150.375 ;
        RECT 14.375 149.305 14.705 149.555 ;
        RECT 14.915 149.275 15.245 149.645 ;
        RECT 15.480 149.570 15.650 149.825 ;
        RECT 15.480 149.240 15.765 149.570 ;
        RECT 13.575 147.995 13.785 149.135 ;
        RECT 13.955 148.165 14.285 149.145 ;
        RECT 14.455 147.995 14.685 149.135 ;
        RECT 15.480 149.095 15.650 149.240 ;
        RECT 14.985 148.925 15.650 149.095 ;
        RECT 15.935 149.070 16.105 149.870 ;
        RECT 14.985 148.165 15.155 148.925 ;
        RECT 15.335 147.995 15.665 148.755 ;
        RECT 15.835 148.165 16.105 149.070 ;
        RECT 16.280 149.805 16.535 150.375 ;
        RECT 16.705 150.145 17.035 150.545 ;
        RECT 17.460 150.010 17.990 150.375 ;
        RECT 17.460 149.975 17.635 150.010 ;
        RECT 16.705 149.805 17.635 149.975 ;
        RECT 18.180 149.865 18.455 150.375 ;
        RECT 16.280 149.135 16.450 149.805 ;
        RECT 16.705 149.635 16.875 149.805 ;
        RECT 16.620 149.305 16.875 149.635 ;
        RECT 17.100 149.305 17.295 149.635 ;
        RECT 16.280 148.165 16.615 149.135 ;
        RECT 16.785 147.995 16.955 149.135 ;
        RECT 17.125 148.335 17.295 149.305 ;
        RECT 17.465 148.675 17.635 149.805 ;
        RECT 17.805 149.015 17.975 149.815 ;
        RECT 18.175 149.695 18.455 149.865 ;
        RECT 18.180 149.215 18.455 149.695 ;
        RECT 18.625 149.015 18.815 150.375 ;
        RECT 18.995 150.010 19.505 150.545 ;
        RECT 19.725 149.735 19.970 150.340 ;
        RECT 20.420 150.000 25.765 150.545 ;
        RECT 25.940 150.000 31.285 150.545 ;
        RECT 19.015 149.565 20.245 149.735 ;
        RECT 17.805 148.845 18.815 149.015 ;
        RECT 18.985 149.000 19.735 149.190 ;
        RECT 17.465 148.505 18.590 148.675 ;
        RECT 18.985 148.335 19.155 149.000 ;
        RECT 19.905 148.755 20.245 149.565 ;
        RECT 17.125 148.165 19.155 148.335 ;
        RECT 19.325 147.995 19.495 148.755 ;
        RECT 19.730 148.345 20.245 148.755 ;
        RECT 22.010 148.430 22.360 149.680 ;
        RECT 23.840 149.170 24.180 150.000 ;
        RECT 27.530 148.430 27.880 149.680 ;
        RECT 29.360 149.170 29.700 150.000 ;
        RECT 31.455 149.745 31.795 150.375 ;
        RECT 31.965 149.745 32.215 150.545 ;
        RECT 32.405 149.895 32.735 150.375 ;
        RECT 32.905 150.085 33.130 150.545 ;
        RECT 33.300 149.895 33.630 150.375 ;
        RECT 31.455 149.135 31.630 149.745 ;
        RECT 32.405 149.725 33.630 149.895 ;
        RECT 34.260 149.765 34.760 150.375 ;
        RECT 35.340 149.765 35.840 150.375 ;
        RECT 31.800 149.385 32.495 149.555 ;
        RECT 32.325 149.135 32.495 149.385 ;
        RECT 32.670 149.355 33.090 149.555 ;
        RECT 33.260 149.355 33.590 149.555 ;
        RECT 33.760 149.355 34.090 149.555 ;
        RECT 34.260 149.135 34.430 149.765 ;
        RECT 34.615 149.305 34.965 149.555 ;
        RECT 35.135 149.305 35.485 149.555 ;
        RECT 35.670 149.135 35.840 149.765 ;
        RECT 36.470 149.895 36.800 150.375 ;
        RECT 36.970 150.085 37.195 150.545 ;
        RECT 37.365 149.895 37.695 150.375 ;
        RECT 36.470 149.725 37.695 149.895 ;
        RECT 37.885 149.745 38.135 150.545 ;
        RECT 38.305 149.745 38.645 150.375 ;
        RECT 38.815 149.820 39.105 150.545 ;
        RECT 40.195 149.775 43.705 150.545 ;
        RECT 36.010 149.355 36.340 149.555 ;
        RECT 36.510 149.355 36.840 149.555 ;
        RECT 37.010 149.355 37.430 149.555 ;
        RECT 37.605 149.385 38.300 149.555 ;
        RECT 37.605 149.135 37.775 149.385 ;
        RECT 38.470 149.135 38.645 149.745 ;
        RECT 20.420 147.995 25.765 148.430 ;
        RECT 25.940 147.995 31.285 148.430 ;
        RECT 31.455 148.165 31.795 149.135 ;
        RECT 31.965 147.995 32.135 149.135 ;
        RECT 32.325 148.965 34.760 149.135 ;
        RECT 32.405 147.995 32.655 148.795 ;
        RECT 33.300 148.165 33.630 148.965 ;
        RECT 33.930 147.995 34.260 148.795 ;
        RECT 34.430 148.165 34.760 148.965 ;
        RECT 35.340 148.965 37.775 149.135 ;
        RECT 35.340 148.165 35.670 148.965 ;
        RECT 35.840 147.995 36.170 148.795 ;
        RECT 36.470 148.165 36.800 148.965 ;
        RECT 37.445 147.995 37.695 148.795 ;
        RECT 37.965 147.995 38.135 149.135 ;
        RECT 38.305 148.165 38.645 149.135 ;
        RECT 38.815 147.995 39.105 149.160 ;
        RECT 40.195 149.085 41.885 149.605 ;
        RECT 42.055 149.255 43.705 149.775 ;
        RECT 43.875 149.870 44.145 150.215 ;
        RECT 44.335 150.145 44.715 150.545 ;
        RECT 44.885 149.975 45.055 150.325 ;
        RECT 45.225 150.145 45.555 150.545 ;
        RECT 45.755 149.975 45.925 150.325 ;
        RECT 46.125 150.045 46.455 150.545 ;
        RECT 43.875 149.135 44.045 149.870 ;
        RECT 44.315 149.805 45.925 149.975 ;
        RECT 44.315 149.635 44.485 149.805 ;
        RECT 44.215 149.305 44.485 149.635 ;
        RECT 44.655 149.305 45.060 149.635 ;
        RECT 44.315 149.135 44.485 149.305 ;
        RECT 40.195 147.995 43.705 149.085 ;
        RECT 43.875 148.165 44.145 149.135 ;
        RECT 44.315 148.965 45.040 149.135 ;
        RECT 45.230 149.015 45.940 149.635 ;
        RECT 46.110 149.305 46.460 149.875 ;
        RECT 46.635 149.870 46.905 150.215 ;
        RECT 47.095 150.145 47.475 150.545 ;
        RECT 47.645 149.975 47.815 150.325 ;
        RECT 47.985 150.145 48.315 150.545 ;
        RECT 48.515 149.975 48.685 150.325 ;
        RECT 48.885 150.045 49.215 150.545 ;
        RECT 46.635 149.135 46.805 149.870 ;
        RECT 47.075 149.805 48.685 149.975 ;
        RECT 47.075 149.635 47.245 149.805 ;
        RECT 46.975 149.305 47.245 149.635 ;
        RECT 47.415 149.305 47.820 149.635 ;
        RECT 47.075 149.135 47.245 149.305 ;
        RECT 44.870 148.845 45.040 148.965 ;
        RECT 46.140 148.845 46.460 149.135 ;
        RECT 44.355 147.995 44.635 148.795 ;
        RECT 44.870 148.675 46.460 148.845 ;
        RECT 44.805 148.215 46.460 148.505 ;
        RECT 46.635 148.165 46.905 149.135 ;
        RECT 47.075 148.965 47.800 149.135 ;
        RECT 47.990 149.015 48.700 149.635 ;
        RECT 48.870 149.305 49.220 149.875 ;
        RECT 49.395 149.775 51.065 150.545 ;
        RECT 47.630 148.845 47.800 148.965 ;
        RECT 48.900 148.845 49.220 149.135 ;
        RECT 47.115 147.995 47.395 148.795 ;
        RECT 47.630 148.675 49.220 148.845 ;
        RECT 49.395 149.085 50.145 149.605 ;
        RECT 50.315 149.255 51.065 149.775 ;
        RECT 51.235 149.745 51.575 150.375 ;
        RECT 51.745 149.745 51.995 150.545 ;
        RECT 52.185 149.895 52.515 150.375 ;
        RECT 52.685 150.085 52.910 150.545 ;
        RECT 53.080 149.895 53.410 150.375 ;
        RECT 51.235 149.135 51.410 149.745 ;
        RECT 52.185 149.725 53.410 149.895 ;
        RECT 54.040 149.765 54.540 150.375 ;
        RECT 55.835 149.775 59.345 150.545 ;
        RECT 51.580 149.385 52.275 149.555 ;
        RECT 52.105 149.135 52.275 149.385 ;
        RECT 52.450 149.355 52.870 149.555 ;
        RECT 53.040 149.355 53.370 149.555 ;
        RECT 53.540 149.355 53.870 149.555 ;
        RECT 54.040 149.135 54.210 149.765 ;
        RECT 54.395 149.305 54.745 149.555 ;
        RECT 47.565 148.215 49.220 148.505 ;
        RECT 49.395 147.995 51.065 149.085 ;
        RECT 51.235 148.165 51.575 149.135 ;
        RECT 51.745 147.995 51.915 149.135 ;
        RECT 52.105 148.965 54.540 149.135 ;
        RECT 52.185 147.995 52.435 148.795 ;
        RECT 53.080 148.165 53.410 148.965 ;
        RECT 53.710 147.995 54.040 148.795 ;
        RECT 54.210 148.165 54.540 148.965 ;
        RECT 55.835 149.085 57.525 149.605 ;
        RECT 57.695 149.255 59.345 149.775 ;
        RECT 59.790 149.735 60.035 150.340 ;
        RECT 60.255 150.010 60.765 150.545 ;
        RECT 59.515 149.565 60.745 149.735 ;
        RECT 55.835 147.995 59.345 149.085 ;
        RECT 59.515 148.755 59.855 149.565 ;
        RECT 60.025 149.000 60.775 149.190 ;
        RECT 59.515 148.345 60.030 148.755 ;
        RECT 60.265 147.995 60.435 148.755 ;
        RECT 60.605 148.335 60.775 149.000 ;
        RECT 60.945 149.015 61.135 150.375 ;
        RECT 61.305 149.525 61.580 150.375 ;
        RECT 61.770 150.010 62.300 150.375 ;
        RECT 62.725 150.145 63.055 150.545 ;
        RECT 62.125 149.975 62.300 150.010 ;
        RECT 61.305 149.355 61.585 149.525 ;
        RECT 61.305 149.215 61.580 149.355 ;
        RECT 61.785 149.015 61.955 149.815 ;
        RECT 60.945 148.845 61.955 149.015 ;
        RECT 62.125 149.805 63.055 149.975 ;
        RECT 63.225 149.805 63.480 150.375 ;
        RECT 64.575 149.820 64.865 150.545 ;
        RECT 62.125 148.675 62.295 149.805 ;
        RECT 62.885 149.635 63.055 149.805 ;
        RECT 61.170 148.505 62.295 148.675 ;
        RECT 62.465 149.305 62.660 149.635 ;
        RECT 62.885 149.305 63.140 149.635 ;
        RECT 62.465 148.335 62.635 149.305 ;
        RECT 63.310 149.135 63.480 149.805 ;
        RECT 65.040 149.705 65.300 150.545 ;
        RECT 65.475 149.800 65.730 150.375 ;
        RECT 65.900 150.165 66.230 150.545 ;
        RECT 66.445 149.995 66.615 150.375 ;
        RECT 65.900 149.825 66.615 149.995 ;
        RECT 60.605 148.165 62.635 148.335 ;
        RECT 62.805 147.995 62.975 149.135 ;
        RECT 63.145 148.165 63.480 149.135 ;
        RECT 64.575 147.995 64.865 149.160 ;
        RECT 65.040 147.995 65.300 149.145 ;
        RECT 65.475 149.070 65.645 149.800 ;
        RECT 65.900 149.635 66.070 149.825 ;
        RECT 66.880 149.705 67.140 150.545 ;
        RECT 67.315 149.800 67.570 150.375 ;
        RECT 67.740 150.165 68.070 150.545 ;
        RECT 68.285 149.995 68.455 150.375 ;
        RECT 68.775 150.065 69.055 150.545 ;
        RECT 67.740 149.825 68.455 149.995 ;
        RECT 69.225 149.895 69.485 150.285 ;
        RECT 69.660 150.065 69.915 150.545 ;
        RECT 70.085 149.895 70.380 150.285 ;
        RECT 70.560 150.065 70.835 150.545 ;
        RECT 71.005 150.045 71.305 150.375 ;
        RECT 65.815 149.305 66.070 149.635 ;
        RECT 65.900 149.095 66.070 149.305 ;
        RECT 66.350 149.275 66.705 149.645 ;
        RECT 65.475 148.165 65.730 149.070 ;
        RECT 65.900 148.925 66.615 149.095 ;
        RECT 65.900 147.995 66.230 148.755 ;
        RECT 66.445 148.165 66.615 148.925 ;
        RECT 66.880 147.995 67.140 149.145 ;
        RECT 67.315 149.070 67.485 149.800 ;
        RECT 67.740 149.635 67.910 149.825 ;
        RECT 68.730 149.725 70.380 149.895 ;
        RECT 67.655 149.305 67.910 149.635 ;
        RECT 67.740 149.095 67.910 149.305 ;
        RECT 68.190 149.275 68.545 149.645 ;
        RECT 68.730 149.215 69.135 149.725 ;
        RECT 69.305 149.385 70.445 149.555 ;
        RECT 67.315 148.165 67.570 149.070 ;
        RECT 67.740 148.925 68.455 149.095 ;
        RECT 68.730 149.045 69.485 149.215 ;
        RECT 67.740 147.995 68.070 148.755 ;
        RECT 68.285 148.165 68.455 148.925 ;
        RECT 68.770 147.995 69.055 148.865 ;
        RECT 69.225 148.795 69.485 149.045 ;
        RECT 70.275 149.135 70.445 149.385 ;
        RECT 70.615 149.305 70.965 149.875 ;
        RECT 71.135 149.135 71.305 150.045 ;
        RECT 71.565 149.995 71.735 150.375 ;
        RECT 71.950 150.165 72.280 150.545 ;
        RECT 71.565 149.825 72.280 149.995 ;
        RECT 71.475 149.275 71.830 149.645 ;
        RECT 72.110 149.635 72.280 149.825 ;
        RECT 72.450 149.800 72.705 150.375 ;
        RECT 72.110 149.305 72.365 149.635 ;
        RECT 70.275 148.965 71.305 149.135 ;
        RECT 72.110 149.095 72.280 149.305 ;
        RECT 69.225 148.625 70.345 148.795 ;
        RECT 69.225 148.165 69.485 148.625 ;
        RECT 69.660 147.995 69.915 148.455 ;
        RECT 70.085 148.165 70.345 148.625 ;
        RECT 70.515 147.995 70.825 148.795 ;
        RECT 70.995 148.165 71.305 148.965 ;
        RECT 71.565 148.925 72.280 149.095 ;
        RECT 72.535 149.070 72.705 149.800 ;
        RECT 72.880 149.705 73.140 150.545 ;
        RECT 73.775 149.775 75.445 150.545 ;
        RECT 71.565 148.165 71.735 148.925 ;
        RECT 71.950 147.995 72.280 148.755 ;
        RECT 72.450 148.165 72.705 149.070 ;
        RECT 72.880 147.995 73.140 149.145 ;
        RECT 73.775 149.085 74.525 149.605 ;
        RECT 74.695 149.255 75.445 149.775 ;
        RECT 75.615 150.045 75.915 150.375 ;
        RECT 76.085 150.065 76.360 150.545 ;
        RECT 75.615 149.135 75.785 150.045 ;
        RECT 76.540 149.895 76.835 150.285 ;
        RECT 77.005 150.065 77.260 150.545 ;
        RECT 77.435 149.895 77.695 150.285 ;
        RECT 77.865 150.065 78.145 150.545 ;
        RECT 75.955 149.305 76.305 149.875 ;
        RECT 76.540 149.725 78.190 149.895 ;
        RECT 76.475 149.385 77.615 149.555 ;
        RECT 76.475 149.135 76.645 149.385 ;
        RECT 77.785 149.215 78.190 149.725 ;
        RECT 73.775 147.995 75.445 149.085 ;
        RECT 75.615 148.965 76.645 149.135 ;
        RECT 77.435 149.045 78.190 149.215 ;
        RECT 78.375 149.745 78.715 150.375 ;
        RECT 78.885 149.745 79.135 150.545 ;
        RECT 79.325 149.895 79.655 150.375 ;
        RECT 79.825 150.085 80.050 150.545 ;
        RECT 80.220 149.895 80.550 150.375 ;
        RECT 78.375 149.135 78.550 149.745 ;
        RECT 79.325 149.725 80.550 149.895 ;
        RECT 81.180 149.765 81.680 150.375 ;
        RECT 82.515 149.775 86.025 150.545 ;
        RECT 78.720 149.385 79.415 149.555 ;
        RECT 79.245 149.135 79.415 149.385 ;
        RECT 79.590 149.355 80.010 149.555 ;
        RECT 80.180 149.355 80.510 149.555 ;
        RECT 80.680 149.355 81.010 149.555 ;
        RECT 81.180 149.135 81.350 149.765 ;
        RECT 81.535 149.305 81.885 149.555 ;
        RECT 75.615 148.165 75.925 148.965 ;
        RECT 77.435 148.795 77.695 149.045 ;
        RECT 76.095 147.995 76.405 148.795 ;
        RECT 76.575 148.625 77.695 148.795 ;
        RECT 76.575 148.165 76.835 148.625 ;
        RECT 77.005 147.995 77.260 148.455 ;
        RECT 77.435 148.165 77.695 148.625 ;
        RECT 77.865 147.995 78.150 148.865 ;
        RECT 78.375 148.165 78.715 149.135 ;
        RECT 78.885 147.995 79.055 149.135 ;
        RECT 79.245 148.965 81.680 149.135 ;
        RECT 79.325 147.995 79.575 148.795 ;
        RECT 80.220 148.165 80.550 148.965 ;
        RECT 80.850 147.995 81.180 148.795 ;
        RECT 81.350 148.165 81.680 148.965 ;
        RECT 82.515 149.085 84.205 149.605 ;
        RECT 84.375 149.255 86.025 149.775 ;
        RECT 86.470 149.735 86.715 150.340 ;
        RECT 86.935 150.010 87.445 150.545 ;
        RECT 86.195 149.565 87.425 149.735 ;
        RECT 82.515 147.995 86.025 149.085 ;
        RECT 86.195 148.755 86.535 149.565 ;
        RECT 86.705 149.000 87.455 149.190 ;
        RECT 86.195 148.345 86.710 148.755 ;
        RECT 86.945 147.995 87.115 148.755 ;
        RECT 87.285 148.335 87.455 149.000 ;
        RECT 87.625 149.015 87.815 150.375 ;
        RECT 87.985 149.525 88.260 150.375 ;
        RECT 88.450 150.010 88.980 150.375 ;
        RECT 89.405 150.145 89.735 150.545 ;
        RECT 88.805 149.975 88.980 150.010 ;
        RECT 87.985 149.355 88.265 149.525 ;
        RECT 87.985 149.215 88.260 149.355 ;
        RECT 88.465 149.015 88.635 149.815 ;
        RECT 87.625 148.845 88.635 149.015 ;
        RECT 88.805 149.805 89.735 149.975 ;
        RECT 89.905 149.805 90.160 150.375 ;
        RECT 90.335 149.820 90.625 150.545 ;
        RECT 88.805 148.675 88.975 149.805 ;
        RECT 89.565 149.635 89.735 149.805 ;
        RECT 87.850 148.505 88.975 148.675 ;
        RECT 89.145 149.305 89.340 149.635 ;
        RECT 89.565 149.305 89.820 149.635 ;
        RECT 89.145 148.335 89.315 149.305 ;
        RECT 89.990 149.135 90.160 149.805 ;
        RECT 90.795 149.775 92.465 150.545 ;
        RECT 87.285 148.165 89.315 148.335 ;
        RECT 89.485 147.995 89.655 149.135 ;
        RECT 89.825 148.165 90.160 149.135 ;
        RECT 90.335 147.995 90.625 149.160 ;
        RECT 90.795 149.085 91.545 149.605 ;
        RECT 91.715 149.255 92.465 149.775 ;
        RECT 92.695 149.725 92.905 150.545 ;
        RECT 93.075 149.745 93.405 150.375 ;
        RECT 93.075 149.145 93.325 149.745 ;
        RECT 93.575 149.725 93.805 150.545 ;
        RECT 94.565 149.995 94.735 150.375 ;
        RECT 94.915 150.165 95.245 150.545 ;
        RECT 94.565 149.825 95.230 149.995 ;
        RECT 95.425 149.870 95.685 150.375 ;
        RECT 93.495 149.305 93.825 149.555 ;
        RECT 94.495 149.275 94.825 149.645 ;
        RECT 95.060 149.570 95.230 149.825 ;
        RECT 95.060 149.240 95.345 149.570 ;
        RECT 90.795 147.995 92.465 149.085 ;
        RECT 92.695 147.995 92.905 149.135 ;
        RECT 93.075 148.165 93.405 149.145 ;
        RECT 93.575 147.995 93.805 149.135 ;
        RECT 95.060 149.095 95.230 149.240 ;
        RECT 94.565 148.925 95.230 149.095 ;
        RECT 95.515 149.070 95.685 149.870 ;
        RECT 95.855 149.795 97.065 150.545 ;
        RECT 97.240 150.000 102.585 150.545 ;
        RECT 94.565 148.165 94.735 148.925 ;
        RECT 94.915 147.995 95.245 148.755 ;
        RECT 95.415 148.165 95.685 149.070 ;
        RECT 95.855 149.085 96.375 149.625 ;
        RECT 96.545 149.255 97.065 149.795 ;
        RECT 95.855 147.995 97.065 149.085 ;
        RECT 98.830 148.430 99.180 149.680 ;
        RECT 100.660 149.170 101.000 150.000 ;
        RECT 102.960 149.765 103.460 150.375 ;
        RECT 102.755 149.305 103.105 149.555 ;
        RECT 103.290 149.135 103.460 149.765 ;
        RECT 104.090 149.895 104.420 150.375 ;
        RECT 104.590 150.085 104.815 150.545 ;
        RECT 104.985 149.895 105.315 150.375 ;
        RECT 104.090 149.725 105.315 149.895 ;
        RECT 105.505 149.745 105.755 150.545 ;
        RECT 105.925 149.745 106.265 150.375 ;
        RECT 103.630 149.355 103.960 149.555 ;
        RECT 104.130 149.355 104.460 149.555 ;
        RECT 104.630 149.355 105.050 149.555 ;
        RECT 105.225 149.385 105.920 149.555 ;
        RECT 105.225 149.135 105.395 149.385 ;
        RECT 106.090 149.135 106.265 149.745 ;
        RECT 102.960 148.965 105.395 149.135 ;
        RECT 97.240 147.995 102.585 148.430 ;
        RECT 102.960 148.165 103.290 148.965 ;
        RECT 103.460 147.995 103.790 148.795 ;
        RECT 104.090 148.165 104.420 148.965 ;
        RECT 105.065 147.995 105.315 148.795 ;
        RECT 105.585 147.995 105.755 149.135 ;
        RECT 105.925 148.165 106.265 149.135 ;
        RECT 106.435 149.745 106.775 150.375 ;
        RECT 106.945 149.745 107.195 150.545 ;
        RECT 107.385 149.895 107.715 150.375 ;
        RECT 107.885 150.085 108.110 150.545 ;
        RECT 108.280 149.895 108.610 150.375 ;
        RECT 106.435 149.135 106.610 149.745 ;
        RECT 107.385 149.725 108.610 149.895 ;
        RECT 109.240 149.765 109.740 150.375 ;
        RECT 110.115 149.775 111.785 150.545 ;
        RECT 106.780 149.385 107.475 149.555 ;
        RECT 107.305 149.135 107.475 149.385 ;
        RECT 107.650 149.355 108.070 149.555 ;
        RECT 108.240 149.355 108.570 149.555 ;
        RECT 108.740 149.355 109.070 149.555 ;
        RECT 109.240 149.135 109.410 149.765 ;
        RECT 109.595 149.305 109.945 149.555 ;
        RECT 106.435 148.165 106.775 149.135 ;
        RECT 106.945 147.995 107.115 149.135 ;
        RECT 107.305 148.965 109.740 149.135 ;
        RECT 107.385 147.995 107.635 148.795 ;
        RECT 108.280 148.165 108.610 148.965 ;
        RECT 108.910 147.995 109.240 148.795 ;
        RECT 109.410 148.165 109.740 148.965 ;
        RECT 110.115 149.085 110.865 149.605 ;
        RECT 111.035 149.255 111.785 149.775 ;
        RECT 112.230 149.735 112.475 150.340 ;
        RECT 112.695 150.010 113.205 150.545 ;
        RECT 111.955 149.565 113.185 149.735 ;
        RECT 110.115 147.995 111.785 149.085 ;
        RECT 111.955 148.755 112.295 149.565 ;
        RECT 112.465 149.000 113.215 149.190 ;
        RECT 111.955 148.345 112.470 148.755 ;
        RECT 112.705 147.995 112.875 148.755 ;
        RECT 113.045 148.335 113.215 149.000 ;
        RECT 113.385 149.015 113.575 150.375 ;
        RECT 113.745 149.525 114.020 150.375 ;
        RECT 114.210 150.010 114.740 150.375 ;
        RECT 115.165 150.145 115.495 150.545 ;
        RECT 114.565 149.975 114.740 150.010 ;
        RECT 113.745 149.355 114.025 149.525 ;
        RECT 113.745 149.215 114.020 149.355 ;
        RECT 114.225 149.015 114.395 149.815 ;
        RECT 113.385 148.845 114.395 149.015 ;
        RECT 114.565 149.805 115.495 149.975 ;
        RECT 115.665 149.805 115.920 150.375 ;
        RECT 116.095 149.820 116.385 150.545 ;
        RECT 114.565 148.675 114.735 149.805 ;
        RECT 115.325 149.635 115.495 149.805 ;
        RECT 113.610 148.505 114.735 148.675 ;
        RECT 114.905 149.305 115.100 149.635 ;
        RECT 115.325 149.305 115.580 149.635 ;
        RECT 114.905 148.335 115.075 149.305 ;
        RECT 115.750 149.135 115.920 149.805 ;
        RECT 117.480 149.805 117.735 150.375 ;
        RECT 117.905 150.145 118.235 150.545 ;
        RECT 118.660 150.010 119.190 150.375 ;
        RECT 118.660 149.975 118.835 150.010 ;
        RECT 117.905 149.805 118.835 149.975 ;
        RECT 113.045 148.165 115.075 148.335 ;
        RECT 115.245 147.995 115.415 149.135 ;
        RECT 115.585 148.165 115.920 149.135 ;
        RECT 116.095 147.995 116.385 149.160 ;
        RECT 117.480 149.135 117.650 149.805 ;
        RECT 117.905 149.635 118.075 149.805 ;
        RECT 117.820 149.305 118.075 149.635 ;
        RECT 118.300 149.305 118.495 149.635 ;
        RECT 117.480 148.165 117.815 149.135 ;
        RECT 117.985 147.995 118.155 149.135 ;
        RECT 118.325 148.335 118.495 149.305 ;
        RECT 118.665 148.675 118.835 149.805 ;
        RECT 119.005 149.015 119.175 149.815 ;
        RECT 119.380 149.525 119.655 150.375 ;
        RECT 119.375 149.355 119.655 149.525 ;
        RECT 119.380 149.215 119.655 149.355 ;
        RECT 119.825 149.015 120.015 150.375 ;
        RECT 120.195 150.010 120.705 150.545 ;
        RECT 120.925 149.735 121.170 150.340 ;
        RECT 121.705 149.995 121.875 150.375 ;
        RECT 122.055 150.165 122.385 150.545 ;
        RECT 121.705 149.825 122.370 149.995 ;
        RECT 122.565 149.870 122.825 150.375 ;
        RECT 120.215 149.565 121.445 149.735 ;
        RECT 119.005 148.845 120.015 149.015 ;
        RECT 120.185 149.000 120.935 149.190 ;
        RECT 118.665 148.505 119.790 148.675 ;
        RECT 120.185 148.335 120.355 149.000 ;
        RECT 121.105 148.755 121.445 149.565 ;
        RECT 121.635 149.275 121.965 149.645 ;
        RECT 122.200 149.570 122.370 149.825 ;
        RECT 122.200 149.240 122.485 149.570 ;
        RECT 122.200 149.095 122.370 149.240 ;
        RECT 118.325 148.165 120.355 148.335 ;
        RECT 120.525 147.995 120.695 148.755 ;
        RECT 120.930 148.345 121.445 148.755 ;
        RECT 121.705 148.925 122.370 149.095 ;
        RECT 122.655 149.070 122.825 149.870 ;
        RECT 122.995 149.795 124.205 150.545 ;
        RECT 121.705 148.165 121.875 148.925 ;
        RECT 122.055 147.995 122.385 148.755 ;
        RECT 122.555 148.165 122.825 149.070 ;
        RECT 122.995 149.085 123.515 149.625 ;
        RECT 123.685 149.255 124.205 149.795 ;
        RECT 124.375 149.775 127.885 150.545 ;
        RECT 128.055 149.795 129.265 150.545 ;
        RECT 124.375 149.085 126.065 149.605 ;
        RECT 126.235 149.255 127.885 149.775 ;
        RECT 128.055 149.085 128.575 149.625 ;
        RECT 128.745 149.255 129.265 149.795 ;
        RECT 122.995 147.995 124.205 149.085 ;
        RECT 124.375 147.995 127.885 149.085 ;
        RECT 128.055 147.995 129.265 149.085 ;
        RECT 9.290 147.825 129.350 147.995 ;
        RECT 9.375 146.735 10.585 147.825 ;
        RECT 11.130 147.485 11.385 147.515 ;
        RECT 11.045 147.315 11.385 147.485 ;
        RECT 9.375 146.025 9.895 146.565 ;
        RECT 10.065 146.195 10.585 146.735 ;
        RECT 11.130 146.845 11.385 147.315 ;
        RECT 11.565 147.025 11.850 147.825 ;
        RECT 12.030 147.105 12.360 147.615 ;
        RECT 9.375 145.275 10.585 146.025 ;
        RECT 11.130 145.985 11.310 146.845 ;
        RECT 12.030 146.515 12.280 147.105 ;
        RECT 12.630 146.955 12.800 147.565 ;
        RECT 12.970 147.135 13.300 147.825 ;
        RECT 13.530 147.275 13.770 147.565 ;
        RECT 13.970 147.445 14.390 147.825 ;
        RECT 14.570 147.355 15.200 147.605 ;
        RECT 15.670 147.445 16.000 147.825 ;
        RECT 14.570 147.275 14.740 147.355 ;
        RECT 16.170 147.275 16.340 147.565 ;
        RECT 16.520 147.445 16.900 147.825 ;
        RECT 17.140 147.440 17.970 147.610 ;
        RECT 13.530 147.105 14.740 147.275 ;
        RECT 11.480 146.185 12.280 146.515 ;
        RECT 11.130 145.455 11.385 145.985 ;
        RECT 11.565 145.275 11.850 145.735 ;
        RECT 12.030 145.535 12.280 146.185 ;
        RECT 12.480 146.935 12.800 146.955 ;
        RECT 12.480 146.765 14.400 146.935 ;
        RECT 12.480 145.870 12.670 146.765 ;
        RECT 14.570 146.595 14.740 147.105 ;
        RECT 14.910 146.845 15.430 147.155 ;
        RECT 12.840 146.425 14.740 146.595 ;
        RECT 12.840 146.365 13.170 146.425 ;
        RECT 13.320 146.195 13.650 146.255 ;
        RECT 12.990 145.925 13.650 146.195 ;
        RECT 12.480 145.540 12.800 145.870 ;
        RECT 12.980 145.275 13.640 145.755 ;
        RECT 13.840 145.665 14.010 146.425 ;
        RECT 14.910 146.255 15.090 146.665 ;
        RECT 14.180 146.085 14.510 146.205 ;
        RECT 15.260 146.085 15.430 146.845 ;
        RECT 14.180 145.915 15.430 146.085 ;
        RECT 15.600 147.025 16.970 147.275 ;
        RECT 15.600 146.255 15.790 147.025 ;
        RECT 16.720 146.765 16.970 147.025 ;
        RECT 15.960 146.595 16.210 146.755 ;
        RECT 17.140 146.595 17.310 147.440 ;
        RECT 18.205 147.155 18.375 147.655 ;
        RECT 18.545 147.325 18.875 147.825 ;
        RECT 17.480 146.765 17.980 147.145 ;
        RECT 18.205 146.985 18.900 147.155 ;
        RECT 15.960 146.425 17.310 146.595 ;
        RECT 16.890 146.385 17.310 146.425 ;
        RECT 15.600 145.915 16.020 146.255 ;
        RECT 16.310 145.925 16.720 146.255 ;
        RECT 13.840 145.495 14.690 145.665 ;
        RECT 15.250 145.275 15.570 145.735 ;
        RECT 15.770 145.485 16.020 145.915 ;
        RECT 16.310 145.275 16.720 145.715 ;
        RECT 16.890 145.655 17.060 146.385 ;
        RECT 17.230 145.835 17.580 146.205 ;
        RECT 17.760 145.895 17.980 146.765 ;
        RECT 18.150 146.195 18.560 146.815 ;
        RECT 18.730 146.015 18.900 146.985 ;
        RECT 18.205 145.825 18.900 146.015 ;
        RECT 16.890 145.455 17.905 145.655 ;
        RECT 18.205 145.495 18.375 145.825 ;
        RECT 18.545 145.275 18.875 145.655 ;
        RECT 19.090 145.535 19.315 147.655 ;
        RECT 19.485 147.325 19.815 147.825 ;
        RECT 19.985 147.155 20.155 147.655 ;
        RECT 19.490 146.985 20.155 147.155 ;
        RECT 19.490 145.995 19.720 146.985 ;
        RECT 19.890 146.165 20.240 146.815 ;
        RECT 20.455 146.685 20.685 147.825 ;
        RECT 20.855 146.675 21.185 147.655 ;
        RECT 21.355 146.685 21.565 147.825 ;
        RECT 21.795 147.065 22.310 147.475 ;
        RECT 22.545 147.065 22.715 147.825 ;
        RECT 22.885 147.485 24.915 147.655 ;
        RECT 20.435 146.265 20.765 146.515 ;
        RECT 19.490 145.825 20.155 145.995 ;
        RECT 19.485 145.275 19.815 145.655 ;
        RECT 19.985 145.535 20.155 145.825 ;
        RECT 20.455 145.275 20.685 146.095 ;
        RECT 20.935 146.075 21.185 146.675 ;
        RECT 21.795 146.255 22.135 147.065 ;
        RECT 22.885 146.820 23.055 147.485 ;
        RECT 23.450 147.145 24.575 147.315 ;
        RECT 22.305 146.630 23.055 146.820 ;
        RECT 23.225 146.805 24.235 146.975 ;
        RECT 20.855 145.445 21.185 146.075 ;
        RECT 21.355 145.275 21.565 146.095 ;
        RECT 21.795 146.085 23.025 146.255 ;
        RECT 22.070 145.480 22.315 146.085 ;
        RECT 22.535 145.275 23.045 145.810 ;
        RECT 23.225 145.445 23.415 146.805 ;
        RECT 23.585 146.465 23.860 146.605 ;
        RECT 23.585 146.295 23.865 146.465 ;
        RECT 23.585 145.445 23.860 146.295 ;
        RECT 24.065 146.005 24.235 146.805 ;
        RECT 24.405 146.015 24.575 147.145 ;
        RECT 24.745 146.515 24.915 147.485 ;
        RECT 25.085 146.685 25.255 147.825 ;
        RECT 25.425 146.685 25.760 147.655 ;
        RECT 24.745 146.185 24.940 146.515 ;
        RECT 25.165 146.185 25.420 146.515 ;
        RECT 25.165 146.015 25.335 146.185 ;
        RECT 25.590 146.015 25.760 146.685 ;
        RECT 25.935 146.660 26.225 147.825 ;
        RECT 26.945 146.895 27.115 147.655 ;
        RECT 27.295 147.065 27.625 147.825 ;
        RECT 26.945 146.725 27.610 146.895 ;
        RECT 27.795 146.750 28.065 147.655 ;
        RECT 27.440 146.580 27.610 146.725 ;
        RECT 26.875 146.175 27.205 146.545 ;
        RECT 27.440 146.250 27.725 146.580 ;
        RECT 24.405 145.845 25.335 146.015 ;
        RECT 24.405 145.810 24.580 145.845 ;
        RECT 24.050 145.445 24.580 145.810 ;
        RECT 25.005 145.275 25.335 145.675 ;
        RECT 25.505 145.445 25.760 146.015 ;
        RECT 25.935 145.275 26.225 146.000 ;
        RECT 27.440 145.995 27.610 146.250 ;
        RECT 26.945 145.825 27.610 145.995 ;
        RECT 27.895 145.950 28.065 146.750 ;
        RECT 28.695 146.735 32.205 147.825 ;
        RECT 28.695 146.215 30.385 146.735 ;
        RECT 32.375 146.685 32.645 147.655 ;
        RECT 32.855 147.025 33.135 147.825 ;
        RECT 33.305 147.315 34.960 147.605 ;
        RECT 33.370 146.975 34.960 147.145 ;
        RECT 33.370 146.855 33.540 146.975 ;
        RECT 32.815 146.685 33.540 146.855 ;
        RECT 30.555 146.045 32.205 146.565 ;
        RECT 26.945 145.445 27.115 145.825 ;
        RECT 27.295 145.275 27.625 145.655 ;
        RECT 27.805 145.445 28.065 145.950 ;
        RECT 28.695 145.275 32.205 146.045 ;
        RECT 32.375 145.950 32.545 146.685 ;
        RECT 32.815 146.515 32.985 146.685 ;
        RECT 32.715 146.185 32.985 146.515 ;
        RECT 33.155 146.185 33.560 146.515 ;
        RECT 33.730 146.185 34.440 146.805 ;
        RECT 34.640 146.685 34.960 146.975 ;
        RECT 35.340 146.855 35.670 147.655 ;
        RECT 35.840 147.025 36.170 147.825 ;
        RECT 36.470 146.855 36.800 147.655 ;
        RECT 37.445 147.025 37.695 147.825 ;
        RECT 35.340 146.685 37.775 146.855 ;
        RECT 37.965 146.685 38.135 147.825 ;
        RECT 38.305 146.685 38.645 147.655 ;
        RECT 32.815 146.015 32.985 146.185 ;
        RECT 32.375 145.605 32.645 145.950 ;
        RECT 32.815 145.845 34.425 146.015 ;
        RECT 34.610 145.945 34.960 146.515 ;
        RECT 35.135 146.265 35.485 146.515 ;
        RECT 35.670 146.055 35.840 146.685 ;
        RECT 36.010 146.265 36.340 146.465 ;
        RECT 36.510 146.265 36.840 146.465 ;
        RECT 37.010 146.265 37.430 146.465 ;
        RECT 37.605 146.435 37.775 146.685 ;
        RECT 37.605 146.265 38.300 146.435 ;
        RECT 32.835 145.275 33.215 145.675 ;
        RECT 33.385 145.495 33.555 145.845 ;
        RECT 33.725 145.275 34.055 145.675 ;
        RECT 34.255 145.495 34.425 145.845 ;
        RECT 34.625 145.275 34.955 145.775 ;
        RECT 35.340 145.445 35.840 146.055 ;
        RECT 36.470 145.925 37.695 146.095 ;
        RECT 38.470 146.075 38.645 146.685 ;
        RECT 38.815 146.735 40.485 147.825 ;
        RECT 40.660 147.390 46.005 147.825 ;
        RECT 38.815 146.215 39.565 146.735 ;
        RECT 36.470 145.445 36.800 145.925 ;
        RECT 36.970 145.275 37.195 145.735 ;
        RECT 37.365 145.445 37.695 145.925 ;
        RECT 37.885 145.275 38.135 146.075 ;
        RECT 38.305 145.445 38.645 146.075 ;
        RECT 39.735 146.045 40.485 146.565 ;
        RECT 42.250 146.140 42.600 147.390 ;
        RECT 46.215 146.685 46.445 147.825 ;
        RECT 46.615 146.675 46.945 147.655 ;
        RECT 47.115 146.685 47.325 147.825 ;
        RECT 47.555 147.065 48.070 147.475 ;
        RECT 48.305 147.065 48.475 147.825 ;
        RECT 48.645 147.485 50.675 147.655 ;
        RECT 38.815 145.275 40.485 146.045 ;
        RECT 44.080 145.820 44.420 146.650 ;
        RECT 46.195 146.265 46.525 146.515 ;
        RECT 40.660 145.275 46.005 145.820 ;
        RECT 46.215 145.275 46.445 146.095 ;
        RECT 46.695 146.075 46.945 146.675 ;
        RECT 47.555 146.255 47.895 147.065 ;
        RECT 48.645 146.820 48.815 147.485 ;
        RECT 49.210 147.145 50.335 147.315 ;
        RECT 48.065 146.630 48.815 146.820 ;
        RECT 48.985 146.805 49.995 146.975 ;
        RECT 46.615 145.445 46.945 146.075 ;
        RECT 47.115 145.275 47.325 146.095 ;
        RECT 47.555 146.085 48.785 146.255 ;
        RECT 47.830 145.480 48.075 146.085 ;
        RECT 48.295 145.275 48.805 145.810 ;
        RECT 48.985 145.445 49.175 146.805 ;
        RECT 49.345 146.125 49.620 146.605 ;
        RECT 49.345 145.955 49.625 146.125 ;
        RECT 49.825 146.005 49.995 146.805 ;
        RECT 50.165 146.015 50.335 147.145 ;
        RECT 50.505 146.515 50.675 147.485 ;
        RECT 50.845 146.685 51.015 147.825 ;
        RECT 51.185 146.685 51.520 147.655 ;
        RECT 50.505 146.185 50.700 146.515 ;
        RECT 50.925 146.185 51.180 146.515 ;
        RECT 50.925 146.015 51.095 146.185 ;
        RECT 51.350 146.015 51.520 146.685 ;
        RECT 51.695 146.660 51.985 147.825 ;
        RECT 52.155 146.685 52.495 147.655 ;
        RECT 52.665 146.685 52.835 147.825 ;
        RECT 53.105 147.025 53.355 147.825 ;
        RECT 54.000 146.855 54.330 147.655 ;
        RECT 54.630 147.025 54.960 147.825 ;
        RECT 55.130 146.855 55.460 147.655 ;
        RECT 53.025 146.685 55.460 146.855 ;
        RECT 56.295 146.735 59.805 147.825 ;
        RECT 60.065 147.080 60.335 147.825 ;
        RECT 60.965 147.820 67.240 147.825 ;
        RECT 60.505 146.910 60.795 147.650 ;
        RECT 60.965 147.095 61.220 147.820 ;
        RECT 61.405 146.925 61.665 147.650 ;
        RECT 61.835 147.095 62.080 147.820 ;
        RECT 62.265 146.925 62.525 147.650 ;
        RECT 62.695 147.095 62.940 147.820 ;
        RECT 63.125 146.925 63.385 147.650 ;
        RECT 63.555 147.095 63.800 147.820 ;
        RECT 63.970 146.925 64.230 147.650 ;
        RECT 64.400 147.095 64.660 147.820 ;
        RECT 64.830 146.925 65.090 147.650 ;
        RECT 65.260 147.095 65.520 147.820 ;
        RECT 65.690 146.925 65.950 147.650 ;
        RECT 66.120 147.095 66.380 147.820 ;
        RECT 66.550 146.925 66.810 147.650 ;
        RECT 66.980 147.025 67.240 147.820 ;
        RECT 61.405 146.910 66.810 146.925 ;
        RECT 49.345 145.445 49.620 145.955 ;
        RECT 50.165 145.845 51.095 146.015 ;
        RECT 50.165 145.810 50.340 145.845 ;
        RECT 49.810 145.445 50.340 145.810 ;
        RECT 50.765 145.275 51.095 145.675 ;
        RECT 51.265 145.445 51.520 146.015 ;
        RECT 52.155 146.075 52.330 146.685 ;
        RECT 53.025 146.435 53.195 146.685 ;
        RECT 52.500 146.265 53.195 146.435 ;
        RECT 53.370 146.265 53.790 146.465 ;
        RECT 53.960 146.265 54.290 146.465 ;
        RECT 54.460 146.265 54.790 146.465 ;
        RECT 51.695 145.275 51.985 146.000 ;
        RECT 52.155 145.445 52.495 146.075 ;
        RECT 52.665 145.275 52.915 146.075 ;
        RECT 53.105 145.925 54.330 146.095 ;
        RECT 53.105 145.445 53.435 145.925 ;
        RECT 53.605 145.275 53.830 145.735 ;
        RECT 54.000 145.445 54.330 145.925 ;
        RECT 54.960 146.055 55.130 146.685 ;
        RECT 55.315 146.265 55.665 146.515 ;
        RECT 56.295 146.215 57.985 146.735 ;
        RECT 60.065 146.685 66.810 146.910 ;
        RECT 54.960 145.445 55.460 146.055 ;
        RECT 58.155 146.045 59.805 146.565 ;
        RECT 56.295 145.275 59.805 146.045 ;
        RECT 60.065 146.095 61.230 146.685 ;
        RECT 67.410 146.515 67.660 147.650 ;
        RECT 67.840 147.015 68.100 147.825 ;
        RECT 68.275 146.515 68.520 147.655 ;
        RECT 68.700 147.015 68.995 147.825 ;
        RECT 69.725 146.895 69.895 147.655 ;
        RECT 70.110 147.065 70.440 147.825 ;
        RECT 69.725 146.725 70.440 146.895 ;
        RECT 70.610 146.750 70.865 147.655 ;
        RECT 61.400 146.265 68.520 146.515 ;
        RECT 60.065 145.925 66.810 146.095 ;
        RECT 60.065 145.275 60.365 145.755 ;
        RECT 60.535 145.470 60.795 145.925 ;
        RECT 60.965 145.275 61.225 145.755 ;
        RECT 61.405 145.470 61.665 145.925 ;
        RECT 61.835 145.275 62.085 145.755 ;
        RECT 62.265 145.470 62.525 145.925 ;
        RECT 62.695 145.275 62.945 145.755 ;
        RECT 63.125 145.470 63.385 145.925 ;
        RECT 63.555 145.275 63.800 145.755 ;
        RECT 63.970 145.470 64.245 145.925 ;
        RECT 64.415 145.275 64.660 145.755 ;
        RECT 64.830 145.470 65.090 145.925 ;
        RECT 65.260 145.275 65.520 145.755 ;
        RECT 65.690 145.470 65.950 145.925 ;
        RECT 66.120 145.275 66.380 145.755 ;
        RECT 66.550 145.470 66.810 145.925 ;
        RECT 66.980 145.275 67.240 145.835 ;
        RECT 67.410 145.455 67.660 146.265 ;
        RECT 67.840 145.275 68.100 145.800 ;
        RECT 68.270 145.455 68.520 146.265 ;
        RECT 68.690 145.955 69.005 146.515 ;
        RECT 69.635 146.175 69.990 146.545 ;
        RECT 70.270 146.515 70.440 146.725 ;
        RECT 70.270 146.185 70.525 146.515 ;
        RECT 70.270 145.995 70.440 146.185 ;
        RECT 70.695 146.020 70.865 146.750 ;
        RECT 71.040 146.675 71.300 147.825 ;
        RECT 71.940 147.390 77.285 147.825 ;
        RECT 73.530 146.140 73.880 147.390 ;
        RECT 77.455 146.660 77.745 147.825 ;
        RECT 77.915 146.685 78.185 147.655 ;
        RECT 78.395 147.025 78.675 147.825 ;
        RECT 78.845 147.315 80.500 147.605 ;
        RECT 78.910 146.975 80.500 147.145 ;
        RECT 78.910 146.855 79.080 146.975 ;
        RECT 78.355 146.685 79.080 146.855 ;
        RECT 69.725 145.825 70.440 145.995 ;
        RECT 68.700 145.275 69.005 145.785 ;
        RECT 69.725 145.445 69.895 145.825 ;
        RECT 70.110 145.275 70.440 145.655 ;
        RECT 70.610 145.445 70.865 146.020 ;
        RECT 71.040 145.275 71.300 146.115 ;
        RECT 75.360 145.820 75.700 146.650 ;
        RECT 71.940 145.275 77.285 145.820 ;
        RECT 77.455 145.275 77.745 146.000 ;
        RECT 77.915 145.950 78.085 146.685 ;
        RECT 78.355 146.515 78.525 146.685 ;
        RECT 78.255 146.185 78.525 146.515 ;
        RECT 78.695 146.185 79.100 146.515 ;
        RECT 79.270 146.185 79.980 146.805 ;
        RECT 80.180 146.685 80.500 146.975 ;
        RECT 81.135 146.735 83.725 147.825 ;
        RECT 78.355 146.015 78.525 146.185 ;
        RECT 77.915 145.605 78.185 145.950 ;
        RECT 78.355 145.845 79.965 146.015 ;
        RECT 80.150 145.945 80.500 146.515 ;
        RECT 81.135 146.215 82.345 146.735 ;
        RECT 83.955 146.685 84.165 147.825 ;
        RECT 84.335 146.675 84.665 147.655 ;
        RECT 84.835 146.685 85.065 147.825 ;
        RECT 85.275 147.065 85.790 147.475 ;
        RECT 86.025 147.065 86.195 147.825 ;
        RECT 86.365 147.485 88.395 147.655 ;
        RECT 82.515 146.045 83.725 146.565 ;
        RECT 78.375 145.275 78.755 145.675 ;
        RECT 78.925 145.495 79.095 145.845 ;
        RECT 79.265 145.275 79.595 145.675 ;
        RECT 79.795 145.495 79.965 145.845 ;
        RECT 80.165 145.275 80.495 145.775 ;
        RECT 81.135 145.275 83.725 146.045 ;
        RECT 83.955 145.275 84.165 146.095 ;
        RECT 84.335 146.075 84.585 146.675 ;
        RECT 84.755 146.265 85.085 146.515 ;
        RECT 85.275 146.255 85.615 147.065 ;
        RECT 86.365 146.820 86.535 147.485 ;
        RECT 86.930 147.145 88.055 147.315 ;
        RECT 85.785 146.630 86.535 146.820 ;
        RECT 86.705 146.805 87.715 146.975 ;
        RECT 84.335 145.445 84.665 146.075 ;
        RECT 84.835 145.275 85.065 146.095 ;
        RECT 85.275 146.085 86.505 146.255 ;
        RECT 85.550 145.480 85.795 146.085 ;
        RECT 86.015 145.275 86.525 145.810 ;
        RECT 86.705 145.445 86.895 146.805 ;
        RECT 87.065 145.785 87.340 146.605 ;
        RECT 87.545 146.005 87.715 146.805 ;
        RECT 87.885 146.015 88.055 147.145 ;
        RECT 88.225 146.515 88.395 147.485 ;
        RECT 88.565 146.685 88.735 147.825 ;
        RECT 88.905 146.685 89.240 147.655 ;
        RECT 88.225 146.185 88.420 146.515 ;
        RECT 88.645 146.185 88.900 146.515 ;
        RECT 88.645 146.015 88.815 146.185 ;
        RECT 89.070 146.015 89.240 146.685 ;
        RECT 87.885 145.845 88.815 146.015 ;
        RECT 87.885 145.810 88.060 145.845 ;
        RECT 87.065 145.615 87.345 145.785 ;
        RECT 87.065 145.445 87.340 145.615 ;
        RECT 87.530 145.445 88.060 145.810 ;
        RECT 88.485 145.275 88.815 145.675 ;
        RECT 88.985 145.445 89.240 146.015 ;
        RECT 89.880 146.635 90.135 147.515 ;
        RECT 90.305 146.685 90.610 147.825 ;
        RECT 90.950 147.445 91.280 147.825 ;
        RECT 91.460 147.275 91.630 147.565 ;
        RECT 91.800 147.365 92.050 147.825 ;
        RECT 90.830 147.105 91.630 147.275 ;
        RECT 92.220 147.315 93.090 147.655 ;
        RECT 89.880 145.985 90.090 146.635 ;
        RECT 90.830 146.515 91.000 147.105 ;
        RECT 92.220 146.935 92.390 147.315 ;
        RECT 93.325 147.195 93.495 147.655 ;
        RECT 93.665 147.365 94.035 147.825 ;
        RECT 94.330 147.225 94.500 147.565 ;
        RECT 94.670 147.395 95.000 147.825 ;
        RECT 95.235 147.225 95.405 147.565 ;
        RECT 91.170 146.765 92.390 146.935 ;
        RECT 92.560 146.855 93.020 147.145 ;
        RECT 93.325 147.025 93.885 147.195 ;
        RECT 94.330 147.055 95.405 147.225 ;
        RECT 95.575 147.325 96.255 147.655 ;
        RECT 96.470 147.325 96.720 147.655 ;
        RECT 96.890 147.365 97.140 147.825 ;
        RECT 93.715 146.885 93.885 147.025 ;
        RECT 92.560 146.845 93.525 146.855 ;
        RECT 92.220 146.675 92.390 146.765 ;
        RECT 92.850 146.685 93.525 146.845 ;
        RECT 90.260 146.485 91.000 146.515 ;
        RECT 90.260 146.185 91.175 146.485 ;
        RECT 90.850 146.010 91.175 146.185 ;
        RECT 89.880 145.455 90.135 145.985 ;
        RECT 90.305 145.275 90.610 145.735 ;
        RECT 90.855 145.655 91.175 146.010 ;
        RECT 91.345 146.225 91.885 146.595 ;
        RECT 92.220 146.505 92.625 146.675 ;
        RECT 91.345 145.825 91.585 146.225 ;
        RECT 92.065 146.055 92.285 146.335 ;
        RECT 91.755 145.885 92.285 146.055 ;
        RECT 91.755 145.655 91.925 145.885 ;
        RECT 92.455 145.725 92.625 146.505 ;
        RECT 92.795 145.895 93.145 146.515 ;
        RECT 93.315 145.895 93.525 146.685 ;
        RECT 93.715 146.715 95.215 146.885 ;
        RECT 93.715 146.025 93.885 146.715 ;
        RECT 95.575 146.545 95.745 147.325 ;
        RECT 96.550 147.195 96.720 147.325 ;
        RECT 94.055 146.375 95.745 146.545 ;
        RECT 95.915 146.765 96.380 147.155 ;
        RECT 96.550 147.025 96.945 147.195 ;
        RECT 94.055 146.195 94.225 146.375 ;
        RECT 90.855 145.485 91.925 145.655 ;
        RECT 92.095 145.275 92.285 145.715 ;
        RECT 92.455 145.445 93.405 145.725 ;
        RECT 93.715 145.635 93.975 146.025 ;
        RECT 94.395 145.955 95.185 146.205 ;
        RECT 93.625 145.465 93.975 145.635 ;
        RECT 94.185 145.275 94.515 145.735 ;
        RECT 95.390 145.665 95.560 146.375 ;
        RECT 95.915 146.175 96.085 146.765 ;
        RECT 95.730 145.955 96.085 146.175 ;
        RECT 96.255 145.955 96.605 146.575 ;
        RECT 96.775 145.665 96.945 147.025 ;
        RECT 97.310 146.855 97.635 147.640 ;
        RECT 97.115 145.805 97.575 146.855 ;
        RECT 95.390 145.495 96.245 145.665 ;
        RECT 96.450 145.495 96.945 145.665 ;
        RECT 97.115 145.275 97.445 145.635 ;
        RECT 97.805 145.535 97.975 147.655 ;
        RECT 98.145 147.325 98.475 147.825 ;
        RECT 98.645 147.155 98.900 147.655 ;
        RECT 98.150 146.985 98.900 147.155 ;
        RECT 98.150 145.995 98.380 146.985 ;
        RECT 98.550 146.165 98.900 146.815 ;
        RECT 99.535 146.735 103.045 147.825 ;
        RECT 99.535 146.215 101.225 146.735 ;
        RECT 103.215 146.660 103.505 147.825 ;
        RECT 103.675 146.685 103.945 147.655 ;
        RECT 104.155 147.025 104.435 147.825 ;
        RECT 104.605 147.315 106.260 147.605 ;
        RECT 104.670 146.975 106.260 147.145 ;
        RECT 104.670 146.855 104.840 146.975 ;
        RECT 104.115 146.685 104.840 146.855 ;
        RECT 101.395 146.045 103.045 146.565 ;
        RECT 98.150 145.825 98.900 145.995 ;
        RECT 98.145 145.275 98.475 145.655 ;
        RECT 98.645 145.535 98.900 145.825 ;
        RECT 99.535 145.275 103.045 146.045 ;
        RECT 103.215 145.275 103.505 146.000 ;
        RECT 103.675 145.950 103.845 146.685 ;
        RECT 104.115 146.515 104.285 146.685 ;
        RECT 105.030 146.635 105.745 146.805 ;
        RECT 105.940 146.685 106.260 146.975 ;
        RECT 106.435 146.685 106.775 147.655 ;
        RECT 106.945 146.685 107.115 147.825 ;
        RECT 107.385 147.025 107.635 147.825 ;
        RECT 108.280 146.855 108.610 147.655 ;
        RECT 108.910 147.025 109.240 147.825 ;
        RECT 109.410 146.855 109.740 147.655 ;
        RECT 107.305 146.685 109.740 146.855 ;
        RECT 110.115 146.685 110.455 147.655 ;
        RECT 110.625 146.685 110.795 147.825 ;
        RECT 111.065 147.025 111.315 147.825 ;
        RECT 111.960 146.855 112.290 147.655 ;
        RECT 112.590 147.025 112.920 147.825 ;
        RECT 113.090 146.855 113.420 147.655 ;
        RECT 110.985 146.685 113.420 146.855 ;
        RECT 114.255 146.735 116.845 147.825 ;
        RECT 117.020 147.390 122.365 147.825 ;
        RECT 122.540 147.390 127.885 147.825 ;
        RECT 104.015 146.185 104.285 146.515 ;
        RECT 104.455 146.185 104.860 146.515 ;
        RECT 105.030 146.185 105.740 146.635 ;
        RECT 104.115 146.015 104.285 146.185 ;
        RECT 103.675 145.605 103.945 145.950 ;
        RECT 104.115 145.845 105.725 146.015 ;
        RECT 105.910 145.945 106.260 146.515 ;
        RECT 106.435 146.075 106.610 146.685 ;
        RECT 107.305 146.435 107.475 146.685 ;
        RECT 106.780 146.265 107.475 146.435 ;
        RECT 107.650 146.265 108.070 146.465 ;
        RECT 108.240 146.265 108.570 146.465 ;
        RECT 108.740 146.265 109.070 146.465 ;
        RECT 104.135 145.275 104.515 145.675 ;
        RECT 104.685 145.495 104.855 145.845 ;
        RECT 105.025 145.275 105.355 145.675 ;
        RECT 105.555 145.495 105.725 145.845 ;
        RECT 105.925 145.275 106.255 145.775 ;
        RECT 106.435 145.445 106.775 146.075 ;
        RECT 106.945 145.275 107.195 146.075 ;
        RECT 107.385 145.925 108.610 146.095 ;
        RECT 107.385 145.445 107.715 145.925 ;
        RECT 107.885 145.275 108.110 145.735 ;
        RECT 108.280 145.445 108.610 145.925 ;
        RECT 109.240 146.055 109.410 146.685 ;
        RECT 109.595 146.265 109.945 146.515 ;
        RECT 110.115 146.125 110.290 146.685 ;
        RECT 110.985 146.435 111.155 146.685 ;
        RECT 110.460 146.265 111.155 146.435 ;
        RECT 111.330 146.265 111.750 146.465 ;
        RECT 111.920 146.265 112.250 146.465 ;
        RECT 112.420 146.265 112.750 146.465 ;
        RECT 110.115 146.075 110.345 146.125 ;
        RECT 109.240 145.445 109.740 146.055 ;
        RECT 110.115 145.445 110.455 146.075 ;
        RECT 110.625 145.275 110.875 146.075 ;
        RECT 111.065 145.925 112.290 146.095 ;
        RECT 111.065 145.445 111.395 145.925 ;
        RECT 111.565 145.275 111.790 145.735 ;
        RECT 111.960 145.445 112.290 145.925 ;
        RECT 112.920 146.055 113.090 146.685 ;
        RECT 113.275 146.265 113.625 146.515 ;
        RECT 114.255 146.215 115.465 146.735 ;
        RECT 112.920 145.445 113.420 146.055 ;
        RECT 115.635 146.045 116.845 146.565 ;
        RECT 118.610 146.140 118.960 147.390 ;
        RECT 114.255 145.275 116.845 146.045 ;
        RECT 120.440 145.820 120.780 146.650 ;
        RECT 124.130 146.140 124.480 147.390 ;
        RECT 128.055 146.735 129.265 147.825 ;
        RECT 125.960 145.820 126.300 146.650 ;
        RECT 128.055 146.195 128.575 146.735 ;
        RECT 128.745 146.025 129.265 146.565 ;
        RECT 117.020 145.275 122.365 145.820 ;
        RECT 122.540 145.275 127.885 145.820 ;
        RECT 128.055 145.275 129.265 146.025 ;
        RECT 9.290 145.105 129.350 145.275 ;
        RECT 9.375 144.355 10.585 145.105 ;
        RECT 9.375 143.815 9.895 144.355 ;
        RECT 11.215 144.335 12.885 145.105 ;
        RECT 13.055 144.380 13.345 145.105 ;
        RECT 13.515 144.355 14.725 145.105 ;
        RECT 14.985 144.555 15.155 144.935 ;
        RECT 15.335 144.725 15.665 145.105 ;
        RECT 14.985 144.385 15.650 144.555 ;
        RECT 15.845 144.430 16.105 144.935 ;
        RECT 10.065 143.645 10.585 144.185 ;
        RECT 9.375 142.555 10.585 143.645 ;
        RECT 11.215 143.645 11.965 144.165 ;
        RECT 12.135 143.815 12.885 144.335 ;
        RECT 11.215 142.555 12.885 143.645 ;
        RECT 13.055 142.555 13.345 143.720 ;
        RECT 13.515 143.645 14.035 144.185 ;
        RECT 14.205 143.815 14.725 144.355 ;
        RECT 14.915 143.835 15.245 144.205 ;
        RECT 15.480 144.130 15.650 144.385 ;
        RECT 15.480 143.800 15.765 144.130 ;
        RECT 15.480 143.655 15.650 143.800 ;
        RECT 13.515 142.555 14.725 143.645 ;
        RECT 14.985 143.485 15.650 143.655 ;
        RECT 15.935 143.630 16.105 144.430 ;
        RECT 14.985 142.725 15.155 143.485 ;
        RECT 15.335 142.555 15.665 143.315 ;
        RECT 15.835 142.725 16.105 143.630 ;
        RECT 16.280 144.365 16.535 144.935 ;
        RECT 16.705 144.705 17.035 145.105 ;
        RECT 17.460 144.570 17.990 144.935 ;
        RECT 17.460 144.535 17.635 144.570 ;
        RECT 16.705 144.365 17.635 144.535 ;
        RECT 18.180 144.425 18.455 144.935 ;
        RECT 16.280 143.695 16.450 144.365 ;
        RECT 16.705 144.195 16.875 144.365 ;
        RECT 16.620 143.865 16.875 144.195 ;
        RECT 17.100 143.865 17.295 144.195 ;
        RECT 16.280 142.725 16.615 143.695 ;
        RECT 16.785 142.555 16.955 143.695 ;
        RECT 17.125 142.895 17.295 143.865 ;
        RECT 17.465 143.235 17.635 144.365 ;
        RECT 17.805 143.575 17.975 144.375 ;
        RECT 18.175 144.255 18.455 144.425 ;
        RECT 18.180 143.775 18.455 144.255 ;
        RECT 18.625 143.575 18.815 144.935 ;
        RECT 18.995 144.570 19.505 145.105 ;
        RECT 19.725 144.295 19.970 144.900 ;
        RECT 20.790 144.425 21.045 144.925 ;
        RECT 21.225 144.645 21.510 145.105 ;
        RECT 20.705 144.395 21.045 144.425 ;
        RECT 19.015 144.125 20.245 144.295 ;
        RECT 20.705 144.255 20.970 144.395 ;
        RECT 17.805 143.405 18.815 143.575 ;
        RECT 18.985 143.560 19.735 143.750 ;
        RECT 17.465 143.065 18.590 143.235 ;
        RECT 18.985 142.895 19.155 143.560 ;
        RECT 19.905 143.315 20.245 144.125 ;
        RECT 17.125 142.725 19.155 142.895 ;
        RECT 19.325 142.555 19.495 143.315 ;
        RECT 19.730 142.905 20.245 143.315 ;
        RECT 20.790 143.535 20.970 144.255 ;
        RECT 21.690 144.195 21.940 144.845 ;
        RECT 21.140 143.865 21.940 144.195 ;
        RECT 20.790 142.865 21.045 143.535 ;
        RECT 21.225 142.555 21.510 143.355 ;
        RECT 21.690 143.275 21.940 143.865 ;
        RECT 22.140 144.510 22.460 144.840 ;
        RECT 22.640 144.625 23.300 145.105 ;
        RECT 23.500 144.715 24.350 144.885 ;
        RECT 22.140 143.615 22.330 144.510 ;
        RECT 22.650 144.185 23.310 144.455 ;
        RECT 22.980 144.125 23.310 144.185 ;
        RECT 22.500 143.955 22.830 144.015 ;
        RECT 23.500 143.955 23.670 144.715 ;
        RECT 24.910 144.645 25.230 145.105 ;
        RECT 25.430 144.465 25.680 144.895 ;
        RECT 25.970 144.665 26.380 145.105 ;
        RECT 26.550 144.725 27.565 144.925 ;
        RECT 23.840 144.295 25.090 144.465 ;
        RECT 23.840 144.175 24.170 144.295 ;
        RECT 22.500 143.785 24.400 143.955 ;
        RECT 22.140 143.445 24.060 143.615 ;
        RECT 22.140 143.425 22.460 143.445 ;
        RECT 21.690 142.765 22.020 143.275 ;
        RECT 22.290 142.815 22.460 143.425 ;
        RECT 24.230 143.275 24.400 143.785 ;
        RECT 24.570 143.715 24.750 144.125 ;
        RECT 24.920 143.535 25.090 144.295 ;
        RECT 22.630 142.555 22.960 143.245 ;
        RECT 23.190 143.105 24.400 143.275 ;
        RECT 24.570 143.225 25.090 143.535 ;
        RECT 25.260 144.125 25.680 144.465 ;
        RECT 25.970 144.125 26.380 144.455 ;
        RECT 25.260 143.355 25.450 144.125 ;
        RECT 26.550 143.995 26.720 144.725 ;
        RECT 27.865 144.555 28.035 144.885 ;
        RECT 28.205 144.725 28.535 145.105 ;
        RECT 26.890 144.175 27.240 144.545 ;
        RECT 26.550 143.955 26.970 143.995 ;
        RECT 25.620 143.785 26.970 143.955 ;
        RECT 25.620 143.625 25.870 143.785 ;
        RECT 26.380 143.355 26.630 143.615 ;
        RECT 25.260 143.105 26.630 143.355 ;
        RECT 23.190 142.815 23.430 143.105 ;
        RECT 24.230 143.025 24.400 143.105 ;
        RECT 23.630 142.555 24.050 142.935 ;
        RECT 24.230 142.775 24.860 143.025 ;
        RECT 25.330 142.555 25.660 142.935 ;
        RECT 25.830 142.815 26.000 143.105 ;
        RECT 26.800 142.940 26.970 143.785 ;
        RECT 27.420 143.615 27.640 144.485 ;
        RECT 27.865 144.365 28.560 144.555 ;
        RECT 27.140 143.235 27.640 143.615 ;
        RECT 27.810 143.565 28.220 144.185 ;
        RECT 28.390 143.395 28.560 144.365 ;
        RECT 27.865 143.225 28.560 143.395 ;
        RECT 26.180 142.555 26.560 142.935 ;
        RECT 26.800 142.770 27.630 142.940 ;
        RECT 27.865 142.725 28.035 143.225 ;
        RECT 28.205 142.555 28.535 143.055 ;
        RECT 28.750 142.725 28.975 144.845 ;
        RECT 29.145 144.725 29.475 145.105 ;
        RECT 29.645 144.555 29.815 144.845 ;
        RECT 29.150 144.385 29.815 144.555 ;
        RECT 29.150 143.395 29.380 144.385 ;
        RECT 30.535 144.335 32.205 145.105 ;
        RECT 29.550 143.565 29.900 144.215 ;
        RECT 30.535 143.645 31.285 144.165 ;
        RECT 31.455 143.815 32.205 144.335 ;
        RECT 32.375 144.305 32.715 144.935 ;
        RECT 32.885 144.305 33.135 145.105 ;
        RECT 33.325 144.455 33.655 144.935 ;
        RECT 33.825 144.645 34.050 145.105 ;
        RECT 34.220 144.455 34.550 144.935 ;
        RECT 32.375 144.255 32.605 144.305 ;
        RECT 33.325 144.285 34.550 144.455 ;
        RECT 35.180 144.325 35.680 144.935 ;
        RECT 36.055 144.335 38.645 145.105 ;
        RECT 38.815 144.380 39.105 145.105 ;
        RECT 39.275 144.335 42.785 145.105 ;
        RECT 32.375 143.695 32.550 144.255 ;
        RECT 32.720 143.945 33.415 144.115 ;
        RECT 33.245 143.695 33.415 143.945 ;
        RECT 33.590 143.915 34.010 144.115 ;
        RECT 34.180 143.915 34.510 144.115 ;
        RECT 34.680 143.915 35.010 144.115 ;
        RECT 35.180 143.695 35.350 144.325 ;
        RECT 35.535 143.865 35.885 144.115 ;
        RECT 29.150 143.225 29.815 143.395 ;
        RECT 29.145 142.555 29.475 143.055 ;
        RECT 29.645 142.725 29.815 143.225 ;
        RECT 30.535 142.555 32.205 143.645 ;
        RECT 32.375 142.725 32.715 143.695 ;
        RECT 32.885 142.555 33.055 143.695 ;
        RECT 33.245 143.525 35.680 143.695 ;
        RECT 33.325 142.555 33.575 143.355 ;
        RECT 34.220 142.725 34.550 143.525 ;
        RECT 34.850 142.555 35.180 143.355 ;
        RECT 35.350 142.725 35.680 143.525 ;
        RECT 36.055 143.645 37.265 144.165 ;
        RECT 37.435 143.815 38.645 144.335 ;
        RECT 36.055 142.555 38.645 143.645 ;
        RECT 38.815 142.555 39.105 143.720 ;
        RECT 39.275 143.645 40.965 144.165 ;
        RECT 41.135 143.815 42.785 144.335 ;
        RECT 42.955 144.430 43.225 144.775 ;
        RECT 43.415 144.705 43.795 145.105 ;
        RECT 43.965 144.535 44.135 144.885 ;
        RECT 44.305 144.705 44.635 145.105 ;
        RECT 44.835 144.535 45.005 144.885 ;
        RECT 45.205 144.605 45.535 145.105 ;
        RECT 42.955 143.695 43.125 144.430 ;
        RECT 43.395 144.365 45.005 144.535 ;
        RECT 43.395 144.195 43.565 144.365 ;
        RECT 43.295 143.865 43.565 144.195 ;
        RECT 43.735 143.865 44.140 144.195 ;
        RECT 43.395 143.695 43.565 143.865 ;
        RECT 39.275 142.555 42.785 143.645 ;
        RECT 42.955 142.725 43.225 143.695 ;
        RECT 43.395 143.525 44.120 143.695 ;
        RECT 44.310 143.575 45.020 144.195 ;
        RECT 45.190 143.865 45.540 144.435 ;
        RECT 46.090 144.395 46.345 144.925 ;
        RECT 46.525 144.645 46.810 145.105 ;
        RECT 43.950 143.405 44.120 143.525 ;
        RECT 45.220 143.405 45.540 143.695 ;
        RECT 43.435 142.555 43.715 143.355 ;
        RECT 43.950 143.235 45.540 143.405 ;
        RECT 46.090 143.535 46.270 144.395 ;
        RECT 46.990 144.195 47.240 144.845 ;
        RECT 46.440 143.865 47.240 144.195 ;
        RECT 46.090 143.065 46.345 143.535 ;
        RECT 43.885 142.775 45.540 143.065 ;
        RECT 46.005 142.895 46.345 143.065 ;
        RECT 46.090 142.865 46.345 142.895 ;
        RECT 46.525 142.555 46.810 143.355 ;
        RECT 46.990 143.275 47.240 143.865 ;
        RECT 47.440 144.510 47.760 144.840 ;
        RECT 47.940 144.625 48.600 145.105 ;
        RECT 48.800 144.715 49.650 144.885 ;
        RECT 47.440 143.615 47.630 144.510 ;
        RECT 47.950 144.185 48.610 144.455 ;
        RECT 48.280 144.125 48.610 144.185 ;
        RECT 47.800 143.955 48.130 144.015 ;
        RECT 48.800 143.955 48.970 144.715 ;
        RECT 50.210 144.645 50.530 145.105 ;
        RECT 50.730 144.465 50.980 144.895 ;
        RECT 51.270 144.665 51.680 145.105 ;
        RECT 51.850 144.725 52.865 144.925 ;
        RECT 49.140 144.295 50.390 144.465 ;
        RECT 49.140 144.175 49.470 144.295 ;
        RECT 47.800 143.785 49.700 143.955 ;
        RECT 47.440 143.445 49.360 143.615 ;
        RECT 47.440 143.425 47.760 143.445 ;
        RECT 46.990 142.765 47.320 143.275 ;
        RECT 47.590 142.815 47.760 143.425 ;
        RECT 49.530 143.275 49.700 143.785 ;
        RECT 49.870 143.715 50.050 144.125 ;
        RECT 50.220 143.535 50.390 144.295 ;
        RECT 47.930 142.555 48.260 143.245 ;
        RECT 48.490 143.105 49.700 143.275 ;
        RECT 49.870 143.225 50.390 143.535 ;
        RECT 50.560 144.125 50.980 144.465 ;
        RECT 51.270 144.125 51.680 144.455 ;
        RECT 50.560 143.355 50.750 144.125 ;
        RECT 51.850 143.995 52.020 144.725 ;
        RECT 53.165 144.555 53.335 144.885 ;
        RECT 53.505 144.725 53.835 145.105 ;
        RECT 52.190 144.175 52.540 144.545 ;
        RECT 51.850 143.955 52.270 143.995 ;
        RECT 50.920 143.785 52.270 143.955 ;
        RECT 50.920 143.625 51.170 143.785 ;
        RECT 51.680 143.355 51.930 143.615 ;
        RECT 50.560 143.105 51.930 143.355 ;
        RECT 48.490 142.815 48.730 143.105 ;
        RECT 49.530 143.025 49.700 143.105 ;
        RECT 48.930 142.555 49.350 142.935 ;
        RECT 49.530 142.775 50.160 143.025 ;
        RECT 50.630 142.555 50.960 142.935 ;
        RECT 51.130 142.815 51.300 143.105 ;
        RECT 52.100 142.940 52.270 143.785 ;
        RECT 52.720 143.615 52.940 144.485 ;
        RECT 53.165 144.365 53.860 144.555 ;
        RECT 52.440 143.235 52.940 143.615 ;
        RECT 53.110 143.565 53.520 144.185 ;
        RECT 53.690 143.395 53.860 144.365 ;
        RECT 53.165 143.225 53.860 143.395 ;
        RECT 51.480 142.555 51.860 142.935 ;
        RECT 52.100 142.770 52.930 142.940 ;
        RECT 53.165 142.725 53.335 143.225 ;
        RECT 53.505 142.555 53.835 143.055 ;
        RECT 54.050 142.725 54.275 144.845 ;
        RECT 54.445 144.725 54.775 145.105 ;
        RECT 54.945 144.555 55.115 144.845 ;
        RECT 54.450 144.385 55.115 144.555 ;
        RECT 54.450 143.395 54.680 144.385 ;
        RECT 55.835 144.335 59.345 145.105 ;
        RECT 54.850 143.565 55.200 144.215 ;
        RECT 55.835 143.645 57.525 144.165 ;
        RECT 57.695 143.815 59.345 144.335 ;
        RECT 59.555 144.285 59.785 145.105 ;
        RECT 59.955 144.305 60.285 144.935 ;
        RECT 59.535 143.865 59.865 144.115 ;
        RECT 60.035 143.705 60.285 144.305 ;
        RECT 60.455 144.285 60.665 145.105 ;
        RECT 60.895 144.305 61.235 144.935 ;
        RECT 61.405 144.305 61.655 145.105 ;
        RECT 61.845 144.455 62.175 144.935 ;
        RECT 62.345 144.645 62.570 145.105 ;
        RECT 62.740 144.455 63.070 144.935 ;
        RECT 54.450 143.225 55.115 143.395 ;
        RECT 54.445 142.555 54.775 143.055 ;
        RECT 54.945 142.725 55.115 143.225 ;
        RECT 55.835 142.555 59.345 143.645 ;
        RECT 59.555 142.555 59.785 143.695 ;
        RECT 59.955 142.725 60.285 143.705 ;
        RECT 60.895 143.695 61.070 144.305 ;
        RECT 61.845 144.285 63.070 144.455 ;
        RECT 63.700 144.325 64.200 144.935 ;
        RECT 64.575 144.380 64.865 145.105 ;
        RECT 65.960 144.560 71.305 145.105 ;
        RECT 71.480 144.560 76.825 145.105 ;
        RECT 61.240 143.945 61.935 144.115 ;
        RECT 61.765 143.695 61.935 143.945 ;
        RECT 62.110 143.915 62.530 144.115 ;
        RECT 62.700 143.915 63.030 144.115 ;
        RECT 63.200 143.915 63.530 144.115 ;
        RECT 63.700 143.695 63.870 144.325 ;
        RECT 64.055 143.865 64.405 144.115 ;
        RECT 60.455 142.555 60.665 143.695 ;
        RECT 60.895 142.725 61.235 143.695 ;
        RECT 61.405 142.555 61.575 143.695 ;
        RECT 61.765 143.525 64.200 143.695 ;
        RECT 61.845 142.555 62.095 143.355 ;
        RECT 62.740 142.725 63.070 143.525 ;
        RECT 63.370 142.555 63.700 143.355 ;
        RECT 63.870 142.725 64.200 143.525 ;
        RECT 64.575 142.555 64.865 143.720 ;
        RECT 67.550 142.990 67.900 144.240 ;
        RECT 69.380 143.730 69.720 144.560 ;
        RECT 73.070 142.990 73.420 144.240 ;
        RECT 74.900 143.730 75.240 144.560 ;
        RECT 77.200 144.325 77.700 144.935 ;
        RECT 76.995 143.865 77.345 144.115 ;
        RECT 77.530 143.695 77.700 144.325 ;
        RECT 78.330 144.455 78.660 144.935 ;
        RECT 78.830 144.645 79.055 145.105 ;
        RECT 79.225 144.455 79.555 144.935 ;
        RECT 78.330 144.285 79.555 144.455 ;
        RECT 79.745 144.305 79.995 145.105 ;
        RECT 80.165 144.305 80.505 144.935 ;
        RECT 80.275 144.255 80.505 144.305 ;
        RECT 77.870 143.915 78.200 144.115 ;
        RECT 78.370 143.915 78.700 144.115 ;
        RECT 78.870 143.915 79.290 144.115 ;
        RECT 79.465 143.945 80.160 144.115 ;
        RECT 79.465 143.695 79.635 143.945 ;
        RECT 80.330 143.695 80.505 144.255 ;
        RECT 77.200 143.525 79.635 143.695 ;
        RECT 65.960 142.555 71.305 142.990 ;
        RECT 71.480 142.555 76.825 142.990 ;
        RECT 77.200 142.725 77.530 143.525 ;
        RECT 77.700 142.555 78.030 143.355 ;
        RECT 78.330 142.725 78.660 143.525 ;
        RECT 79.305 142.555 79.555 143.355 ;
        RECT 79.825 142.555 79.995 143.695 ;
        RECT 80.165 142.725 80.505 143.695 ;
        RECT 81.050 144.395 81.305 144.925 ;
        RECT 81.485 144.645 81.770 145.105 ;
        RECT 81.050 143.535 81.230 144.395 ;
        RECT 81.950 144.195 82.200 144.845 ;
        RECT 81.400 143.865 82.200 144.195 ;
        RECT 81.050 143.065 81.305 143.535 ;
        RECT 80.965 142.895 81.305 143.065 ;
        RECT 81.050 142.865 81.305 142.895 ;
        RECT 81.485 142.555 81.770 143.355 ;
        RECT 81.950 143.275 82.200 143.865 ;
        RECT 82.400 144.510 82.720 144.840 ;
        RECT 82.900 144.625 83.560 145.105 ;
        RECT 83.760 144.715 84.610 144.885 ;
        RECT 82.400 143.615 82.590 144.510 ;
        RECT 82.910 144.185 83.570 144.455 ;
        RECT 83.240 144.125 83.570 144.185 ;
        RECT 82.760 143.955 83.090 144.015 ;
        RECT 83.760 143.955 83.930 144.715 ;
        RECT 85.170 144.645 85.490 145.105 ;
        RECT 85.690 144.465 85.940 144.895 ;
        RECT 86.230 144.665 86.640 145.105 ;
        RECT 86.810 144.725 87.825 144.925 ;
        RECT 84.100 144.295 85.350 144.465 ;
        RECT 84.100 144.175 84.430 144.295 ;
        RECT 82.760 143.785 84.660 143.955 ;
        RECT 82.400 143.445 84.320 143.615 ;
        RECT 82.400 143.425 82.720 143.445 ;
        RECT 81.950 142.765 82.280 143.275 ;
        RECT 82.550 142.815 82.720 143.425 ;
        RECT 84.490 143.275 84.660 143.785 ;
        RECT 84.830 143.715 85.010 144.125 ;
        RECT 85.180 143.535 85.350 144.295 ;
        RECT 82.890 142.555 83.220 143.245 ;
        RECT 83.450 143.105 84.660 143.275 ;
        RECT 84.830 143.225 85.350 143.535 ;
        RECT 85.520 144.125 85.940 144.465 ;
        RECT 86.230 144.125 86.640 144.455 ;
        RECT 85.520 143.355 85.710 144.125 ;
        RECT 86.810 143.995 86.980 144.725 ;
        RECT 88.125 144.555 88.295 144.885 ;
        RECT 88.465 144.725 88.795 145.105 ;
        RECT 87.150 144.175 87.500 144.545 ;
        RECT 86.810 143.955 87.230 143.995 ;
        RECT 85.880 143.785 87.230 143.955 ;
        RECT 85.880 143.625 86.130 143.785 ;
        RECT 86.640 143.355 86.890 143.615 ;
        RECT 85.520 143.105 86.890 143.355 ;
        RECT 83.450 142.815 83.690 143.105 ;
        RECT 84.490 143.025 84.660 143.105 ;
        RECT 83.890 142.555 84.310 142.935 ;
        RECT 84.490 142.775 85.120 143.025 ;
        RECT 85.590 142.555 85.920 142.935 ;
        RECT 86.090 142.815 86.260 143.105 ;
        RECT 87.060 142.940 87.230 143.785 ;
        RECT 87.680 143.615 87.900 144.485 ;
        RECT 88.125 144.365 88.820 144.555 ;
        RECT 87.400 143.235 87.900 143.615 ;
        RECT 88.070 143.565 88.480 144.185 ;
        RECT 88.650 143.395 88.820 144.365 ;
        RECT 88.125 143.225 88.820 143.395 ;
        RECT 86.440 142.555 86.820 142.935 ;
        RECT 87.060 142.770 87.890 142.940 ;
        RECT 88.125 142.725 88.295 143.225 ;
        RECT 88.465 142.555 88.795 143.055 ;
        RECT 89.010 142.725 89.235 144.845 ;
        RECT 89.405 144.725 89.735 145.105 ;
        RECT 89.905 144.555 90.075 144.845 ;
        RECT 89.410 144.385 90.075 144.555 ;
        RECT 89.410 143.395 89.640 144.385 ;
        RECT 90.335 144.380 90.625 145.105 ;
        RECT 90.795 144.430 91.055 144.935 ;
        RECT 91.235 144.725 91.565 145.105 ;
        RECT 91.745 144.555 91.915 144.935 ;
        RECT 89.810 143.565 90.160 144.215 ;
        RECT 89.410 143.225 90.075 143.395 ;
        RECT 89.405 142.555 89.735 143.055 ;
        RECT 89.905 142.725 90.075 143.225 ;
        RECT 90.335 142.555 90.625 143.720 ;
        RECT 90.795 143.630 90.965 144.430 ;
        RECT 91.250 144.385 91.915 144.555 ;
        RECT 91.250 144.130 91.420 144.385 ;
        RECT 92.175 144.335 93.845 145.105 ;
        RECT 94.020 144.560 99.365 145.105 ;
        RECT 99.540 144.560 104.885 145.105 ;
        RECT 105.065 144.605 105.395 145.105 ;
        RECT 91.135 143.800 91.420 144.130 ;
        RECT 91.655 143.835 91.985 144.205 ;
        RECT 91.250 143.655 91.420 143.800 ;
        RECT 90.795 142.725 91.065 143.630 ;
        RECT 91.250 143.485 91.915 143.655 ;
        RECT 91.235 142.555 91.565 143.315 ;
        RECT 91.745 142.725 91.915 143.485 ;
        RECT 92.175 143.645 92.925 144.165 ;
        RECT 93.095 143.815 93.845 144.335 ;
        RECT 92.175 142.555 93.845 143.645 ;
        RECT 95.610 142.990 95.960 144.240 ;
        RECT 97.440 143.730 97.780 144.560 ;
        RECT 101.130 142.990 101.480 144.240 ;
        RECT 102.960 143.730 103.300 144.560 ;
        RECT 105.595 144.535 105.765 144.885 ;
        RECT 105.965 144.705 106.295 145.105 ;
        RECT 106.465 144.535 106.635 144.885 ;
        RECT 106.805 144.705 107.185 145.105 ;
        RECT 105.060 143.865 105.410 144.435 ;
        RECT 105.595 144.365 107.205 144.535 ;
        RECT 107.375 144.430 107.645 144.775 ;
        RECT 107.035 144.195 107.205 144.365 ;
        RECT 105.580 143.745 106.290 144.195 ;
        RECT 106.460 143.865 106.865 144.195 ;
        RECT 107.035 143.865 107.305 144.195 ;
        RECT 105.060 143.405 105.380 143.695 ;
        RECT 105.575 143.575 106.290 143.745 ;
        RECT 107.035 143.695 107.205 143.865 ;
        RECT 107.475 143.695 107.645 144.430 ;
        RECT 107.815 144.355 109.025 145.105 ;
        RECT 106.480 143.525 107.205 143.695 ;
        RECT 106.480 143.405 106.650 143.525 ;
        RECT 105.060 143.235 106.650 143.405 ;
        RECT 94.020 142.555 99.365 142.990 ;
        RECT 99.540 142.555 104.885 142.990 ;
        RECT 105.060 142.775 106.715 143.065 ;
        RECT 106.885 142.555 107.165 143.355 ;
        RECT 107.375 142.725 107.645 143.695 ;
        RECT 107.815 143.645 108.335 144.185 ;
        RECT 108.505 143.815 109.025 144.355 ;
        RECT 109.400 144.325 109.900 144.935 ;
        RECT 109.195 143.865 109.545 144.115 ;
        RECT 109.730 143.695 109.900 144.325 ;
        RECT 110.530 144.455 110.860 144.935 ;
        RECT 111.030 144.645 111.255 145.105 ;
        RECT 111.425 144.455 111.755 144.935 ;
        RECT 110.530 144.285 111.755 144.455 ;
        RECT 111.945 144.305 112.195 145.105 ;
        RECT 112.365 144.305 112.705 144.935 ;
        RECT 112.885 144.605 113.215 145.105 ;
        RECT 113.415 144.535 113.585 144.885 ;
        RECT 113.785 144.705 114.115 145.105 ;
        RECT 114.285 144.535 114.455 144.885 ;
        RECT 114.625 144.705 115.005 145.105 ;
        RECT 112.475 144.255 112.705 144.305 ;
        RECT 110.070 143.915 110.400 144.115 ;
        RECT 110.570 143.915 110.900 144.115 ;
        RECT 111.070 143.915 111.490 144.115 ;
        RECT 111.665 143.945 112.360 144.115 ;
        RECT 111.665 143.695 111.835 143.945 ;
        RECT 112.530 143.695 112.705 144.255 ;
        RECT 112.880 143.865 113.230 144.435 ;
        RECT 113.415 144.365 115.025 144.535 ;
        RECT 115.195 144.430 115.465 144.775 ;
        RECT 114.855 144.195 115.025 144.365 ;
        RECT 113.400 143.745 114.110 144.195 ;
        RECT 114.280 143.865 114.685 144.195 ;
        RECT 114.855 143.865 115.125 144.195 ;
        RECT 107.815 142.555 109.025 143.645 ;
        RECT 109.400 143.525 111.835 143.695 ;
        RECT 109.400 142.725 109.730 143.525 ;
        RECT 109.900 142.555 110.230 143.355 ;
        RECT 110.530 142.725 110.860 143.525 ;
        RECT 111.505 142.555 111.755 143.355 ;
        RECT 112.025 142.555 112.195 143.695 ;
        RECT 112.365 142.725 112.705 143.695 ;
        RECT 112.880 143.405 113.200 143.695 ;
        RECT 113.395 143.575 114.110 143.745 ;
        RECT 114.855 143.695 115.025 143.865 ;
        RECT 115.295 143.695 115.465 144.430 ;
        RECT 116.095 144.380 116.385 145.105 ;
        RECT 117.020 144.560 122.365 145.105 ;
        RECT 122.540 144.560 127.885 145.105 ;
        RECT 114.300 143.525 115.025 143.695 ;
        RECT 114.300 143.405 114.470 143.525 ;
        RECT 112.880 143.235 114.470 143.405 ;
        RECT 112.880 142.775 114.535 143.065 ;
        RECT 114.705 142.555 114.985 143.355 ;
        RECT 115.195 142.725 115.465 143.695 ;
        RECT 116.095 142.555 116.385 143.720 ;
        RECT 118.610 142.990 118.960 144.240 ;
        RECT 120.440 143.730 120.780 144.560 ;
        RECT 124.130 142.990 124.480 144.240 ;
        RECT 125.960 143.730 126.300 144.560 ;
        RECT 128.055 144.355 129.265 145.105 ;
        RECT 128.055 143.645 128.575 144.185 ;
        RECT 128.745 143.815 129.265 144.355 ;
        RECT 117.020 142.555 122.365 142.990 ;
        RECT 122.540 142.555 127.885 142.990 ;
        RECT 128.055 142.555 129.265 143.645 ;
        RECT 9.290 142.385 129.350 142.555 ;
        RECT 9.375 141.295 10.585 142.385 ;
        RECT 9.375 140.585 9.895 141.125 ;
        RECT 10.065 140.755 10.585 141.295 ;
        RECT 10.755 141.295 14.265 142.385 ;
        RECT 14.525 141.715 14.695 142.215 ;
        RECT 14.865 141.885 15.195 142.385 ;
        RECT 14.525 141.545 15.190 141.715 ;
        RECT 10.755 140.775 12.445 141.295 ;
        RECT 12.615 140.605 14.265 141.125 ;
        RECT 14.440 140.725 14.790 141.375 ;
        RECT 9.375 139.835 10.585 140.585 ;
        RECT 10.755 139.835 14.265 140.605 ;
        RECT 14.960 140.555 15.190 141.545 ;
        RECT 14.525 140.385 15.190 140.555 ;
        RECT 14.525 140.095 14.695 140.385 ;
        RECT 14.865 139.835 15.195 140.215 ;
        RECT 15.365 140.095 15.590 142.215 ;
        RECT 15.805 141.885 16.135 142.385 ;
        RECT 16.305 141.715 16.475 142.215 ;
        RECT 16.710 142.000 17.540 142.170 ;
        RECT 17.780 142.005 18.160 142.385 ;
        RECT 15.780 141.545 16.475 141.715 ;
        RECT 15.780 140.575 15.950 141.545 ;
        RECT 16.120 140.755 16.530 141.375 ;
        RECT 16.700 141.325 17.200 141.705 ;
        RECT 15.780 140.385 16.475 140.575 ;
        RECT 16.700 140.455 16.920 141.325 ;
        RECT 17.370 141.155 17.540 142.000 ;
        RECT 18.340 141.835 18.510 142.125 ;
        RECT 18.680 142.005 19.010 142.385 ;
        RECT 19.480 141.915 20.110 142.165 ;
        RECT 20.290 142.005 20.710 142.385 ;
        RECT 19.940 141.835 20.110 141.915 ;
        RECT 20.910 141.835 21.150 142.125 ;
        RECT 17.710 141.585 19.080 141.835 ;
        RECT 17.710 141.325 17.960 141.585 ;
        RECT 18.470 141.155 18.720 141.315 ;
        RECT 17.370 140.985 18.720 141.155 ;
        RECT 17.370 140.945 17.790 140.985 ;
        RECT 17.100 140.395 17.450 140.765 ;
        RECT 15.805 139.835 16.135 140.215 ;
        RECT 16.305 140.055 16.475 140.385 ;
        RECT 17.620 140.215 17.790 140.945 ;
        RECT 18.890 140.815 19.080 141.585 ;
        RECT 17.960 140.485 18.370 140.815 ;
        RECT 18.660 140.475 19.080 140.815 ;
        RECT 19.250 141.405 19.770 141.715 ;
        RECT 19.940 141.665 21.150 141.835 ;
        RECT 21.380 141.695 21.710 142.385 ;
        RECT 19.250 140.645 19.420 141.405 ;
        RECT 19.590 140.815 19.770 141.225 ;
        RECT 19.940 141.155 20.110 141.665 ;
        RECT 21.880 141.515 22.050 142.125 ;
        RECT 22.320 141.665 22.650 142.175 ;
        RECT 21.880 141.495 22.200 141.515 ;
        RECT 20.280 141.325 22.200 141.495 ;
        RECT 19.940 140.985 21.840 141.155 ;
        RECT 20.170 140.645 20.500 140.765 ;
        RECT 19.250 140.475 20.500 140.645 ;
        RECT 16.775 140.015 17.790 140.215 ;
        RECT 17.960 139.835 18.370 140.275 ;
        RECT 18.660 140.045 18.910 140.475 ;
        RECT 19.110 139.835 19.430 140.295 ;
        RECT 20.670 140.225 20.840 140.985 ;
        RECT 21.510 140.925 21.840 140.985 ;
        RECT 21.030 140.755 21.360 140.815 ;
        RECT 21.030 140.485 21.690 140.755 ;
        RECT 22.010 140.430 22.200 141.325 ;
        RECT 19.990 140.055 20.840 140.225 ;
        RECT 21.040 139.835 21.700 140.315 ;
        RECT 21.880 140.100 22.200 140.430 ;
        RECT 22.400 141.075 22.650 141.665 ;
        RECT 22.830 141.585 23.115 142.385 ;
        RECT 23.295 142.045 23.550 142.075 ;
        RECT 23.295 141.875 23.635 142.045 ;
        RECT 23.295 141.405 23.550 141.875 ;
        RECT 22.400 140.745 23.200 141.075 ;
        RECT 22.400 140.095 22.650 140.745 ;
        RECT 23.370 140.545 23.550 141.405 ;
        RECT 24.095 141.295 25.765 142.385 ;
        RECT 24.095 140.775 24.845 141.295 ;
        RECT 25.935 141.220 26.225 142.385 ;
        RECT 26.860 141.950 32.205 142.385 ;
        RECT 25.015 140.605 25.765 141.125 ;
        RECT 28.450 140.700 28.800 141.950 ;
        RECT 32.375 141.245 32.715 142.215 ;
        RECT 32.885 141.245 33.055 142.385 ;
        RECT 33.325 141.585 33.575 142.385 ;
        RECT 34.220 141.415 34.550 142.215 ;
        RECT 34.850 141.585 35.180 142.385 ;
        RECT 35.350 141.415 35.680 142.215 ;
        RECT 33.245 141.245 35.680 141.415 ;
        RECT 36.055 141.295 37.265 142.385 ;
        RECT 37.435 141.295 40.945 142.385 ;
        RECT 41.120 141.950 46.465 142.385 ;
        RECT 22.830 139.835 23.115 140.295 ;
        RECT 23.295 140.015 23.550 140.545 ;
        RECT 24.095 139.835 25.765 140.605 ;
        RECT 25.935 139.835 26.225 140.560 ;
        RECT 30.280 140.380 30.620 141.210 ;
        RECT 32.375 140.635 32.550 141.245 ;
        RECT 33.245 140.995 33.415 141.245 ;
        RECT 32.720 140.825 33.415 140.995 ;
        RECT 33.590 140.825 34.010 141.025 ;
        RECT 34.180 140.825 34.510 141.025 ;
        RECT 34.680 140.825 35.010 141.025 ;
        RECT 26.860 139.835 32.205 140.380 ;
        RECT 32.375 140.005 32.715 140.635 ;
        RECT 32.885 139.835 33.135 140.635 ;
        RECT 33.325 140.485 34.550 140.655 ;
        RECT 33.325 140.005 33.655 140.485 ;
        RECT 33.825 139.835 34.050 140.295 ;
        RECT 34.220 140.005 34.550 140.485 ;
        RECT 35.180 140.615 35.350 141.245 ;
        RECT 35.535 140.825 35.885 141.075 ;
        RECT 36.055 140.755 36.575 141.295 ;
        RECT 35.180 140.005 35.680 140.615 ;
        RECT 36.745 140.585 37.265 141.125 ;
        RECT 37.435 140.775 39.125 141.295 ;
        RECT 39.295 140.605 40.945 141.125 ;
        RECT 42.710 140.700 43.060 141.950 ;
        RECT 46.635 141.245 46.975 142.215 ;
        RECT 47.145 141.245 47.315 142.385 ;
        RECT 47.585 141.585 47.835 142.385 ;
        RECT 48.480 141.415 48.810 142.215 ;
        RECT 49.110 141.585 49.440 142.385 ;
        RECT 49.610 141.415 49.940 142.215 ;
        RECT 47.505 141.245 49.940 141.415 ;
        RECT 50.315 141.295 51.525 142.385 ;
        RECT 36.055 139.835 37.265 140.585 ;
        RECT 37.435 139.835 40.945 140.605 ;
        RECT 44.540 140.380 44.880 141.210 ;
        RECT 46.635 140.635 46.810 141.245 ;
        RECT 47.505 140.995 47.675 141.245 ;
        RECT 46.980 140.825 47.675 140.995 ;
        RECT 47.850 140.825 48.270 141.025 ;
        RECT 48.440 140.825 48.770 141.025 ;
        RECT 48.940 140.825 49.270 141.025 ;
        RECT 41.120 139.835 46.465 140.380 ;
        RECT 46.635 140.005 46.975 140.635 ;
        RECT 47.145 139.835 47.395 140.635 ;
        RECT 47.585 140.485 48.810 140.655 ;
        RECT 47.585 140.005 47.915 140.485 ;
        RECT 48.085 139.835 48.310 140.295 ;
        RECT 48.480 140.005 48.810 140.485 ;
        RECT 49.440 140.615 49.610 141.245 ;
        RECT 49.795 140.825 50.145 141.075 ;
        RECT 50.315 140.755 50.835 141.295 ;
        RECT 51.695 141.220 51.985 142.385 ;
        RECT 52.705 141.455 52.875 142.215 ;
        RECT 53.055 141.625 53.385 142.385 ;
        RECT 52.705 141.285 53.370 141.455 ;
        RECT 53.555 141.310 53.825 142.215 ;
        RECT 53.200 141.140 53.370 141.285 ;
        RECT 49.440 140.005 49.940 140.615 ;
        RECT 51.005 140.585 51.525 141.125 ;
        RECT 52.635 140.735 52.965 141.105 ;
        RECT 53.200 140.810 53.485 141.140 ;
        RECT 50.315 139.835 51.525 140.585 ;
        RECT 51.695 139.835 51.985 140.560 ;
        RECT 53.200 140.555 53.370 140.810 ;
        RECT 52.705 140.385 53.370 140.555 ;
        RECT 53.655 140.510 53.825 141.310 ;
        RECT 53.995 141.295 55.665 142.385 ;
        RECT 55.840 141.995 56.175 142.215 ;
        RECT 57.180 142.005 57.535 142.385 ;
        RECT 55.840 141.375 56.095 141.995 ;
        RECT 56.345 141.835 56.575 141.875 ;
        RECT 57.705 141.835 57.955 142.215 ;
        RECT 56.345 141.635 57.955 141.835 ;
        RECT 56.345 141.545 56.530 141.635 ;
        RECT 57.120 141.625 57.955 141.635 ;
        RECT 58.205 141.605 58.455 142.385 ;
        RECT 58.625 141.535 58.885 142.215 ;
        RECT 59.145 141.715 59.315 142.215 ;
        RECT 59.485 141.885 59.815 142.385 ;
        RECT 59.145 141.545 59.810 141.715 ;
        RECT 56.685 141.435 57.015 141.465 ;
        RECT 56.685 141.375 58.485 141.435 ;
        RECT 53.995 140.775 54.745 141.295 ;
        RECT 55.840 141.265 58.545 141.375 ;
        RECT 55.840 141.205 57.015 141.265 ;
        RECT 58.345 141.230 58.545 141.265 ;
        RECT 54.915 140.605 55.665 141.125 ;
        RECT 55.835 140.825 56.325 141.025 ;
        RECT 56.515 140.825 56.990 141.035 ;
        RECT 52.705 140.005 52.875 140.385 ;
        RECT 53.055 139.835 53.385 140.215 ;
        RECT 53.565 140.005 53.825 140.510 ;
        RECT 53.995 139.835 55.665 140.605 ;
        RECT 55.840 139.835 56.295 140.600 ;
        RECT 56.770 140.425 56.990 140.825 ;
        RECT 57.235 140.825 57.565 141.035 ;
        RECT 57.235 140.425 57.445 140.825 ;
        RECT 57.735 140.790 58.145 141.095 ;
        RECT 58.375 140.655 58.545 141.230 ;
        RECT 58.275 140.535 58.545 140.655 ;
        RECT 57.700 140.490 58.545 140.535 ;
        RECT 57.700 140.365 58.455 140.490 ;
        RECT 57.700 140.215 57.870 140.365 ;
        RECT 58.715 140.335 58.885 141.535 ;
        RECT 59.060 140.725 59.410 141.375 ;
        RECT 59.580 140.555 59.810 141.545 ;
        RECT 56.570 140.005 57.870 140.215 ;
        RECT 58.125 139.835 58.455 140.195 ;
        RECT 58.625 140.005 58.885 140.335 ;
        RECT 59.145 140.385 59.810 140.555 ;
        RECT 59.145 140.095 59.315 140.385 ;
        RECT 59.485 139.835 59.815 140.215 ;
        RECT 59.985 140.095 60.210 142.215 ;
        RECT 60.425 141.885 60.755 142.385 ;
        RECT 60.925 141.715 61.095 142.215 ;
        RECT 61.330 142.000 62.160 142.170 ;
        RECT 62.400 142.005 62.780 142.385 ;
        RECT 60.400 141.545 61.095 141.715 ;
        RECT 60.400 140.575 60.570 141.545 ;
        RECT 60.740 140.755 61.150 141.375 ;
        RECT 61.320 141.325 61.820 141.705 ;
        RECT 60.400 140.385 61.095 140.575 ;
        RECT 61.320 140.455 61.540 141.325 ;
        RECT 61.990 141.155 62.160 142.000 ;
        RECT 62.960 141.835 63.130 142.125 ;
        RECT 63.300 142.005 63.630 142.385 ;
        RECT 64.100 141.915 64.730 142.165 ;
        RECT 64.910 142.005 65.330 142.385 ;
        RECT 64.560 141.835 64.730 141.915 ;
        RECT 65.530 141.835 65.770 142.125 ;
        RECT 62.330 141.585 63.700 141.835 ;
        RECT 62.330 141.325 62.580 141.585 ;
        RECT 63.090 141.155 63.340 141.315 ;
        RECT 61.990 140.985 63.340 141.155 ;
        RECT 61.990 140.945 62.410 140.985 ;
        RECT 61.720 140.395 62.070 140.765 ;
        RECT 60.425 139.835 60.755 140.215 ;
        RECT 60.925 140.055 61.095 140.385 ;
        RECT 62.240 140.215 62.410 140.945 ;
        RECT 63.510 140.815 63.700 141.585 ;
        RECT 62.580 140.485 62.990 140.815 ;
        RECT 63.280 140.475 63.700 140.815 ;
        RECT 63.870 141.405 64.390 141.715 ;
        RECT 64.560 141.665 65.770 141.835 ;
        RECT 66.000 141.695 66.330 142.385 ;
        RECT 63.870 140.645 64.040 141.405 ;
        RECT 64.210 140.815 64.390 141.225 ;
        RECT 64.560 141.155 64.730 141.665 ;
        RECT 66.500 141.515 66.670 142.125 ;
        RECT 66.940 141.665 67.270 142.175 ;
        RECT 66.500 141.495 66.820 141.515 ;
        RECT 64.900 141.325 66.820 141.495 ;
        RECT 64.560 140.985 66.460 141.155 ;
        RECT 64.790 140.645 65.120 140.765 ;
        RECT 63.870 140.475 65.120 140.645 ;
        RECT 61.395 140.015 62.410 140.215 ;
        RECT 62.580 139.835 62.990 140.275 ;
        RECT 63.280 140.045 63.530 140.475 ;
        RECT 63.730 139.835 64.050 140.295 ;
        RECT 65.290 140.225 65.460 140.985 ;
        RECT 66.130 140.925 66.460 140.985 ;
        RECT 65.650 140.755 65.980 140.815 ;
        RECT 65.650 140.485 66.310 140.755 ;
        RECT 66.630 140.430 66.820 141.325 ;
        RECT 64.610 140.055 65.460 140.225 ;
        RECT 65.660 139.835 66.320 140.315 ;
        RECT 66.500 140.100 66.820 140.430 ;
        RECT 67.020 141.075 67.270 141.665 ;
        RECT 67.450 141.585 67.735 142.385 ;
        RECT 67.915 142.045 68.170 142.075 ;
        RECT 67.915 141.875 68.255 142.045 ;
        RECT 67.915 141.405 68.170 141.875 ;
        RECT 67.020 140.745 67.820 141.075 ;
        RECT 67.020 140.095 67.270 140.745 ;
        RECT 67.990 140.545 68.170 141.405 ;
        RECT 67.450 139.835 67.735 140.295 ;
        RECT 67.915 140.015 68.170 140.545 ;
        RECT 68.715 141.245 69.055 142.215 ;
        RECT 69.225 141.245 69.395 142.385 ;
        RECT 69.665 141.585 69.915 142.385 ;
        RECT 70.560 141.415 70.890 142.215 ;
        RECT 71.190 141.585 71.520 142.385 ;
        RECT 71.690 141.415 72.020 142.215 ;
        RECT 69.585 141.245 72.020 141.415 ;
        RECT 72.455 141.245 72.665 142.385 ;
        RECT 68.715 140.635 68.890 141.245 ;
        RECT 69.585 140.995 69.755 141.245 ;
        RECT 69.060 140.825 69.755 140.995 ;
        RECT 69.930 140.825 70.350 141.025 ;
        RECT 70.520 140.825 70.850 141.025 ;
        RECT 71.020 140.825 71.350 141.025 ;
        RECT 68.715 140.005 69.055 140.635 ;
        RECT 69.225 139.835 69.475 140.635 ;
        RECT 69.665 140.485 70.890 140.655 ;
        RECT 69.665 140.005 69.995 140.485 ;
        RECT 70.165 139.835 70.390 140.295 ;
        RECT 70.560 140.005 70.890 140.485 ;
        RECT 71.520 140.615 71.690 141.245 ;
        RECT 72.835 141.235 73.165 142.215 ;
        RECT 73.335 141.245 73.565 142.385 ;
        RECT 73.775 141.295 77.285 142.385 ;
        RECT 71.875 140.825 72.225 141.075 ;
        RECT 71.520 140.005 72.020 140.615 ;
        RECT 72.455 139.835 72.665 140.655 ;
        RECT 72.835 140.635 73.085 141.235 ;
        RECT 73.255 140.825 73.585 141.075 ;
        RECT 73.775 140.775 75.465 141.295 ;
        RECT 77.455 141.220 77.745 142.385 ;
        RECT 77.915 141.245 78.185 142.215 ;
        RECT 78.395 141.585 78.675 142.385 ;
        RECT 78.845 141.875 80.500 142.165 ;
        RECT 81.140 141.950 86.485 142.385 ;
        RECT 86.660 141.950 92.005 142.385 ;
        RECT 92.180 141.950 97.525 142.385 ;
        RECT 97.700 141.950 103.045 142.385 ;
        RECT 78.910 141.535 80.500 141.705 ;
        RECT 78.910 141.415 79.080 141.535 ;
        RECT 78.355 141.245 79.080 141.415 ;
        RECT 72.835 140.005 73.165 140.635 ;
        RECT 73.335 139.835 73.565 140.655 ;
        RECT 75.635 140.605 77.285 141.125 ;
        RECT 73.775 139.835 77.285 140.605 ;
        RECT 77.455 139.835 77.745 140.560 ;
        RECT 77.915 140.510 78.085 141.245 ;
        RECT 78.355 141.075 78.525 141.245 ;
        RECT 78.255 140.745 78.525 141.075 ;
        RECT 78.695 140.745 79.100 141.075 ;
        RECT 79.270 140.745 79.980 141.365 ;
        RECT 80.180 141.245 80.500 141.535 ;
        RECT 78.355 140.575 78.525 140.745 ;
        RECT 77.915 140.165 78.185 140.510 ;
        RECT 78.355 140.405 79.965 140.575 ;
        RECT 80.150 140.505 80.500 141.075 ;
        RECT 82.730 140.700 83.080 141.950 ;
        RECT 78.375 139.835 78.755 140.235 ;
        RECT 78.925 140.055 79.095 140.405 ;
        RECT 79.265 139.835 79.595 140.235 ;
        RECT 79.795 140.055 79.965 140.405 ;
        RECT 84.560 140.380 84.900 141.210 ;
        RECT 88.250 140.700 88.600 141.950 ;
        RECT 90.080 140.380 90.420 141.210 ;
        RECT 93.770 140.700 94.120 141.950 ;
        RECT 95.600 140.380 95.940 141.210 ;
        RECT 99.290 140.700 99.640 141.950 ;
        RECT 103.215 141.220 103.505 142.385 ;
        RECT 103.675 141.295 104.885 142.385 ;
        RECT 105.055 141.295 108.565 142.385 ;
        RECT 101.120 140.380 101.460 141.210 ;
        RECT 103.675 140.755 104.195 141.295 ;
        RECT 104.365 140.585 104.885 141.125 ;
        RECT 105.055 140.775 106.745 141.295 ;
        RECT 108.735 141.245 109.075 142.215 ;
        RECT 109.245 141.245 109.415 142.385 ;
        RECT 109.685 141.585 109.935 142.385 ;
        RECT 110.580 141.415 110.910 142.215 ;
        RECT 111.210 141.585 111.540 142.385 ;
        RECT 111.710 141.415 112.040 142.215 ;
        RECT 109.605 141.245 112.040 141.415 ;
        RECT 112.875 141.295 116.385 142.385 ;
        RECT 106.915 140.605 108.565 141.125 ;
        RECT 80.165 139.835 80.495 140.335 ;
        RECT 81.140 139.835 86.485 140.380 ;
        RECT 86.660 139.835 92.005 140.380 ;
        RECT 92.180 139.835 97.525 140.380 ;
        RECT 97.700 139.835 103.045 140.380 ;
        RECT 103.215 139.835 103.505 140.560 ;
        RECT 103.675 139.835 104.885 140.585 ;
        RECT 105.055 139.835 108.565 140.605 ;
        RECT 108.735 140.635 108.910 141.245 ;
        RECT 109.605 140.995 109.775 141.245 ;
        RECT 109.080 140.825 109.775 140.995 ;
        RECT 109.950 140.825 110.370 141.025 ;
        RECT 110.540 140.825 110.870 141.025 ;
        RECT 111.040 140.825 111.370 141.025 ;
        RECT 108.735 140.005 109.075 140.635 ;
        RECT 109.245 139.835 109.495 140.635 ;
        RECT 109.685 140.485 110.910 140.655 ;
        RECT 109.685 140.005 110.015 140.485 ;
        RECT 110.185 139.835 110.410 140.295 ;
        RECT 110.580 140.005 110.910 140.485 ;
        RECT 111.540 140.615 111.710 141.245 ;
        RECT 111.895 140.825 112.245 141.075 ;
        RECT 112.875 140.775 114.565 141.295 ;
        RECT 116.595 141.245 116.825 142.385 ;
        RECT 116.995 141.235 117.325 142.215 ;
        RECT 117.495 141.245 117.705 142.385 ;
        RECT 117.935 141.625 118.450 142.035 ;
        RECT 118.685 141.625 118.855 142.385 ;
        RECT 119.025 142.045 121.055 142.215 ;
        RECT 111.540 140.005 112.040 140.615 ;
        RECT 114.735 140.605 116.385 141.125 ;
        RECT 116.575 140.825 116.905 141.075 ;
        RECT 112.875 139.835 116.385 140.605 ;
        RECT 116.595 139.835 116.825 140.655 ;
        RECT 117.075 140.635 117.325 141.235 ;
        RECT 117.935 140.815 118.275 141.625 ;
        RECT 119.025 141.380 119.195 142.045 ;
        RECT 119.590 141.705 120.715 141.875 ;
        RECT 118.445 141.190 119.195 141.380 ;
        RECT 119.365 141.365 120.375 141.535 ;
        RECT 116.995 140.005 117.325 140.635 ;
        RECT 117.495 139.835 117.705 140.655 ;
        RECT 117.935 140.645 119.165 140.815 ;
        RECT 118.210 140.040 118.455 140.645 ;
        RECT 118.675 139.835 119.185 140.370 ;
        RECT 119.365 140.005 119.555 141.365 ;
        RECT 119.725 141.025 120.000 141.165 ;
        RECT 119.725 140.855 120.005 141.025 ;
        RECT 119.725 140.005 120.000 140.855 ;
        RECT 120.205 140.565 120.375 141.365 ;
        RECT 120.545 140.575 120.715 141.705 ;
        RECT 120.885 141.075 121.055 142.045 ;
        RECT 121.225 141.245 121.395 142.385 ;
        RECT 121.565 141.245 121.900 142.215 ;
        RECT 123.085 141.455 123.255 142.215 ;
        RECT 123.435 141.625 123.765 142.385 ;
        RECT 123.085 141.285 123.750 141.455 ;
        RECT 123.935 141.310 124.205 142.215 ;
        RECT 120.885 140.745 121.080 141.075 ;
        RECT 121.305 140.745 121.560 141.075 ;
        RECT 121.305 140.575 121.475 140.745 ;
        RECT 121.730 140.575 121.900 141.245 ;
        RECT 123.580 141.140 123.750 141.285 ;
        RECT 123.015 140.735 123.345 141.105 ;
        RECT 123.580 140.810 123.865 141.140 ;
        RECT 120.545 140.405 121.475 140.575 ;
        RECT 120.545 140.370 120.720 140.405 ;
        RECT 120.190 140.005 120.720 140.370 ;
        RECT 121.145 139.835 121.475 140.235 ;
        RECT 121.645 140.005 121.900 140.575 ;
        RECT 123.580 140.555 123.750 140.810 ;
        RECT 123.085 140.385 123.750 140.555 ;
        RECT 124.035 140.510 124.205 141.310 ;
        RECT 124.375 141.295 127.885 142.385 ;
        RECT 128.055 141.295 129.265 142.385 ;
        RECT 124.375 140.775 126.065 141.295 ;
        RECT 126.235 140.605 127.885 141.125 ;
        RECT 128.055 140.755 128.575 141.295 ;
        RECT 123.085 140.005 123.255 140.385 ;
        RECT 123.435 139.835 123.765 140.215 ;
        RECT 123.945 140.005 124.205 140.510 ;
        RECT 124.375 139.835 127.885 140.605 ;
        RECT 128.745 140.585 129.265 141.125 ;
        RECT 128.055 139.835 129.265 140.585 ;
        RECT 9.290 139.665 129.350 139.835 ;
        RECT 9.375 138.915 10.585 139.665 ;
        RECT 9.375 138.375 9.895 138.915 ;
        RECT 11.215 138.895 12.885 139.665 ;
        RECT 13.055 138.940 13.345 139.665 ;
        RECT 13.975 138.895 17.485 139.665 ;
        RECT 10.065 138.205 10.585 138.745 ;
        RECT 9.375 137.115 10.585 138.205 ;
        RECT 11.215 138.205 11.965 138.725 ;
        RECT 12.135 138.375 12.885 138.895 ;
        RECT 11.215 137.115 12.885 138.205 ;
        RECT 13.055 137.115 13.345 138.280 ;
        RECT 13.975 138.205 15.665 138.725 ;
        RECT 15.835 138.375 17.485 138.895 ;
        RECT 17.695 138.845 17.925 139.665 ;
        RECT 18.095 138.865 18.425 139.495 ;
        RECT 17.675 138.425 18.005 138.675 ;
        RECT 18.175 138.265 18.425 138.865 ;
        RECT 18.595 138.845 18.805 139.665 ;
        RECT 19.035 138.895 21.625 139.665 ;
        RECT 21.800 139.120 27.145 139.665 ;
        RECT 13.975 137.115 17.485 138.205 ;
        RECT 17.695 137.115 17.925 138.255 ;
        RECT 18.095 137.285 18.425 138.265 ;
        RECT 18.595 137.115 18.805 138.255 ;
        RECT 19.035 138.205 20.245 138.725 ;
        RECT 20.415 138.375 21.625 138.895 ;
        RECT 19.035 137.115 21.625 138.205 ;
        RECT 23.390 137.550 23.740 138.800 ;
        RECT 25.220 138.290 25.560 139.120 ;
        RECT 27.315 138.990 27.585 139.335 ;
        RECT 27.775 139.265 28.155 139.665 ;
        RECT 28.325 139.095 28.495 139.445 ;
        RECT 28.665 139.265 28.995 139.665 ;
        RECT 29.195 139.095 29.365 139.445 ;
        RECT 29.565 139.165 29.895 139.665 ;
        RECT 27.315 138.255 27.485 138.990 ;
        RECT 27.755 138.925 29.365 139.095 ;
        RECT 27.755 138.755 27.925 138.925 ;
        RECT 27.655 138.425 27.925 138.755 ;
        RECT 28.095 138.425 28.500 138.755 ;
        RECT 27.755 138.255 27.925 138.425 ;
        RECT 28.670 138.305 29.380 138.755 ;
        RECT 29.550 138.425 29.900 138.995 ;
        RECT 30.075 138.990 30.345 139.335 ;
        RECT 30.535 139.265 30.915 139.665 ;
        RECT 31.085 139.095 31.255 139.445 ;
        RECT 31.425 139.265 31.755 139.665 ;
        RECT 31.955 139.095 32.125 139.445 ;
        RECT 32.325 139.165 32.655 139.665 ;
        RECT 21.800 137.115 27.145 137.550 ;
        RECT 27.315 137.285 27.585 138.255 ;
        RECT 27.755 138.085 28.480 138.255 ;
        RECT 28.670 138.135 29.385 138.305 ;
        RECT 30.075 138.255 30.245 138.990 ;
        RECT 30.515 138.925 32.125 139.095 ;
        RECT 30.515 138.755 30.685 138.925 ;
        RECT 30.415 138.425 30.685 138.755 ;
        RECT 30.855 138.425 31.260 138.755 ;
        RECT 30.515 138.255 30.685 138.425 ;
        RECT 31.430 138.305 32.140 138.755 ;
        RECT 32.310 138.425 32.660 138.995 ;
        RECT 32.835 138.990 33.105 139.335 ;
        RECT 33.295 139.265 33.675 139.665 ;
        RECT 33.845 139.095 34.015 139.445 ;
        RECT 34.185 139.265 34.515 139.665 ;
        RECT 34.715 139.095 34.885 139.445 ;
        RECT 35.085 139.165 35.415 139.665 ;
        RECT 28.310 137.965 28.480 138.085 ;
        RECT 29.580 137.965 29.900 138.255 ;
        RECT 27.795 137.115 28.075 137.915 ;
        RECT 28.310 137.795 29.900 137.965 ;
        RECT 28.245 137.335 29.900 137.625 ;
        RECT 30.075 137.285 30.345 138.255 ;
        RECT 30.515 138.085 31.240 138.255 ;
        RECT 31.430 138.135 32.145 138.305 ;
        RECT 32.835 138.255 33.005 138.990 ;
        RECT 33.275 138.925 34.885 139.095 ;
        RECT 33.275 138.755 33.445 138.925 ;
        RECT 33.175 138.425 33.445 138.755 ;
        RECT 33.615 138.425 34.020 138.755 ;
        RECT 33.275 138.255 33.445 138.425 ;
        RECT 34.190 138.305 34.900 138.755 ;
        RECT 35.070 138.425 35.420 138.995 ;
        RECT 36.055 138.895 38.645 139.665 ;
        RECT 38.815 138.940 39.105 139.665 ;
        RECT 39.735 138.895 42.325 139.665 ;
        RECT 42.500 139.120 47.845 139.665 ;
        RECT 31.070 137.965 31.240 138.085 ;
        RECT 32.340 137.965 32.660 138.255 ;
        RECT 30.555 137.115 30.835 137.915 ;
        RECT 31.070 137.795 32.660 137.965 ;
        RECT 31.005 137.335 32.660 137.625 ;
        RECT 32.835 137.285 33.105 138.255 ;
        RECT 33.275 138.085 34.000 138.255 ;
        RECT 34.190 138.135 34.905 138.305 ;
        RECT 33.830 137.965 34.000 138.085 ;
        RECT 35.100 137.965 35.420 138.255 ;
        RECT 33.315 137.115 33.595 137.915 ;
        RECT 33.830 137.795 35.420 137.965 ;
        RECT 36.055 138.205 37.265 138.725 ;
        RECT 37.435 138.375 38.645 138.895 ;
        RECT 33.765 137.335 35.420 137.625 ;
        RECT 36.055 137.115 38.645 138.205 ;
        RECT 38.815 137.115 39.105 138.280 ;
        RECT 39.735 138.205 40.945 138.725 ;
        RECT 41.115 138.375 42.325 138.895 ;
        RECT 39.735 137.115 42.325 138.205 ;
        RECT 44.090 137.550 44.440 138.800 ;
        RECT 45.920 138.290 46.260 139.120 ;
        RECT 48.020 138.925 48.275 139.495 ;
        RECT 48.445 139.265 48.775 139.665 ;
        RECT 49.200 139.130 49.730 139.495 ;
        RECT 49.920 139.325 50.195 139.495 ;
        RECT 49.915 139.155 50.195 139.325 ;
        RECT 49.200 139.095 49.375 139.130 ;
        RECT 48.445 138.925 49.375 139.095 ;
        RECT 48.020 138.255 48.190 138.925 ;
        RECT 48.445 138.755 48.615 138.925 ;
        RECT 48.360 138.425 48.615 138.755 ;
        RECT 48.840 138.425 49.035 138.755 ;
        RECT 42.500 137.115 47.845 137.550 ;
        RECT 48.020 137.285 48.355 138.255 ;
        RECT 48.525 137.115 48.695 138.255 ;
        RECT 48.865 137.455 49.035 138.425 ;
        RECT 49.205 137.795 49.375 138.925 ;
        RECT 49.545 138.135 49.715 138.935 ;
        RECT 49.920 138.335 50.195 139.155 ;
        RECT 50.365 138.135 50.555 139.495 ;
        RECT 50.735 139.130 51.245 139.665 ;
        RECT 51.465 138.855 51.710 139.460 ;
        RECT 52.615 138.895 55.205 139.665 ;
        RECT 55.380 139.120 60.725 139.665 ;
        RECT 50.755 138.685 51.985 138.855 ;
        RECT 49.545 137.965 50.555 138.135 ;
        RECT 50.725 138.120 51.475 138.310 ;
        RECT 49.205 137.625 50.330 137.795 ;
        RECT 50.725 137.455 50.895 138.120 ;
        RECT 51.645 137.875 51.985 138.685 ;
        RECT 48.865 137.285 50.895 137.455 ;
        RECT 51.065 137.115 51.235 137.875 ;
        RECT 51.470 137.465 51.985 137.875 ;
        RECT 52.615 138.205 53.825 138.725 ;
        RECT 53.995 138.375 55.205 138.895 ;
        RECT 52.615 137.115 55.205 138.205 ;
        RECT 56.970 137.550 57.320 138.800 ;
        RECT 58.800 138.290 59.140 139.120 ;
        RECT 60.895 138.865 61.235 139.495 ;
        RECT 61.405 138.865 61.655 139.665 ;
        RECT 61.845 139.015 62.175 139.495 ;
        RECT 62.345 139.205 62.570 139.665 ;
        RECT 62.740 139.015 63.070 139.495 ;
        RECT 60.895 138.255 61.070 138.865 ;
        RECT 61.845 138.845 63.070 139.015 ;
        RECT 63.700 138.885 64.200 139.495 ;
        RECT 64.575 138.940 64.865 139.665 ;
        RECT 65.495 138.895 68.085 139.665 ;
        RECT 61.240 138.505 61.935 138.675 ;
        RECT 61.765 138.255 61.935 138.505 ;
        RECT 62.110 138.475 62.530 138.675 ;
        RECT 62.700 138.475 63.030 138.675 ;
        RECT 63.200 138.475 63.530 138.675 ;
        RECT 63.700 138.255 63.870 138.885 ;
        RECT 64.055 138.425 64.405 138.675 ;
        RECT 55.380 137.115 60.725 137.550 ;
        RECT 60.895 137.285 61.235 138.255 ;
        RECT 61.405 137.115 61.575 138.255 ;
        RECT 61.765 138.085 64.200 138.255 ;
        RECT 61.845 137.115 62.095 137.915 ;
        RECT 62.740 137.285 63.070 138.085 ;
        RECT 63.370 137.115 63.700 137.915 ;
        RECT 63.870 137.285 64.200 138.085 ;
        RECT 64.575 137.115 64.865 138.280 ;
        RECT 65.495 138.205 66.705 138.725 ;
        RECT 66.875 138.375 68.085 138.895 ;
        RECT 68.630 138.955 68.885 139.485 ;
        RECT 69.065 139.205 69.350 139.665 ;
        RECT 65.495 137.115 68.085 138.205 ;
        RECT 68.630 138.095 68.810 138.955 ;
        RECT 69.530 138.755 69.780 139.405 ;
        RECT 68.980 138.425 69.780 138.755 ;
        RECT 68.630 137.625 68.885 138.095 ;
        RECT 68.545 137.455 68.885 137.625 ;
        RECT 68.630 137.425 68.885 137.455 ;
        RECT 69.065 137.115 69.350 137.915 ;
        RECT 69.530 137.835 69.780 138.425 ;
        RECT 69.980 139.070 70.300 139.400 ;
        RECT 70.480 139.185 71.140 139.665 ;
        RECT 71.340 139.275 72.190 139.445 ;
        RECT 69.980 138.175 70.170 139.070 ;
        RECT 70.490 138.745 71.150 139.015 ;
        RECT 70.820 138.685 71.150 138.745 ;
        RECT 70.340 138.515 70.670 138.575 ;
        RECT 71.340 138.515 71.510 139.275 ;
        RECT 72.750 139.205 73.070 139.665 ;
        RECT 73.270 139.025 73.520 139.455 ;
        RECT 73.810 139.225 74.220 139.665 ;
        RECT 74.390 139.285 75.405 139.485 ;
        RECT 71.680 138.855 72.930 139.025 ;
        RECT 71.680 138.735 72.010 138.855 ;
        RECT 70.340 138.345 72.240 138.515 ;
        RECT 69.980 138.005 71.900 138.175 ;
        RECT 69.980 137.985 70.300 138.005 ;
        RECT 69.530 137.325 69.860 137.835 ;
        RECT 70.130 137.375 70.300 137.985 ;
        RECT 72.070 137.835 72.240 138.345 ;
        RECT 72.410 138.275 72.590 138.685 ;
        RECT 72.760 138.095 72.930 138.855 ;
        RECT 70.470 137.115 70.800 137.805 ;
        RECT 71.030 137.665 72.240 137.835 ;
        RECT 72.410 137.785 72.930 138.095 ;
        RECT 73.100 138.685 73.520 139.025 ;
        RECT 73.810 138.685 74.220 139.015 ;
        RECT 73.100 137.915 73.290 138.685 ;
        RECT 74.390 138.555 74.560 139.285 ;
        RECT 75.705 139.115 75.875 139.445 ;
        RECT 76.045 139.285 76.375 139.665 ;
        RECT 74.730 138.735 75.080 139.105 ;
        RECT 74.390 138.515 74.810 138.555 ;
        RECT 73.460 138.345 74.810 138.515 ;
        RECT 73.460 138.185 73.710 138.345 ;
        RECT 74.220 137.915 74.470 138.175 ;
        RECT 73.100 137.665 74.470 137.915 ;
        RECT 71.030 137.375 71.270 137.665 ;
        RECT 72.070 137.585 72.240 137.665 ;
        RECT 71.470 137.115 71.890 137.495 ;
        RECT 72.070 137.335 72.700 137.585 ;
        RECT 73.170 137.115 73.500 137.495 ;
        RECT 73.670 137.375 73.840 137.665 ;
        RECT 74.640 137.500 74.810 138.345 ;
        RECT 75.260 138.175 75.480 139.045 ;
        RECT 75.705 138.925 76.400 139.115 ;
        RECT 74.980 137.795 75.480 138.175 ;
        RECT 75.650 138.125 76.060 138.745 ;
        RECT 76.230 137.955 76.400 138.925 ;
        RECT 75.705 137.785 76.400 137.955 ;
        RECT 74.020 137.115 74.400 137.495 ;
        RECT 74.640 137.330 75.470 137.500 ;
        RECT 75.705 137.285 75.875 137.785 ;
        RECT 76.045 137.115 76.375 137.615 ;
        RECT 76.590 137.285 76.815 139.405 ;
        RECT 76.985 139.285 77.315 139.665 ;
        RECT 77.485 139.115 77.655 139.405 ;
        RECT 76.990 138.945 77.655 139.115 ;
        RECT 76.990 137.955 77.220 138.945 ;
        RECT 77.915 138.915 79.125 139.665 ;
        RECT 77.390 138.125 77.740 138.775 ;
        RECT 77.915 138.205 78.435 138.745 ;
        RECT 78.605 138.375 79.125 138.915 ;
        RECT 79.295 138.865 79.635 139.495 ;
        RECT 79.805 138.865 80.055 139.665 ;
        RECT 80.245 139.015 80.575 139.495 ;
        RECT 80.745 139.205 80.970 139.665 ;
        RECT 81.140 139.015 81.470 139.495 ;
        RECT 79.295 138.255 79.470 138.865 ;
        RECT 80.245 138.845 81.470 139.015 ;
        RECT 82.100 138.885 82.600 139.495 ;
        RECT 83.440 139.120 88.785 139.665 ;
        RECT 79.640 138.505 80.335 138.675 ;
        RECT 80.165 138.255 80.335 138.505 ;
        RECT 80.510 138.475 80.930 138.675 ;
        RECT 81.100 138.475 81.430 138.675 ;
        RECT 81.600 138.475 81.930 138.675 ;
        RECT 82.100 138.255 82.270 138.885 ;
        RECT 82.455 138.425 82.805 138.675 ;
        RECT 76.990 137.785 77.655 137.955 ;
        RECT 76.985 137.115 77.315 137.615 ;
        RECT 77.485 137.285 77.655 137.785 ;
        RECT 77.915 137.115 79.125 138.205 ;
        RECT 79.295 137.285 79.635 138.255 ;
        RECT 79.805 137.115 79.975 138.255 ;
        RECT 80.165 138.085 82.600 138.255 ;
        RECT 80.245 137.115 80.495 137.915 ;
        RECT 81.140 137.285 81.470 138.085 ;
        RECT 81.770 137.115 82.100 137.915 ;
        RECT 82.270 137.285 82.600 138.085 ;
        RECT 85.030 137.550 85.380 138.800 ;
        RECT 86.860 138.290 87.200 139.120 ;
        RECT 89.015 138.845 89.225 139.665 ;
        RECT 89.395 138.865 89.725 139.495 ;
        RECT 89.395 138.265 89.645 138.865 ;
        RECT 89.895 138.845 90.125 139.665 ;
        RECT 90.335 138.940 90.625 139.665 ;
        RECT 91.260 139.120 96.605 139.665 ;
        RECT 89.815 138.425 90.145 138.675 ;
        RECT 83.440 137.115 88.785 137.550 ;
        RECT 89.015 137.115 89.225 138.255 ;
        RECT 89.395 137.285 89.725 138.265 ;
        RECT 89.895 137.115 90.125 138.255 ;
        RECT 90.335 137.115 90.625 138.280 ;
        RECT 92.850 137.550 93.200 138.800 ;
        RECT 94.680 138.290 95.020 139.120 ;
        RECT 96.775 138.990 97.045 139.335 ;
        RECT 97.235 139.265 97.615 139.665 ;
        RECT 97.785 139.095 97.955 139.445 ;
        RECT 98.125 139.265 98.455 139.665 ;
        RECT 98.655 139.095 98.825 139.445 ;
        RECT 99.025 139.165 99.355 139.665 ;
        RECT 96.775 138.255 96.945 138.990 ;
        RECT 97.215 138.925 98.825 139.095 ;
        RECT 97.215 138.755 97.385 138.925 ;
        RECT 97.115 138.425 97.385 138.755 ;
        RECT 97.555 138.425 97.960 138.755 ;
        RECT 97.215 138.255 97.385 138.425 ;
        RECT 98.130 138.305 98.840 138.755 ;
        RECT 99.010 138.425 99.360 138.995 ;
        RECT 99.535 138.865 99.875 139.495 ;
        RECT 100.045 138.865 100.295 139.665 ;
        RECT 100.485 139.015 100.815 139.495 ;
        RECT 100.985 139.205 101.210 139.665 ;
        RECT 101.380 139.015 101.710 139.495 ;
        RECT 99.535 138.815 99.765 138.865 ;
        RECT 100.485 138.845 101.710 139.015 ;
        RECT 102.340 138.885 102.840 139.495 ;
        RECT 103.675 138.990 103.945 139.335 ;
        RECT 104.135 139.265 104.515 139.665 ;
        RECT 104.685 139.095 104.855 139.445 ;
        RECT 105.025 139.265 105.355 139.665 ;
        RECT 105.555 139.095 105.725 139.445 ;
        RECT 105.925 139.165 106.255 139.665 ;
        RECT 91.260 137.115 96.605 137.550 ;
        RECT 96.775 137.285 97.045 138.255 ;
        RECT 97.215 138.085 97.940 138.255 ;
        RECT 98.130 138.135 98.845 138.305 ;
        RECT 99.535 138.255 99.710 138.815 ;
        RECT 99.880 138.505 100.575 138.675 ;
        RECT 100.405 138.255 100.575 138.505 ;
        RECT 100.750 138.475 101.170 138.675 ;
        RECT 101.340 138.475 101.670 138.675 ;
        RECT 101.840 138.475 102.170 138.675 ;
        RECT 102.340 138.255 102.510 138.885 ;
        RECT 102.695 138.425 103.045 138.675 ;
        RECT 103.675 138.255 103.845 138.990 ;
        RECT 104.115 138.925 105.725 139.095 ;
        RECT 104.115 138.755 104.285 138.925 ;
        RECT 104.015 138.425 104.285 138.755 ;
        RECT 104.455 138.425 104.860 138.755 ;
        RECT 104.115 138.255 104.285 138.425 ;
        RECT 97.770 137.965 97.940 138.085 ;
        RECT 99.040 137.965 99.360 138.255 ;
        RECT 97.255 137.115 97.535 137.915 ;
        RECT 97.770 137.795 99.360 137.965 ;
        RECT 97.705 137.335 99.360 137.625 ;
        RECT 99.535 137.285 99.875 138.255 ;
        RECT 100.045 137.115 100.215 138.255 ;
        RECT 100.405 138.085 102.840 138.255 ;
        RECT 100.485 137.115 100.735 137.915 ;
        RECT 101.380 137.285 101.710 138.085 ;
        RECT 102.010 137.115 102.340 137.915 ;
        RECT 102.510 137.285 102.840 138.085 ;
        RECT 103.675 137.285 103.945 138.255 ;
        RECT 104.115 138.085 104.840 138.255 ;
        RECT 105.030 138.135 105.740 138.755 ;
        RECT 105.910 138.425 106.260 138.995 ;
        RECT 106.435 138.865 106.775 139.495 ;
        RECT 106.945 138.865 107.195 139.665 ;
        RECT 107.385 139.015 107.715 139.495 ;
        RECT 107.885 139.205 108.110 139.665 ;
        RECT 108.280 139.015 108.610 139.495 ;
        RECT 106.435 138.815 106.665 138.865 ;
        RECT 107.385 138.845 108.610 139.015 ;
        RECT 109.240 138.885 109.740 139.495 ;
        RECT 110.115 138.895 111.785 139.665 ;
        RECT 106.435 138.255 106.610 138.815 ;
        RECT 106.780 138.505 107.475 138.675 ;
        RECT 107.305 138.255 107.475 138.505 ;
        RECT 107.650 138.475 108.070 138.675 ;
        RECT 108.240 138.475 108.570 138.675 ;
        RECT 108.740 138.475 109.070 138.675 ;
        RECT 109.240 138.255 109.410 138.885 ;
        RECT 109.595 138.425 109.945 138.675 ;
        RECT 104.670 137.965 104.840 138.085 ;
        RECT 105.940 137.965 106.260 138.255 ;
        RECT 104.155 137.115 104.435 137.915 ;
        RECT 104.670 137.795 106.260 137.965 ;
        RECT 104.605 137.335 106.260 137.625 ;
        RECT 106.435 137.285 106.775 138.255 ;
        RECT 106.945 137.115 107.115 138.255 ;
        RECT 107.305 138.085 109.740 138.255 ;
        RECT 107.385 137.115 107.635 137.915 ;
        RECT 108.280 137.285 108.610 138.085 ;
        RECT 108.910 137.115 109.240 137.915 ;
        RECT 109.410 137.285 109.740 138.085 ;
        RECT 110.115 138.205 110.865 138.725 ;
        RECT 111.035 138.375 111.785 138.895 ;
        RECT 112.230 138.855 112.475 139.460 ;
        RECT 112.695 139.130 113.205 139.665 ;
        RECT 111.955 138.685 113.185 138.855 ;
        RECT 110.115 137.115 111.785 138.205 ;
        RECT 111.955 137.875 112.295 138.685 ;
        RECT 112.465 138.120 113.215 138.310 ;
        RECT 111.955 137.465 112.470 137.875 ;
        RECT 112.705 137.115 112.875 137.875 ;
        RECT 113.045 137.455 113.215 138.120 ;
        RECT 113.385 138.135 113.575 139.495 ;
        RECT 113.745 138.985 114.020 139.495 ;
        RECT 114.210 139.130 114.740 139.495 ;
        RECT 115.165 139.265 115.495 139.665 ;
        RECT 114.565 139.095 114.740 139.130 ;
        RECT 113.745 138.815 114.025 138.985 ;
        RECT 113.745 138.335 114.020 138.815 ;
        RECT 114.225 138.135 114.395 138.935 ;
        RECT 113.385 137.965 114.395 138.135 ;
        RECT 114.565 138.925 115.495 139.095 ;
        RECT 115.665 138.925 115.920 139.495 ;
        RECT 116.095 138.940 116.385 139.665 ;
        RECT 114.565 137.795 114.735 138.925 ;
        RECT 115.325 138.755 115.495 138.925 ;
        RECT 113.610 137.625 114.735 137.795 ;
        RECT 114.905 138.425 115.100 138.755 ;
        RECT 115.325 138.425 115.580 138.755 ;
        RECT 114.905 137.455 115.075 138.425 ;
        RECT 115.750 138.255 115.920 138.925 ;
        RECT 116.595 138.845 116.825 139.665 ;
        RECT 116.995 138.865 117.325 139.495 ;
        RECT 116.575 138.425 116.905 138.675 ;
        RECT 113.045 137.285 115.075 137.455 ;
        RECT 115.245 137.115 115.415 138.255 ;
        RECT 115.585 137.285 115.920 138.255 ;
        RECT 116.095 137.115 116.385 138.280 ;
        RECT 117.075 138.265 117.325 138.865 ;
        RECT 117.495 138.845 117.705 139.665 ;
        RECT 118.310 139.325 118.565 139.485 ;
        RECT 118.225 139.155 118.565 139.325 ;
        RECT 118.745 139.205 119.030 139.665 ;
        RECT 118.310 138.955 118.565 139.155 ;
        RECT 116.595 137.115 116.825 138.255 ;
        RECT 116.995 137.285 117.325 138.265 ;
        RECT 117.495 137.115 117.705 138.255 ;
        RECT 118.310 138.095 118.490 138.955 ;
        RECT 119.210 138.755 119.460 139.405 ;
        RECT 118.660 138.425 119.460 138.755 ;
        RECT 118.310 137.425 118.565 138.095 ;
        RECT 118.745 137.115 119.030 137.915 ;
        RECT 119.210 137.835 119.460 138.425 ;
        RECT 119.660 139.070 119.980 139.400 ;
        RECT 120.160 139.185 120.820 139.665 ;
        RECT 121.020 139.275 121.870 139.445 ;
        RECT 119.660 138.175 119.850 139.070 ;
        RECT 120.170 138.745 120.830 139.015 ;
        RECT 120.500 138.685 120.830 138.745 ;
        RECT 120.020 138.515 120.350 138.575 ;
        RECT 121.020 138.515 121.190 139.275 ;
        RECT 122.430 139.205 122.750 139.665 ;
        RECT 122.950 139.025 123.200 139.455 ;
        RECT 123.490 139.225 123.900 139.665 ;
        RECT 124.070 139.285 125.085 139.485 ;
        RECT 121.360 138.855 122.610 139.025 ;
        RECT 121.360 138.735 121.690 138.855 ;
        RECT 120.020 138.345 121.920 138.515 ;
        RECT 119.660 138.005 121.580 138.175 ;
        RECT 119.660 137.985 119.980 138.005 ;
        RECT 119.210 137.325 119.540 137.835 ;
        RECT 119.810 137.375 119.980 137.985 ;
        RECT 121.750 137.835 121.920 138.345 ;
        RECT 122.090 138.275 122.270 138.685 ;
        RECT 122.440 138.095 122.610 138.855 ;
        RECT 120.150 137.115 120.480 137.805 ;
        RECT 120.710 137.665 121.920 137.835 ;
        RECT 122.090 137.785 122.610 138.095 ;
        RECT 122.780 138.685 123.200 139.025 ;
        RECT 123.490 138.685 123.900 139.015 ;
        RECT 122.780 137.915 122.970 138.685 ;
        RECT 124.070 138.555 124.240 139.285 ;
        RECT 125.385 139.115 125.555 139.445 ;
        RECT 125.725 139.285 126.055 139.665 ;
        RECT 124.410 138.735 124.760 139.105 ;
        RECT 124.070 138.515 124.490 138.555 ;
        RECT 123.140 138.345 124.490 138.515 ;
        RECT 123.140 138.185 123.390 138.345 ;
        RECT 123.900 137.915 124.150 138.175 ;
        RECT 122.780 137.665 124.150 137.915 ;
        RECT 120.710 137.375 120.950 137.665 ;
        RECT 121.750 137.585 121.920 137.665 ;
        RECT 121.150 137.115 121.570 137.495 ;
        RECT 121.750 137.335 122.380 137.585 ;
        RECT 122.850 137.115 123.180 137.495 ;
        RECT 123.350 137.375 123.520 137.665 ;
        RECT 124.320 137.500 124.490 138.345 ;
        RECT 124.940 138.175 125.160 139.045 ;
        RECT 125.385 138.925 126.080 139.115 ;
        RECT 124.660 137.795 125.160 138.175 ;
        RECT 125.330 138.125 125.740 138.745 ;
        RECT 125.910 137.955 126.080 138.925 ;
        RECT 125.385 137.785 126.080 137.955 ;
        RECT 123.700 137.115 124.080 137.495 ;
        RECT 124.320 137.330 125.150 137.500 ;
        RECT 125.385 137.285 125.555 137.785 ;
        RECT 125.725 137.115 126.055 137.615 ;
        RECT 126.270 137.285 126.495 139.405 ;
        RECT 126.665 139.285 126.995 139.665 ;
        RECT 127.165 139.115 127.335 139.405 ;
        RECT 126.670 138.945 127.335 139.115 ;
        RECT 126.670 137.955 126.900 138.945 ;
        RECT 128.055 138.915 129.265 139.665 ;
        RECT 127.070 138.125 127.420 138.775 ;
        RECT 128.055 138.205 128.575 138.745 ;
        RECT 128.745 138.375 129.265 138.915 ;
        RECT 126.670 137.785 127.335 137.955 ;
        RECT 126.665 137.115 126.995 137.615 ;
        RECT 127.165 137.285 127.335 137.785 ;
        RECT 128.055 137.115 129.265 138.205 ;
        RECT 9.290 136.945 129.350 137.115 ;
        RECT 9.375 135.855 10.585 136.945 ;
        RECT 9.375 135.145 9.895 135.685 ;
        RECT 10.065 135.315 10.585 135.855 ;
        RECT 11.215 135.855 14.725 136.945 ;
        RECT 14.900 136.510 20.245 136.945 ;
        RECT 20.420 136.510 25.765 136.945 ;
        RECT 11.215 135.335 12.905 135.855 ;
        RECT 13.075 135.165 14.725 135.685 ;
        RECT 16.490 135.260 16.840 136.510 ;
        RECT 9.375 134.395 10.585 135.145 ;
        RECT 11.215 134.395 14.725 135.165 ;
        RECT 18.320 134.940 18.660 135.770 ;
        RECT 22.010 135.260 22.360 136.510 ;
        RECT 25.935 135.780 26.225 136.945 ;
        RECT 26.855 135.855 28.525 136.945 ;
        RECT 28.700 136.510 34.045 136.945 ;
        RECT 34.220 136.510 39.565 136.945 ;
        RECT 23.840 134.940 24.180 135.770 ;
        RECT 26.855 135.335 27.605 135.855 ;
        RECT 27.775 135.165 28.525 135.685 ;
        RECT 30.290 135.260 30.640 136.510 ;
        RECT 14.900 134.395 20.245 134.940 ;
        RECT 20.420 134.395 25.765 134.940 ;
        RECT 25.935 134.395 26.225 135.120 ;
        RECT 26.855 134.395 28.525 135.165 ;
        RECT 32.120 134.940 32.460 135.770 ;
        RECT 35.810 135.260 36.160 136.510 ;
        RECT 39.775 135.805 40.005 136.945 ;
        RECT 40.175 135.795 40.505 136.775 ;
        RECT 40.675 135.805 40.885 136.945 ;
        RECT 41.490 135.965 41.745 136.635 ;
        RECT 41.925 136.145 42.210 136.945 ;
        RECT 42.390 136.225 42.720 136.735 ;
        RECT 37.640 134.940 37.980 135.770 ;
        RECT 39.755 135.385 40.085 135.635 ;
        RECT 28.700 134.395 34.045 134.940 ;
        RECT 34.220 134.395 39.565 134.940 ;
        RECT 39.775 134.395 40.005 135.215 ;
        RECT 40.255 135.195 40.505 135.795 ;
        RECT 40.175 134.565 40.505 135.195 ;
        RECT 40.675 134.395 40.885 135.215 ;
        RECT 41.490 135.105 41.670 135.965 ;
        RECT 42.390 135.635 42.640 136.225 ;
        RECT 42.990 136.075 43.160 136.685 ;
        RECT 43.330 136.255 43.660 136.945 ;
        RECT 43.890 136.395 44.130 136.685 ;
        RECT 44.330 136.565 44.750 136.945 ;
        RECT 44.930 136.475 45.560 136.725 ;
        RECT 46.030 136.565 46.360 136.945 ;
        RECT 44.930 136.395 45.100 136.475 ;
        RECT 46.530 136.395 46.700 136.685 ;
        RECT 46.880 136.565 47.260 136.945 ;
        RECT 47.500 136.560 48.330 136.730 ;
        RECT 43.890 136.225 45.100 136.395 ;
        RECT 41.840 135.305 42.640 135.635 ;
        RECT 41.490 134.905 41.745 135.105 ;
        RECT 41.405 134.735 41.745 134.905 ;
        RECT 41.490 134.575 41.745 134.735 ;
        RECT 41.925 134.395 42.210 134.855 ;
        RECT 42.390 134.655 42.640 135.305 ;
        RECT 42.840 136.055 43.160 136.075 ;
        RECT 42.840 135.885 44.760 136.055 ;
        RECT 42.840 134.990 43.030 135.885 ;
        RECT 44.930 135.715 45.100 136.225 ;
        RECT 45.270 135.965 45.790 136.275 ;
        RECT 43.200 135.545 45.100 135.715 ;
        RECT 43.200 135.485 43.530 135.545 ;
        RECT 43.680 135.315 44.010 135.375 ;
        RECT 43.350 135.045 44.010 135.315 ;
        RECT 42.840 134.660 43.160 134.990 ;
        RECT 43.340 134.395 44.000 134.875 ;
        RECT 44.200 134.785 44.370 135.545 ;
        RECT 45.270 135.375 45.450 135.785 ;
        RECT 44.540 135.205 44.870 135.325 ;
        RECT 45.620 135.205 45.790 135.965 ;
        RECT 44.540 135.035 45.790 135.205 ;
        RECT 45.960 136.145 47.330 136.395 ;
        RECT 45.960 135.375 46.150 136.145 ;
        RECT 47.080 135.885 47.330 136.145 ;
        RECT 46.320 135.715 46.570 135.875 ;
        RECT 47.500 135.715 47.670 136.560 ;
        RECT 48.565 136.275 48.735 136.775 ;
        RECT 48.905 136.445 49.235 136.945 ;
        RECT 47.840 135.885 48.340 136.265 ;
        RECT 48.565 136.105 49.260 136.275 ;
        RECT 46.320 135.545 47.670 135.715 ;
        RECT 47.250 135.505 47.670 135.545 ;
        RECT 45.960 135.035 46.380 135.375 ;
        RECT 46.670 135.045 47.080 135.375 ;
        RECT 44.200 134.615 45.050 134.785 ;
        RECT 45.610 134.395 45.930 134.855 ;
        RECT 46.130 134.605 46.380 135.035 ;
        RECT 46.670 134.395 47.080 134.835 ;
        RECT 47.250 134.775 47.420 135.505 ;
        RECT 47.590 134.955 47.940 135.325 ;
        RECT 48.120 135.015 48.340 135.885 ;
        RECT 48.510 135.315 48.920 135.935 ;
        RECT 49.090 135.135 49.260 136.105 ;
        RECT 48.565 134.945 49.260 135.135 ;
        RECT 47.250 134.575 48.265 134.775 ;
        RECT 48.565 134.615 48.735 134.945 ;
        RECT 48.905 134.395 49.235 134.775 ;
        RECT 49.450 134.655 49.675 136.775 ;
        RECT 49.845 136.445 50.175 136.945 ;
        RECT 50.345 136.275 50.515 136.775 ;
        RECT 49.850 136.105 50.515 136.275 ;
        RECT 49.850 135.115 50.080 136.105 ;
        RECT 50.250 135.285 50.600 135.935 ;
        RECT 51.695 135.780 51.985 136.945 ;
        RECT 53.080 136.510 58.425 136.945 ;
        RECT 58.600 136.510 63.945 136.945 ;
        RECT 54.670 135.260 55.020 136.510 ;
        RECT 49.850 134.945 50.515 135.115 ;
        RECT 49.845 134.395 50.175 134.775 ;
        RECT 50.345 134.655 50.515 134.945 ;
        RECT 51.695 134.395 51.985 135.120 ;
        RECT 56.500 134.940 56.840 135.770 ;
        RECT 60.190 135.260 60.540 136.510 ;
        RECT 64.115 135.805 64.455 136.775 ;
        RECT 64.625 135.805 64.795 136.945 ;
        RECT 65.065 136.145 65.315 136.945 ;
        RECT 65.960 135.975 66.290 136.775 ;
        RECT 66.590 136.145 66.920 136.945 ;
        RECT 67.090 135.975 67.420 136.775 ;
        RECT 64.985 135.805 67.420 135.975 ;
        RECT 67.795 136.185 68.310 136.595 ;
        RECT 68.545 136.185 68.715 136.945 ;
        RECT 68.885 136.605 70.915 136.775 ;
        RECT 62.020 134.940 62.360 135.770 ;
        RECT 64.115 135.195 64.290 135.805 ;
        RECT 64.985 135.555 65.155 135.805 ;
        RECT 64.460 135.385 65.155 135.555 ;
        RECT 65.330 135.385 65.750 135.585 ;
        RECT 65.920 135.385 66.250 135.585 ;
        RECT 66.420 135.385 66.750 135.585 ;
        RECT 53.080 134.395 58.425 134.940 ;
        RECT 58.600 134.395 63.945 134.940 ;
        RECT 64.115 134.565 64.455 135.195 ;
        RECT 64.625 134.395 64.875 135.195 ;
        RECT 65.065 135.045 66.290 135.215 ;
        RECT 65.065 134.565 65.395 135.045 ;
        RECT 65.565 134.395 65.790 134.855 ;
        RECT 65.960 134.565 66.290 135.045 ;
        RECT 66.920 135.175 67.090 135.805 ;
        RECT 67.275 135.385 67.625 135.635 ;
        RECT 67.795 135.375 68.135 136.185 ;
        RECT 68.885 135.940 69.055 136.605 ;
        RECT 69.450 136.265 70.575 136.435 ;
        RECT 68.305 135.750 69.055 135.940 ;
        RECT 69.225 135.925 70.235 136.095 ;
        RECT 67.795 135.205 69.025 135.375 ;
        RECT 66.920 134.565 67.420 135.175 ;
        RECT 68.070 134.600 68.315 135.205 ;
        RECT 68.535 134.395 69.045 134.930 ;
        RECT 69.225 134.565 69.415 135.925 ;
        RECT 69.585 135.245 69.860 135.725 ;
        RECT 69.585 135.075 69.865 135.245 ;
        RECT 70.065 135.125 70.235 135.925 ;
        RECT 70.405 135.135 70.575 136.265 ;
        RECT 70.745 135.635 70.915 136.605 ;
        RECT 71.085 135.805 71.255 136.945 ;
        RECT 71.425 135.805 71.760 136.775 ;
        RECT 70.745 135.305 70.940 135.635 ;
        RECT 71.165 135.305 71.420 135.635 ;
        RECT 71.165 135.135 71.335 135.305 ;
        RECT 71.590 135.135 71.760 135.805 ;
        RECT 71.935 135.855 73.145 136.945 ;
        RECT 73.405 136.015 73.575 136.775 ;
        RECT 73.755 136.185 74.085 136.945 ;
        RECT 71.935 135.315 72.455 135.855 ;
        RECT 73.405 135.845 74.070 136.015 ;
        RECT 74.255 135.870 74.525 136.775 ;
        RECT 73.900 135.700 74.070 135.845 ;
        RECT 72.625 135.145 73.145 135.685 ;
        RECT 73.335 135.295 73.665 135.665 ;
        RECT 73.900 135.370 74.185 135.700 ;
        RECT 69.585 134.565 69.860 135.075 ;
        RECT 70.405 134.965 71.335 135.135 ;
        RECT 70.405 134.930 70.580 134.965 ;
        RECT 70.050 134.565 70.580 134.930 ;
        RECT 71.005 134.395 71.335 134.795 ;
        RECT 71.505 134.565 71.760 135.135 ;
        RECT 71.935 134.395 73.145 135.145 ;
        RECT 73.900 135.115 74.070 135.370 ;
        RECT 73.405 134.945 74.070 135.115 ;
        RECT 74.355 135.070 74.525 135.870 ;
        RECT 74.695 135.855 77.285 136.945 ;
        RECT 74.695 135.335 75.905 135.855 ;
        RECT 77.455 135.780 77.745 136.945 ;
        RECT 78.840 136.510 84.185 136.945 ;
        RECT 84.730 136.605 84.985 136.635 ;
        RECT 76.075 135.165 77.285 135.685 ;
        RECT 80.430 135.260 80.780 136.510 ;
        RECT 84.645 136.435 84.985 136.605 ;
        RECT 84.730 135.965 84.985 136.435 ;
        RECT 85.165 136.145 85.450 136.945 ;
        RECT 85.630 136.225 85.960 136.735 ;
        RECT 73.405 134.565 73.575 134.945 ;
        RECT 73.755 134.395 74.085 134.775 ;
        RECT 74.265 134.565 74.525 135.070 ;
        RECT 74.695 134.395 77.285 135.165 ;
        RECT 77.455 134.395 77.745 135.120 ;
        RECT 82.260 134.940 82.600 135.770 ;
        RECT 84.730 135.105 84.910 135.965 ;
        RECT 85.630 135.635 85.880 136.225 ;
        RECT 86.230 136.075 86.400 136.685 ;
        RECT 86.570 136.255 86.900 136.945 ;
        RECT 87.130 136.395 87.370 136.685 ;
        RECT 87.570 136.565 87.990 136.945 ;
        RECT 88.170 136.475 88.800 136.725 ;
        RECT 89.270 136.565 89.600 136.945 ;
        RECT 88.170 136.395 88.340 136.475 ;
        RECT 89.770 136.395 89.940 136.685 ;
        RECT 90.120 136.565 90.500 136.945 ;
        RECT 90.740 136.560 91.570 136.730 ;
        RECT 87.130 136.225 88.340 136.395 ;
        RECT 85.080 135.305 85.880 135.635 ;
        RECT 78.840 134.395 84.185 134.940 ;
        RECT 84.730 134.575 84.985 135.105 ;
        RECT 85.165 134.395 85.450 134.855 ;
        RECT 85.630 134.655 85.880 135.305 ;
        RECT 86.080 136.055 86.400 136.075 ;
        RECT 86.080 135.885 88.000 136.055 ;
        RECT 86.080 134.990 86.270 135.885 ;
        RECT 88.170 135.715 88.340 136.225 ;
        RECT 88.510 135.965 89.030 136.275 ;
        RECT 86.440 135.545 88.340 135.715 ;
        RECT 86.440 135.485 86.770 135.545 ;
        RECT 86.920 135.315 87.250 135.375 ;
        RECT 86.590 135.045 87.250 135.315 ;
        RECT 86.080 134.660 86.400 134.990 ;
        RECT 86.580 134.395 87.240 134.875 ;
        RECT 87.440 134.785 87.610 135.545 ;
        RECT 88.510 135.375 88.690 135.785 ;
        RECT 87.780 135.205 88.110 135.325 ;
        RECT 88.860 135.205 89.030 135.965 ;
        RECT 87.780 135.035 89.030 135.205 ;
        RECT 89.200 136.145 90.570 136.395 ;
        RECT 89.200 135.375 89.390 136.145 ;
        RECT 90.320 135.885 90.570 136.145 ;
        RECT 89.560 135.715 89.810 135.875 ;
        RECT 90.740 135.715 90.910 136.560 ;
        RECT 91.805 136.275 91.975 136.775 ;
        RECT 92.145 136.445 92.475 136.945 ;
        RECT 91.080 135.885 91.580 136.265 ;
        RECT 91.805 136.105 92.500 136.275 ;
        RECT 89.560 135.545 90.910 135.715 ;
        RECT 90.490 135.505 90.910 135.545 ;
        RECT 89.200 135.035 89.620 135.375 ;
        RECT 89.910 135.045 90.320 135.375 ;
        RECT 87.440 134.615 88.290 134.785 ;
        RECT 88.850 134.395 89.170 134.855 ;
        RECT 89.370 134.605 89.620 135.035 ;
        RECT 89.910 134.395 90.320 134.835 ;
        RECT 90.490 134.775 90.660 135.505 ;
        RECT 90.830 134.955 91.180 135.325 ;
        RECT 91.360 135.015 91.580 135.885 ;
        RECT 91.750 135.315 92.160 135.935 ;
        RECT 92.330 135.135 92.500 136.105 ;
        RECT 91.805 134.945 92.500 135.135 ;
        RECT 90.490 134.575 91.505 134.775 ;
        RECT 91.805 134.615 91.975 134.945 ;
        RECT 92.145 134.395 92.475 134.775 ;
        RECT 92.690 134.655 92.915 136.775 ;
        RECT 93.085 136.445 93.415 136.945 ;
        RECT 93.585 136.275 93.755 136.775 ;
        RECT 93.090 136.105 93.755 136.275 ;
        RECT 93.090 135.115 93.320 136.105 ;
        RECT 93.490 135.285 93.840 135.935 ;
        RECT 94.015 135.855 97.525 136.945 ;
        RECT 97.700 136.510 103.045 136.945 ;
        RECT 94.015 135.335 95.705 135.855 ;
        RECT 95.875 135.165 97.525 135.685 ;
        RECT 99.290 135.260 99.640 136.510 ;
        RECT 103.215 135.780 103.505 136.945 ;
        RECT 104.135 135.855 106.725 136.945 ;
        RECT 93.090 134.945 93.755 135.115 ;
        RECT 93.085 134.395 93.415 134.775 ;
        RECT 93.585 134.655 93.755 134.945 ;
        RECT 94.015 134.395 97.525 135.165 ;
        RECT 101.120 134.940 101.460 135.770 ;
        RECT 104.135 135.335 105.345 135.855 ;
        RECT 106.895 135.805 107.165 136.775 ;
        RECT 107.375 136.145 107.655 136.945 ;
        RECT 107.825 136.435 109.480 136.725 ;
        RECT 107.890 136.095 109.480 136.265 ;
        RECT 107.890 135.975 108.060 136.095 ;
        RECT 107.335 135.805 108.060 135.975 ;
        RECT 105.515 135.165 106.725 135.685 ;
        RECT 97.700 134.395 103.045 134.940 ;
        RECT 103.215 134.395 103.505 135.120 ;
        RECT 104.135 134.395 106.725 135.165 ;
        RECT 106.895 135.070 107.065 135.805 ;
        RECT 107.335 135.635 107.505 135.805 ;
        RECT 107.235 135.305 107.505 135.635 ;
        RECT 107.675 135.305 108.080 135.635 ;
        RECT 108.250 135.305 108.960 135.925 ;
        RECT 109.160 135.805 109.480 136.095 ;
        RECT 109.655 135.855 111.325 136.945 ;
        RECT 111.500 136.510 116.845 136.945 ;
        RECT 117.390 136.605 117.645 136.635 ;
        RECT 107.335 135.135 107.505 135.305 ;
        RECT 106.895 134.725 107.165 135.070 ;
        RECT 107.335 134.965 108.945 135.135 ;
        RECT 109.130 135.065 109.480 135.635 ;
        RECT 109.655 135.335 110.405 135.855 ;
        RECT 110.575 135.165 111.325 135.685 ;
        RECT 113.090 135.260 113.440 136.510 ;
        RECT 117.305 136.435 117.645 136.605 ;
        RECT 117.390 135.965 117.645 136.435 ;
        RECT 117.825 136.145 118.110 136.945 ;
        RECT 118.290 136.225 118.620 136.735 ;
        RECT 107.355 134.395 107.735 134.795 ;
        RECT 107.905 134.615 108.075 134.965 ;
        RECT 108.245 134.395 108.575 134.795 ;
        RECT 108.775 134.615 108.945 134.965 ;
        RECT 109.145 134.395 109.475 134.895 ;
        RECT 109.655 134.395 111.325 135.165 ;
        RECT 114.920 134.940 115.260 135.770 ;
        RECT 117.390 135.105 117.570 135.965 ;
        RECT 118.290 135.635 118.540 136.225 ;
        RECT 118.890 136.075 119.060 136.685 ;
        RECT 119.230 136.255 119.560 136.945 ;
        RECT 119.790 136.395 120.030 136.685 ;
        RECT 120.230 136.565 120.650 136.945 ;
        RECT 120.830 136.475 121.460 136.725 ;
        RECT 121.930 136.565 122.260 136.945 ;
        RECT 120.830 136.395 121.000 136.475 ;
        RECT 122.430 136.395 122.600 136.685 ;
        RECT 122.780 136.565 123.160 136.945 ;
        RECT 123.400 136.560 124.230 136.730 ;
        RECT 119.790 136.225 121.000 136.395 ;
        RECT 117.740 135.305 118.540 135.635 ;
        RECT 111.500 134.395 116.845 134.940 ;
        RECT 117.390 134.575 117.645 135.105 ;
        RECT 117.825 134.395 118.110 134.855 ;
        RECT 118.290 134.655 118.540 135.305 ;
        RECT 118.740 136.055 119.060 136.075 ;
        RECT 118.740 135.885 120.660 136.055 ;
        RECT 118.740 134.990 118.930 135.885 ;
        RECT 120.830 135.715 121.000 136.225 ;
        RECT 121.170 135.965 121.690 136.275 ;
        RECT 119.100 135.545 121.000 135.715 ;
        RECT 119.100 135.485 119.430 135.545 ;
        RECT 119.580 135.315 119.910 135.375 ;
        RECT 119.250 135.045 119.910 135.315 ;
        RECT 118.740 134.660 119.060 134.990 ;
        RECT 119.240 134.395 119.900 134.875 ;
        RECT 120.100 134.785 120.270 135.545 ;
        RECT 121.170 135.375 121.350 135.785 ;
        RECT 120.440 135.205 120.770 135.325 ;
        RECT 121.520 135.205 121.690 135.965 ;
        RECT 120.440 135.035 121.690 135.205 ;
        RECT 121.860 136.145 123.230 136.395 ;
        RECT 121.860 135.375 122.050 136.145 ;
        RECT 122.980 135.885 123.230 136.145 ;
        RECT 122.220 135.715 122.470 135.875 ;
        RECT 123.400 135.715 123.570 136.560 ;
        RECT 124.465 136.275 124.635 136.775 ;
        RECT 124.805 136.445 125.135 136.945 ;
        RECT 123.740 135.885 124.240 136.265 ;
        RECT 124.465 136.105 125.160 136.275 ;
        RECT 122.220 135.545 123.570 135.715 ;
        RECT 123.150 135.505 123.570 135.545 ;
        RECT 121.860 135.035 122.280 135.375 ;
        RECT 122.570 135.045 122.980 135.375 ;
        RECT 120.100 134.615 120.950 134.785 ;
        RECT 121.510 134.395 121.830 134.855 ;
        RECT 122.030 134.605 122.280 135.035 ;
        RECT 122.570 134.395 122.980 134.835 ;
        RECT 123.150 134.775 123.320 135.505 ;
        RECT 123.490 134.955 123.840 135.325 ;
        RECT 124.020 135.015 124.240 135.885 ;
        RECT 124.410 135.315 124.820 135.935 ;
        RECT 124.990 135.135 125.160 136.105 ;
        RECT 124.465 134.945 125.160 135.135 ;
        RECT 123.150 134.575 124.165 134.775 ;
        RECT 124.465 134.615 124.635 134.945 ;
        RECT 124.805 134.395 125.135 134.775 ;
        RECT 125.350 134.655 125.575 136.775 ;
        RECT 125.745 136.445 126.075 136.945 ;
        RECT 126.245 136.275 126.415 136.775 ;
        RECT 125.750 136.105 126.415 136.275 ;
        RECT 125.750 135.115 125.980 136.105 ;
        RECT 126.150 135.285 126.500 135.935 ;
        RECT 126.675 135.855 127.885 136.945 ;
        RECT 128.055 135.855 129.265 136.945 ;
        RECT 126.675 135.315 127.195 135.855 ;
        RECT 127.365 135.145 127.885 135.685 ;
        RECT 128.055 135.315 128.575 135.855 ;
        RECT 128.745 135.145 129.265 135.685 ;
        RECT 125.750 134.945 126.415 135.115 ;
        RECT 125.745 134.395 126.075 134.775 ;
        RECT 126.245 134.655 126.415 134.945 ;
        RECT 126.675 134.395 127.885 135.145 ;
        RECT 128.055 134.395 129.265 135.145 ;
        RECT 9.290 134.225 129.350 134.395 ;
        RECT 9.375 133.475 10.585 134.225 ;
        RECT 9.375 132.935 9.895 133.475 ;
        RECT 11.215 133.455 12.885 134.225 ;
        RECT 13.055 133.500 13.345 134.225 ;
        RECT 13.515 133.455 16.105 134.225 ;
        RECT 10.065 132.765 10.585 133.305 ;
        RECT 9.375 131.675 10.585 132.765 ;
        RECT 11.215 132.765 11.965 133.285 ;
        RECT 12.135 132.935 12.885 133.455 ;
        RECT 11.215 131.675 12.885 132.765 ;
        RECT 13.055 131.675 13.345 132.840 ;
        RECT 13.515 132.765 14.725 133.285 ;
        RECT 14.895 132.935 16.105 133.455 ;
        RECT 16.550 133.415 16.795 134.020 ;
        RECT 17.015 133.690 17.525 134.225 ;
        RECT 16.275 133.245 17.505 133.415 ;
        RECT 13.515 131.675 16.105 132.765 ;
        RECT 16.275 132.435 16.615 133.245 ;
        RECT 16.785 132.680 17.535 132.870 ;
        RECT 16.275 132.025 16.790 132.435 ;
        RECT 17.025 131.675 17.195 132.435 ;
        RECT 17.365 132.015 17.535 132.680 ;
        RECT 17.705 132.695 17.895 134.055 ;
        RECT 18.065 133.205 18.340 134.055 ;
        RECT 18.530 133.690 19.060 134.055 ;
        RECT 19.485 133.825 19.815 134.225 ;
        RECT 18.885 133.655 19.060 133.690 ;
        RECT 18.065 133.035 18.345 133.205 ;
        RECT 18.065 132.895 18.340 133.035 ;
        RECT 18.545 132.695 18.715 133.495 ;
        RECT 17.705 132.525 18.715 132.695 ;
        RECT 18.885 133.485 19.815 133.655 ;
        RECT 19.985 133.485 20.240 134.055 ;
        RECT 20.420 133.680 25.765 134.225 ;
        RECT 18.885 132.355 19.055 133.485 ;
        RECT 19.645 133.315 19.815 133.485 ;
        RECT 17.930 132.185 19.055 132.355 ;
        RECT 19.225 132.985 19.420 133.315 ;
        RECT 19.645 132.985 19.900 133.315 ;
        RECT 19.225 132.015 19.395 132.985 ;
        RECT 20.070 132.815 20.240 133.485 ;
        RECT 17.365 131.845 19.395 132.015 ;
        RECT 19.565 131.675 19.735 132.815 ;
        RECT 19.905 131.845 20.240 132.815 ;
        RECT 22.010 132.110 22.360 133.360 ;
        RECT 23.840 132.850 24.180 133.680 ;
        RECT 26.135 133.595 26.465 133.955 ;
        RECT 27.085 133.765 27.335 134.225 ;
        RECT 27.505 133.765 28.065 134.055 ;
        RECT 26.135 133.405 27.525 133.595 ;
        RECT 27.355 133.315 27.525 133.405 ;
        RECT 25.950 132.985 26.625 133.235 ;
        RECT 26.845 132.985 27.185 133.235 ;
        RECT 27.355 132.985 27.645 133.315 ;
        RECT 25.950 132.625 26.215 132.985 ;
        RECT 27.355 132.735 27.525 132.985 ;
        RECT 26.585 132.565 27.525 132.735 ;
        RECT 20.420 131.675 25.765 132.110 ;
        RECT 26.135 131.675 26.415 132.345 ;
        RECT 26.585 132.015 26.885 132.565 ;
        RECT 27.815 132.395 28.065 133.765 ;
        RECT 28.435 133.595 28.765 133.955 ;
        RECT 29.385 133.765 29.635 134.225 ;
        RECT 29.805 133.765 30.365 134.055 ;
        RECT 28.435 133.405 29.825 133.595 ;
        RECT 29.655 133.315 29.825 133.405 ;
        RECT 28.250 132.985 28.925 133.235 ;
        RECT 29.145 132.985 29.485 133.235 ;
        RECT 29.655 132.985 29.945 133.315 ;
        RECT 28.250 132.625 28.515 132.985 ;
        RECT 29.655 132.735 29.825 132.985 ;
        RECT 27.085 131.675 27.415 132.395 ;
        RECT 27.605 131.845 28.065 132.395 ;
        RECT 28.885 132.565 29.825 132.735 ;
        RECT 28.435 131.675 28.715 132.345 ;
        RECT 28.885 132.015 29.185 132.565 ;
        RECT 30.115 132.395 30.365 133.765 ;
        RECT 30.735 133.595 31.065 133.955 ;
        RECT 31.685 133.765 31.935 134.225 ;
        RECT 32.105 133.765 32.665 134.055 ;
        RECT 30.735 133.405 32.125 133.595 ;
        RECT 31.955 133.315 32.125 133.405 ;
        RECT 30.550 132.985 31.225 133.235 ;
        RECT 31.445 132.985 31.785 133.235 ;
        RECT 31.955 132.985 32.245 133.315 ;
        RECT 30.550 132.625 30.815 132.985 ;
        RECT 31.955 132.735 32.125 132.985 ;
        RECT 29.385 131.675 29.715 132.395 ;
        RECT 29.905 131.845 30.365 132.395 ;
        RECT 31.185 132.565 32.125 132.735 ;
        RECT 30.735 131.675 31.015 132.345 ;
        RECT 31.185 132.015 31.485 132.565 ;
        RECT 32.415 132.395 32.665 133.765 ;
        RECT 33.300 133.680 38.645 134.225 ;
        RECT 31.685 131.675 32.015 132.395 ;
        RECT 32.205 131.845 32.665 132.395 ;
        RECT 34.890 132.110 35.240 133.360 ;
        RECT 36.720 132.850 37.060 133.680 ;
        RECT 38.815 133.500 39.105 134.225 ;
        RECT 39.275 133.455 40.945 134.225 ;
        RECT 33.300 131.675 38.645 132.110 ;
        RECT 38.815 131.675 39.105 132.840 ;
        RECT 39.275 132.765 40.025 133.285 ;
        RECT 40.195 132.935 40.945 133.455 ;
        RECT 41.115 133.550 41.385 133.895 ;
        RECT 41.575 133.825 41.955 134.225 ;
        RECT 42.125 133.655 42.295 134.005 ;
        RECT 42.465 133.825 42.795 134.225 ;
        RECT 42.995 133.655 43.165 134.005 ;
        RECT 43.365 133.725 43.695 134.225 ;
        RECT 41.115 132.815 41.285 133.550 ;
        RECT 41.555 133.485 43.165 133.655 ;
        RECT 41.555 133.315 41.725 133.485 ;
        RECT 41.455 132.985 41.725 133.315 ;
        RECT 41.895 132.985 42.300 133.315 ;
        RECT 41.555 132.815 41.725 132.985 ;
        RECT 42.470 132.865 43.180 133.315 ;
        RECT 43.350 132.985 43.700 133.555 ;
        RECT 43.875 133.455 45.545 134.225 ;
        RECT 39.275 131.675 40.945 132.765 ;
        RECT 41.115 131.845 41.385 132.815 ;
        RECT 41.555 132.645 42.280 132.815 ;
        RECT 42.470 132.695 43.185 132.865 ;
        RECT 42.110 132.525 42.280 132.645 ;
        RECT 43.380 132.525 43.700 132.815 ;
        RECT 41.595 131.675 41.875 132.475 ;
        RECT 42.110 132.355 43.700 132.525 ;
        RECT 43.875 132.765 44.625 133.285 ;
        RECT 44.795 132.935 45.545 133.455 ;
        RECT 45.715 133.425 46.055 134.055 ;
        RECT 46.225 133.425 46.475 134.225 ;
        RECT 46.665 133.575 46.995 134.055 ;
        RECT 47.165 133.765 47.390 134.225 ;
        RECT 47.560 133.575 47.890 134.055 ;
        RECT 45.715 133.375 45.945 133.425 ;
        RECT 46.665 133.405 47.890 133.575 ;
        RECT 48.520 133.445 49.020 134.055 ;
        RECT 49.395 133.550 49.655 134.055 ;
        RECT 49.835 133.845 50.165 134.225 ;
        RECT 50.345 133.675 50.515 134.055 ;
        RECT 45.715 132.815 45.890 133.375 ;
        RECT 46.060 133.065 46.755 133.235 ;
        RECT 46.585 132.815 46.755 133.065 ;
        RECT 46.930 133.035 47.350 133.235 ;
        RECT 47.520 133.035 47.850 133.235 ;
        RECT 48.020 133.035 48.350 133.235 ;
        RECT 48.520 132.815 48.690 133.445 ;
        RECT 48.875 132.985 49.225 133.235 ;
        RECT 42.045 131.895 43.700 132.185 ;
        RECT 43.875 131.675 45.545 132.765 ;
        RECT 45.715 131.845 46.055 132.815 ;
        RECT 46.225 131.675 46.395 132.815 ;
        RECT 46.585 132.645 49.020 132.815 ;
        RECT 46.665 131.675 46.915 132.475 ;
        RECT 47.560 131.845 47.890 132.645 ;
        RECT 48.190 131.675 48.520 132.475 ;
        RECT 48.690 131.845 49.020 132.645 ;
        RECT 49.395 132.750 49.565 133.550 ;
        RECT 49.850 133.505 50.515 133.675 ;
        RECT 49.850 133.250 50.020 133.505 ;
        RECT 51.695 133.455 55.205 134.225 ;
        RECT 49.735 132.920 50.020 133.250 ;
        RECT 50.255 132.955 50.585 133.325 ;
        RECT 49.850 132.775 50.020 132.920 ;
        RECT 49.395 131.845 49.665 132.750 ;
        RECT 49.850 132.605 50.515 132.775 ;
        RECT 49.835 131.675 50.165 132.435 ;
        RECT 50.345 131.845 50.515 132.605 ;
        RECT 51.695 132.765 53.385 133.285 ;
        RECT 53.555 132.935 55.205 133.455 ;
        RECT 55.415 133.405 55.645 134.225 ;
        RECT 55.815 133.425 56.145 134.055 ;
        RECT 55.395 132.985 55.725 133.235 ;
        RECT 55.895 132.825 56.145 133.425 ;
        RECT 56.315 133.405 56.525 134.225 ;
        RECT 56.845 133.675 57.015 134.055 ;
        RECT 57.195 133.845 57.525 134.225 ;
        RECT 56.845 133.505 57.510 133.675 ;
        RECT 57.705 133.550 57.965 134.055 ;
        RECT 59.060 133.680 64.405 134.225 ;
        RECT 56.775 132.955 57.105 133.325 ;
        RECT 57.340 133.250 57.510 133.505 ;
        RECT 51.695 131.675 55.205 132.765 ;
        RECT 55.415 131.675 55.645 132.815 ;
        RECT 55.815 131.845 56.145 132.825 ;
        RECT 57.340 132.920 57.625 133.250 ;
        RECT 56.315 131.675 56.525 132.815 ;
        RECT 57.340 132.775 57.510 132.920 ;
        RECT 56.845 132.605 57.510 132.775 ;
        RECT 57.795 132.750 57.965 133.550 ;
        RECT 56.845 131.845 57.015 132.605 ;
        RECT 57.195 131.675 57.525 132.435 ;
        RECT 57.695 131.845 57.965 132.750 ;
        RECT 60.650 132.110 61.000 133.360 ;
        RECT 62.480 132.850 62.820 133.680 ;
        RECT 64.575 133.500 64.865 134.225 ;
        RECT 65.495 133.455 69.005 134.225 ;
        RECT 69.180 133.680 74.525 134.225 ;
        RECT 74.700 133.680 80.045 134.225 ;
        RECT 59.060 131.675 64.405 132.110 ;
        RECT 64.575 131.675 64.865 132.840 ;
        RECT 65.495 132.765 67.185 133.285 ;
        RECT 67.355 132.935 69.005 133.455 ;
        RECT 65.495 131.675 69.005 132.765 ;
        RECT 70.770 132.110 71.120 133.360 ;
        RECT 72.600 132.850 72.940 133.680 ;
        RECT 76.290 132.110 76.640 133.360 ;
        RECT 78.120 132.850 78.460 133.680 ;
        RECT 80.215 133.425 80.555 134.055 ;
        RECT 80.725 133.425 80.975 134.225 ;
        RECT 81.165 133.575 81.495 134.055 ;
        RECT 81.665 133.765 81.890 134.225 ;
        RECT 82.060 133.575 82.390 134.055 ;
        RECT 80.215 132.815 80.390 133.425 ;
        RECT 81.165 133.405 82.390 133.575 ;
        RECT 83.020 133.445 83.520 134.055 ;
        RECT 80.560 133.065 81.255 133.235 ;
        RECT 81.085 132.815 81.255 133.065 ;
        RECT 81.430 133.035 81.850 133.235 ;
        RECT 82.020 133.035 82.350 133.235 ;
        RECT 82.520 133.035 82.850 133.235 ;
        RECT 83.020 132.815 83.190 133.445 ;
        RECT 84.630 133.415 84.875 134.020 ;
        RECT 85.095 133.690 85.605 134.225 ;
        RECT 84.355 133.245 85.585 133.415 ;
        RECT 83.375 132.985 83.725 133.235 ;
        RECT 69.180 131.675 74.525 132.110 ;
        RECT 74.700 131.675 80.045 132.110 ;
        RECT 80.215 131.845 80.555 132.815 ;
        RECT 80.725 131.675 80.895 132.815 ;
        RECT 81.085 132.645 83.520 132.815 ;
        RECT 81.165 131.675 81.415 132.475 ;
        RECT 82.060 131.845 82.390 132.645 ;
        RECT 82.690 131.675 83.020 132.475 ;
        RECT 83.190 131.845 83.520 132.645 ;
        RECT 84.355 132.435 84.695 133.245 ;
        RECT 84.865 132.680 85.615 132.870 ;
        RECT 84.355 132.025 84.870 132.435 ;
        RECT 85.105 131.675 85.275 132.435 ;
        RECT 85.445 132.015 85.615 132.680 ;
        RECT 85.785 132.695 85.975 134.055 ;
        RECT 86.145 133.205 86.420 134.055 ;
        RECT 86.610 133.690 87.140 134.055 ;
        RECT 87.565 133.825 87.895 134.225 ;
        RECT 86.965 133.655 87.140 133.690 ;
        RECT 86.145 133.035 86.425 133.205 ;
        RECT 86.145 132.895 86.420 133.035 ;
        RECT 86.625 132.695 86.795 133.495 ;
        RECT 85.785 132.525 86.795 132.695 ;
        RECT 86.965 133.485 87.895 133.655 ;
        RECT 88.065 133.485 88.320 134.055 ;
        RECT 89.045 133.675 89.215 134.055 ;
        RECT 89.395 133.845 89.725 134.225 ;
        RECT 89.045 133.505 89.710 133.675 ;
        RECT 89.905 133.550 90.165 134.055 ;
        RECT 86.965 132.355 87.135 133.485 ;
        RECT 87.725 133.315 87.895 133.485 ;
        RECT 86.010 132.185 87.135 132.355 ;
        RECT 87.305 132.985 87.500 133.315 ;
        RECT 87.725 132.985 87.980 133.315 ;
        RECT 87.305 132.015 87.475 132.985 ;
        RECT 88.150 132.815 88.320 133.485 ;
        RECT 88.975 132.955 89.305 133.325 ;
        RECT 89.540 133.250 89.710 133.505 ;
        RECT 85.445 131.845 87.475 132.015 ;
        RECT 87.645 131.675 87.815 132.815 ;
        RECT 87.985 131.845 88.320 132.815 ;
        RECT 89.540 132.920 89.825 133.250 ;
        RECT 89.540 132.775 89.710 132.920 ;
        RECT 89.045 132.605 89.710 132.775 ;
        RECT 89.995 132.750 90.165 133.550 ;
        RECT 90.335 133.500 90.625 134.225 ;
        RECT 90.800 133.680 96.145 134.225 ;
        RECT 89.045 131.845 89.215 132.605 ;
        RECT 89.395 131.675 89.725 132.435 ;
        RECT 89.895 131.845 90.165 132.750 ;
        RECT 90.335 131.675 90.625 132.840 ;
        RECT 92.390 132.110 92.740 133.360 ;
        RECT 94.220 132.850 94.560 133.680 ;
        RECT 96.355 133.405 96.585 134.225 ;
        RECT 96.755 133.425 97.085 134.055 ;
        RECT 96.335 132.985 96.665 133.235 ;
        RECT 96.835 132.825 97.085 133.425 ;
        RECT 97.255 133.405 97.465 134.225 ;
        RECT 97.970 133.415 98.215 134.020 ;
        RECT 98.435 133.690 98.945 134.225 ;
        RECT 90.800 131.675 96.145 132.110 ;
        RECT 96.355 131.675 96.585 132.815 ;
        RECT 96.755 131.845 97.085 132.825 ;
        RECT 97.695 133.245 98.925 133.415 ;
        RECT 97.255 131.675 97.465 132.815 ;
        RECT 97.695 132.435 98.035 133.245 ;
        RECT 98.205 132.680 98.955 132.870 ;
        RECT 97.695 132.025 98.210 132.435 ;
        RECT 98.445 131.675 98.615 132.435 ;
        RECT 98.785 132.015 98.955 132.680 ;
        RECT 99.125 132.695 99.315 134.055 ;
        RECT 99.485 133.205 99.760 134.055 ;
        RECT 99.950 133.690 100.480 134.055 ;
        RECT 100.905 133.825 101.235 134.225 ;
        RECT 100.305 133.655 100.480 133.690 ;
        RECT 99.485 133.035 99.765 133.205 ;
        RECT 99.485 132.895 99.760 133.035 ;
        RECT 99.965 132.695 100.135 133.495 ;
        RECT 99.125 132.525 100.135 132.695 ;
        RECT 100.305 133.485 101.235 133.655 ;
        RECT 101.405 133.485 101.660 134.055 ;
        RECT 102.760 133.680 108.105 134.225 ;
        RECT 100.305 132.355 100.475 133.485 ;
        RECT 101.065 133.315 101.235 133.485 ;
        RECT 99.350 132.185 100.475 132.355 ;
        RECT 100.645 132.985 100.840 133.315 ;
        RECT 101.065 132.985 101.320 133.315 ;
        RECT 100.645 132.015 100.815 132.985 ;
        RECT 101.490 132.815 101.660 133.485 ;
        RECT 98.785 131.845 100.815 132.015 ;
        RECT 100.985 131.675 101.155 132.815 ;
        RECT 101.325 131.845 101.660 132.815 ;
        RECT 104.350 132.110 104.700 133.360 ;
        RECT 106.180 132.850 106.520 133.680 ;
        RECT 108.550 133.415 108.795 134.020 ;
        RECT 109.015 133.690 109.525 134.225 ;
        RECT 108.275 133.245 109.505 133.415 ;
        RECT 108.275 132.435 108.615 133.245 ;
        RECT 108.785 132.680 109.535 132.870 ;
        RECT 102.760 131.675 108.105 132.110 ;
        RECT 108.275 132.025 108.790 132.435 ;
        RECT 109.025 131.675 109.195 132.435 ;
        RECT 109.365 132.015 109.535 132.680 ;
        RECT 109.705 132.695 109.895 134.055 ;
        RECT 110.065 133.885 110.340 134.055 ;
        RECT 110.065 133.715 110.345 133.885 ;
        RECT 110.065 132.895 110.340 133.715 ;
        RECT 110.530 133.690 111.060 134.055 ;
        RECT 111.485 133.825 111.815 134.225 ;
        RECT 110.885 133.655 111.060 133.690 ;
        RECT 110.545 132.695 110.715 133.495 ;
        RECT 109.705 132.525 110.715 132.695 ;
        RECT 110.885 133.485 111.815 133.655 ;
        RECT 111.985 133.485 112.240 134.055 ;
        RECT 112.505 133.675 112.675 134.055 ;
        RECT 112.855 133.845 113.185 134.225 ;
        RECT 112.505 133.505 113.170 133.675 ;
        RECT 113.365 133.550 113.625 134.055 ;
        RECT 110.885 132.355 111.055 133.485 ;
        RECT 111.645 133.315 111.815 133.485 ;
        RECT 109.930 132.185 111.055 132.355 ;
        RECT 111.225 132.985 111.420 133.315 ;
        RECT 111.645 132.985 111.900 133.315 ;
        RECT 111.225 132.015 111.395 132.985 ;
        RECT 112.070 132.815 112.240 133.485 ;
        RECT 112.435 132.955 112.765 133.325 ;
        RECT 113.000 133.250 113.170 133.505 ;
        RECT 109.365 131.845 111.395 132.015 ;
        RECT 111.565 131.675 111.735 132.815 ;
        RECT 111.905 131.845 112.240 132.815 ;
        RECT 113.000 132.920 113.285 133.250 ;
        RECT 113.000 132.775 113.170 132.920 ;
        RECT 112.505 132.605 113.170 132.775 ;
        RECT 113.455 132.750 113.625 133.550 ;
        RECT 114.255 133.455 115.925 134.225 ;
        RECT 116.095 133.500 116.385 134.225 ;
        RECT 117.020 133.680 122.365 134.225 ;
        RECT 112.505 131.845 112.675 132.605 ;
        RECT 112.855 131.675 113.185 132.435 ;
        RECT 113.355 131.845 113.625 132.750 ;
        RECT 114.255 132.765 115.005 133.285 ;
        RECT 115.175 132.935 115.925 133.455 ;
        RECT 114.255 131.675 115.925 132.765 ;
        RECT 116.095 131.675 116.385 132.840 ;
        RECT 118.610 132.110 118.960 133.360 ;
        RECT 120.440 132.850 120.780 133.680 ;
        RECT 122.625 133.675 122.795 134.055 ;
        RECT 122.975 133.845 123.305 134.225 ;
        RECT 122.625 133.505 123.290 133.675 ;
        RECT 123.485 133.550 123.745 134.055 ;
        RECT 122.555 132.955 122.885 133.325 ;
        RECT 123.120 133.250 123.290 133.505 ;
        RECT 123.120 132.920 123.405 133.250 ;
        RECT 123.120 132.775 123.290 132.920 ;
        RECT 122.625 132.605 123.290 132.775 ;
        RECT 123.575 132.750 123.745 133.550 ;
        RECT 124.375 133.455 127.885 134.225 ;
        RECT 128.055 133.475 129.265 134.225 ;
        RECT 117.020 131.675 122.365 132.110 ;
        RECT 122.625 131.845 122.795 132.605 ;
        RECT 122.975 131.675 123.305 132.435 ;
        RECT 123.475 131.845 123.745 132.750 ;
        RECT 124.375 132.765 126.065 133.285 ;
        RECT 126.235 132.935 127.885 133.455 ;
        RECT 128.055 132.765 128.575 133.305 ;
        RECT 128.745 132.935 129.265 133.475 ;
        RECT 124.375 131.675 127.885 132.765 ;
        RECT 128.055 131.675 129.265 132.765 ;
        RECT 9.290 131.505 129.350 131.675 ;
        RECT 9.375 130.415 10.585 131.505 ;
        RECT 12.050 130.525 12.305 131.195 ;
        RECT 12.485 130.705 12.770 131.505 ;
        RECT 12.950 130.785 13.280 131.295 ;
        RECT 12.050 130.485 12.230 130.525 ;
        RECT 9.375 129.705 9.895 130.245 ;
        RECT 10.065 129.875 10.585 130.415 ;
        RECT 11.965 130.315 12.230 130.485 ;
        RECT 9.375 128.955 10.585 129.705 ;
        RECT 12.050 129.665 12.230 130.315 ;
        RECT 12.950 130.195 13.200 130.785 ;
        RECT 13.550 130.635 13.720 131.245 ;
        RECT 13.890 130.815 14.220 131.505 ;
        RECT 14.450 130.955 14.690 131.245 ;
        RECT 14.890 131.125 15.310 131.505 ;
        RECT 15.490 131.035 16.120 131.285 ;
        RECT 16.590 131.125 16.920 131.505 ;
        RECT 15.490 130.955 15.660 131.035 ;
        RECT 17.090 130.955 17.260 131.245 ;
        RECT 17.440 131.125 17.820 131.505 ;
        RECT 18.060 131.120 18.890 131.290 ;
        RECT 14.450 130.785 15.660 130.955 ;
        RECT 12.400 129.865 13.200 130.195 ;
        RECT 12.050 129.135 12.305 129.665 ;
        RECT 12.485 128.955 12.770 129.415 ;
        RECT 12.950 129.215 13.200 129.865 ;
        RECT 13.400 130.615 13.720 130.635 ;
        RECT 13.400 130.445 15.320 130.615 ;
        RECT 13.400 129.550 13.590 130.445 ;
        RECT 15.490 130.275 15.660 130.785 ;
        RECT 15.830 130.525 16.350 130.835 ;
        RECT 13.760 130.105 15.660 130.275 ;
        RECT 13.760 130.045 14.090 130.105 ;
        RECT 14.240 129.875 14.570 129.935 ;
        RECT 13.910 129.605 14.570 129.875 ;
        RECT 13.400 129.220 13.720 129.550 ;
        RECT 13.900 128.955 14.560 129.435 ;
        RECT 14.760 129.345 14.930 130.105 ;
        RECT 15.830 129.935 16.010 130.345 ;
        RECT 15.100 129.765 15.430 129.885 ;
        RECT 16.180 129.765 16.350 130.525 ;
        RECT 15.100 129.595 16.350 129.765 ;
        RECT 16.520 130.705 17.890 130.955 ;
        RECT 16.520 129.935 16.710 130.705 ;
        RECT 17.640 130.445 17.890 130.705 ;
        RECT 16.880 130.275 17.130 130.435 ;
        RECT 18.060 130.275 18.230 131.120 ;
        RECT 19.125 130.835 19.295 131.335 ;
        RECT 19.465 131.005 19.795 131.505 ;
        RECT 18.400 130.445 18.900 130.825 ;
        RECT 19.125 130.665 19.820 130.835 ;
        RECT 16.880 130.105 18.230 130.275 ;
        RECT 17.810 130.065 18.230 130.105 ;
        RECT 16.520 129.595 16.940 129.935 ;
        RECT 17.230 129.605 17.640 129.935 ;
        RECT 14.760 129.175 15.610 129.345 ;
        RECT 16.170 128.955 16.490 129.415 ;
        RECT 16.690 129.165 16.940 129.595 ;
        RECT 17.230 128.955 17.640 129.395 ;
        RECT 17.810 129.335 17.980 130.065 ;
        RECT 18.150 129.515 18.500 129.885 ;
        RECT 18.680 129.575 18.900 130.445 ;
        RECT 19.070 129.875 19.480 130.495 ;
        RECT 19.650 129.695 19.820 130.665 ;
        RECT 19.125 129.505 19.820 129.695 ;
        RECT 17.810 129.135 18.825 129.335 ;
        RECT 19.125 129.175 19.295 129.505 ;
        RECT 19.465 128.955 19.795 129.335 ;
        RECT 20.010 129.215 20.235 131.335 ;
        RECT 20.405 131.005 20.735 131.505 ;
        RECT 20.905 130.835 21.075 131.335 ;
        RECT 20.410 130.665 21.075 130.835 ;
        RECT 20.410 129.675 20.640 130.665 ;
        RECT 20.810 129.845 21.160 130.495 ;
        RECT 21.335 130.430 21.605 131.335 ;
        RECT 21.775 130.745 22.105 131.505 ;
        RECT 22.285 130.575 22.455 131.335 ;
        RECT 20.410 129.505 21.075 129.675 ;
        RECT 20.405 128.955 20.735 129.335 ;
        RECT 20.905 129.215 21.075 129.505 ;
        RECT 21.335 129.630 21.505 130.430 ;
        RECT 21.790 130.405 22.455 130.575 ;
        RECT 23.175 130.430 23.445 131.335 ;
        RECT 23.615 130.745 23.945 131.505 ;
        RECT 24.125 130.575 24.295 131.335 ;
        RECT 21.790 130.260 21.960 130.405 ;
        RECT 21.675 129.930 21.960 130.260 ;
        RECT 21.790 129.675 21.960 129.930 ;
        RECT 22.195 129.855 22.525 130.225 ;
        RECT 21.335 129.125 21.595 129.630 ;
        RECT 21.790 129.505 22.455 129.675 ;
        RECT 21.775 128.955 22.105 129.335 ;
        RECT 22.285 129.125 22.455 129.505 ;
        RECT 23.175 129.630 23.345 130.430 ;
        RECT 23.630 130.405 24.295 130.575 ;
        RECT 24.555 130.415 25.765 131.505 ;
        RECT 23.630 130.260 23.800 130.405 ;
        RECT 23.515 129.930 23.800 130.260 ;
        RECT 23.630 129.675 23.800 129.930 ;
        RECT 24.035 129.855 24.365 130.225 ;
        RECT 24.555 129.875 25.075 130.415 ;
        RECT 25.935 130.340 26.225 131.505 ;
        RECT 27.315 130.415 30.825 131.505 ;
        RECT 31.085 130.575 31.255 131.335 ;
        RECT 31.435 130.745 31.765 131.505 ;
        RECT 25.245 129.705 25.765 130.245 ;
        RECT 27.315 129.895 29.005 130.415 ;
        RECT 31.085 130.405 31.750 130.575 ;
        RECT 31.935 130.430 32.205 131.335 ;
        RECT 32.575 130.835 32.855 131.505 ;
        RECT 33.025 130.615 33.325 131.165 ;
        RECT 33.525 130.785 33.855 131.505 ;
        RECT 34.045 130.785 34.505 131.335 ;
        RECT 31.580 130.260 31.750 130.405 ;
        RECT 29.175 129.725 30.825 130.245 ;
        RECT 31.015 129.855 31.345 130.225 ;
        RECT 31.580 129.930 31.865 130.260 ;
        RECT 23.175 129.125 23.435 129.630 ;
        RECT 23.630 129.505 24.295 129.675 ;
        RECT 23.615 128.955 23.945 129.335 ;
        RECT 24.125 129.125 24.295 129.505 ;
        RECT 24.555 128.955 25.765 129.705 ;
        RECT 25.935 128.955 26.225 129.680 ;
        RECT 27.315 128.955 30.825 129.725 ;
        RECT 31.580 129.675 31.750 129.930 ;
        RECT 31.085 129.505 31.750 129.675 ;
        RECT 32.035 129.630 32.205 130.430 ;
        RECT 32.390 130.195 32.655 130.555 ;
        RECT 33.025 130.445 33.965 130.615 ;
        RECT 33.795 130.195 33.965 130.445 ;
        RECT 32.390 129.945 33.065 130.195 ;
        RECT 33.285 129.945 33.625 130.195 ;
        RECT 33.795 129.865 34.085 130.195 ;
        RECT 33.795 129.775 33.965 129.865 ;
        RECT 31.085 129.125 31.255 129.505 ;
        RECT 31.435 128.955 31.765 129.335 ;
        RECT 31.945 129.125 32.205 129.630 ;
        RECT 32.575 129.585 33.965 129.775 ;
        RECT 32.575 129.225 32.905 129.585 ;
        RECT 34.255 129.415 34.505 130.785 ;
        RECT 34.675 130.415 36.345 131.505 ;
        RECT 34.675 129.895 35.425 130.415 ;
        RECT 36.515 130.365 36.785 131.335 ;
        RECT 36.995 130.705 37.275 131.505 ;
        RECT 37.445 130.995 39.100 131.285 ;
        RECT 37.510 130.655 39.100 130.825 ;
        RECT 37.510 130.535 37.680 130.655 ;
        RECT 36.955 130.365 37.680 130.535 ;
        RECT 35.595 129.725 36.345 130.245 ;
        RECT 33.525 128.955 33.775 129.415 ;
        RECT 33.945 129.125 34.505 129.415 ;
        RECT 34.675 128.955 36.345 129.725 ;
        RECT 36.515 129.630 36.685 130.365 ;
        RECT 36.955 130.195 37.125 130.365 ;
        RECT 36.855 129.865 37.125 130.195 ;
        RECT 37.295 129.865 37.700 130.195 ;
        RECT 37.870 129.865 38.580 130.485 ;
        RECT 38.780 130.365 39.100 130.655 ;
        RECT 39.275 130.365 39.545 131.335 ;
        RECT 39.755 130.705 40.035 131.505 ;
        RECT 40.205 130.995 41.860 131.285 ;
        RECT 40.270 130.655 41.860 130.825 ;
        RECT 40.270 130.535 40.440 130.655 ;
        RECT 39.715 130.365 40.440 130.535 ;
        RECT 36.955 129.695 37.125 129.865 ;
        RECT 36.515 129.285 36.785 129.630 ;
        RECT 36.955 129.525 38.565 129.695 ;
        RECT 38.750 129.625 39.100 130.195 ;
        RECT 39.275 129.630 39.445 130.365 ;
        RECT 39.715 130.195 39.885 130.365 ;
        RECT 39.615 129.865 39.885 130.195 ;
        RECT 40.055 129.865 40.460 130.195 ;
        RECT 40.630 129.865 41.340 130.485 ;
        RECT 41.540 130.365 41.860 130.655 ;
        RECT 42.035 130.415 43.705 131.505 ;
        RECT 39.715 129.695 39.885 129.865 ;
        RECT 36.975 128.955 37.355 129.355 ;
        RECT 37.525 129.175 37.695 129.525 ;
        RECT 37.865 128.955 38.195 129.355 ;
        RECT 38.395 129.175 38.565 129.525 ;
        RECT 38.765 128.955 39.095 129.455 ;
        RECT 39.275 129.285 39.545 129.630 ;
        RECT 39.715 129.525 41.325 129.695 ;
        RECT 41.510 129.625 41.860 130.195 ;
        RECT 42.035 129.895 42.785 130.415 ;
        RECT 43.875 130.365 44.215 131.335 ;
        RECT 44.385 130.365 44.555 131.505 ;
        RECT 44.825 130.705 45.075 131.505 ;
        RECT 45.720 130.535 46.050 131.335 ;
        RECT 46.350 130.705 46.680 131.505 ;
        RECT 46.850 130.535 47.180 131.335 ;
        RECT 44.745 130.365 47.180 130.535 ;
        RECT 47.555 130.745 48.070 131.155 ;
        RECT 48.305 130.745 48.475 131.505 ;
        RECT 48.645 131.165 50.675 131.335 ;
        RECT 42.955 129.725 43.705 130.245 ;
        RECT 39.735 128.955 40.115 129.355 ;
        RECT 40.285 129.175 40.455 129.525 ;
        RECT 40.625 128.955 40.955 129.355 ;
        RECT 41.155 129.175 41.325 129.525 ;
        RECT 41.525 128.955 41.855 129.455 ;
        RECT 42.035 128.955 43.705 129.725 ;
        RECT 43.875 129.805 44.050 130.365 ;
        RECT 44.745 130.115 44.915 130.365 ;
        RECT 44.220 129.945 44.915 130.115 ;
        RECT 45.090 129.945 45.510 130.145 ;
        RECT 45.680 129.945 46.010 130.145 ;
        RECT 46.180 129.945 46.510 130.145 ;
        RECT 43.875 129.755 44.105 129.805 ;
        RECT 43.875 129.125 44.215 129.755 ;
        RECT 44.385 128.955 44.635 129.755 ;
        RECT 44.825 129.605 46.050 129.775 ;
        RECT 44.825 129.125 45.155 129.605 ;
        RECT 45.325 128.955 45.550 129.415 ;
        RECT 45.720 129.125 46.050 129.605 ;
        RECT 46.680 129.735 46.850 130.365 ;
        RECT 47.035 129.945 47.385 130.195 ;
        RECT 47.555 129.935 47.895 130.745 ;
        RECT 48.645 130.500 48.815 131.165 ;
        RECT 49.210 130.825 50.335 130.995 ;
        RECT 48.065 130.310 48.815 130.500 ;
        RECT 48.985 130.485 49.995 130.655 ;
        RECT 47.555 129.765 48.785 129.935 ;
        RECT 46.680 129.125 47.180 129.735 ;
        RECT 47.830 129.160 48.075 129.765 ;
        RECT 48.295 128.955 48.805 129.490 ;
        RECT 48.985 129.125 49.175 130.485 ;
        RECT 49.345 130.145 49.620 130.285 ;
        RECT 49.345 129.975 49.625 130.145 ;
        RECT 49.345 129.125 49.620 129.975 ;
        RECT 49.825 129.685 49.995 130.485 ;
        RECT 50.165 129.695 50.335 130.825 ;
        RECT 50.505 130.195 50.675 131.165 ;
        RECT 50.845 130.365 51.015 131.505 ;
        RECT 51.185 130.365 51.520 131.335 ;
        RECT 50.505 129.865 50.700 130.195 ;
        RECT 50.925 129.865 51.180 130.195 ;
        RECT 50.925 129.695 51.095 129.865 ;
        RECT 51.350 129.695 51.520 130.365 ;
        RECT 51.695 130.340 51.985 131.505 ;
        RECT 52.530 130.525 52.785 131.195 ;
        RECT 52.965 130.705 53.250 131.505 ;
        RECT 53.430 130.785 53.760 131.295 ;
        RECT 50.165 129.525 51.095 129.695 ;
        RECT 50.165 129.490 50.340 129.525 ;
        RECT 49.810 129.125 50.340 129.490 ;
        RECT 50.765 128.955 51.095 129.355 ;
        RECT 51.265 129.125 51.520 129.695 ;
        RECT 51.695 128.955 51.985 129.680 ;
        RECT 52.530 129.665 52.710 130.525 ;
        RECT 53.430 130.195 53.680 130.785 ;
        RECT 54.030 130.635 54.200 131.245 ;
        RECT 54.370 130.815 54.700 131.505 ;
        RECT 54.930 130.955 55.170 131.245 ;
        RECT 55.370 131.125 55.790 131.505 ;
        RECT 55.970 131.035 56.600 131.285 ;
        RECT 57.070 131.125 57.400 131.505 ;
        RECT 55.970 130.955 56.140 131.035 ;
        RECT 57.570 130.955 57.740 131.245 ;
        RECT 57.920 131.125 58.300 131.505 ;
        RECT 58.540 131.120 59.370 131.290 ;
        RECT 54.930 130.785 56.140 130.955 ;
        RECT 52.880 129.865 53.680 130.195 ;
        RECT 52.530 129.465 52.785 129.665 ;
        RECT 52.445 129.295 52.785 129.465 ;
        RECT 52.530 129.135 52.785 129.295 ;
        RECT 52.965 128.955 53.250 129.415 ;
        RECT 53.430 129.215 53.680 129.865 ;
        RECT 53.880 130.615 54.200 130.635 ;
        RECT 53.880 130.445 55.800 130.615 ;
        RECT 53.880 129.550 54.070 130.445 ;
        RECT 55.970 130.275 56.140 130.785 ;
        RECT 56.310 130.525 56.830 130.835 ;
        RECT 54.240 130.105 56.140 130.275 ;
        RECT 54.240 130.045 54.570 130.105 ;
        RECT 54.720 129.875 55.050 129.935 ;
        RECT 54.390 129.605 55.050 129.875 ;
        RECT 53.880 129.220 54.200 129.550 ;
        RECT 54.380 128.955 55.040 129.435 ;
        RECT 55.240 129.345 55.410 130.105 ;
        RECT 56.310 129.935 56.490 130.345 ;
        RECT 55.580 129.765 55.910 129.885 ;
        RECT 56.660 129.765 56.830 130.525 ;
        RECT 55.580 129.595 56.830 129.765 ;
        RECT 57.000 130.705 58.370 130.955 ;
        RECT 57.000 129.935 57.190 130.705 ;
        RECT 58.120 130.445 58.370 130.705 ;
        RECT 57.360 130.275 57.610 130.435 ;
        RECT 58.540 130.275 58.710 131.120 ;
        RECT 59.605 130.835 59.775 131.335 ;
        RECT 59.945 131.005 60.275 131.505 ;
        RECT 58.880 130.445 59.380 130.825 ;
        RECT 59.605 130.665 60.300 130.835 ;
        RECT 57.360 130.105 58.710 130.275 ;
        RECT 58.290 130.065 58.710 130.105 ;
        RECT 57.000 129.595 57.420 129.935 ;
        RECT 57.710 129.605 58.120 129.935 ;
        RECT 55.240 129.175 56.090 129.345 ;
        RECT 56.650 128.955 56.970 129.415 ;
        RECT 57.170 129.165 57.420 129.595 ;
        RECT 57.710 128.955 58.120 129.395 ;
        RECT 58.290 129.335 58.460 130.065 ;
        RECT 58.630 129.515 58.980 129.885 ;
        RECT 59.160 129.575 59.380 130.445 ;
        RECT 59.550 129.875 59.960 130.495 ;
        RECT 60.130 129.695 60.300 130.665 ;
        RECT 59.605 129.505 60.300 129.695 ;
        RECT 58.290 129.135 59.305 129.335 ;
        RECT 59.605 129.175 59.775 129.505 ;
        RECT 59.945 128.955 60.275 129.335 ;
        RECT 60.490 129.215 60.715 131.335 ;
        RECT 60.885 131.005 61.215 131.505 ;
        RECT 61.385 130.835 61.555 131.335 ;
        RECT 60.890 130.665 61.555 130.835 ;
        RECT 60.890 129.675 61.120 130.665 ;
        RECT 61.290 129.845 61.640 130.495 ;
        RECT 62.275 130.415 65.785 131.505 ;
        RECT 65.955 130.745 66.470 131.155 ;
        RECT 66.705 130.745 66.875 131.505 ;
        RECT 67.045 131.165 69.075 131.335 ;
        RECT 62.275 129.895 63.965 130.415 ;
        RECT 64.135 129.725 65.785 130.245 ;
        RECT 65.955 129.935 66.295 130.745 ;
        RECT 67.045 130.500 67.215 131.165 ;
        RECT 67.610 130.825 68.735 130.995 ;
        RECT 66.465 130.310 67.215 130.500 ;
        RECT 67.385 130.485 68.395 130.655 ;
        RECT 65.955 129.765 67.185 129.935 ;
        RECT 60.890 129.505 61.555 129.675 ;
        RECT 60.885 128.955 61.215 129.335 ;
        RECT 61.385 129.215 61.555 129.505 ;
        RECT 62.275 128.955 65.785 129.725 ;
        RECT 66.230 129.160 66.475 129.765 ;
        RECT 66.695 128.955 67.205 129.490 ;
        RECT 67.385 129.125 67.575 130.485 ;
        RECT 67.745 129.805 68.020 130.285 ;
        RECT 67.745 129.635 68.025 129.805 ;
        RECT 68.225 129.685 68.395 130.485 ;
        RECT 68.565 129.695 68.735 130.825 ;
        RECT 68.905 130.195 69.075 131.165 ;
        RECT 69.245 130.365 69.415 131.505 ;
        RECT 69.585 130.365 69.920 131.335 ;
        RECT 70.645 130.575 70.815 131.335 ;
        RECT 70.995 130.745 71.325 131.505 ;
        RECT 70.645 130.405 71.310 130.575 ;
        RECT 71.495 130.430 71.765 131.335 ;
        RECT 68.905 129.865 69.100 130.195 ;
        RECT 69.325 129.865 69.580 130.195 ;
        RECT 69.325 129.695 69.495 129.865 ;
        RECT 69.750 129.695 69.920 130.365 ;
        RECT 71.140 130.260 71.310 130.405 ;
        RECT 70.575 129.855 70.905 130.225 ;
        RECT 71.140 129.930 71.425 130.260 ;
        RECT 67.745 129.125 68.020 129.635 ;
        RECT 68.565 129.525 69.495 129.695 ;
        RECT 68.565 129.490 68.740 129.525 ;
        RECT 68.210 129.125 68.740 129.490 ;
        RECT 69.165 128.955 69.495 129.355 ;
        RECT 69.665 129.125 69.920 129.695 ;
        RECT 71.140 129.675 71.310 129.930 ;
        RECT 70.645 129.505 71.310 129.675 ;
        RECT 71.595 129.630 71.765 130.430 ;
        RECT 71.935 130.415 74.525 131.505 ;
        RECT 71.935 129.895 73.145 130.415 ;
        RECT 74.695 130.365 74.965 131.335 ;
        RECT 75.175 130.705 75.455 131.505 ;
        RECT 75.625 130.995 77.280 131.285 ;
        RECT 75.690 130.655 77.280 130.825 ;
        RECT 75.690 130.535 75.860 130.655 ;
        RECT 75.135 130.365 75.860 130.535 ;
        RECT 73.315 129.725 74.525 130.245 ;
        RECT 70.645 129.125 70.815 129.505 ;
        RECT 70.995 128.955 71.325 129.335 ;
        RECT 71.505 129.125 71.765 129.630 ;
        RECT 71.935 128.955 74.525 129.725 ;
        RECT 74.695 129.630 74.865 130.365 ;
        RECT 75.135 130.195 75.305 130.365 ;
        RECT 75.035 129.865 75.305 130.195 ;
        RECT 75.475 129.865 75.880 130.195 ;
        RECT 76.050 129.865 76.760 130.485 ;
        RECT 76.960 130.365 77.280 130.655 ;
        RECT 77.455 130.340 77.745 131.505 ;
        RECT 77.915 130.415 79.585 131.505 ;
        RECT 75.135 129.695 75.305 129.865 ;
        RECT 74.695 129.285 74.965 129.630 ;
        RECT 75.135 129.525 76.745 129.695 ;
        RECT 76.930 129.625 77.280 130.195 ;
        RECT 77.915 129.895 78.665 130.415 ;
        RECT 79.755 130.365 80.095 131.335 ;
        RECT 80.265 130.365 80.435 131.505 ;
        RECT 80.705 130.705 80.955 131.505 ;
        RECT 81.600 130.535 81.930 131.335 ;
        RECT 82.230 130.705 82.560 131.505 ;
        RECT 82.730 130.535 83.060 131.335 ;
        RECT 80.625 130.365 83.060 130.535 ;
        RECT 83.435 130.415 85.105 131.505 ;
        RECT 85.275 130.745 85.790 131.155 ;
        RECT 86.025 130.745 86.195 131.505 ;
        RECT 86.365 131.165 88.395 131.335 ;
        RECT 78.835 129.725 79.585 130.245 ;
        RECT 75.155 128.955 75.535 129.355 ;
        RECT 75.705 129.175 75.875 129.525 ;
        RECT 76.045 128.955 76.375 129.355 ;
        RECT 76.575 129.175 76.745 129.525 ;
        RECT 76.945 128.955 77.275 129.455 ;
        RECT 77.455 128.955 77.745 129.680 ;
        RECT 77.915 128.955 79.585 129.725 ;
        RECT 79.755 129.805 79.930 130.365 ;
        RECT 80.625 130.115 80.795 130.365 ;
        RECT 80.100 129.945 80.795 130.115 ;
        RECT 80.970 129.945 81.390 130.145 ;
        RECT 81.560 129.945 81.890 130.145 ;
        RECT 82.060 129.945 82.390 130.145 ;
        RECT 79.755 129.755 79.985 129.805 ;
        RECT 79.755 129.125 80.095 129.755 ;
        RECT 80.265 128.955 80.515 129.755 ;
        RECT 80.705 129.605 81.930 129.775 ;
        RECT 80.705 129.125 81.035 129.605 ;
        RECT 81.205 128.955 81.430 129.415 ;
        RECT 81.600 129.125 81.930 129.605 ;
        RECT 82.560 129.735 82.730 130.365 ;
        RECT 82.915 129.945 83.265 130.195 ;
        RECT 83.435 129.895 84.185 130.415 ;
        RECT 82.560 129.125 83.060 129.735 ;
        RECT 84.355 129.725 85.105 130.245 ;
        RECT 85.275 129.935 85.615 130.745 ;
        RECT 86.365 130.500 86.535 131.165 ;
        RECT 86.930 130.825 88.055 130.995 ;
        RECT 85.785 130.310 86.535 130.500 ;
        RECT 86.705 130.485 87.715 130.655 ;
        RECT 85.275 129.765 86.505 129.935 ;
        RECT 83.435 128.955 85.105 129.725 ;
        RECT 85.550 129.160 85.795 129.765 ;
        RECT 86.015 128.955 86.525 129.490 ;
        RECT 86.705 129.125 86.895 130.485 ;
        RECT 87.065 130.145 87.340 130.285 ;
        RECT 87.065 129.975 87.345 130.145 ;
        RECT 87.065 129.125 87.340 129.975 ;
        RECT 87.545 129.685 87.715 130.485 ;
        RECT 87.885 129.695 88.055 130.825 ;
        RECT 88.225 130.195 88.395 131.165 ;
        RECT 88.565 130.365 88.735 131.505 ;
        RECT 88.905 130.365 89.240 131.335 ;
        RECT 88.225 129.865 88.420 130.195 ;
        RECT 88.645 129.865 88.900 130.195 ;
        RECT 88.645 129.695 88.815 129.865 ;
        RECT 89.070 129.695 89.240 130.365 ;
        RECT 87.885 129.525 88.815 129.695 ;
        RECT 87.885 129.490 88.060 129.525 ;
        RECT 87.530 129.125 88.060 129.490 ;
        RECT 88.485 128.955 88.815 129.355 ;
        RECT 88.985 129.125 89.240 129.695 ;
        RECT 89.415 130.430 89.685 131.335 ;
        RECT 89.855 130.745 90.185 131.505 ;
        RECT 90.365 130.575 90.535 131.335 ;
        RECT 89.415 129.630 89.585 130.430 ;
        RECT 89.870 130.405 90.535 130.575 ;
        RECT 90.795 130.415 93.385 131.505 ;
        RECT 93.930 131.165 94.185 131.195 ;
        RECT 93.845 130.995 94.185 131.165 ;
        RECT 93.930 130.525 94.185 130.995 ;
        RECT 94.365 130.705 94.650 131.505 ;
        RECT 94.830 130.785 95.160 131.295 ;
        RECT 89.870 130.260 90.040 130.405 ;
        RECT 89.755 129.930 90.040 130.260 ;
        RECT 89.870 129.675 90.040 129.930 ;
        RECT 90.275 129.855 90.605 130.225 ;
        RECT 90.795 129.895 92.005 130.415 ;
        RECT 92.175 129.725 93.385 130.245 ;
        RECT 89.415 129.125 89.675 129.630 ;
        RECT 89.870 129.505 90.535 129.675 ;
        RECT 89.855 128.955 90.185 129.335 ;
        RECT 90.365 129.125 90.535 129.505 ;
        RECT 90.795 128.955 93.385 129.725 ;
        RECT 93.930 129.665 94.110 130.525 ;
        RECT 94.830 130.195 95.080 130.785 ;
        RECT 95.430 130.635 95.600 131.245 ;
        RECT 95.770 130.815 96.100 131.505 ;
        RECT 96.330 130.955 96.570 131.245 ;
        RECT 96.770 131.125 97.190 131.505 ;
        RECT 97.370 131.035 98.000 131.285 ;
        RECT 98.470 131.125 98.800 131.505 ;
        RECT 97.370 130.955 97.540 131.035 ;
        RECT 98.970 130.955 99.140 131.245 ;
        RECT 99.320 131.125 99.700 131.505 ;
        RECT 99.940 131.120 100.770 131.290 ;
        RECT 96.330 130.785 97.540 130.955 ;
        RECT 94.280 129.865 95.080 130.195 ;
        RECT 93.930 129.135 94.185 129.665 ;
        RECT 94.365 128.955 94.650 129.415 ;
        RECT 94.830 129.215 95.080 129.865 ;
        RECT 95.280 130.615 95.600 130.635 ;
        RECT 95.280 130.445 97.200 130.615 ;
        RECT 95.280 129.550 95.470 130.445 ;
        RECT 97.370 130.275 97.540 130.785 ;
        RECT 97.710 130.525 98.230 130.835 ;
        RECT 95.640 130.105 97.540 130.275 ;
        RECT 95.640 130.045 95.970 130.105 ;
        RECT 96.120 129.875 96.450 129.935 ;
        RECT 95.790 129.605 96.450 129.875 ;
        RECT 95.280 129.220 95.600 129.550 ;
        RECT 95.780 128.955 96.440 129.435 ;
        RECT 96.640 129.345 96.810 130.105 ;
        RECT 97.710 129.935 97.890 130.345 ;
        RECT 96.980 129.765 97.310 129.885 ;
        RECT 98.060 129.765 98.230 130.525 ;
        RECT 96.980 129.595 98.230 129.765 ;
        RECT 98.400 130.705 99.770 130.955 ;
        RECT 98.400 129.935 98.590 130.705 ;
        RECT 99.520 130.445 99.770 130.705 ;
        RECT 98.760 130.275 99.010 130.435 ;
        RECT 99.940 130.275 100.110 131.120 ;
        RECT 101.005 130.835 101.175 131.335 ;
        RECT 101.345 131.005 101.675 131.505 ;
        RECT 100.280 130.445 100.780 130.825 ;
        RECT 101.005 130.665 101.700 130.835 ;
        RECT 98.760 130.105 100.110 130.275 ;
        RECT 99.690 130.065 100.110 130.105 ;
        RECT 98.400 129.595 98.820 129.935 ;
        RECT 99.110 129.605 99.520 129.935 ;
        RECT 96.640 129.175 97.490 129.345 ;
        RECT 98.050 128.955 98.370 129.415 ;
        RECT 98.570 129.165 98.820 129.595 ;
        RECT 99.110 128.955 99.520 129.395 ;
        RECT 99.690 129.335 99.860 130.065 ;
        RECT 100.030 129.515 100.380 129.885 ;
        RECT 100.560 129.575 100.780 130.445 ;
        RECT 100.950 129.875 101.360 130.495 ;
        RECT 101.530 129.695 101.700 130.665 ;
        RECT 101.005 129.505 101.700 129.695 ;
        RECT 99.690 129.135 100.705 129.335 ;
        RECT 101.005 129.175 101.175 129.505 ;
        RECT 101.345 128.955 101.675 129.335 ;
        RECT 101.890 129.215 102.115 131.335 ;
        RECT 102.285 131.005 102.615 131.505 ;
        RECT 102.785 130.835 102.955 131.335 ;
        RECT 102.290 130.665 102.955 130.835 ;
        RECT 102.290 129.675 102.520 130.665 ;
        RECT 102.690 129.845 103.040 130.495 ;
        RECT 103.215 130.340 103.505 131.505 ;
        RECT 104.135 130.415 105.805 131.505 ;
        RECT 106.350 130.525 106.605 131.195 ;
        RECT 106.785 130.705 107.070 131.505 ;
        RECT 107.250 130.785 107.580 131.295 ;
        RECT 104.135 129.895 104.885 130.415 ;
        RECT 105.055 129.725 105.805 130.245 ;
        RECT 106.350 130.145 106.530 130.525 ;
        RECT 107.250 130.195 107.500 130.785 ;
        RECT 107.850 130.635 108.020 131.245 ;
        RECT 108.190 130.815 108.520 131.505 ;
        RECT 108.750 130.955 108.990 131.245 ;
        RECT 109.190 131.125 109.610 131.505 ;
        RECT 109.790 131.035 110.420 131.285 ;
        RECT 110.890 131.125 111.220 131.505 ;
        RECT 109.790 130.955 109.960 131.035 ;
        RECT 111.390 130.955 111.560 131.245 ;
        RECT 111.740 131.125 112.120 131.505 ;
        RECT 112.360 131.120 113.190 131.290 ;
        RECT 108.750 130.785 109.960 130.955 ;
        RECT 106.265 129.975 106.530 130.145 ;
        RECT 102.290 129.505 102.955 129.675 ;
        RECT 102.285 128.955 102.615 129.335 ;
        RECT 102.785 129.215 102.955 129.505 ;
        RECT 103.215 128.955 103.505 129.680 ;
        RECT 104.135 128.955 105.805 129.725 ;
        RECT 106.350 129.665 106.530 129.975 ;
        RECT 106.700 129.865 107.500 130.195 ;
        RECT 106.350 129.135 106.605 129.665 ;
        RECT 106.785 128.955 107.070 129.415 ;
        RECT 107.250 129.215 107.500 129.865 ;
        RECT 107.700 130.615 108.020 130.635 ;
        RECT 107.700 130.445 109.620 130.615 ;
        RECT 107.700 129.550 107.890 130.445 ;
        RECT 109.790 130.275 109.960 130.785 ;
        RECT 110.130 130.525 110.650 130.835 ;
        RECT 108.060 130.105 109.960 130.275 ;
        RECT 108.060 130.045 108.390 130.105 ;
        RECT 108.540 129.875 108.870 129.935 ;
        RECT 108.210 129.605 108.870 129.875 ;
        RECT 107.700 129.220 108.020 129.550 ;
        RECT 108.200 128.955 108.860 129.435 ;
        RECT 109.060 129.345 109.230 130.105 ;
        RECT 110.130 129.935 110.310 130.345 ;
        RECT 109.400 129.765 109.730 129.885 ;
        RECT 110.480 129.765 110.650 130.525 ;
        RECT 109.400 129.595 110.650 129.765 ;
        RECT 110.820 130.705 112.190 130.955 ;
        RECT 110.820 129.935 111.010 130.705 ;
        RECT 111.940 130.445 112.190 130.705 ;
        RECT 111.180 130.275 111.430 130.435 ;
        RECT 112.360 130.275 112.530 131.120 ;
        RECT 113.425 130.835 113.595 131.335 ;
        RECT 113.765 131.005 114.095 131.505 ;
        RECT 112.700 130.445 113.200 130.825 ;
        RECT 113.425 130.665 114.120 130.835 ;
        RECT 111.180 130.105 112.530 130.275 ;
        RECT 112.110 130.065 112.530 130.105 ;
        RECT 110.820 129.595 111.240 129.935 ;
        RECT 111.530 129.605 111.940 129.935 ;
        RECT 109.060 129.175 109.910 129.345 ;
        RECT 110.470 128.955 110.790 129.415 ;
        RECT 110.990 129.165 111.240 129.595 ;
        RECT 111.530 128.955 111.940 129.395 ;
        RECT 112.110 129.335 112.280 130.065 ;
        RECT 112.450 129.515 112.800 129.885 ;
        RECT 112.980 129.575 113.200 130.445 ;
        RECT 113.370 129.875 113.780 130.495 ;
        RECT 113.950 129.695 114.120 130.665 ;
        RECT 113.425 129.505 114.120 129.695 ;
        RECT 112.110 129.135 113.125 129.335 ;
        RECT 113.425 129.175 113.595 129.505 ;
        RECT 113.765 128.955 114.095 129.335 ;
        RECT 114.310 129.215 114.535 131.335 ;
        RECT 114.705 131.005 115.035 131.505 ;
        RECT 115.205 130.835 115.375 131.335 ;
        RECT 114.710 130.665 115.375 130.835 ;
        RECT 114.710 129.675 114.940 130.665 ;
        RECT 115.110 129.845 115.460 130.495 ;
        RECT 115.635 130.415 116.845 131.505 ;
        RECT 117.020 131.070 122.365 131.505 ;
        RECT 122.540 131.070 127.885 131.505 ;
        RECT 115.635 129.875 116.155 130.415 ;
        RECT 116.325 129.705 116.845 130.245 ;
        RECT 118.610 129.820 118.960 131.070 ;
        RECT 114.710 129.505 115.375 129.675 ;
        RECT 114.705 128.955 115.035 129.335 ;
        RECT 115.205 129.215 115.375 129.505 ;
        RECT 115.635 128.955 116.845 129.705 ;
        RECT 120.440 129.500 120.780 130.330 ;
        RECT 124.130 129.820 124.480 131.070 ;
        RECT 128.055 130.415 129.265 131.505 ;
        RECT 125.960 129.500 126.300 130.330 ;
        RECT 128.055 129.875 128.575 130.415 ;
        RECT 128.745 129.705 129.265 130.245 ;
        RECT 117.020 128.955 122.365 129.500 ;
        RECT 122.540 128.955 127.885 129.500 ;
        RECT 128.055 128.955 129.265 129.705 ;
        RECT 9.290 128.785 129.350 128.955 ;
        RECT 9.375 128.035 10.585 128.785 ;
        RECT 9.375 127.495 9.895 128.035 ;
        RECT 11.735 127.965 11.945 128.785 ;
        RECT 12.115 127.985 12.445 128.615 ;
        RECT 10.065 127.325 10.585 127.865 ;
        RECT 12.115 127.385 12.365 127.985 ;
        RECT 12.615 127.965 12.845 128.785 ;
        RECT 13.055 128.060 13.345 128.785 ;
        RECT 13.890 128.445 14.145 128.605 ;
        RECT 13.805 128.275 14.145 128.445 ;
        RECT 14.325 128.325 14.610 128.785 ;
        RECT 13.890 128.075 14.145 128.275 ;
        RECT 12.535 127.545 12.865 127.795 ;
        RECT 9.375 126.235 10.585 127.325 ;
        RECT 11.735 126.235 11.945 127.375 ;
        RECT 12.115 126.405 12.445 127.385 ;
        RECT 12.615 126.235 12.845 127.375 ;
        RECT 13.055 126.235 13.345 127.400 ;
        RECT 13.890 127.215 14.070 128.075 ;
        RECT 14.790 127.875 15.040 128.525 ;
        RECT 14.240 127.545 15.040 127.875 ;
        RECT 13.890 126.545 14.145 127.215 ;
        RECT 14.325 126.235 14.610 127.035 ;
        RECT 14.790 126.955 15.040 127.545 ;
        RECT 15.240 128.190 15.560 128.520 ;
        RECT 15.740 128.305 16.400 128.785 ;
        RECT 16.600 128.395 17.450 128.565 ;
        RECT 15.240 127.295 15.430 128.190 ;
        RECT 15.750 127.865 16.410 128.135 ;
        RECT 16.080 127.805 16.410 127.865 ;
        RECT 15.600 127.635 15.930 127.695 ;
        RECT 16.600 127.635 16.770 128.395 ;
        RECT 18.010 128.325 18.330 128.785 ;
        RECT 18.530 128.145 18.780 128.575 ;
        RECT 19.070 128.345 19.480 128.785 ;
        RECT 19.650 128.405 20.665 128.605 ;
        RECT 16.940 127.975 18.190 128.145 ;
        RECT 16.940 127.855 17.270 127.975 ;
        RECT 15.600 127.465 17.500 127.635 ;
        RECT 15.240 127.125 17.160 127.295 ;
        RECT 15.240 127.105 15.560 127.125 ;
        RECT 14.790 126.445 15.120 126.955 ;
        RECT 15.390 126.495 15.560 127.105 ;
        RECT 17.330 126.955 17.500 127.465 ;
        RECT 17.670 127.395 17.850 127.805 ;
        RECT 18.020 127.215 18.190 127.975 ;
        RECT 15.730 126.235 16.060 126.925 ;
        RECT 16.290 126.785 17.500 126.955 ;
        RECT 17.670 126.905 18.190 127.215 ;
        RECT 18.360 127.805 18.780 128.145 ;
        RECT 19.070 127.805 19.480 128.135 ;
        RECT 18.360 127.035 18.550 127.805 ;
        RECT 19.650 127.675 19.820 128.405 ;
        RECT 20.965 128.235 21.135 128.565 ;
        RECT 21.305 128.405 21.635 128.785 ;
        RECT 19.990 127.855 20.340 128.225 ;
        RECT 19.650 127.635 20.070 127.675 ;
        RECT 18.720 127.465 20.070 127.635 ;
        RECT 18.720 127.305 18.970 127.465 ;
        RECT 19.480 127.035 19.730 127.295 ;
        RECT 18.360 126.785 19.730 127.035 ;
        RECT 16.290 126.495 16.530 126.785 ;
        RECT 17.330 126.705 17.500 126.785 ;
        RECT 16.730 126.235 17.150 126.615 ;
        RECT 17.330 126.455 17.960 126.705 ;
        RECT 18.430 126.235 18.760 126.615 ;
        RECT 18.930 126.495 19.100 126.785 ;
        RECT 19.900 126.620 20.070 127.465 ;
        RECT 20.520 127.295 20.740 128.165 ;
        RECT 20.965 128.045 21.660 128.235 ;
        RECT 20.240 126.915 20.740 127.295 ;
        RECT 20.910 127.245 21.320 127.865 ;
        RECT 21.490 127.075 21.660 128.045 ;
        RECT 20.965 126.905 21.660 127.075 ;
        RECT 19.280 126.235 19.660 126.615 ;
        RECT 19.900 126.450 20.730 126.620 ;
        RECT 20.965 126.405 21.135 126.905 ;
        RECT 21.305 126.235 21.635 126.735 ;
        RECT 21.850 126.405 22.075 128.525 ;
        RECT 22.245 128.405 22.575 128.785 ;
        RECT 22.745 128.235 22.915 128.525 ;
        RECT 22.250 128.065 22.915 128.235 ;
        RECT 22.250 127.075 22.480 128.065 ;
        RECT 23.450 127.975 23.695 128.580 ;
        RECT 23.915 128.250 24.425 128.785 ;
        RECT 22.650 127.245 23.000 127.895 ;
        RECT 23.175 127.805 24.405 127.975 ;
        RECT 22.250 126.905 22.915 127.075 ;
        RECT 22.245 126.235 22.575 126.735 ;
        RECT 22.745 126.405 22.915 126.905 ;
        RECT 23.175 126.995 23.515 127.805 ;
        RECT 23.685 127.240 24.435 127.430 ;
        RECT 23.175 126.585 23.690 126.995 ;
        RECT 23.925 126.235 24.095 126.995 ;
        RECT 24.265 126.575 24.435 127.240 ;
        RECT 24.605 127.255 24.795 128.615 ;
        RECT 24.965 128.105 25.240 128.615 ;
        RECT 25.430 128.250 25.960 128.615 ;
        RECT 26.385 128.385 26.715 128.785 ;
        RECT 25.785 128.215 25.960 128.250 ;
        RECT 24.965 127.935 25.245 128.105 ;
        RECT 24.965 127.455 25.240 127.935 ;
        RECT 25.445 127.255 25.615 128.055 ;
        RECT 24.605 127.085 25.615 127.255 ;
        RECT 25.785 128.045 26.715 128.215 ;
        RECT 26.885 128.045 27.140 128.615 ;
        RECT 27.405 128.305 27.705 128.785 ;
        RECT 27.875 128.135 28.135 128.590 ;
        RECT 28.305 128.305 28.565 128.785 ;
        RECT 28.745 128.135 29.005 128.590 ;
        RECT 29.175 128.305 29.425 128.785 ;
        RECT 29.605 128.135 29.865 128.590 ;
        RECT 30.035 128.305 30.285 128.785 ;
        RECT 30.465 128.135 30.725 128.590 ;
        RECT 30.895 128.305 31.140 128.785 ;
        RECT 31.310 128.135 31.585 128.590 ;
        RECT 31.755 128.305 32.000 128.785 ;
        RECT 32.170 128.135 32.430 128.590 ;
        RECT 32.600 128.305 32.860 128.785 ;
        RECT 33.030 128.135 33.290 128.590 ;
        RECT 33.460 128.305 33.720 128.785 ;
        RECT 33.890 128.135 34.150 128.590 ;
        RECT 34.320 128.225 34.580 128.785 ;
        RECT 25.785 126.915 25.955 128.045 ;
        RECT 26.545 127.875 26.715 128.045 ;
        RECT 24.830 126.745 25.955 126.915 ;
        RECT 26.125 127.545 26.320 127.875 ;
        RECT 26.545 127.545 26.800 127.875 ;
        RECT 26.125 126.575 26.295 127.545 ;
        RECT 26.970 127.375 27.140 128.045 ;
        RECT 24.265 126.405 26.295 126.575 ;
        RECT 26.465 126.235 26.635 127.375 ;
        RECT 26.805 126.405 27.140 127.375 ;
        RECT 27.405 127.965 34.150 128.135 ;
        RECT 27.405 127.375 28.570 127.965 ;
        RECT 34.750 127.795 35.000 128.605 ;
        RECT 35.180 128.260 35.440 128.785 ;
        RECT 35.610 127.795 35.860 128.605 ;
        RECT 36.040 128.275 36.345 128.785 ;
        RECT 28.740 127.545 35.860 127.795 ;
        RECT 36.030 127.545 36.345 128.105 ;
        RECT 36.975 128.015 38.645 128.785 ;
        RECT 38.815 128.060 39.105 128.785 ;
        RECT 40.200 128.240 45.545 128.785 ;
        RECT 45.715 128.325 46.275 128.615 ;
        RECT 46.445 128.325 46.695 128.785 ;
        RECT 27.405 127.150 34.150 127.375 ;
        RECT 27.405 126.235 27.675 126.980 ;
        RECT 27.845 126.410 28.135 127.150 ;
        RECT 28.745 127.135 34.150 127.150 ;
        RECT 28.305 126.240 28.560 126.965 ;
        RECT 28.745 126.410 29.005 127.135 ;
        RECT 29.175 126.240 29.420 126.965 ;
        RECT 29.605 126.410 29.865 127.135 ;
        RECT 30.035 126.240 30.280 126.965 ;
        RECT 30.465 126.410 30.725 127.135 ;
        RECT 30.895 126.240 31.140 126.965 ;
        RECT 31.310 126.410 31.570 127.135 ;
        RECT 31.740 126.240 32.000 126.965 ;
        RECT 32.170 126.410 32.430 127.135 ;
        RECT 32.600 126.240 32.860 126.965 ;
        RECT 33.030 126.410 33.290 127.135 ;
        RECT 33.460 126.240 33.720 126.965 ;
        RECT 33.890 126.410 34.150 127.135 ;
        RECT 34.320 126.240 34.580 127.035 ;
        RECT 34.750 126.410 35.000 127.545 ;
        RECT 28.305 126.235 34.580 126.240 ;
        RECT 35.180 126.235 35.440 127.045 ;
        RECT 35.615 126.405 35.860 127.545 ;
        RECT 36.975 127.325 37.725 127.845 ;
        RECT 37.895 127.495 38.645 128.015 ;
        RECT 36.040 126.235 36.335 127.045 ;
        RECT 36.975 126.235 38.645 127.325 ;
        RECT 38.815 126.235 39.105 127.400 ;
        RECT 41.790 126.670 42.140 127.920 ;
        RECT 43.620 127.410 43.960 128.240 ;
        RECT 45.715 126.955 45.965 128.325 ;
        RECT 47.315 128.155 47.645 128.515 ;
        RECT 46.255 127.965 47.645 128.155 ;
        RECT 48.015 127.985 48.355 128.615 ;
        RECT 48.525 127.985 48.775 128.785 ;
        RECT 48.965 128.135 49.295 128.615 ;
        RECT 49.465 128.325 49.690 128.785 ;
        RECT 49.860 128.135 50.190 128.615 ;
        RECT 46.255 127.875 46.425 127.965 ;
        RECT 46.135 127.545 46.425 127.875 ;
        RECT 46.595 127.545 46.935 127.795 ;
        RECT 47.155 127.545 47.830 127.795 ;
        RECT 46.255 127.295 46.425 127.545 ;
        RECT 46.255 127.125 47.195 127.295 ;
        RECT 47.565 127.185 47.830 127.545 ;
        RECT 48.015 127.375 48.190 127.985 ;
        RECT 48.965 127.965 50.190 128.135 ;
        RECT 50.820 128.005 51.320 128.615 ;
        RECT 52.155 128.015 53.825 128.785 ;
        RECT 48.360 127.625 49.055 127.795 ;
        RECT 48.885 127.375 49.055 127.625 ;
        RECT 49.230 127.595 49.650 127.795 ;
        RECT 49.820 127.595 50.150 127.795 ;
        RECT 50.320 127.595 50.650 127.795 ;
        RECT 50.820 127.375 50.990 128.005 ;
        RECT 51.175 127.545 51.525 127.795 ;
        RECT 40.200 126.235 45.545 126.670 ;
        RECT 45.715 126.405 46.175 126.955 ;
        RECT 46.365 126.235 46.695 126.955 ;
        RECT 46.895 126.575 47.195 127.125 ;
        RECT 47.365 126.235 47.645 126.905 ;
        RECT 48.015 126.405 48.355 127.375 ;
        RECT 48.525 126.235 48.695 127.375 ;
        RECT 48.885 127.205 51.320 127.375 ;
        RECT 48.965 126.235 49.215 127.035 ;
        RECT 49.860 126.405 50.190 127.205 ;
        RECT 50.490 126.235 50.820 127.035 ;
        RECT 50.990 126.405 51.320 127.205 ;
        RECT 52.155 127.325 52.905 127.845 ;
        RECT 53.075 127.495 53.825 128.015 ;
        RECT 54.270 127.975 54.515 128.580 ;
        RECT 54.735 128.250 55.245 128.785 ;
        RECT 53.995 127.805 55.225 127.975 ;
        RECT 52.155 126.235 53.825 127.325 ;
        RECT 53.995 126.995 54.335 127.805 ;
        RECT 54.505 127.240 55.255 127.430 ;
        RECT 53.995 126.585 54.510 126.995 ;
        RECT 54.745 126.235 54.915 126.995 ;
        RECT 55.085 126.575 55.255 127.240 ;
        RECT 55.425 127.255 55.615 128.615 ;
        RECT 55.785 128.105 56.060 128.615 ;
        RECT 56.250 128.250 56.780 128.615 ;
        RECT 57.205 128.385 57.535 128.785 ;
        RECT 56.605 128.215 56.780 128.250 ;
        RECT 55.785 127.935 56.065 128.105 ;
        RECT 55.785 127.455 56.060 127.935 ;
        RECT 56.265 127.255 56.435 128.055 ;
        RECT 55.425 127.085 56.435 127.255 ;
        RECT 56.605 128.045 57.535 128.215 ;
        RECT 57.705 128.045 57.960 128.615 ;
        RECT 56.605 126.915 56.775 128.045 ;
        RECT 57.365 127.875 57.535 128.045 ;
        RECT 55.650 126.745 56.775 126.915 ;
        RECT 56.945 127.545 57.140 127.875 ;
        RECT 57.365 127.545 57.620 127.875 ;
        RECT 56.945 126.575 57.115 127.545 ;
        RECT 57.790 127.375 57.960 128.045 ;
        RECT 58.135 128.035 59.345 128.785 ;
        RECT 55.085 126.405 57.115 126.575 ;
        RECT 57.285 126.235 57.455 127.375 ;
        RECT 57.625 126.405 57.960 127.375 ;
        RECT 58.135 127.325 58.655 127.865 ;
        RECT 58.825 127.495 59.345 128.035 ;
        RECT 59.515 128.015 63.025 128.785 ;
        RECT 59.515 127.325 61.205 127.845 ;
        RECT 61.375 127.495 63.025 128.015 ;
        RECT 63.235 127.965 63.465 128.785 ;
        RECT 63.635 127.985 63.965 128.615 ;
        RECT 63.215 127.545 63.545 127.795 ;
        RECT 63.715 127.385 63.965 127.985 ;
        RECT 64.135 127.965 64.345 128.785 ;
        RECT 64.575 128.060 64.865 128.785 ;
        RECT 65.870 128.445 66.125 128.605 ;
        RECT 65.785 128.275 66.125 128.445 ;
        RECT 66.305 128.325 66.590 128.785 ;
        RECT 65.870 128.075 66.125 128.275 ;
        RECT 58.135 126.235 59.345 127.325 ;
        RECT 59.515 126.235 63.025 127.325 ;
        RECT 63.235 126.235 63.465 127.375 ;
        RECT 63.635 126.405 63.965 127.385 ;
        RECT 64.135 126.235 64.345 127.375 ;
        RECT 64.575 126.235 64.865 127.400 ;
        RECT 65.870 127.215 66.050 128.075 ;
        RECT 66.770 127.875 67.020 128.525 ;
        RECT 66.220 127.545 67.020 127.875 ;
        RECT 65.870 126.545 66.125 127.215 ;
        RECT 66.305 126.235 66.590 127.035 ;
        RECT 66.770 126.955 67.020 127.545 ;
        RECT 67.220 128.190 67.540 128.520 ;
        RECT 67.720 128.305 68.380 128.785 ;
        RECT 68.580 128.395 69.430 128.565 ;
        RECT 67.220 127.295 67.410 128.190 ;
        RECT 67.730 127.865 68.390 128.135 ;
        RECT 68.060 127.805 68.390 127.865 ;
        RECT 67.580 127.635 67.910 127.695 ;
        RECT 68.580 127.635 68.750 128.395 ;
        RECT 69.990 128.325 70.310 128.785 ;
        RECT 70.510 128.145 70.760 128.575 ;
        RECT 71.050 128.345 71.460 128.785 ;
        RECT 71.630 128.405 72.645 128.605 ;
        RECT 68.920 127.975 70.170 128.145 ;
        RECT 68.920 127.855 69.250 127.975 ;
        RECT 67.580 127.465 69.480 127.635 ;
        RECT 67.220 127.125 69.140 127.295 ;
        RECT 67.220 127.105 67.540 127.125 ;
        RECT 66.770 126.445 67.100 126.955 ;
        RECT 67.370 126.495 67.540 127.105 ;
        RECT 69.310 126.955 69.480 127.465 ;
        RECT 69.650 127.395 69.830 127.805 ;
        RECT 70.000 127.215 70.170 127.975 ;
        RECT 67.710 126.235 68.040 126.925 ;
        RECT 68.270 126.785 69.480 126.955 ;
        RECT 69.650 126.905 70.170 127.215 ;
        RECT 70.340 127.805 70.760 128.145 ;
        RECT 71.050 127.805 71.460 128.135 ;
        RECT 70.340 127.035 70.530 127.805 ;
        RECT 71.630 127.675 71.800 128.405 ;
        RECT 72.945 128.235 73.115 128.565 ;
        RECT 73.285 128.405 73.615 128.785 ;
        RECT 71.970 127.855 72.320 128.225 ;
        RECT 71.630 127.635 72.050 127.675 ;
        RECT 70.700 127.465 72.050 127.635 ;
        RECT 70.700 127.305 70.950 127.465 ;
        RECT 71.460 127.035 71.710 127.295 ;
        RECT 70.340 126.785 71.710 127.035 ;
        RECT 68.270 126.495 68.510 126.785 ;
        RECT 69.310 126.705 69.480 126.785 ;
        RECT 68.710 126.235 69.130 126.615 ;
        RECT 69.310 126.455 69.940 126.705 ;
        RECT 70.410 126.235 70.740 126.615 ;
        RECT 70.910 126.495 71.080 126.785 ;
        RECT 71.880 126.620 72.050 127.465 ;
        RECT 72.500 127.295 72.720 128.165 ;
        RECT 72.945 128.045 73.640 128.235 ;
        RECT 72.220 126.915 72.720 127.295 ;
        RECT 72.890 127.245 73.300 127.865 ;
        RECT 73.470 127.075 73.640 128.045 ;
        RECT 72.945 126.905 73.640 127.075 ;
        RECT 71.260 126.235 71.640 126.615 ;
        RECT 71.880 126.450 72.710 126.620 ;
        RECT 72.945 126.405 73.115 126.905 ;
        RECT 73.285 126.235 73.615 126.735 ;
        RECT 73.830 126.405 74.055 128.525 ;
        RECT 74.225 128.405 74.555 128.785 ;
        RECT 74.725 128.235 74.895 128.525 ;
        RECT 74.230 128.065 74.895 128.235 ;
        RECT 74.230 127.075 74.460 128.065 ;
        RECT 75.155 128.015 77.745 128.785 ;
        RECT 74.630 127.245 74.980 127.895 ;
        RECT 75.155 127.325 76.365 127.845 ;
        RECT 76.535 127.495 77.745 128.015 ;
        RECT 77.915 128.110 78.185 128.455 ;
        RECT 78.375 128.385 78.755 128.785 ;
        RECT 78.925 128.215 79.095 128.565 ;
        RECT 79.265 128.385 79.595 128.785 ;
        RECT 79.795 128.215 79.965 128.565 ;
        RECT 80.165 128.285 80.495 128.785 ;
        RECT 81.050 128.445 81.305 128.605 ;
        RECT 80.965 128.275 81.305 128.445 ;
        RECT 81.485 128.325 81.770 128.785 ;
        RECT 77.915 127.375 78.085 128.110 ;
        RECT 78.355 128.045 79.965 128.215 ;
        RECT 78.355 127.875 78.525 128.045 ;
        RECT 78.255 127.545 78.525 127.875 ;
        RECT 78.695 127.545 79.100 127.875 ;
        RECT 78.355 127.375 78.525 127.545 ;
        RECT 74.230 126.905 74.895 127.075 ;
        RECT 74.225 126.235 74.555 126.735 ;
        RECT 74.725 126.405 74.895 126.905 ;
        RECT 75.155 126.235 77.745 127.325 ;
        RECT 77.915 126.405 78.185 127.375 ;
        RECT 78.355 127.205 79.080 127.375 ;
        RECT 79.270 127.255 79.980 127.875 ;
        RECT 80.150 127.545 80.500 128.115 ;
        RECT 81.050 128.075 81.305 128.275 ;
        RECT 78.910 127.085 79.080 127.205 ;
        RECT 80.180 127.085 80.500 127.375 ;
        RECT 78.395 126.235 78.675 127.035 ;
        RECT 78.910 126.915 80.500 127.085 ;
        RECT 81.050 127.215 81.230 128.075 ;
        RECT 81.950 127.875 82.200 128.525 ;
        RECT 81.400 127.545 82.200 127.875 ;
        RECT 78.845 126.455 80.500 126.745 ;
        RECT 81.050 126.545 81.305 127.215 ;
        RECT 81.485 126.235 81.770 127.035 ;
        RECT 81.950 126.955 82.200 127.545 ;
        RECT 82.400 128.190 82.720 128.520 ;
        RECT 82.900 128.305 83.560 128.785 ;
        RECT 83.760 128.395 84.610 128.565 ;
        RECT 82.400 127.295 82.590 128.190 ;
        RECT 82.910 127.865 83.570 128.135 ;
        RECT 83.240 127.805 83.570 127.865 ;
        RECT 82.760 127.635 83.090 127.695 ;
        RECT 83.760 127.635 83.930 128.395 ;
        RECT 85.170 128.325 85.490 128.785 ;
        RECT 85.690 128.145 85.940 128.575 ;
        RECT 86.230 128.345 86.640 128.785 ;
        RECT 86.810 128.405 87.825 128.605 ;
        RECT 84.100 127.975 85.350 128.145 ;
        RECT 84.100 127.855 84.430 127.975 ;
        RECT 82.760 127.465 84.660 127.635 ;
        RECT 82.400 127.125 84.320 127.295 ;
        RECT 82.400 127.105 82.720 127.125 ;
        RECT 81.950 126.445 82.280 126.955 ;
        RECT 82.550 126.495 82.720 127.105 ;
        RECT 84.490 126.955 84.660 127.465 ;
        RECT 84.830 127.395 85.010 127.805 ;
        RECT 85.180 127.215 85.350 127.975 ;
        RECT 82.890 126.235 83.220 126.925 ;
        RECT 83.450 126.785 84.660 126.955 ;
        RECT 84.830 126.905 85.350 127.215 ;
        RECT 85.520 127.805 85.940 128.145 ;
        RECT 86.230 127.805 86.640 128.135 ;
        RECT 85.520 127.035 85.710 127.805 ;
        RECT 86.810 127.675 86.980 128.405 ;
        RECT 88.125 128.235 88.295 128.565 ;
        RECT 88.465 128.405 88.795 128.785 ;
        RECT 87.150 127.855 87.500 128.225 ;
        RECT 86.810 127.635 87.230 127.675 ;
        RECT 85.880 127.465 87.230 127.635 ;
        RECT 85.880 127.305 86.130 127.465 ;
        RECT 86.640 127.035 86.890 127.295 ;
        RECT 85.520 126.785 86.890 127.035 ;
        RECT 83.450 126.495 83.690 126.785 ;
        RECT 84.490 126.705 84.660 126.785 ;
        RECT 83.890 126.235 84.310 126.615 ;
        RECT 84.490 126.455 85.120 126.705 ;
        RECT 85.590 126.235 85.920 126.615 ;
        RECT 86.090 126.495 86.260 126.785 ;
        RECT 87.060 126.620 87.230 127.465 ;
        RECT 87.680 127.295 87.900 128.165 ;
        RECT 88.125 128.045 88.820 128.235 ;
        RECT 87.400 126.915 87.900 127.295 ;
        RECT 88.070 127.245 88.480 127.865 ;
        RECT 88.650 127.075 88.820 128.045 ;
        RECT 88.125 126.905 88.820 127.075 ;
        RECT 86.440 126.235 86.820 126.615 ;
        RECT 87.060 126.450 87.890 126.620 ;
        RECT 88.125 126.405 88.295 126.905 ;
        RECT 88.465 126.235 88.795 126.735 ;
        RECT 89.010 126.405 89.235 128.525 ;
        RECT 89.405 128.405 89.735 128.785 ;
        RECT 89.905 128.235 90.075 128.525 ;
        RECT 89.410 128.065 90.075 128.235 ;
        RECT 89.410 127.075 89.640 128.065 ;
        RECT 90.335 128.060 90.625 128.785 ;
        RECT 90.855 127.965 91.065 128.785 ;
        RECT 91.235 127.985 91.565 128.615 ;
        RECT 89.810 127.245 90.160 127.895 ;
        RECT 89.410 126.905 90.075 127.075 ;
        RECT 89.405 126.235 89.735 126.735 ;
        RECT 89.905 126.405 90.075 126.905 ;
        RECT 90.335 126.235 90.625 127.400 ;
        RECT 91.235 127.385 91.485 127.985 ;
        RECT 91.735 127.965 91.965 128.785 ;
        RECT 92.175 128.035 93.385 128.785 ;
        RECT 91.655 127.545 91.985 127.795 ;
        RECT 90.855 126.235 91.065 127.375 ;
        RECT 91.235 126.405 91.565 127.385 ;
        RECT 91.735 126.235 91.965 127.375 ;
        RECT 92.175 127.325 92.695 127.865 ;
        RECT 92.865 127.495 93.385 128.035 ;
        RECT 93.555 128.015 97.065 128.785 ;
        RECT 93.555 127.325 95.245 127.845 ;
        RECT 95.415 127.495 97.065 128.015 ;
        RECT 97.435 128.155 97.765 128.515 ;
        RECT 98.385 128.325 98.635 128.785 ;
        RECT 98.805 128.325 99.365 128.615 ;
        RECT 97.435 127.965 98.825 128.155 ;
        RECT 98.655 127.875 98.825 127.965 ;
        RECT 97.250 127.545 97.925 127.795 ;
        RECT 98.145 127.545 98.485 127.795 ;
        RECT 98.655 127.545 98.945 127.875 ;
        RECT 92.175 126.235 93.385 127.325 ;
        RECT 93.555 126.235 97.065 127.325 ;
        RECT 97.250 127.185 97.515 127.545 ;
        RECT 98.655 127.295 98.825 127.545 ;
        RECT 97.885 127.125 98.825 127.295 ;
        RECT 97.435 126.235 97.715 126.905 ;
        RECT 97.885 126.575 98.185 127.125 ;
        RECT 99.115 126.955 99.365 128.325 ;
        RECT 98.385 126.235 98.715 126.955 ;
        RECT 98.905 126.405 99.365 126.955 ;
        RECT 100.455 128.110 100.715 128.615 ;
        RECT 100.895 128.405 101.225 128.785 ;
        RECT 101.405 128.235 101.575 128.615 ;
        RECT 100.455 127.310 100.625 128.110 ;
        RECT 100.910 128.065 101.575 128.235 ;
        RECT 100.910 127.810 101.080 128.065 ;
        RECT 102.295 128.015 103.965 128.785 ;
        RECT 100.795 127.480 101.080 127.810 ;
        RECT 101.315 127.515 101.645 127.885 ;
        RECT 100.910 127.335 101.080 127.480 ;
        RECT 100.455 126.405 100.725 127.310 ;
        RECT 100.910 127.165 101.575 127.335 ;
        RECT 100.895 126.235 101.225 126.995 ;
        RECT 101.405 126.405 101.575 127.165 ;
        RECT 102.295 127.325 103.045 127.845 ;
        RECT 103.215 127.495 103.965 128.015 ;
        RECT 104.335 128.155 104.665 128.515 ;
        RECT 105.285 128.325 105.535 128.785 ;
        RECT 105.705 128.325 106.265 128.615 ;
        RECT 104.335 127.965 105.725 128.155 ;
        RECT 105.555 127.875 105.725 127.965 ;
        RECT 104.150 127.545 104.825 127.795 ;
        RECT 105.045 127.545 105.385 127.795 ;
        RECT 105.555 127.545 105.845 127.875 ;
        RECT 102.295 126.235 103.965 127.325 ;
        RECT 104.150 127.185 104.415 127.545 ;
        RECT 105.555 127.295 105.725 127.545 ;
        RECT 104.785 127.125 105.725 127.295 ;
        RECT 104.335 126.235 104.615 126.905 ;
        RECT 104.785 126.575 105.085 127.125 ;
        RECT 106.015 126.955 106.265 128.325 ;
        RECT 107.395 127.965 107.625 128.785 ;
        RECT 107.795 127.985 108.125 128.615 ;
        RECT 107.375 127.545 107.705 127.795 ;
        RECT 107.875 127.385 108.125 127.985 ;
        RECT 108.295 127.965 108.505 128.785 ;
        RECT 108.735 128.325 109.295 128.615 ;
        RECT 109.465 128.325 109.715 128.785 ;
        RECT 105.285 126.235 105.615 126.955 ;
        RECT 105.805 126.405 106.265 126.955 ;
        RECT 107.395 126.235 107.625 127.375 ;
        RECT 107.795 126.405 108.125 127.385 ;
        RECT 108.295 126.235 108.505 127.375 ;
        RECT 108.735 126.955 108.985 128.325 ;
        RECT 110.335 128.155 110.665 128.515 ;
        RECT 109.275 127.965 110.665 128.155 ;
        RECT 112.155 128.155 112.485 128.515 ;
        RECT 113.105 128.325 113.355 128.785 ;
        RECT 113.525 128.325 114.085 128.615 ;
        RECT 112.155 127.965 113.545 128.155 ;
        RECT 109.275 127.875 109.445 127.965 ;
        RECT 109.155 127.545 109.445 127.875 ;
        RECT 113.375 127.875 113.545 127.965 ;
        RECT 109.615 127.545 109.955 127.795 ;
        RECT 110.175 127.545 110.850 127.795 ;
        RECT 109.275 127.295 109.445 127.545 ;
        RECT 109.275 127.125 110.215 127.295 ;
        RECT 110.585 127.185 110.850 127.545 ;
        RECT 111.970 127.545 112.645 127.795 ;
        RECT 112.865 127.545 113.205 127.795 ;
        RECT 113.375 127.545 113.665 127.875 ;
        RECT 111.970 127.185 112.235 127.545 ;
        RECT 113.375 127.295 113.545 127.545 ;
        RECT 108.735 126.405 109.195 126.955 ;
        RECT 109.385 126.235 109.715 126.955 ;
        RECT 109.915 126.575 110.215 127.125 ;
        RECT 112.605 127.125 113.545 127.295 ;
        RECT 110.385 126.235 110.665 126.905 ;
        RECT 112.155 126.235 112.435 126.905 ;
        RECT 112.605 126.575 112.905 127.125 ;
        RECT 113.835 126.955 114.085 128.325 ;
        RECT 114.255 128.015 115.925 128.785 ;
        RECT 116.095 128.060 116.385 128.785 ;
        RECT 117.020 128.240 122.365 128.785 ;
        RECT 122.540 128.240 127.885 128.785 ;
        RECT 113.105 126.235 113.435 126.955 ;
        RECT 113.625 126.405 114.085 126.955 ;
        RECT 114.255 127.325 115.005 127.845 ;
        RECT 115.175 127.495 115.925 128.015 ;
        RECT 114.255 126.235 115.925 127.325 ;
        RECT 116.095 126.235 116.385 127.400 ;
        RECT 118.610 126.670 118.960 127.920 ;
        RECT 120.440 127.410 120.780 128.240 ;
        RECT 124.130 126.670 124.480 127.920 ;
        RECT 125.960 127.410 126.300 128.240 ;
        RECT 128.055 128.035 129.265 128.785 ;
        RECT 128.055 127.325 128.575 127.865 ;
        RECT 128.745 127.495 129.265 128.035 ;
        RECT 117.020 126.235 122.365 126.670 ;
        RECT 122.540 126.235 127.885 126.670 ;
        RECT 128.055 126.235 129.265 127.325 ;
        RECT 9.290 126.065 129.350 126.235 ;
        RECT 9.375 124.975 10.585 126.065 ;
        RECT 9.375 124.265 9.895 124.805 ;
        RECT 10.065 124.435 10.585 124.975 ;
        RECT 11.675 124.975 15.185 126.065 ;
        RECT 11.675 124.455 13.365 124.975 ;
        RECT 15.395 124.925 15.625 126.065 ;
        RECT 15.795 124.915 16.125 125.895 ;
        RECT 16.295 124.925 16.505 126.065 ;
        RECT 16.735 125.305 17.250 125.715 ;
        RECT 17.485 125.305 17.655 126.065 ;
        RECT 17.825 125.725 19.855 125.895 ;
        RECT 13.535 124.285 15.185 124.805 ;
        RECT 15.375 124.505 15.705 124.755 ;
        RECT 9.375 123.515 10.585 124.265 ;
        RECT 11.675 123.515 15.185 124.285 ;
        RECT 15.395 123.515 15.625 124.335 ;
        RECT 15.875 124.315 16.125 124.915 ;
        RECT 16.735 124.495 17.075 125.305 ;
        RECT 17.825 125.060 17.995 125.725 ;
        RECT 18.390 125.385 19.515 125.555 ;
        RECT 17.245 124.870 17.995 125.060 ;
        RECT 18.165 125.045 19.175 125.215 ;
        RECT 15.795 123.685 16.125 124.315 ;
        RECT 16.295 123.515 16.505 124.335 ;
        RECT 16.735 124.325 17.965 124.495 ;
        RECT 17.010 123.720 17.255 124.325 ;
        RECT 17.475 123.515 17.985 124.050 ;
        RECT 18.165 123.685 18.355 125.045 ;
        RECT 18.525 124.025 18.800 124.845 ;
        RECT 19.005 124.245 19.175 125.045 ;
        RECT 19.345 124.255 19.515 125.385 ;
        RECT 19.685 124.755 19.855 125.725 ;
        RECT 20.025 124.925 20.195 126.065 ;
        RECT 20.365 124.925 20.700 125.895 ;
        RECT 19.685 124.425 19.880 124.755 ;
        RECT 20.105 124.425 20.360 124.755 ;
        RECT 20.105 124.255 20.275 124.425 ;
        RECT 20.530 124.255 20.700 124.925 ;
        RECT 20.875 124.975 24.385 126.065 ;
        RECT 20.875 124.455 22.565 124.975 ;
        RECT 24.595 124.925 24.825 126.065 ;
        RECT 24.995 124.915 25.325 125.895 ;
        RECT 25.495 124.925 25.705 126.065 ;
        RECT 22.735 124.285 24.385 124.805 ;
        RECT 24.575 124.505 24.905 124.755 ;
        RECT 19.345 124.085 20.275 124.255 ;
        RECT 19.345 124.050 19.520 124.085 ;
        RECT 18.525 123.855 18.805 124.025 ;
        RECT 18.525 123.685 18.800 123.855 ;
        RECT 18.990 123.685 19.520 124.050 ;
        RECT 19.945 123.515 20.275 123.915 ;
        RECT 20.445 123.685 20.700 124.255 ;
        RECT 20.875 123.515 24.385 124.285 ;
        RECT 24.595 123.515 24.825 124.335 ;
        RECT 25.075 124.315 25.325 124.915 ;
        RECT 25.935 124.900 26.225 126.065 ;
        RECT 26.770 125.725 27.025 125.755 ;
        RECT 26.685 125.555 27.025 125.725 ;
        RECT 26.770 125.085 27.025 125.555 ;
        RECT 27.205 125.265 27.490 126.065 ;
        RECT 27.670 125.345 28.000 125.855 ;
        RECT 24.995 123.685 25.325 124.315 ;
        RECT 25.495 123.515 25.705 124.335 ;
        RECT 25.935 123.515 26.225 124.240 ;
        RECT 26.770 124.225 26.950 125.085 ;
        RECT 27.670 124.755 27.920 125.345 ;
        RECT 28.270 125.195 28.440 125.805 ;
        RECT 28.610 125.375 28.940 126.065 ;
        RECT 29.170 125.515 29.410 125.805 ;
        RECT 29.610 125.685 30.030 126.065 ;
        RECT 30.210 125.595 30.840 125.845 ;
        RECT 31.310 125.685 31.640 126.065 ;
        RECT 30.210 125.515 30.380 125.595 ;
        RECT 31.810 125.515 31.980 125.805 ;
        RECT 32.160 125.685 32.540 126.065 ;
        RECT 32.780 125.680 33.610 125.850 ;
        RECT 29.170 125.345 30.380 125.515 ;
        RECT 27.120 124.425 27.920 124.755 ;
        RECT 26.770 123.695 27.025 124.225 ;
        RECT 27.205 123.515 27.490 123.975 ;
        RECT 27.670 123.775 27.920 124.425 ;
        RECT 28.120 125.175 28.440 125.195 ;
        RECT 28.120 125.005 30.040 125.175 ;
        RECT 28.120 124.110 28.310 125.005 ;
        RECT 30.210 124.835 30.380 125.345 ;
        RECT 30.550 125.085 31.070 125.395 ;
        RECT 28.480 124.665 30.380 124.835 ;
        RECT 28.480 124.605 28.810 124.665 ;
        RECT 28.960 124.435 29.290 124.495 ;
        RECT 28.630 124.165 29.290 124.435 ;
        RECT 28.120 123.780 28.440 124.110 ;
        RECT 28.620 123.515 29.280 123.995 ;
        RECT 29.480 123.905 29.650 124.665 ;
        RECT 30.550 124.495 30.730 124.905 ;
        RECT 29.820 124.325 30.150 124.445 ;
        RECT 30.900 124.325 31.070 125.085 ;
        RECT 29.820 124.155 31.070 124.325 ;
        RECT 31.240 125.265 32.610 125.515 ;
        RECT 31.240 124.495 31.430 125.265 ;
        RECT 32.360 125.005 32.610 125.265 ;
        RECT 31.600 124.835 31.850 124.995 ;
        RECT 32.780 124.835 32.950 125.680 ;
        RECT 33.845 125.395 34.015 125.895 ;
        RECT 34.185 125.565 34.515 126.065 ;
        RECT 33.120 125.005 33.620 125.385 ;
        RECT 33.845 125.225 34.540 125.395 ;
        RECT 31.600 124.665 32.950 124.835 ;
        RECT 32.530 124.625 32.950 124.665 ;
        RECT 31.240 124.155 31.660 124.495 ;
        RECT 31.950 124.165 32.360 124.495 ;
        RECT 29.480 123.735 30.330 123.905 ;
        RECT 30.890 123.515 31.210 123.975 ;
        RECT 31.410 123.725 31.660 124.155 ;
        RECT 31.950 123.515 32.360 123.955 ;
        RECT 32.530 123.895 32.700 124.625 ;
        RECT 32.870 124.075 33.220 124.445 ;
        RECT 33.400 124.135 33.620 125.005 ;
        RECT 33.790 124.435 34.200 125.055 ;
        RECT 34.370 124.255 34.540 125.225 ;
        RECT 33.845 124.065 34.540 124.255 ;
        RECT 32.530 123.695 33.545 123.895 ;
        RECT 33.845 123.735 34.015 124.065 ;
        RECT 34.185 123.515 34.515 123.895 ;
        RECT 34.730 123.775 34.955 125.895 ;
        RECT 35.125 125.565 35.455 126.065 ;
        RECT 35.625 125.395 35.795 125.895 ;
        RECT 35.130 125.225 35.795 125.395 ;
        RECT 36.115 125.230 36.370 126.065 ;
        RECT 35.130 124.235 35.360 125.225 ;
        RECT 36.540 125.060 36.800 125.865 ;
        RECT 36.970 125.230 37.230 126.065 ;
        RECT 37.400 125.060 37.655 125.865 ;
        RECT 35.530 124.405 35.880 125.055 ;
        RECT 36.055 124.890 37.655 125.060 ;
        RECT 38.855 124.925 39.085 126.065 ;
        RECT 39.255 124.915 39.585 125.895 ;
        RECT 39.755 124.925 39.965 126.065 ;
        RECT 41.125 125.255 41.420 126.065 ;
        RECT 36.055 124.325 36.335 124.890 ;
        RECT 36.505 124.495 37.725 124.720 ;
        RECT 38.835 124.505 39.165 124.755 ;
        RECT 35.130 124.065 35.795 124.235 ;
        RECT 36.055 124.155 36.785 124.325 ;
        RECT 35.125 123.515 35.455 123.895 ;
        RECT 35.625 123.775 35.795 124.065 ;
        RECT 36.060 123.515 36.390 123.985 ;
        RECT 36.560 123.710 36.785 124.155 ;
        RECT 36.955 123.515 37.250 124.040 ;
        RECT 38.855 123.515 39.085 124.335 ;
        RECT 39.335 124.315 39.585 124.915 ;
        RECT 41.600 124.755 41.845 125.895 ;
        RECT 42.020 125.255 42.280 126.065 ;
        RECT 42.880 126.060 49.155 126.065 ;
        RECT 42.460 124.755 42.710 125.890 ;
        RECT 42.880 125.265 43.140 126.060 ;
        RECT 43.310 125.165 43.570 125.890 ;
        RECT 43.740 125.335 44.000 126.060 ;
        RECT 44.170 125.165 44.430 125.890 ;
        RECT 44.600 125.335 44.860 126.060 ;
        RECT 45.030 125.165 45.290 125.890 ;
        RECT 45.460 125.335 45.720 126.060 ;
        RECT 45.890 125.165 46.150 125.890 ;
        RECT 46.320 125.335 46.565 126.060 ;
        RECT 46.735 125.165 46.995 125.890 ;
        RECT 47.180 125.335 47.425 126.060 ;
        RECT 47.595 125.165 47.855 125.890 ;
        RECT 48.040 125.335 48.285 126.060 ;
        RECT 48.455 125.165 48.715 125.890 ;
        RECT 48.900 125.335 49.155 126.060 ;
        RECT 43.310 125.150 48.715 125.165 ;
        RECT 49.325 125.150 49.615 125.890 ;
        RECT 49.785 125.320 50.055 126.065 ;
        RECT 43.310 125.045 50.055 125.150 ;
        RECT 43.310 124.925 50.085 125.045 ;
        RECT 48.890 124.875 50.085 124.925 ;
        RECT 50.315 124.975 51.525 126.065 ;
        RECT 39.255 123.685 39.585 124.315 ;
        RECT 39.755 123.515 39.965 124.335 ;
        RECT 41.115 124.195 41.430 124.755 ;
        RECT 41.600 124.505 48.720 124.755 ;
        RECT 41.115 123.515 41.420 124.025 ;
        RECT 41.600 123.695 41.850 124.505 ;
        RECT 42.020 123.515 42.280 124.040 ;
        RECT 42.460 123.695 42.710 124.505 ;
        RECT 48.890 124.335 50.055 124.875 ;
        RECT 50.315 124.435 50.835 124.975 ;
        RECT 51.695 124.900 51.985 126.065 ;
        RECT 52.620 125.630 57.965 126.065 ;
        RECT 43.310 124.165 50.055 124.335 ;
        RECT 51.005 124.265 51.525 124.805 ;
        RECT 54.210 124.380 54.560 125.630 ;
        RECT 58.225 125.135 58.395 125.895 ;
        RECT 58.575 125.305 58.905 126.065 ;
        RECT 58.225 124.965 58.890 125.135 ;
        RECT 59.075 124.990 59.345 125.895 ;
        RECT 42.880 123.515 43.140 124.075 ;
        RECT 43.310 123.710 43.570 124.165 ;
        RECT 43.740 123.515 44.000 123.995 ;
        RECT 44.170 123.710 44.430 124.165 ;
        RECT 44.600 123.515 44.860 123.995 ;
        RECT 45.030 123.710 45.290 124.165 ;
        RECT 45.460 123.515 45.705 123.995 ;
        RECT 45.875 123.710 46.150 124.165 ;
        RECT 46.320 123.515 46.565 123.995 ;
        RECT 46.735 123.710 46.995 124.165 ;
        RECT 47.175 123.515 47.425 123.995 ;
        RECT 47.595 123.710 47.855 124.165 ;
        RECT 48.035 123.515 48.285 123.995 ;
        RECT 48.455 123.710 48.715 124.165 ;
        RECT 48.895 123.515 49.155 123.995 ;
        RECT 49.325 123.710 49.585 124.165 ;
        RECT 49.755 123.515 50.055 123.995 ;
        RECT 50.315 123.515 51.525 124.265 ;
        RECT 51.695 123.515 51.985 124.240 ;
        RECT 56.040 124.060 56.380 124.890 ;
        RECT 58.720 124.820 58.890 124.965 ;
        RECT 58.155 124.415 58.485 124.785 ;
        RECT 58.720 124.490 59.005 124.820 ;
        RECT 58.720 124.235 58.890 124.490 ;
        RECT 58.225 124.065 58.890 124.235 ;
        RECT 59.175 124.190 59.345 124.990 ;
        RECT 59.515 125.305 60.030 125.715 ;
        RECT 60.265 125.305 60.435 126.065 ;
        RECT 60.605 125.725 62.635 125.895 ;
        RECT 59.515 124.495 59.855 125.305 ;
        RECT 60.605 125.060 60.775 125.725 ;
        RECT 61.170 125.385 62.295 125.555 ;
        RECT 60.025 124.870 60.775 125.060 ;
        RECT 60.945 125.045 61.955 125.215 ;
        RECT 59.515 124.325 60.745 124.495 ;
        RECT 52.620 123.515 57.965 124.060 ;
        RECT 58.225 123.685 58.395 124.065 ;
        RECT 58.575 123.515 58.905 123.895 ;
        RECT 59.085 123.685 59.345 124.190 ;
        RECT 59.790 123.720 60.035 124.325 ;
        RECT 60.255 123.515 60.765 124.050 ;
        RECT 60.945 123.685 61.135 125.045 ;
        RECT 61.305 124.705 61.580 124.845 ;
        RECT 61.305 124.535 61.585 124.705 ;
        RECT 61.305 123.685 61.580 124.535 ;
        RECT 61.785 124.245 61.955 125.045 ;
        RECT 62.125 124.255 62.295 125.385 ;
        RECT 62.465 124.755 62.635 125.725 ;
        RECT 62.805 124.925 62.975 126.065 ;
        RECT 63.145 124.925 63.480 125.895 ;
        RECT 64.580 125.640 64.915 126.065 ;
        RECT 65.085 125.460 65.270 125.865 ;
        RECT 62.465 124.425 62.660 124.755 ;
        RECT 62.885 124.425 63.140 124.755 ;
        RECT 62.885 124.255 63.055 124.425 ;
        RECT 63.310 124.255 63.480 124.925 ;
        RECT 62.125 124.085 63.055 124.255 ;
        RECT 62.125 124.050 62.300 124.085 ;
        RECT 61.770 123.685 62.300 124.050 ;
        RECT 62.725 123.515 63.055 123.915 ;
        RECT 63.225 123.685 63.480 124.255 ;
        RECT 64.605 125.285 65.270 125.460 ;
        RECT 65.475 125.285 65.805 126.065 ;
        RECT 64.605 124.255 64.945 125.285 ;
        RECT 65.975 125.095 66.245 125.865 ;
        RECT 65.115 124.925 66.245 125.095 ;
        RECT 65.115 124.425 65.365 124.925 ;
        RECT 64.605 124.085 65.290 124.255 ;
        RECT 65.545 124.175 65.905 124.755 ;
        RECT 64.580 123.515 64.915 123.915 ;
        RECT 65.085 123.685 65.290 124.085 ;
        RECT 66.075 124.015 66.245 124.925 ;
        RECT 65.500 123.515 65.775 123.995 ;
        RECT 65.985 123.685 66.245 124.015 ;
        RECT 66.415 125.095 66.685 125.865 ;
        RECT 66.855 125.285 67.185 126.065 ;
        RECT 67.390 125.460 67.575 125.865 ;
        RECT 67.745 125.640 68.080 126.065 ;
        RECT 67.390 125.285 68.055 125.460 ;
        RECT 66.415 124.925 67.545 125.095 ;
        RECT 66.415 124.015 66.585 124.925 ;
        RECT 66.755 124.175 67.115 124.755 ;
        RECT 67.295 124.425 67.545 124.925 ;
        RECT 67.715 124.255 68.055 125.285 ;
        RECT 67.370 124.085 68.055 124.255 ;
        RECT 68.255 125.345 68.715 125.895 ;
        RECT 68.905 125.345 69.235 126.065 ;
        RECT 66.415 123.685 66.675 124.015 ;
        RECT 66.885 123.515 67.160 123.995 ;
        RECT 67.370 123.685 67.575 124.085 ;
        RECT 68.255 123.975 68.505 125.345 ;
        RECT 69.435 125.175 69.735 125.725 ;
        RECT 69.905 125.395 70.185 126.065 ;
        RECT 68.795 125.005 69.735 125.175 ;
        RECT 68.795 124.755 68.965 125.005 ;
        RECT 70.105 124.755 70.370 125.115 ;
        RECT 68.675 124.425 68.965 124.755 ;
        RECT 69.135 124.505 69.475 124.755 ;
        RECT 69.695 124.505 70.370 124.755 ;
        RECT 70.555 124.975 71.765 126.065 ;
        RECT 71.940 125.630 77.285 126.065 ;
        RECT 70.555 124.435 71.075 124.975 ;
        RECT 68.795 124.335 68.965 124.425 ;
        RECT 68.795 124.145 70.185 124.335 ;
        RECT 71.245 124.265 71.765 124.805 ;
        RECT 73.530 124.380 73.880 125.630 ;
        RECT 77.455 124.900 77.745 126.065 ;
        RECT 77.915 124.975 80.505 126.065 ;
        RECT 80.685 125.255 80.980 126.065 ;
        RECT 67.745 123.515 68.080 123.915 ;
        RECT 68.255 123.685 68.815 123.975 ;
        RECT 68.985 123.515 69.235 123.975 ;
        RECT 69.855 123.785 70.185 124.145 ;
        RECT 70.555 123.515 71.765 124.265 ;
        RECT 75.360 124.060 75.700 124.890 ;
        RECT 77.915 124.455 79.125 124.975 ;
        RECT 79.295 124.285 80.505 124.805 ;
        RECT 81.160 124.755 81.405 125.895 ;
        RECT 81.580 125.255 81.840 126.065 ;
        RECT 82.440 126.060 88.715 126.065 ;
        RECT 82.020 124.755 82.270 125.890 ;
        RECT 82.440 125.265 82.700 126.060 ;
        RECT 82.870 125.165 83.130 125.890 ;
        RECT 83.300 125.335 83.560 126.060 ;
        RECT 83.730 125.165 83.990 125.890 ;
        RECT 84.160 125.335 84.420 126.060 ;
        RECT 84.590 125.165 84.850 125.890 ;
        RECT 85.020 125.335 85.280 126.060 ;
        RECT 85.450 125.165 85.710 125.890 ;
        RECT 85.880 125.335 86.125 126.060 ;
        RECT 86.295 125.165 86.555 125.890 ;
        RECT 86.740 125.335 86.985 126.060 ;
        RECT 87.155 125.165 87.415 125.890 ;
        RECT 87.600 125.335 87.845 126.060 ;
        RECT 88.015 125.165 88.275 125.890 ;
        RECT 88.460 125.335 88.715 126.060 ;
        RECT 82.870 125.150 88.275 125.165 ;
        RECT 88.885 125.150 89.175 125.890 ;
        RECT 89.345 125.320 89.615 126.065 ;
        RECT 82.870 125.045 89.615 125.150 ;
        RECT 82.870 124.925 89.645 125.045 ;
        RECT 88.450 124.875 89.645 124.925 ;
        RECT 90.335 124.975 93.845 126.065 ;
        RECT 94.025 125.255 94.320 126.065 ;
        RECT 71.940 123.515 77.285 124.060 ;
        RECT 77.455 123.515 77.745 124.240 ;
        RECT 77.915 123.515 80.505 124.285 ;
        RECT 80.675 124.195 80.990 124.755 ;
        RECT 81.160 124.505 88.280 124.755 ;
        RECT 80.675 123.515 80.980 124.025 ;
        RECT 81.160 123.695 81.410 124.505 ;
        RECT 81.580 123.515 81.840 124.040 ;
        RECT 82.020 123.695 82.270 124.505 ;
        RECT 88.450 124.335 89.615 124.875 ;
        RECT 90.335 124.455 92.025 124.975 ;
        RECT 82.870 124.165 89.615 124.335 ;
        RECT 92.195 124.285 93.845 124.805 ;
        RECT 94.500 124.755 94.745 125.895 ;
        RECT 94.920 125.255 95.180 126.065 ;
        RECT 95.780 126.060 102.055 126.065 ;
        RECT 95.360 124.755 95.610 125.890 ;
        RECT 95.780 125.265 96.040 126.060 ;
        RECT 96.210 125.165 96.470 125.890 ;
        RECT 96.640 125.335 96.900 126.060 ;
        RECT 97.070 125.165 97.330 125.890 ;
        RECT 97.500 125.335 97.760 126.060 ;
        RECT 97.930 125.165 98.190 125.890 ;
        RECT 98.360 125.335 98.620 126.060 ;
        RECT 98.790 125.165 99.050 125.890 ;
        RECT 99.220 125.335 99.465 126.060 ;
        RECT 99.635 125.165 99.895 125.890 ;
        RECT 100.080 125.335 100.325 126.060 ;
        RECT 100.495 125.165 100.755 125.890 ;
        RECT 100.940 125.335 101.185 126.060 ;
        RECT 101.355 125.165 101.615 125.890 ;
        RECT 101.800 125.335 102.055 126.060 ;
        RECT 96.210 125.150 101.615 125.165 ;
        RECT 102.225 125.150 102.515 125.890 ;
        RECT 102.685 125.320 102.955 126.065 ;
        RECT 96.210 125.045 102.955 125.150 ;
        RECT 96.210 124.925 102.985 125.045 ;
        RECT 101.790 124.875 102.985 124.925 ;
        RECT 103.215 124.900 103.505 126.065 ;
        RECT 104.135 124.975 106.725 126.065 ;
        RECT 106.895 125.345 107.355 125.895 ;
        RECT 107.545 125.345 107.875 126.065 ;
        RECT 82.440 123.515 82.700 124.075 ;
        RECT 82.870 123.710 83.130 124.165 ;
        RECT 83.300 123.515 83.560 123.995 ;
        RECT 83.730 123.710 83.990 124.165 ;
        RECT 84.160 123.515 84.420 123.995 ;
        RECT 84.590 123.710 84.850 124.165 ;
        RECT 85.020 123.515 85.265 123.995 ;
        RECT 85.435 123.710 85.710 124.165 ;
        RECT 85.880 123.515 86.125 123.995 ;
        RECT 86.295 123.710 86.555 124.165 ;
        RECT 86.735 123.515 86.985 123.995 ;
        RECT 87.155 123.710 87.415 124.165 ;
        RECT 87.595 123.515 87.845 123.995 ;
        RECT 88.015 123.710 88.275 124.165 ;
        RECT 88.455 123.515 88.715 123.995 ;
        RECT 88.885 123.710 89.145 124.165 ;
        RECT 89.315 123.515 89.615 123.995 ;
        RECT 90.335 123.515 93.845 124.285 ;
        RECT 94.015 124.195 94.330 124.755 ;
        RECT 94.500 124.505 101.620 124.755 ;
        RECT 94.015 123.515 94.320 124.025 ;
        RECT 94.500 123.695 94.750 124.505 ;
        RECT 94.920 123.515 95.180 124.040 ;
        RECT 95.360 123.695 95.610 124.505 ;
        RECT 101.790 124.335 102.955 124.875 ;
        RECT 104.135 124.455 105.345 124.975 ;
        RECT 96.210 124.165 102.955 124.335 ;
        RECT 105.515 124.285 106.725 124.805 ;
        RECT 95.780 123.515 96.040 124.075 ;
        RECT 96.210 123.710 96.470 124.165 ;
        RECT 96.640 123.515 96.900 123.995 ;
        RECT 97.070 123.710 97.330 124.165 ;
        RECT 97.500 123.515 97.760 123.995 ;
        RECT 97.930 123.710 98.190 124.165 ;
        RECT 98.360 123.515 98.605 123.995 ;
        RECT 98.775 123.710 99.050 124.165 ;
        RECT 99.220 123.515 99.465 123.995 ;
        RECT 99.635 123.710 99.895 124.165 ;
        RECT 100.075 123.515 100.325 123.995 ;
        RECT 100.495 123.710 100.755 124.165 ;
        RECT 100.935 123.515 101.185 123.995 ;
        RECT 101.355 123.710 101.615 124.165 ;
        RECT 101.795 123.515 102.055 123.995 ;
        RECT 102.225 123.710 102.485 124.165 ;
        RECT 102.655 123.515 102.955 123.995 ;
        RECT 103.215 123.515 103.505 124.240 ;
        RECT 104.135 123.515 106.725 124.285 ;
        RECT 106.895 123.975 107.145 125.345 ;
        RECT 108.075 125.175 108.375 125.725 ;
        RECT 108.545 125.395 108.825 126.065 ;
        RECT 107.435 125.005 108.375 125.175 ;
        RECT 107.435 124.755 107.605 125.005 ;
        RECT 108.745 124.755 109.010 125.115 ;
        RECT 107.315 124.425 107.605 124.755 ;
        RECT 107.775 124.505 108.115 124.755 ;
        RECT 108.335 124.505 109.010 124.755 ;
        RECT 109.195 124.975 110.865 126.065 ;
        RECT 111.035 125.345 111.495 125.895 ;
        RECT 111.685 125.345 112.015 126.065 ;
        RECT 109.195 124.455 109.945 124.975 ;
        RECT 107.435 124.335 107.605 124.425 ;
        RECT 107.435 124.145 108.825 124.335 ;
        RECT 110.115 124.285 110.865 124.805 ;
        RECT 106.895 123.685 107.455 123.975 ;
        RECT 107.625 123.515 107.875 123.975 ;
        RECT 108.495 123.785 108.825 124.145 ;
        RECT 109.195 123.515 110.865 124.285 ;
        RECT 111.035 123.975 111.285 125.345 ;
        RECT 112.215 125.175 112.515 125.725 ;
        RECT 112.685 125.395 112.965 126.065 ;
        RECT 111.575 125.005 112.515 125.175 ;
        RECT 111.575 124.755 111.745 125.005 ;
        RECT 112.885 124.755 113.150 125.115 ;
        RECT 111.455 124.425 111.745 124.755 ;
        RECT 111.915 124.505 112.255 124.755 ;
        RECT 112.475 124.505 113.150 124.755 ;
        RECT 113.335 124.975 115.925 126.065 ;
        RECT 113.335 124.455 114.545 124.975 ;
        RECT 116.135 124.925 116.365 126.065 ;
        RECT 116.535 124.915 116.865 125.895 ;
        RECT 117.035 124.925 117.245 126.065 ;
        RECT 117.850 125.085 118.105 125.755 ;
        RECT 118.285 125.265 118.570 126.065 ;
        RECT 118.750 125.345 119.080 125.855 ;
        RECT 111.575 124.335 111.745 124.425 ;
        RECT 111.575 124.145 112.965 124.335 ;
        RECT 114.715 124.285 115.925 124.805 ;
        RECT 116.115 124.505 116.445 124.755 ;
        RECT 111.035 123.685 111.595 123.975 ;
        RECT 111.765 123.515 112.015 123.975 ;
        RECT 112.635 123.785 112.965 124.145 ;
        RECT 113.335 123.515 115.925 124.285 ;
        RECT 116.135 123.515 116.365 124.335 ;
        RECT 116.615 124.315 116.865 124.915 ;
        RECT 117.850 124.365 118.030 125.085 ;
        RECT 118.750 124.755 119.000 125.345 ;
        RECT 119.350 125.195 119.520 125.805 ;
        RECT 119.690 125.375 120.020 126.065 ;
        RECT 120.250 125.515 120.490 125.805 ;
        RECT 120.690 125.685 121.110 126.065 ;
        RECT 121.290 125.595 121.920 125.845 ;
        RECT 122.390 125.685 122.720 126.065 ;
        RECT 121.290 125.515 121.460 125.595 ;
        RECT 122.890 125.515 123.060 125.805 ;
        RECT 123.240 125.685 123.620 126.065 ;
        RECT 123.860 125.680 124.690 125.850 ;
        RECT 120.250 125.345 121.460 125.515 ;
        RECT 118.200 124.425 119.000 124.755 ;
        RECT 116.535 123.685 116.865 124.315 ;
        RECT 117.035 123.515 117.245 124.335 ;
        RECT 117.765 124.225 118.030 124.365 ;
        RECT 117.765 124.195 118.105 124.225 ;
        RECT 117.850 123.695 118.105 124.195 ;
        RECT 118.285 123.515 118.570 123.975 ;
        RECT 118.750 123.775 119.000 124.425 ;
        RECT 119.200 125.175 119.520 125.195 ;
        RECT 119.200 125.005 121.120 125.175 ;
        RECT 119.200 124.110 119.390 125.005 ;
        RECT 121.290 124.835 121.460 125.345 ;
        RECT 121.630 125.085 122.150 125.395 ;
        RECT 119.560 124.665 121.460 124.835 ;
        RECT 119.560 124.605 119.890 124.665 ;
        RECT 120.040 124.435 120.370 124.495 ;
        RECT 119.710 124.165 120.370 124.435 ;
        RECT 119.200 123.780 119.520 124.110 ;
        RECT 119.700 123.515 120.360 123.995 ;
        RECT 120.560 123.905 120.730 124.665 ;
        RECT 121.630 124.495 121.810 124.905 ;
        RECT 120.900 124.325 121.230 124.445 ;
        RECT 121.980 124.325 122.150 125.085 ;
        RECT 120.900 124.155 122.150 124.325 ;
        RECT 122.320 125.265 123.690 125.515 ;
        RECT 122.320 124.495 122.510 125.265 ;
        RECT 123.440 125.005 123.690 125.265 ;
        RECT 122.680 124.835 122.930 124.995 ;
        RECT 123.860 124.835 124.030 125.680 ;
        RECT 124.925 125.395 125.095 125.895 ;
        RECT 125.265 125.565 125.595 126.065 ;
        RECT 124.200 125.005 124.700 125.385 ;
        RECT 124.925 125.225 125.620 125.395 ;
        RECT 122.680 124.665 124.030 124.835 ;
        RECT 123.610 124.625 124.030 124.665 ;
        RECT 122.320 124.155 122.740 124.495 ;
        RECT 123.030 124.165 123.440 124.495 ;
        RECT 120.560 123.735 121.410 123.905 ;
        RECT 121.970 123.515 122.290 123.975 ;
        RECT 122.490 123.725 122.740 124.155 ;
        RECT 123.030 123.515 123.440 123.955 ;
        RECT 123.610 123.895 123.780 124.625 ;
        RECT 123.950 124.075 124.300 124.445 ;
        RECT 124.480 124.135 124.700 125.005 ;
        RECT 124.870 124.435 125.280 125.055 ;
        RECT 125.450 124.255 125.620 125.225 ;
        RECT 124.925 124.065 125.620 124.255 ;
        RECT 123.610 123.695 124.625 123.895 ;
        RECT 124.925 123.735 125.095 124.065 ;
        RECT 125.265 123.515 125.595 123.895 ;
        RECT 125.810 123.775 126.035 125.895 ;
        RECT 126.205 125.565 126.535 126.065 ;
        RECT 126.705 125.395 126.875 125.895 ;
        RECT 126.210 125.225 126.875 125.395 ;
        RECT 126.210 124.235 126.440 125.225 ;
        RECT 126.610 124.405 126.960 125.055 ;
        RECT 128.055 124.975 129.265 126.065 ;
        RECT 128.055 124.435 128.575 124.975 ;
        RECT 128.745 124.265 129.265 124.805 ;
        RECT 126.210 124.065 126.875 124.235 ;
        RECT 126.205 123.515 126.535 123.895 ;
        RECT 126.705 123.775 126.875 124.065 ;
        RECT 128.055 123.515 129.265 124.265 ;
        RECT 9.290 123.345 129.350 123.515 ;
        RECT 9.375 122.595 10.585 123.345 ;
        RECT 9.375 122.055 9.895 122.595 ;
        RECT 11.215 122.575 12.885 123.345 ;
        RECT 13.055 122.620 13.345 123.345 ;
        RECT 13.520 122.800 18.865 123.345 ;
        RECT 19.040 122.800 24.385 123.345 ;
        RECT 24.560 122.800 29.905 123.345 ;
        RECT 10.065 121.885 10.585 122.425 ;
        RECT 9.375 120.795 10.585 121.885 ;
        RECT 11.215 121.885 11.965 122.405 ;
        RECT 12.135 122.055 12.885 122.575 ;
        RECT 11.215 120.795 12.885 121.885 ;
        RECT 13.055 120.795 13.345 121.960 ;
        RECT 15.110 121.230 15.460 122.480 ;
        RECT 16.940 121.970 17.280 122.800 ;
        RECT 20.630 121.230 20.980 122.480 ;
        RECT 22.460 121.970 22.800 122.800 ;
        RECT 26.150 121.230 26.500 122.480 ;
        RECT 27.980 121.970 28.320 122.800 ;
        RECT 30.275 122.715 30.605 123.075 ;
        RECT 31.225 122.885 31.475 123.345 ;
        RECT 31.645 122.885 32.205 123.175 ;
        RECT 30.275 122.525 31.665 122.715 ;
        RECT 31.495 122.435 31.665 122.525 ;
        RECT 30.090 122.105 30.765 122.355 ;
        RECT 30.985 122.105 31.325 122.355 ;
        RECT 31.495 122.105 31.785 122.435 ;
        RECT 30.090 121.745 30.355 122.105 ;
        RECT 31.495 121.855 31.665 122.105 ;
        RECT 30.725 121.685 31.665 121.855 ;
        RECT 13.520 120.795 18.865 121.230 ;
        RECT 19.040 120.795 24.385 121.230 ;
        RECT 24.560 120.795 29.905 121.230 ;
        RECT 30.275 120.795 30.555 121.465 ;
        RECT 30.725 121.135 31.025 121.685 ;
        RECT 31.955 121.515 32.205 122.885 ;
        RECT 32.575 122.715 32.905 123.075 ;
        RECT 33.525 122.885 33.775 123.345 ;
        RECT 33.945 122.885 34.505 123.175 ;
        RECT 32.575 122.525 33.965 122.715 ;
        RECT 33.795 122.435 33.965 122.525 ;
        RECT 32.390 122.105 33.065 122.355 ;
        RECT 33.285 122.105 33.625 122.355 ;
        RECT 33.795 122.105 34.085 122.435 ;
        RECT 32.390 121.745 32.655 122.105 ;
        RECT 33.795 121.855 33.965 122.105 ;
        RECT 31.225 120.795 31.555 121.515 ;
        RECT 31.745 120.965 32.205 121.515 ;
        RECT 33.025 121.685 33.965 121.855 ;
        RECT 32.575 120.795 32.855 121.465 ;
        RECT 33.025 121.135 33.325 121.685 ;
        RECT 34.255 121.515 34.505 122.885 ;
        RECT 34.950 122.535 35.195 123.140 ;
        RECT 35.415 122.810 35.925 123.345 ;
        RECT 33.525 120.795 33.855 121.515 ;
        RECT 34.045 120.965 34.505 121.515 ;
        RECT 34.675 122.365 35.905 122.535 ;
        RECT 34.675 121.555 35.015 122.365 ;
        RECT 35.185 121.800 35.935 121.990 ;
        RECT 34.675 121.145 35.190 121.555 ;
        RECT 35.425 120.795 35.595 121.555 ;
        RECT 35.765 121.135 35.935 121.800 ;
        RECT 36.105 121.815 36.295 123.175 ;
        RECT 36.465 123.005 36.740 123.175 ;
        RECT 36.465 122.835 36.745 123.005 ;
        RECT 36.465 122.015 36.740 122.835 ;
        RECT 36.930 122.810 37.460 123.175 ;
        RECT 37.885 122.945 38.215 123.345 ;
        RECT 37.285 122.775 37.460 122.810 ;
        RECT 36.945 121.815 37.115 122.615 ;
        RECT 36.105 121.645 37.115 121.815 ;
        RECT 37.285 122.605 38.215 122.775 ;
        RECT 38.385 122.605 38.640 123.175 ;
        RECT 38.815 122.620 39.105 123.345 ;
        RECT 39.935 122.715 40.265 123.075 ;
        RECT 40.885 122.885 41.135 123.345 ;
        RECT 41.305 122.885 41.865 123.175 ;
        RECT 37.285 121.475 37.455 122.605 ;
        RECT 38.045 122.435 38.215 122.605 ;
        RECT 36.330 121.305 37.455 121.475 ;
        RECT 37.625 122.105 37.820 122.435 ;
        RECT 38.045 122.105 38.300 122.435 ;
        RECT 37.625 121.135 37.795 122.105 ;
        RECT 38.470 121.935 38.640 122.605 ;
        RECT 39.935 122.525 41.325 122.715 ;
        RECT 41.155 122.435 41.325 122.525 ;
        RECT 39.750 122.105 40.425 122.355 ;
        RECT 40.645 122.105 40.985 122.355 ;
        RECT 41.155 122.105 41.445 122.435 ;
        RECT 35.765 120.965 37.795 121.135 ;
        RECT 37.965 120.795 38.135 121.935 ;
        RECT 38.305 120.965 38.640 121.935 ;
        RECT 38.815 120.795 39.105 121.960 ;
        RECT 39.750 121.745 40.015 122.105 ;
        RECT 41.155 121.855 41.325 122.105 ;
        RECT 40.385 121.685 41.325 121.855 ;
        RECT 39.935 120.795 40.215 121.465 ;
        RECT 40.385 121.135 40.685 121.685 ;
        RECT 41.615 121.515 41.865 122.885 ;
        RECT 42.125 122.795 42.295 123.175 ;
        RECT 42.475 122.965 42.805 123.345 ;
        RECT 42.125 122.625 42.790 122.795 ;
        RECT 42.985 122.670 43.245 123.175 ;
        RECT 42.055 122.075 42.385 122.445 ;
        RECT 42.620 122.370 42.790 122.625 ;
        RECT 42.620 122.040 42.905 122.370 ;
        RECT 42.620 121.895 42.790 122.040 ;
        RECT 40.885 120.795 41.215 121.515 ;
        RECT 41.405 120.965 41.865 121.515 ;
        RECT 42.125 121.725 42.790 121.895 ;
        RECT 43.075 121.870 43.245 122.670 ;
        RECT 43.415 122.575 46.925 123.345 ;
        RECT 47.615 122.875 47.915 123.345 ;
        RECT 48.085 122.705 48.340 123.150 ;
        RECT 48.510 122.875 48.770 123.345 ;
        RECT 48.940 122.705 49.200 123.150 ;
        RECT 49.370 122.875 49.665 123.345 ;
        RECT 42.125 120.965 42.295 121.725 ;
        RECT 42.475 120.795 42.805 121.555 ;
        RECT 42.975 120.965 43.245 121.870 ;
        RECT 43.415 121.885 45.105 122.405 ;
        RECT 45.275 122.055 46.925 122.575 ;
        RECT 47.095 122.535 50.125 122.705 ;
        RECT 50.315 122.575 53.825 123.345 ;
        RECT 54.370 123.005 54.625 123.165 ;
        RECT 54.285 122.835 54.625 123.005 ;
        RECT 54.805 122.885 55.090 123.345 ;
        RECT 47.095 121.970 47.395 122.535 ;
        RECT 47.570 122.140 49.785 122.365 ;
        RECT 49.955 121.970 50.125 122.535 ;
        RECT 43.415 120.795 46.925 121.885 ;
        RECT 47.095 121.800 50.125 121.970 ;
        RECT 50.315 121.885 52.005 122.405 ;
        RECT 52.175 122.055 53.825 122.575 ;
        RECT 54.370 122.635 54.625 122.835 ;
        RECT 47.095 120.795 47.480 121.630 ;
        RECT 47.650 120.995 47.910 121.800 ;
        RECT 48.080 120.795 48.340 121.630 ;
        RECT 48.510 120.995 48.765 121.800 ;
        RECT 48.940 120.795 49.200 121.630 ;
        RECT 49.370 120.995 49.625 121.800 ;
        RECT 49.800 120.795 50.145 121.630 ;
        RECT 50.315 120.795 53.825 121.885 ;
        RECT 54.370 121.775 54.550 122.635 ;
        RECT 55.270 122.435 55.520 123.085 ;
        RECT 54.720 122.105 55.520 122.435 ;
        RECT 54.370 121.105 54.625 121.775 ;
        RECT 54.805 120.795 55.090 121.595 ;
        RECT 55.270 121.515 55.520 122.105 ;
        RECT 55.720 122.750 56.040 123.080 ;
        RECT 56.220 122.865 56.880 123.345 ;
        RECT 57.080 122.955 57.930 123.125 ;
        RECT 55.720 121.855 55.910 122.750 ;
        RECT 56.230 122.425 56.890 122.695 ;
        RECT 56.560 122.365 56.890 122.425 ;
        RECT 56.080 122.195 56.410 122.255 ;
        RECT 57.080 122.195 57.250 122.955 ;
        RECT 58.490 122.885 58.810 123.345 ;
        RECT 59.010 122.705 59.260 123.135 ;
        RECT 59.550 122.905 59.960 123.345 ;
        RECT 60.130 122.965 61.145 123.165 ;
        RECT 57.420 122.535 58.670 122.705 ;
        RECT 57.420 122.415 57.750 122.535 ;
        RECT 56.080 122.025 57.980 122.195 ;
        RECT 55.720 121.685 57.640 121.855 ;
        RECT 55.720 121.665 56.040 121.685 ;
        RECT 55.270 121.005 55.600 121.515 ;
        RECT 55.870 121.055 56.040 121.665 ;
        RECT 57.810 121.515 57.980 122.025 ;
        RECT 58.150 121.955 58.330 122.365 ;
        RECT 58.500 121.775 58.670 122.535 ;
        RECT 56.210 120.795 56.540 121.485 ;
        RECT 56.770 121.345 57.980 121.515 ;
        RECT 58.150 121.465 58.670 121.775 ;
        RECT 58.840 122.365 59.260 122.705 ;
        RECT 59.550 122.365 59.960 122.695 ;
        RECT 58.840 121.595 59.030 122.365 ;
        RECT 60.130 122.235 60.300 122.965 ;
        RECT 61.445 122.795 61.615 123.125 ;
        RECT 61.785 122.965 62.115 123.345 ;
        RECT 60.470 122.415 60.820 122.785 ;
        RECT 60.130 122.195 60.550 122.235 ;
        RECT 59.200 122.025 60.550 122.195 ;
        RECT 59.200 121.865 59.450 122.025 ;
        RECT 59.960 121.595 60.210 121.855 ;
        RECT 58.840 121.345 60.210 121.595 ;
        RECT 56.770 121.055 57.010 121.345 ;
        RECT 57.810 121.265 57.980 121.345 ;
        RECT 57.210 120.795 57.630 121.175 ;
        RECT 57.810 121.015 58.440 121.265 ;
        RECT 58.910 120.795 59.240 121.175 ;
        RECT 59.410 121.055 59.580 121.345 ;
        RECT 60.380 121.180 60.550 122.025 ;
        RECT 61.000 121.855 61.220 122.725 ;
        RECT 61.445 122.605 62.140 122.795 ;
        RECT 60.720 121.475 61.220 121.855 ;
        RECT 61.390 121.805 61.800 122.425 ;
        RECT 61.970 121.635 62.140 122.605 ;
        RECT 61.445 121.465 62.140 121.635 ;
        RECT 59.760 120.795 60.140 121.175 ;
        RECT 60.380 121.010 61.210 121.180 ;
        RECT 61.445 120.965 61.615 121.465 ;
        RECT 61.785 120.795 62.115 121.295 ;
        RECT 62.330 120.965 62.555 123.085 ;
        RECT 62.725 122.965 63.055 123.345 ;
        RECT 63.225 122.795 63.395 123.085 ;
        RECT 62.730 122.625 63.395 122.795 ;
        RECT 62.730 121.635 62.960 122.625 ;
        RECT 64.575 122.620 64.865 123.345 ;
        RECT 65.095 122.865 65.375 123.345 ;
        RECT 65.545 122.695 65.805 123.085 ;
        RECT 65.980 122.865 66.235 123.345 ;
        RECT 66.405 122.695 66.700 123.085 ;
        RECT 66.880 122.865 67.155 123.345 ;
        RECT 67.325 122.845 67.625 123.175 ;
        RECT 65.050 122.525 66.700 122.695 ;
        RECT 63.130 121.805 63.480 122.455 ;
        RECT 65.050 122.015 65.455 122.525 ;
        RECT 65.625 122.185 66.765 122.355 ;
        RECT 62.730 121.465 63.395 121.635 ;
        RECT 62.725 120.795 63.055 121.295 ;
        RECT 63.225 120.965 63.395 121.465 ;
        RECT 64.575 120.795 64.865 121.960 ;
        RECT 65.050 121.845 65.805 122.015 ;
        RECT 65.090 120.795 65.375 121.665 ;
        RECT 65.545 121.595 65.805 121.845 ;
        RECT 66.595 121.935 66.765 122.185 ;
        RECT 66.935 122.105 67.285 122.675 ;
        RECT 67.455 121.935 67.625 122.845 ;
        RECT 67.795 122.595 69.005 123.345 ;
        RECT 66.595 121.765 67.625 121.935 ;
        RECT 65.545 121.425 66.665 121.595 ;
        RECT 65.545 120.965 65.805 121.425 ;
        RECT 65.980 120.795 66.235 121.255 ;
        RECT 66.405 120.965 66.665 121.425 ;
        RECT 66.835 120.795 67.145 121.595 ;
        RECT 67.315 120.965 67.625 121.765 ;
        RECT 67.795 121.885 68.315 122.425 ;
        RECT 68.485 122.055 69.005 122.595 ;
        RECT 69.175 122.845 69.475 123.175 ;
        RECT 69.645 122.865 69.920 123.345 ;
        RECT 69.175 121.935 69.345 122.845 ;
        RECT 70.100 122.695 70.395 123.085 ;
        RECT 70.565 122.865 70.820 123.345 ;
        RECT 70.995 122.695 71.255 123.085 ;
        RECT 71.425 122.865 71.705 123.345 ;
        RECT 69.515 122.105 69.865 122.675 ;
        RECT 70.100 122.525 71.750 122.695 ;
        RECT 71.935 122.575 74.525 123.345 ;
        RECT 70.035 122.185 71.175 122.355 ;
        RECT 70.035 121.935 70.205 122.185 ;
        RECT 71.345 122.015 71.750 122.525 ;
        RECT 67.795 120.795 69.005 121.885 ;
        RECT 69.175 121.765 70.205 121.935 ;
        RECT 70.995 121.845 71.750 122.015 ;
        RECT 71.935 121.885 73.145 122.405 ;
        RECT 73.315 122.055 74.525 122.575 ;
        RECT 74.895 122.715 75.225 123.075 ;
        RECT 75.845 122.885 76.095 123.345 ;
        RECT 76.265 122.885 76.825 123.175 ;
        RECT 74.895 122.525 76.285 122.715 ;
        RECT 76.115 122.435 76.285 122.525 ;
        RECT 74.710 122.105 75.385 122.355 ;
        RECT 75.605 122.105 75.945 122.355 ;
        RECT 76.115 122.105 76.405 122.435 ;
        RECT 69.175 120.965 69.485 121.765 ;
        RECT 70.995 121.595 71.255 121.845 ;
        RECT 69.655 120.795 69.965 121.595 ;
        RECT 70.135 121.425 71.255 121.595 ;
        RECT 70.135 120.965 70.395 121.425 ;
        RECT 70.565 120.795 70.820 121.255 ;
        RECT 70.995 120.965 71.255 121.425 ;
        RECT 71.425 120.795 71.710 121.665 ;
        RECT 71.935 120.795 74.525 121.885 ;
        RECT 74.710 121.745 74.975 122.105 ;
        RECT 76.115 121.855 76.285 122.105 ;
        RECT 75.345 121.685 76.285 121.855 ;
        RECT 74.895 120.795 75.175 121.465 ;
        RECT 75.345 121.135 75.645 121.685 ;
        RECT 76.575 121.515 76.825 122.885 ;
        RECT 75.845 120.795 76.175 121.515 ;
        RECT 76.365 120.965 76.825 121.515 ;
        RECT 76.995 122.885 77.555 123.175 ;
        RECT 77.725 122.885 77.975 123.345 ;
        RECT 76.995 121.515 77.245 122.885 ;
        RECT 78.595 122.715 78.925 123.075 ;
        RECT 77.535 122.525 78.925 122.715 ;
        RECT 79.755 122.885 80.315 123.175 ;
        RECT 80.485 122.885 80.735 123.345 ;
        RECT 77.535 122.435 77.705 122.525 ;
        RECT 77.415 122.105 77.705 122.435 ;
        RECT 77.875 122.105 78.215 122.355 ;
        RECT 78.435 122.105 79.110 122.355 ;
        RECT 77.535 121.855 77.705 122.105 ;
        RECT 77.535 121.685 78.475 121.855 ;
        RECT 78.845 121.745 79.110 122.105 ;
        RECT 76.995 120.965 77.455 121.515 ;
        RECT 77.645 120.795 77.975 121.515 ;
        RECT 78.175 121.135 78.475 121.685 ;
        RECT 79.755 121.515 80.005 122.885 ;
        RECT 81.355 122.715 81.685 123.075 ;
        RECT 80.295 122.525 81.685 122.715 ;
        RECT 82.055 122.885 82.615 123.175 ;
        RECT 82.785 122.885 83.035 123.345 ;
        RECT 80.295 122.435 80.465 122.525 ;
        RECT 80.175 122.105 80.465 122.435 ;
        RECT 80.635 122.105 80.975 122.355 ;
        RECT 81.195 122.105 81.870 122.355 ;
        RECT 80.295 121.855 80.465 122.105 ;
        RECT 80.295 121.685 81.235 121.855 ;
        RECT 81.605 121.745 81.870 122.105 ;
        RECT 78.645 120.795 78.925 121.465 ;
        RECT 79.755 120.965 80.215 121.515 ;
        RECT 80.405 120.795 80.735 121.515 ;
        RECT 80.935 121.135 81.235 121.685 ;
        RECT 82.055 121.515 82.305 122.885 ;
        RECT 83.655 122.715 83.985 123.075 ;
        RECT 82.595 122.525 83.985 122.715 ;
        RECT 84.815 122.575 86.485 123.345 ;
        RECT 87.175 122.875 87.475 123.345 ;
        RECT 87.645 122.705 87.900 123.150 ;
        RECT 88.070 122.875 88.330 123.345 ;
        RECT 88.500 122.705 88.760 123.150 ;
        RECT 88.930 122.875 89.225 123.345 ;
        RECT 82.595 122.435 82.765 122.525 ;
        RECT 82.475 122.105 82.765 122.435 ;
        RECT 82.935 122.105 83.275 122.355 ;
        RECT 83.495 122.105 84.170 122.355 ;
        RECT 82.595 121.855 82.765 122.105 ;
        RECT 82.595 121.685 83.535 121.855 ;
        RECT 83.905 121.745 84.170 122.105 ;
        RECT 84.815 121.885 85.565 122.405 ;
        RECT 85.735 122.055 86.485 122.575 ;
        RECT 86.655 122.535 89.685 122.705 ;
        RECT 90.335 122.620 90.625 123.345 ;
        RECT 90.795 122.575 93.385 123.345 ;
        RECT 93.560 122.800 98.905 123.345 ;
        RECT 99.080 122.800 104.425 123.345 ;
        RECT 86.655 121.970 86.955 122.535 ;
        RECT 87.130 122.140 89.345 122.365 ;
        RECT 89.515 121.970 89.685 122.535 ;
        RECT 81.405 120.795 81.685 121.465 ;
        RECT 82.055 120.965 82.515 121.515 ;
        RECT 82.705 120.795 83.035 121.515 ;
        RECT 83.235 121.135 83.535 121.685 ;
        RECT 83.705 120.795 83.985 121.465 ;
        RECT 84.815 120.795 86.485 121.885 ;
        RECT 86.655 121.800 89.685 121.970 ;
        RECT 86.655 120.795 87.040 121.630 ;
        RECT 87.210 120.995 87.470 121.800 ;
        RECT 87.640 120.795 87.900 121.630 ;
        RECT 88.070 120.995 88.325 121.800 ;
        RECT 88.500 120.795 88.760 121.630 ;
        RECT 88.930 120.995 89.185 121.800 ;
        RECT 89.360 120.795 89.705 121.630 ;
        RECT 90.335 120.795 90.625 121.960 ;
        RECT 90.795 121.885 92.005 122.405 ;
        RECT 92.175 122.055 93.385 122.575 ;
        RECT 90.795 120.795 93.385 121.885 ;
        RECT 95.150 121.230 95.500 122.480 ;
        RECT 96.980 121.970 97.320 122.800 ;
        RECT 100.670 121.230 101.020 122.480 ;
        RECT 102.500 121.970 102.840 122.800 ;
        RECT 104.635 122.525 104.865 123.345 ;
        RECT 105.035 122.545 105.365 123.175 ;
        RECT 104.615 122.105 104.945 122.355 ;
        RECT 105.115 121.945 105.365 122.545 ;
        RECT 105.535 122.525 105.745 123.345 ;
        RECT 106.710 122.535 106.955 123.140 ;
        RECT 107.175 122.810 107.685 123.345 ;
        RECT 93.560 120.795 98.905 121.230 ;
        RECT 99.080 120.795 104.425 121.230 ;
        RECT 104.635 120.795 104.865 121.935 ;
        RECT 105.035 120.965 105.365 121.945 ;
        RECT 106.435 122.365 107.665 122.535 ;
        RECT 105.535 120.795 105.745 121.935 ;
        RECT 106.435 121.555 106.775 122.365 ;
        RECT 106.945 121.800 107.695 121.990 ;
        RECT 106.435 121.145 106.950 121.555 ;
        RECT 107.185 120.795 107.355 121.555 ;
        RECT 107.525 121.135 107.695 121.800 ;
        RECT 107.865 121.815 108.055 123.175 ;
        RECT 108.225 122.325 108.500 123.175 ;
        RECT 108.690 122.810 109.220 123.175 ;
        RECT 109.645 122.945 109.975 123.345 ;
        RECT 109.045 122.775 109.220 122.810 ;
        RECT 108.225 122.155 108.505 122.325 ;
        RECT 108.225 122.015 108.500 122.155 ;
        RECT 108.705 121.815 108.875 122.615 ;
        RECT 107.865 121.645 108.875 121.815 ;
        RECT 109.045 122.605 109.975 122.775 ;
        RECT 110.145 122.605 110.400 123.175 ;
        RECT 109.045 121.475 109.215 122.605 ;
        RECT 109.805 122.435 109.975 122.605 ;
        RECT 108.090 121.305 109.215 121.475 ;
        RECT 109.385 122.105 109.580 122.435 ;
        RECT 109.805 122.105 110.060 122.435 ;
        RECT 109.385 121.135 109.555 122.105 ;
        RECT 110.230 121.935 110.400 122.605 ;
        RECT 110.575 122.595 111.785 123.345 ;
        RECT 107.525 120.965 109.555 121.135 ;
        RECT 109.725 120.795 109.895 121.935 ;
        RECT 110.065 120.965 110.400 121.935 ;
        RECT 110.575 121.885 111.095 122.425 ;
        RECT 111.265 122.055 111.785 122.595 ;
        RECT 112.230 122.535 112.475 123.140 ;
        RECT 112.695 122.810 113.205 123.345 ;
        RECT 111.955 122.365 113.185 122.535 ;
        RECT 110.575 120.795 111.785 121.885 ;
        RECT 111.955 121.555 112.295 122.365 ;
        RECT 112.465 121.800 113.215 121.990 ;
        RECT 111.955 121.145 112.470 121.555 ;
        RECT 112.705 120.795 112.875 121.555 ;
        RECT 113.045 121.135 113.215 121.800 ;
        RECT 113.385 121.815 113.575 123.175 ;
        RECT 113.745 123.005 114.020 123.175 ;
        RECT 113.745 122.835 114.025 123.005 ;
        RECT 113.745 122.015 114.020 122.835 ;
        RECT 114.210 122.810 114.740 123.175 ;
        RECT 115.165 122.945 115.495 123.345 ;
        RECT 114.565 122.775 114.740 122.810 ;
        RECT 114.225 121.815 114.395 122.615 ;
        RECT 113.385 121.645 114.395 121.815 ;
        RECT 114.565 122.605 115.495 122.775 ;
        RECT 115.665 122.605 115.920 123.175 ;
        RECT 116.095 122.620 116.385 123.345 ;
        RECT 116.930 123.005 117.185 123.165 ;
        RECT 116.845 122.835 117.185 123.005 ;
        RECT 117.365 122.885 117.650 123.345 ;
        RECT 116.930 122.635 117.185 122.835 ;
        RECT 114.565 121.475 114.735 122.605 ;
        RECT 115.325 122.435 115.495 122.605 ;
        RECT 113.610 121.305 114.735 121.475 ;
        RECT 114.905 122.105 115.100 122.435 ;
        RECT 115.325 122.105 115.580 122.435 ;
        RECT 114.905 121.135 115.075 122.105 ;
        RECT 115.750 121.935 115.920 122.605 ;
        RECT 113.045 120.965 115.075 121.135 ;
        RECT 115.245 120.795 115.415 121.935 ;
        RECT 115.585 120.965 115.920 121.935 ;
        RECT 116.095 120.795 116.385 121.960 ;
        RECT 116.930 121.775 117.110 122.635 ;
        RECT 117.830 122.435 118.080 123.085 ;
        RECT 117.280 122.105 118.080 122.435 ;
        RECT 116.930 121.105 117.185 121.775 ;
        RECT 117.365 120.795 117.650 121.595 ;
        RECT 117.830 121.515 118.080 122.105 ;
        RECT 118.280 122.750 118.600 123.080 ;
        RECT 118.780 122.865 119.440 123.345 ;
        RECT 119.640 122.955 120.490 123.125 ;
        RECT 118.280 121.855 118.470 122.750 ;
        RECT 118.790 122.425 119.450 122.695 ;
        RECT 119.120 122.365 119.450 122.425 ;
        RECT 118.640 122.195 118.970 122.255 ;
        RECT 119.640 122.195 119.810 122.955 ;
        RECT 121.050 122.885 121.370 123.345 ;
        RECT 121.570 122.705 121.820 123.135 ;
        RECT 122.110 122.905 122.520 123.345 ;
        RECT 122.690 122.965 123.705 123.165 ;
        RECT 119.980 122.535 121.230 122.705 ;
        RECT 119.980 122.415 120.310 122.535 ;
        RECT 118.640 122.025 120.540 122.195 ;
        RECT 118.280 121.685 120.200 121.855 ;
        RECT 118.280 121.665 118.600 121.685 ;
        RECT 117.830 121.005 118.160 121.515 ;
        RECT 118.430 121.055 118.600 121.665 ;
        RECT 120.370 121.515 120.540 122.025 ;
        RECT 120.710 121.955 120.890 122.365 ;
        RECT 121.060 121.775 121.230 122.535 ;
        RECT 118.770 120.795 119.100 121.485 ;
        RECT 119.330 121.345 120.540 121.515 ;
        RECT 120.710 121.465 121.230 121.775 ;
        RECT 121.400 122.365 121.820 122.705 ;
        RECT 122.110 122.365 122.520 122.695 ;
        RECT 121.400 121.595 121.590 122.365 ;
        RECT 122.690 122.235 122.860 122.965 ;
        RECT 124.005 122.795 124.175 123.125 ;
        RECT 124.345 122.965 124.675 123.345 ;
        RECT 123.030 122.415 123.380 122.785 ;
        RECT 122.690 122.195 123.110 122.235 ;
        RECT 121.760 122.025 123.110 122.195 ;
        RECT 121.760 121.865 122.010 122.025 ;
        RECT 122.520 121.595 122.770 121.855 ;
        RECT 121.400 121.345 122.770 121.595 ;
        RECT 119.330 121.055 119.570 121.345 ;
        RECT 120.370 121.265 120.540 121.345 ;
        RECT 119.770 120.795 120.190 121.175 ;
        RECT 120.370 121.015 121.000 121.265 ;
        RECT 121.470 120.795 121.800 121.175 ;
        RECT 121.970 121.055 122.140 121.345 ;
        RECT 122.940 121.180 123.110 122.025 ;
        RECT 123.560 121.855 123.780 122.725 ;
        RECT 124.005 122.605 124.700 122.795 ;
        RECT 123.280 121.475 123.780 121.855 ;
        RECT 123.950 121.805 124.360 122.425 ;
        RECT 124.530 121.635 124.700 122.605 ;
        RECT 124.005 121.465 124.700 121.635 ;
        RECT 122.320 120.795 122.700 121.175 ;
        RECT 122.940 121.010 123.770 121.180 ;
        RECT 124.005 120.965 124.175 121.465 ;
        RECT 124.345 120.795 124.675 121.295 ;
        RECT 124.890 120.965 125.115 123.085 ;
        RECT 125.285 122.965 125.615 123.345 ;
        RECT 125.785 122.795 125.955 123.085 ;
        RECT 125.290 122.625 125.955 122.795 ;
        RECT 126.215 122.670 126.475 123.175 ;
        RECT 126.655 122.965 126.985 123.345 ;
        RECT 127.165 122.795 127.335 123.175 ;
        RECT 125.290 121.635 125.520 122.625 ;
        RECT 125.690 121.805 126.040 122.455 ;
        RECT 126.215 121.870 126.385 122.670 ;
        RECT 126.670 122.625 127.335 122.795 ;
        RECT 126.670 122.370 126.840 122.625 ;
        RECT 128.055 122.595 129.265 123.345 ;
        RECT 126.555 122.040 126.840 122.370 ;
        RECT 127.075 122.075 127.405 122.445 ;
        RECT 126.670 121.895 126.840 122.040 ;
        RECT 125.290 121.465 125.955 121.635 ;
        RECT 125.285 120.795 125.615 121.295 ;
        RECT 125.785 120.965 125.955 121.465 ;
        RECT 126.215 120.965 126.485 121.870 ;
        RECT 126.670 121.725 127.335 121.895 ;
        RECT 126.655 120.795 126.985 121.555 ;
        RECT 127.165 120.965 127.335 121.725 ;
        RECT 128.055 121.885 128.575 122.425 ;
        RECT 128.745 122.055 129.265 122.595 ;
        RECT 128.055 120.795 129.265 121.885 ;
        RECT 9.290 120.625 129.350 120.795 ;
        RECT 9.375 119.535 10.585 120.625 ;
        RECT 11.220 120.190 16.565 120.625 ;
        RECT 9.375 118.825 9.895 119.365 ;
        RECT 10.065 118.995 10.585 119.535 ;
        RECT 12.810 118.940 13.160 120.190 ;
        RECT 16.735 119.865 17.250 120.275 ;
        RECT 17.485 119.865 17.655 120.625 ;
        RECT 17.825 120.285 19.855 120.455 ;
        RECT 9.375 118.075 10.585 118.825 ;
        RECT 14.640 118.620 14.980 119.450 ;
        RECT 16.735 119.055 17.075 119.865 ;
        RECT 17.825 119.620 17.995 120.285 ;
        RECT 18.390 119.945 19.515 120.115 ;
        RECT 17.245 119.430 17.995 119.620 ;
        RECT 18.165 119.605 19.175 119.775 ;
        RECT 16.735 118.885 17.965 119.055 ;
        RECT 11.220 118.075 16.565 118.620 ;
        RECT 17.010 118.280 17.255 118.885 ;
        RECT 17.475 118.075 17.985 118.610 ;
        RECT 18.165 118.245 18.355 119.605 ;
        RECT 18.525 119.265 18.800 119.405 ;
        RECT 18.525 119.095 18.805 119.265 ;
        RECT 18.525 118.245 18.800 119.095 ;
        RECT 19.005 118.805 19.175 119.605 ;
        RECT 19.345 118.815 19.515 119.945 ;
        RECT 19.685 119.315 19.855 120.285 ;
        RECT 20.025 119.485 20.195 120.625 ;
        RECT 20.365 119.485 20.700 120.455 ;
        RECT 19.685 118.985 19.880 119.315 ;
        RECT 20.105 118.985 20.360 119.315 ;
        RECT 20.105 118.815 20.275 118.985 ;
        RECT 20.530 118.815 20.700 119.485 ;
        RECT 19.345 118.645 20.275 118.815 ;
        RECT 19.345 118.610 19.520 118.645 ;
        RECT 18.990 118.245 19.520 118.610 ;
        RECT 19.945 118.075 20.275 118.475 ;
        RECT 20.445 118.245 20.700 118.815 ;
        RECT 21.800 119.485 22.135 120.455 ;
        RECT 22.305 119.485 22.475 120.625 ;
        RECT 22.645 120.285 24.675 120.455 ;
        RECT 21.800 118.815 21.970 119.485 ;
        RECT 22.645 119.315 22.815 120.285 ;
        RECT 22.140 118.985 22.395 119.315 ;
        RECT 22.620 118.985 22.815 119.315 ;
        RECT 22.985 119.945 24.110 120.115 ;
        RECT 22.225 118.815 22.395 118.985 ;
        RECT 22.985 118.815 23.155 119.945 ;
        RECT 21.800 118.245 22.055 118.815 ;
        RECT 22.225 118.645 23.155 118.815 ;
        RECT 23.325 119.605 24.335 119.775 ;
        RECT 23.325 118.805 23.495 119.605 ;
        RECT 23.700 118.925 23.975 119.405 ;
        RECT 23.695 118.755 23.975 118.925 ;
        RECT 22.980 118.610 23.155 118.645 ;
        RECT 22.225 118.075 22.555 118.475 ;
        RECT 22.980 118.245 23.510 118.610 ;
        RECT 23.700 118.245 23.975 118.755 ;
        RECT 24.145 118.245 24.335 119.605 ;
        RECT 24.505 119.620 24.675 120.285 ;
        RECT 24.845 119.865 25.015 120.625 ;
        RECT 25.250 119.865 25.765 120.275 ;
        RECT 24.505 119.430 25.255 119.620 ;
        RECT 25.425 119.055 25.765 119.865 ;
        RECT 25.935 119.460 26.225 120.625 ;
        RECT 27.315 119.535 30.825 120.625 ;
        RECT 24.535 118.885 25.765 119.055 ;
        RECT 27.315 119.015 29.005 119.535 ;
        RECT 31.000 119.485 31.335 120.455 ;
        RECT 31.505 119.485 31.675 120.625 ;
        RECT 31.845 120.285 33.875 120.455 ;
        RECT 24.515 118.075 25.025 118.610 ;
        RECT 25.245 118.280 25.490 118.885 ;
        RECT 29.175 118.845 30.825 119.365 ;
        RECT 25.935 118.075 26.225 118.800 ;
        RECT 27.315 118.075 30.825 118.845 ;
        RECT 31.000 118.815 31.170 119.485 ;
        RECT 31.845 119.315 32.015 120.285 ;
        RECT 31.340 118.985 31.595 119.315 ;
        RECT 31.820 118.985 32.015 119.315 ;
        RECT 32.185 119.945 33.310 120.115 ;
        RECT 31.425 118.815 31.595 118.985 ;
        RECT 32.185 118.815 32.355 119.945 ;
        RECT 31.000 118.245 31.255 118.815 ;
        RECT 31.425 118.645 32.355 118.815 ;
        RECT 32.525 119.605 33.535 119.775 ;
        RECT 32.525 118.805 32.695 119.605 ;
        RECT 32.900 119.265 33.175 119.405 ;
        RECT 32.895 119.095 33.175 119.265 ;
        RECT 32.180 118.610 32.355 118.645 ;
        RECT 31.425 118.075 31.755 118.475 ;
        RECT 32.180 118.245 32.710 118.610 ;
        RECT 32.900 118.245 33.175 119.095 ;
        RECT 33.345 118.245 33.535 119.605 ;
        RECT 33.705 119.620 33.875 120.285 ;
        RECT 34.045 119.865 34.215 120.625 ;
        RECT 34.450 119.865 34.965 120.275 ;
        RECT 33.705 119.430 34.455 119.620 ;
        RECT 34.625 119.055 34.965 119.865 ;
        RECT 33.735 118.885 34.965 119.055 ;
        RECT 35.970 119.645 36.225 120.315 ;
        RECT 36.405 119.825 36.690 120.625 ;
        RECT 36.870 119.905 37.200 120.415 ;
        RECT 33.715 118.075 34.225 118.610 ;
        RECT 34.445 118.280 34.690 118.885 ;
        RECT 35.970 118.785 36.150 119.645 ;
        RECT 36.870 119.315 37.120 119.905 ;
        RECT 37.470 119.755 37.640 120.365 ;
        RECT 37.810 119.935 38.140 120.625 ;
        RECT 38.370 120.075 38.610 120.365 ;
        RECT 38.810 120.245 39.230 120.625 ;
        RECT 39.410 120.155 40.040 120.405 ;
        RECT 40.510 120.245 40.840 120.625 ;
        RECT 39.410 120.075 39.580 120.155 ;
        RECT 41.010 120.075 41.180 120.365 ;
        RECT 41.360 120.245 41.740 120.625 ;
        RECT 41.980 120.240 42.810 120.410 ;
        RECT 38.370 119.905 39.580 120.075 ;
        RECT 36.320 118.985 37.120 119.315 ;
        RECT 35.970 118.585 36.225 118.785 ;
        RECT 35.885 118.415 36.225 118.585 ;
        RECT 35.970 118.255 36.225 118.415 ;
        RECT 36.405 118.075 36.690 118.535 ;
        RECT 36.870 118.335 37.120 118.985 ;
        RECT 37.320 119.735 37.640 119.755 ;
        RECT 37.320 119.565 39.240 119.735 ;
        RECT 37.320 118.670 37.510 119.565 ;
        RECT 39.410 119.395 39.580 119.905 ;
        RECT 39.750 119.645 40.270 119.955 ;
        RECT 37.680 119.225 39.580 119.395 ;
        RECT 37.680 119.165 38.010 119.225 ;
        RECT 38.160 118.995 38.490 119.055 ;
        RECT 37.830 118.725 38.490 118.995 ;
        RECT 37.320 118.340 37.640 118.670 ;
        RECT 37.820 118.075 38.480 118.555 ;
        RECT 38.680 118.465 38.850 119.225 ;
        RECT 39.750 119.055 39.930 119.465 ;
        RECT 39.020 118.885 39.350 119.005 ;
        RECT 40.100 118.885 40.270 119.645 ;
        RECT 39.020 118.715 40.270 118.885 ;
        RECT 40.440 119.825 41.810 120.075 ;
        RECT 40.440 119.055 40.630 119.825 ;
        RECT 41.560 119.565 41.810 119.825 ;
        RECT 40.800 119.395 41.050 119.555 ;
        RECT 41.980 119.395 42.150 120.240 ;
        RECT 43.045 119.955 43.215 120.455 ;
        RECT 43.385 120.125 43.715 120.625 ;
        RECT 42.320 119.565 42.820 119.945 ;
        RECT 43.045 119.785 43.740 119.955 ;
        RECT 40.800 119.225 42.150 119.395 ;
        RECT 41.730 119.185 42.150 119.225 ;
        RECT 40.440 118.715 40.860 119.055 ;
        RECT 41.150 118.725 41.560 119.055 ;
        RECT 38.680 118.295 39.530 118.465 ;
        RECT 40.090 118.075 40.410 118.535 ;
        RECT 40.610 118.285 40.860 118.715 ;
        RECT 41.150 118.075 41.560 118.515 ;
        RECT 41.730 118.455 41.900 119.185 ;
        RECT 42.070 118.635 42.420 119.005 ;
        RECT 42.600 118.695 42.820 119.565 ;
        RECT 42.990 118.995 43.400 119.615 ;
        RECT 43.570 118.815 43.740 119.785 ;
        RECT 43.045 118.625 43.740 118.815 ;
        RECT 41.730 118.255 42.745 118.455 ;
        RECT 43.045 118.295 43.215 118.625 ;
        RECT 43.385 118.075 43.715 118.455 ;
        RECT 43.930 118.335 44.155 120.455 ;
        RECT 44.325 120.125 44.655 120.625 ;
        RECT 44.825 119.955 44.995 120.455 ;
        RECT 44.330 119.785 44.995 119.955 ;
        RECT 45.255 119.905 45.715 120.455 ;
        RECT 45.905 119.905 46.235 120.625 ;
        RECT 44.330 118.795 44.560 119.785 ;
        RECT 44.730 118.965 45.080 119.615 ;
        RECT 44.330 118.625 44.995 118.795 ;
        RECT 44.325 118.075 44.655 118.455 ;
        RECT 44.825 118.335 44.995 118.625 ;
        RECT 45.255 118.535 45.505 119.905 ;
        RECT 46.435 119.735 46.735 120.285 ;
        RECT 46.905 119.955 47.185 120.625 ;
        RECT 45.795 119.565 46.735 119.735 ;
        RECT 48.475 119.905 48.935 120.455 ;
        RECT 49.125 119.905 49.455 120.625 ;
        RECT 45.795 119.315 45.965 119.565 ;
        RECT 47.105 119.315 47.370 119.675 ;
        RECT 45.675 118.985 45.965 119.315 ;
        RECT 46.135 119.065 46.475 119.315 ;
        RECT 46.695 119.065 47.370 119.315 ;
        RECT 45.795 118.895 45.965 118.985 ;
        RECT 45.795 118.705 47.185 118.895 ;
        RECT 45.255 118.245 45.815 118.535 ;
        RECT 45.985 118.075 46.235 118.535 ;
        RECT 46.855 118.345 47.185 118.705 ;
        RECT 48.475 118.535 48.725 119.905 ;
        RECT 49.655 119.735 49.955 120.285 ;
        RECT 50.125 119.955 50.405 120.625 ;
        RECT 49.015 119.565 49.955 119.735 ;
        RECT 49.015 119.315 49.185 119.565 ;
        RECT 50.325 119.315 50.590 119.675 ;
        RECT 51.695 119.460 51.985 120.625 ;
        RECT 53.080 120.190 58.425 120.625 ;
        RECT 48.895 118.985 49.185 119.315 ;
        RECT 49.355 119.065 49.695 119.315 ;
        RECT 49.915 119.065 50.590 119.315 ;
        RECT 49.015 118.895 49.185 118.985 ;
        RECT 54.670 118.940 55.020 120.190 ;
        RECT 58.655 119.485 58.865 120.625 ;
        RECT 59.035 119.475 59.365 120.455 ;
        RECT 59.535 119.485 59.765 120.625 ;
        RECT 60.895 119.535 64.405 120.625 ;
        RECT 64.665 119.695 64.835 120.455 ;
        RECT 65.015 119.865 65.345 120.625 ;
        RECT 49.015 118.705 50.405 118.895 ;
        RECT 48.475 118.245 49.035 118.535 ;
        RECT 49.205 118.075 49.455 118.535 ;
        RECT 50.075 118.345 50.405 118.705 ;
        RECT 51.695 118.075 51.985 118.800 ;
        RECT 56.500 118.620 56.840 119.450 ;
        RECT 53.080 118.075 58.425 118.620 ;
        RECT 58.655 118.075 58.865 118.895 ;
        RECT 59.035 118.875 59.285 119.475 ;
        RECT 59.455 119.065 59.785 119.315 ;
        RECT 60.895 119.015 62.585 119.535 ;
        RECT 64.665 119.525 65.330 119.695 ;
        RECT 65.515 119.550 65.785 120.455 ;
        RECT 66.420 120.190 71.765 120.625 ;
        RECT 71.940 120.190 77.285 120.625 ;
        RECT 65.160 119.380 65.330 119.525 ;
        RECT 59.035 118.245 59.365 118.875 ;
        RECT 59.535 118.075 59.765 118.895 ;
        RECT 62.755 118.845 64.405 119.365 ;
        RECT 64.595 118.975 64.925 119.345 ;
        RECT 65.160 119.050 65.445 119.380 ;
        RECT 60.895 118.075 64.405 118.845 ;
        RECT 65.160 118.795 65.330 119.050 ;
        RECT 64.665 118.625 65.330 118.795 ;
        RECT 65.615 118.750 65.785 119.550 ;
        RECT 68.010 118.940 68.360 120.190 ;
        RECT 64.665 118.245 64.835 118.625 ;
        RECT 65.015 118.075 65.345 118.455 ;
        RECT 65.525 118.245 65.785 118.750 ;
        RECT 69.840 118.620 70.180 119.450 ;
        RECT 73.530 118.940 73.880 120.190 ;
        RECT 77.455 119.460 77.745 120.625 ;
        RECT 77.915 119.535 79.125 120.625 ;
        RECT 79.295 119.550 79.565 120.455 ;
        RECT 79.735 119.865 80.065 120.625 ;
        RECT 80.245 119.695 80.415 120.455 ;
        RECT 75.360 118.620 75.700 119.450 ;
        RECT 77.915 118.995 78.435 119.535 ;
        RECT 78.605 118.825 79.125 119.365 ;
        RECT 66.420 118.075 71.765 118.620 ;
        RECT 71.940 118.075 77.285 118.620 ;
        RECT 77.455 118.075 77.745 118.800 ;
        RECT 77.915 118.075 79.125 118.825 ;
        RECT 79.295 118.750 79.465 119.550 ;
        RECT 79.750 119.525 80.415 119.695 ;
        RECT 81.595 119.865 82.110 120.275 ;
        RECT 82.345 119.865 82.515 120.625 ;
        RECT 82.685 120.285 84.715 120.455 ;
        RECT 79.750 119.380 79.920 119.525 ;
        RECT 79.635 119.050 79.920 119.380 ;
        RECT 79.750 118.795 79.920 119.050 ;
        RECT 80.155 118.975 80.485 119.345 ;
        RECT 81.595 119.055 81.935 119.865 ;
        RECT 82.685 119.620 82.855 120.285 ;
        RECT 83.250 119.945 84.375 120.115 ;
        RECT 82.105 119.430 82.855 119.620 ;
        RECT 83.025 119.605 84.035 119.775 ;
        RECT 81.595 118.885 82.825 119.055 ;
        RECT 79.295 118.245 79.555 118.750 ;
        RECT 79.750 118.625 80.415 118.795 ;
        RECT 79.735 118.075 80.065 118.455 ;
        RECT 80.245 118.245 80.415 118.625 ;
        RECT 81.870 118.280 82.115 118.885 ;
        RECT 82.335 118.075 82.845 118.610 ;
        RECT 83.025 118.245 83.215 119.605 ;
        RECT 83.385 118.585 83.660 119.405 ;
        RECT 83.865 118.805 84.035 119.605 ;
        RECT 84.205 118.815 84.375 119.945 ;
        RECT 84.545 119.315 84.715 120.285 ;
        RECT 84.885 119.485 85.055 120.625 ;
        RECT 85.225 119.485 85.560 120.455 ;
        RECT 84.545 118.985 84.740 119.315 ;
        RECT 84.965 118.985 85.220 119.315 ;
        RECT 84.965 118.815 85.135 118.985 ;
        RECT 85.390 118.815 85.560 119.485 ;
        RECT 85.735 119.535 86.945 120.625 ;
        RECT 87.490 119.645 87.745 120.315 ;
        RECT 87.925 119.825 88.210 120.625 ;
        RECT 88.390 119.905 88.720 120.415 ;
        RECT 85.735 118.995 86.255 119.535 ;
        RECT 86.425 118.825 86.945 119.365 ;
        RECT 87.490 119.265 87.670 119.645 ;
        RECT 88.390 119.315 88.640 119.905 ;
        RECT 88.990 119.755 89.160 120.365 ;
        RECT 89.330 119.935 89.660 120.625 ;
        RECT 89.890 120.075 90.130 120.365 ;
        RECT 90.330 120.245 90.750 120.625 ;
        RECT 90.930 120.155 91.560 120.405 ;
        RECT 92.030 120.245 92.360 120.625 ;
        RECT 90.930 120.075 91.100 120.155 ;
        RECT 92.530 120.075 92.700 120.365 ;
        RECT 92.880 120.245 93.260 120.625 ;
        RECT 93.500 120.240 94.330 120.410 ;
        RECT 89.890 119.905 91.100 120.075 ;
        RECT 87.405 119.095 87.670 119.265 ;
        RECT 84.205 118.645 85.135 118.815 ;
        RECT 84.205 118.610 84.380 118.645 ;
        RECT 83.385 118.415 83.665 118.585 ;
        RECT 83.385 118.245 83.660 118.415 ;
        RECT 83.850 118.245 84.380 118.610 ;
        RECT 84.805 118.075 85.135 118.475 ;
        RECT 85.305 118.245 85.560 118.815 ;
        RECT 85.735 118.075 86.945 118.825 ;
        RECT 87.490 118.785 87.670 119.095 ;
        RECT 87.840 118.985 88.640 119.315 ;
        RECT 87.490 118.255 87.745 118.785 ;
        RECT 87.925 118.075 88.210 118.535 ;
        RECT 88.390 118.335 88.640 118.985 ;
        RECT 88.840 119.735 89.160 119.755 ;
        RECT 88.840 119.565 90.760 119.735 ;
        RECT 88.840 118.670 89.030 119.565 ;
        RECT 90.930 119.395 91.100 119.905 ;
        RECT 91.270 119.645 91.790 119.955 ;
        RECT 89.200 119.225 91.100 119.395 ;
        RECT 89.200 119.165 89.530 119.225 ;
        RECT 89.680 118.995 90.010 119.055 ;
        RECT 89.350 118.725 90.010 118.995 ;
        RECT 88.840 118.340 89.160 118.670 ;
        RECT 89.340 118.075 90.000 118.555 ;
        RECT 90.200 118.465 90.370 119.225 ;
        RECT 91.270 119.055 91.450 119.465 ;
        RECT 90.540 118.885 90.870 119.005 ;
        RECT 91.620 118.885 91.790 119.645 ;
        RECT 90.540 118.715 91.790 118.885 ;
        RECT 91.960 119.825 93.330 120.075 ;
        RECT 91.960 119.055 92.150 119.825 ;
        RECT 93.080 119.565 93.330 119.825 ;
        RECT 92.320 119.395 92.570 119.555 ;
        RECT 93.500 119.395 93.670 120.240 ;
        RECT 94.565 119.955 94.735 120.455 ;
        RECT 94.905 120.125 95.235 120.625 ;
        RECT 93.840 119.565 94.340 119.945 ;
        RECT 94.565 119.785 95.260 119.955 ;
        RECT 92.320 119.225 93.670 119.395 ;
        RECT 93.250 119.185 93.670 119.225 ;
        RECT 91.960 118.715 92.380 119.055 ;
        RECT 92.670 118.725 93.080 119.055 ;
        RECT 90.200 118.295 91.050 118.465 ;
        RECT 91.610 118.075 91.930 118.535 ;
        RECT 92.130 118.285 92.380 118.715 ;
        RECT 92.670 118.075 93.080 118.515 ;
        RECT 93.250 118.455 93.420 119.185 ;
        RECT 93.590 118.635 93.940 119.005 ;
        RECT 94.120 118.695 94.340 119.565 ;
        RECT 94.510 118.995 94.920 119.615 ;
        RECT 95.090 118.815 95.260 119.785 ;
        RECT 94.565 118.625 95.260 118.815 ;
        RECT 93.250 118.255 94.265 118.455 ;
        RECT 94.565 118.295 94.735 118.625 ;
        RECT 94.905 118.075 95.235 118.455 ;
        RECT 95.450 118.335 95.675 120.455 ;
        RECT 95.845 120.125 96.175 120.625 ;
        RECT 96.345 119.955 96.515 120.455 ;
        RECT 95.850 119.785 96.515 119.955 ;
        RECT 95.850 118.795 96.080 119.785 ;
        RECT 96.250 118.965 96.600 119.615 ;
        RECT 96.775 119.535 97.985 120.625 ;
        RECT 98.155 119.865 98.670 120.275 ;
        RECT 98.905 119.865 99.075 120.625 ;
        RECT 99.245 120.285 101.275 120.455 ;
        RECT 96.775 118.995 97.295 119.535 ;
        RECT 97.465 118.825 97.985 119.365 ;
        RECT 98.155 119.055 98.495 119.865 ;
        RECT 99.245 119.620 99.415 120.285 ;
        RECT 99.810 119.945 100.935 120.115 ;
        RECT 98.665 119.430 99.415 119.620 ;
        RECT 99.585 119.605 100.595 119.775 ;
        RECT 98.155 118.885 99.385 119.055 ;
        RECT 95.850 118.625 96.515 118.795 ;
        RECT 95.845 118.075 96.175 118.455 ;
        RECT 96.345 118.335 96.515 118.625 ;
        RECT 96.775 118.075 97.985 118.825 ;
        RECT 98.430 118.280 98.675 118.885 ;
        RECT 98.895 118.075 99.405 118.610 ;
        RECT 99.585 118.245 99.775 119.605 ;
        RECT 99.945 119.265 100.220 119.405 ;
        RECT 99.945 119.095 100.225 119.265 ;
        RECT 99.945 118.245 100.220 119.095 ;
        RECT 100.425 118.805 100.595 119.605 ;
        RECT 100.765 118.815 100.935 119.945 ;
        RECT 101.105 119.315 101.275 120.285 ;
        RECT 101.445 119.485 101.615 120.625 ;
        RECT 101.785 119.485 102.120 120.455 ;
        RECT 101.105 118.985 101.300 119.315 ;
        RECT 101.525 118.985 101.780 119.315 ;
        RECT 101.525 118.815 101.695 118.985 ;
        RECT 101.950 118.815 102.120 119.485 ;
        RECT 103.215 119.460 103.505 120.625 ;
        RECT 104.050 119.645 104.305 120.315 ;
        RECT 104.485 119.825 104.770 120.625 ;
        RECT 104.950 119.905 105.280 120.415 ;
        RECT 104.050 119.605 104.230 119.645 ;
        RECT 103.965 119.435 104.230 119.605 ;
        RECT 100.765 118.645 101.695 118.815 ;
        RECT 100.765 118.610 100.940 118.645 ;
        RECT 100.410 118.245 100.940 118.610 ;
        RECT 101.365 118.075 101.695 118.475 ;
        RECT 101.865 118.245 102.120 118.815 ;
        RECT 103.215 118.075 103.505 118.800 ;
        RECT 104.050 118.785 104.230 119.435 ;
        RECT 104.950 119.315 105.200 119.905 ;
        RECT 105.550 119.755 105.720 120.365 ;
        RECT 105.890 119.935 106.220 120.625 ;
        RECT 106.450 120.075 106.690 120.365 ;
        RECT 106.890 120.245 107.310 120.625 ;
        RECT 107.490 120.155 108.120 120.405 ;
        RECT 108.590 120.245 108.920 120.625 ;
        RECT 107.490 120.075 107.660 120.155 ;
        RECT 109.090 120.075 109.260 120.365 ;
        RECT 109.440 120.245 109.820 120.625 ;
        RECT 110.060 120.240 110.890 120.410 ;
        RECT 106.450 119.905 107.660 120.075 ;
        RECT 104.400 118.985 105.200 119.315 ;
        RECT 104.050 118.255 104.305 118.785 ;
        RECT 104.485 118.075 104.770 118.535 ;
        RECT 104.950 118.335 105.200 118.985 ;
        RECT 105.400 119.735 105.720 119.755 ;
        RECT 105.400 119.565 107.320 119.735 ;
        RECT 105.400 118.670 105.590 119.565 ;
        RECT 107.490 119.395 107.660 119.905 ;
        RECT 107.830 119.645 108.350 119.955 ;
        RECT 105.760 119.225 107.660 119.395 ;
        RECT 105.760 119.165 106.090 119.225 ;
        RECT 106.240 118.995 106.570 119.055 ;
        RECT 105.910 118.725 106.570 118.995 ;
        RECT 105.400 118.340 105.720 118.670 ;
        RECT 105.900 118.075 106.560 118.555 ;
        RECT 106.760 118.465 106.930 119.225 ;
        RECT 107.830 119.055 108.010 119.465 ;
        RECT 107.100 118.885 107.430 119.005 ;
        RECT 108.180 118.885 108.350 119.645 ;
        RECT 107.100 118.715 108.350 118.885 ;
        RECT 108.520 119.825 109.890 120.075 ;
        RECT 108.520 119.055 108.710 119.825 ;
        RECT 109.640 119.565 109.890 119.825 ;
        RECT 108.880 119.395 109.130 119.555 ;
        RECT 110.060 119.395 110.230 120.240 ;
        RECT 111.125 119.955 111.295 120.455 ;
        RECT 111.465 120.125 111.795 120.625 ;
        RECT 110.400 119.565 110.900 119.945 ;
        RECT 111.125 119.785 111.820 119.955 ;
        RECT 108.880 119.225 110.230 119.395 ;
        RECT 109.810 119.185 110.230 119.225 ;
        RECT 108.520 118.715 108.940 119.055 ;
        RECT 109.230 118.725 109.640 119.055 ;
        RECT 106.760 118.295 107.610 118.465 ;
        RECT 108.170 118.075 108.490 118.535 ;
        RECT 108.690 118.285 108.940 118.715 ;
        RECT 109.230 118.075 109.640 118.515 ;
        RECT 109.810 118.455 109.980 119.185 ;
        RECT 110.150 118.635 110.500 119.005 ;
        RECT 110.680 118.695 110.900 119.565 ;
        RECT 111.070 118.995 111.480 119.615 ;
        RECT 111.650 118.815 111.820 119.785 ;
        RECT 111.125 118.625 111.820 118.815 ;
        RECT 109.810 118.255 110.825 118.455 ;
        RECT 111.125 118.295 111.295 118.625 ;
        RECT 111.465 118.075 111.795 118.455 ;
        RECT 112.010 118.335 112.235 120.455 ;
        RECT 112.405 120.125 112.735 120.625 ;
        RECT 112.905 119.955 113.075 120.455 ;
        RECT 112.410 119.785 113.075 119.955 ;
        RECT 112.410 118.795 112.640 119.785 ;
        RECT 112.810 118.965 113.160 119.615 ;
        RECT 113.795 119.535 115.465 120.625 ;
        RECT 115.635 119.865 116.150 120.275 ;
        RECT 116.385 119.865 116.555 120.625 ;
        RECT 116.725 120.285 118.755 120.455 ;
        RECT 113.795 119.015 114.545 119.535 ;
        RECT 114.715 118.845 115.465 119.365 ;
        RECT 115.635 119.055 115.975 119.865 ;
        RECT 116.725 119.620 116.895 120.285 ;
        RECT 117.290 119.945 118.415 120.115 ;
        RECT 116.145 119.430 116.895 119.620 ;
        RECT 117.065 119.605 118.075 119.775 ;
        RECT 115.635 118.885 116.865 119.055 ;
        RECT 112.410 118.625 113.075 118.795 ;
        RECT 112.405 118.075 112.735 118.455 ;
        RECT 112.905 118.335 113.075 118.625 ;
        RECT 113.795 118.075 115.465 118.845 ;
        RECT 115.910 118.280 116.155 118.885 ;
        RECT 116.375 118.075 116.885 118.610 ;
        RECT 117.065 118.245 117.255 119.605 ;
        RECT 117.425 119.265 117.700 119.405 ;
        RECT 117.425 119.095 117.705 119.265 ;
        RECT 117.425 118.245 117.700 119.095 ;
        RECT 117.905 118.805 118.075 119.605 ;
        RECT 118.245 118.815 118.415 119.945 ;
        RECT 118.585 119.315 118.755 120.285 ;
        RECT 118.925 119.485 119.095 120.625 ;
        RECT 119.265 119.485 119.600 120.455 ;
        RECT 120.275 119.485 120.505 120.625 ;
        RECT 118.585 118.985 118.780 119.315 ;
        RECT 119.005 118.985 119.260 119.315 ;
        RECT 119.005 118.815 119.175 118.985 ;
        RECT 119.430 118.815 119.600 119.485 ;
        RECT 120.675 119.475 121.005 120.455 ;
        RECT 121.175 119.485 121.385 120.625 ;
        RECT 121.705 119.695 121.875 120.455 ;
        RECT 122.055 119.865 122.385 120.625 ;
        RECT 121.705 119.525 122.370 119.695 ;
        RECT 122.555 119.550 122.825 120.455 ;
        RECT 120.255 119.065 120.585 119.315 ;
        RECT 118.245 118.645 119.175 118.815 ;
        RECT 118.245 118.610 118.420 118.645 ;
        RECT 117.890 118.245 118.420 118.610 ;
        RECT 118.845 118.075 119.175 118.475 ;
        RECT 119.345 118.245 119.600 118.815 ;
        RECT 120.275 118.075 120.505 118.895 ;
        RECT 120.755 118.875 121.005 119.475 ;
        RECT 122.200 119.380 122.370 119.525 ;
        RECT 121.635 118.975 121.965 119.345 ;
        RECT 122.200 119.050 122.485 119.380 ;
        RECT 120.675 118.245 121.005 118.875 ;
        RECT 121.175 118.075 121.385 118.895 ;
        RECT 122.200 118.795 122.370 119.050 ;
        RECT 121.705 118.625 122.370 118.795 ;
        RECT 122.655 118.750 122.825 119.550 ;
        RECT 122.995 119.535 124.205 120.625 ;
        RECT 124.375 119.535 127.885 120.625 ;
        RECT 128.055 119.535 129.265 120.625 ;
        RECT 122.995 118.995 123.515 119.535 ;
        RECT 123.685 118.825 124.205 119.365 ;
        RECT 124.375 119.015 126.065 119.535 ;
        RECT 126.235 118.845 127.885 119.365 ;
        RECT 128.055 118.995 128.575 119.535 ;
        RECT 121.705 118.245 121.875 118.625 ;
        RECT 122.055 118.075 122.385 118.455 ;
        RECT 122.565 118.245 122.825 118.750 ;
        RECT 122.995 118.075 124.205 118.825 ;
        RECT 124.375 118.075 127.885 118.845 ;
        RECT 128.745 118.825 129.265 119.365 ;
        RECT 128.055 118.075 129.265 118.825 ;
        RECT 9.290 117.905 129.350 118.075 ;
        RECT 9.375 117.155 10.585 117.905 ;
        RECT 9.375 116.615 9.895 117.155 ;
        RECT 11.215 117.135 12.885 117.905 ;
        RECT 13.055 117.180 13.345 117.905 ;
        RECT 10.065 116.445 10.585 116.985 ;
        RECT 9.375 115.355 10.585 116.445 ;
        RECT 11.215 116.445 11.965 116.965 ;
        RECT 12.135 116.615 12.885 117.135 ;
        RECT 13.555 117.085 13.785 117.905 ;
        RECT 13.955 117.105 14.285 117.735 ;
        RECT 13.535 116.665 13.865 116.915 ;
        RECT 11.215 115.355 12.885 116.445 ;
        RECT 13.055 115.355 13.345 116.520 ;
        RECT 14.035 116.505 14.285 117.105 ;
        RECT 14.455 117.085 14.665 117.905 ;
        RECT 15.270 117.565 15.525 117.725 ;
        RECT 15.185 117.395 15.525 117.565 ;
        RECT 15.705 117.445 15.990 117.905 ;
        RECT 15.270 117.195 15.525 117.395 ;
        RECT 13.555 115.355 13.785 116.495 ;
        RECT 13.955 115.525 14.285 116.505 ;
        RECT 14.455 115.355 14.665 116.495 ;
        RECT 15.270 116.335 15.450 117.195 ;
        RECT 16.170 116.995 16.420 117.645 ;
        RECT 15.620 116.665 16.420 116.995 ;
        RECT 15.270 115.665 15.525 116.335 ;
        RECT 15.705 115.355 15.990 116.155 ;
        RECT 16.170 116.075 16.420 116.665 ;
        RECT 16.620 117.310 16.940 117.640 ;
        RECT 17.120 117.425 17.780 117.905 ;
        RECT 17.980 117.515 18.830 117.685 ;
        RECT 16.620 116.415 16.810 117.310 ;
        RECT 17.130 116.985 17.790 117.255 ;
        RECT 17.460 116.925 17.790 116.985 ;
        RECT 16.980 116.755 17.310 116.815 ;
        RECT 17.980 116.755 18.150 117.515 ;
        RECT 19.390 117.445 19.710 117.905 ;
        RECT 19.910 117.265 20.160 117.695 ;
        RECT 20.450 117.465 20.860 117.905 ;
        RECT 21.030 117.525 22.045 117.725 ;
        RECT 18.320 117.095 19.570 117.265 ;
        RECT 18.320 116.975 18.650 117.095 ;
        RECT 16.980 116.585 18.880 116.755 ;
        RECT 16.620 116.245 18.540 116.415 ;
        RECT 16.620 116.225 16.940 116.245 ;
        RECT 16.170 115.565 16.500 116.075 ;
        RECT 16.770 115.615 16.940 116.225 ;
        RECT 18.710 116.075 18.880 116.585 ;
        RECT 19.050 116.515 19.230 116.925 ;
        RECT 19.400 116.335 19.570 117.095 ;
        RECT 17.110 115.355 17.440 116.045 ;
        RECT 17.670 115.905 18.880 116.075 ;
        RECT 19.050 116.025 19.570 116.335 ;
        RECT 19.740 116.925 20.160 117.265 ;
        RECT 20.450 116.925 20.860 117.255 ;
        RECT 19.740 116.155 19.930 116.925 ;
        RECT 21.030 116.795 21.200 117.525 ;
        RECT 22.345 117.355 22.515 117.685 ;
        RECT 22.685 117.525 23.015 117.905 ;
        RECT 21.370 116.975 21.720 117.345 ;
        RECT 21.030 116.755 21.450 116.795 ;
        RECT 20.100 116.585 21.450 116.755 ;
        RECT 20.100 116.425 20.350 116.585 ;
        RECT 20.860 116.155 21.110 116.415 ;
        RECT 19.740 115.905 21.110 116.155 ;
        RECT 17.670 115.615 17.910 115.905 ;
        RECT 18.710 115.825 18.880 115.905 ;
        RECT 18.110 115.355 18.530 115.735 ;
        RECT 18.710 115.575 19.340 115.825 ;
        RECT 19.810 115.355 20.140 115.735 ;
        RECT 20.310 115.615 20.480 115.905 ;
        RECT 21.280 115.740 21.450 116.585 ;
        RECT 21.900 116.415 22.120 117.285 ;
        RECT 22.345 117.165 23.040 117.355 ;
        RECT 21.620 116.035 22.120 116.415 ;
        RECT 22.290 116.365 22.700 116.985 ;
        RECT 22.870 116.195 23.040 117.165 ;
        RECT 22.345 116.025 23.040 116.195 ;
        RECT 20.660 115.355 21.040 115.735 ;
        RECT 21.280 115.570 22.110 115.740 ;
        RECT 22.345 115.525 22.515 116.025 ;
        RECT 22.685 115.355 23.015 115.855 ;
        RECT 23.230 115.525 23.455 117.645 ;
        RECT 23.625 117.525 23.955 117.905 ;
        RECT 24.125 117.355 24.295 117.645 ;
        RECT 24.930 117.565 25.185 117.725 ;
        RECT 24.845 117.395 25.185 117.565 ;
        RECT 25.365 117.445 25.650 117.905 ;
        RECT 23.630 117.185 24.295 117.355 ;
        RECT 24.930 117.195 25.185 117.395 ;
        RECT 23.630 116.195 23.860 117.185 ;
        RECT 24.030 116.365 24.380 117.015 ;
        RECT 24.930 116.335 25.110 117.195 ;
        RECT 25.830 116.995 26.080 117.645 ;
        RECT 25.280 116.665 26.080 116.995 ;
        RECT 23.630 116.025 24.295 116.195 ;
        RECT 23.625 115.355 23.955 115.855 ;
        RECT 24.125 115.525 24.295 116.025 ;
        RECT 24.930 115.665 25.185 116.335 ;
        RECT 25.365 115.355 25.650 116.155 ;
        RECT 25.830 116.075 26.080 116.665 ;
        RECT 26.280 117.310 26.600 117.640 ;
        RECT 26.780 117.425 27.440 117.905 ;
        RECT 27.640 117.515 28.490 117.685 ;
        RECT 26.280 116.415 26.470 117.310 ;
        RECT 26.790 116.985 27.450 117.255 ;
        RECT 27.120 116.925 27.450 116.985 ;
        RECT 26.640 116.755 26.970 116.815 ;
        RECT 27.640 116.755 27.810 117.515 ;
        RECT 29.050 117.445 29.370 117.905 ;
        RECT 29.570 117.265 29.820 117.695 ;
        RECT 30.110 117.465 30.520 117.905 ;
        RECT 30.690 117.525 31.705 117.725 ;
        RECT 27.980 117.095 29.230 117.265 ;
        RECT 27.980 116.975 28.310 117.095 ;
        RECT 26.640 116.585 28.540 116.755 ;
        RECT 26.280 116.245 28.200 116.415 ;
        RECT 26.280 116.225 26.600 116.245 ;
        RECT 25.830 115.565 26.160 116.075 ;
        RECT 26.430 115.615 26.600 116.225 ;
        RECT 28.370 116.075 28.540 116.585 ;
        RECT 28.710 116.515 28.890 116.925 ;
        RECT 29.060 116.335 29.230 117.095 ;
        RECT 26.770 115.355 27.100 116.045 ;
        RECT 27.330 115.905 28.540 116.075 ;
        RECT 28.710 116.025 29.230 116.335 ;
        RECT 29.400 116.925 29.820 117.265 ;
        RECT 30.110 116.925 30.520 117.255 ;
        RECT 29.400 116.155 29.590 116.925 ;
        RECT 30.690 116.795 30.860 117.525 ;
        RECT 32.005 117.355 32.175 117.685 ;
        RECT 32.345 117.525 32.675 117.905 ;
        RECT 31.030 116.975 31.380 117.345 ;
        RECT 30.690 116.755 31.110 116.795 ;
        RECT 29.760 116.585 31.110 116.755 ;
        RECT 29.760 116.425 30.010 116.585 ;
        RECT 30.520 116.155 30.770 116.415 ;
        RECT 29.400 115.905 30.770 116.155 ;
        RECT 27.330 115.615 27.570 115.905 ;
        RECT 28.370 115.825 28.540 115.905 ;
        RECT 27.770 115.355 28.190 115.735 ;
        RECT 28.370 115.575 29.000 115.825 ;
        RECT 29.470 115.355 29.800 115.735 ;
        RECT 29.970 115.615 30.140 115.905 ;
        RECT 30.940 115.740 31.110 116.585 ;
        RECT 31.560 116.415 31.780 117.285 ;
        RECT 32.005 117.165 32.700 117.355 ;
        RECT 31.280 116.035 31.780 116.415 ;
        RECT 31.950 116.365 32.360 116.985 ;
        RECT 32.530 116.195 32.700 117.165 ;
        RECT 32.005 116.025 32.700 116.195 ;
        RECT 30.320 115.355 30.700 115.735 ;
        RECT 30.940 115.570 31.770 115.740 ;
        RECT 32.005 115.525 32.175 116.025 ;
        RECT 32.345 115.355 32.675 115.855 ;
        RECT 32.890 115.525 33.115 117.645 ;
        RECT 33.285 117.525 33.615 117.905 ;
        RECT 33.785 117.355 33.955 117.645 ;
        RECT 33.290 117.185 33.955 117.355 ;
        RECT 33.290 116.195 33.520 117.185 ;
        RECT 35.175 117.085 35.405 117.905 ;
        RECT 35.575 117.105 35.905 117.735 ;
        RECT 33.690 116.365 34.040 117.015 ;
        RECT 35.155 116.665 35.485 116.915 ;
        RECT 35.655 116.505 35.905 117.105 ;
        RECT 36.075 117.085 36.285 117.905 ;
        RECT 36.975 117.135 38.645 117.905 ;
        RECT 38.815 117.180 39.105 117.905 ;
        RECT 39.275 117.155 40.485 117.905 ;
        RECT 33.290 116.025 33.955 116.195 ;
        RECT 33.285 115.355 33.615 115.855 ;
        RECT 33.785 115.525 33.955 116.025 ;
        RECT 35.175 115.355 35.405 116.495 ;
        RECT 35.575 115.525 35.905 116.505 ;
        RECT 36.075 115.355 36.285 116.495 ;
        RECT 36.975 116.445 37.725 116.965 ;
        RECT 37.895 116.615 38.645 117.135 ;
        RECT 36.975 115.355 38.645 116.445 ;
        RECT 38.815 115.355 39.105 116.520 ;
        RECT 39.275 116.445 39.795 116.985 ;
        RECT 39.965 116.615 40.485 117.155 ;
        RECT 40.655 117.230 40.915 117.735 ;
        RECT 41.095 117.525 41.425 117.905 ;
        RECT 41.605 117.355 41.775 117.735 ;
        RECT 42.960 117.360 48.305 117.905 ;
        RECT 39.275 115.355 40.485 116.445 ;
        RECT 40.655 116.430 40.825 117.230 ;
        RECT 41.110 117.185 41.775 117.355 ;
        RECT 41.110 116.930 41.280 117.185 ;
        RECT 40.995 116.600 41.280 116.930 ;
        RECT 41.515 116.635 41.845 117.005 ;
        RECT 41.110 116.455 41.280 116.600 ;
        RECT 40.655 115.525 40.925 116.430 ;
        RECT 41.110 116.285 41.775 116.455 ;
        RECT 41.095 115.355 41.425 116.115 ;
        RECT 41.605 115.525 41.775 116.285 ;
        RECT 44.550 115.790 44.900 117.040 ;
        RECT 46.380 116.530 46.720 117.360 ;
        RECT 48.515 117.085 48.745 117.905 ;
        RECT 48.915 117.105 49.245 117.735 ;
        RECT 48.495 116.665 48.825 116.915 ;
        RECT 48.995 116.505 49.245 117.105 ;
        RECT 49.415 117.085 49.625 117.905 ;
        RECT 50.130 117.095 50.375 117.700 ;
        RECT 50.595 117.370 51.105 117.905 ;
        RECT 42.960 115.355 48.305 115.790 ;
        RECT 48.515 115.355 48.745 116.495 ;
        RECT 48.915 115.525 49.245 116.505 ;
        RECT 49.855 116.925 51.085 117.095 ;
        RECT 49.415 115.355 49.625 116.495 ;
        RECT 49.855 116.115 50.195 116.925 ;
        RECT 50.365 116.360 51.115 116.550 ;
        RECT 49.855 115.705 50.370 116.115 ;
        RECT 50.605 115.355 50.775 116.115 ;
        RECT 50.945 115.695 51.115 116.360 ;
        RECT 51.285 116.375 51.475 117.735 ;
        RECT 51.645 116.885 51.920 117.735 ;
        RECT 52.110 117.370 52.640 117.735 ;
        RECT 53.065 117.505 53.395 117.905 ;
        RECT 52.465 117.335 52.640 117.370 ;
        RECT 51.645 116.715 51.925 116.885 ;
        RECT 51.645 116.575 51.920 116.715 ;
        RECT 52.125 116.375 52.295 117.175 ;
        RECT 51.285 116.205 52.295 116.375 ;
        RECT 52.465 117.165 53.395 117.335 ;
        RECT 53.565 117.165 53.820 117.735 ;
        RECT 54.085 117.355 54.255 117.735 ;
        RECT 54.435 117.525 54.765 117.905 ;
        RECT 54.085 117.185 54.750 117.355 ;
        RECT 54.945 117.230 55.205 117.735 ;
        RECT 52.465 116.035 52.635 117.165 ;
        RECT 53.225 116.995 53.395 117.165 ;
        RECT 51.510 115.865 52.635 116.035 ;
        RECT 52.805 116.665 53.000 116.995 ;
        RECT 53.225 116.665 53.480 116.995 ;
        RECT 52.805 115.695 52.975 116.665 ;
        RECT 53.650 116.495 53.820 117.165 ;
        RECT 54.015 116.635 54.345 117.005 ;
        RECT 54.580 116.930 54.750 117.185 ;
        RECT 50.945 115.525 52.975 115.695 ;
        RECT 53.145 115.355 53.315 116.495 ;
        RECT 53.485 115.525 53.820 116.495 ;
        RECT 54.580 116.600 54.865 116.930 ;
        RECT 54.580 116.455 54.750 116.600 ;
        RECT 54.085 116.285 54.750 116.455 ;
        RECT 55.035 116.430 55.205 117.230 ;
        RECT 55.525 117.105 55.855 117.905 ;
        RECT 56.025 117.255 56.195 117.735 ;
        RECT 56.365 117.425 56.695 117.905 ;
        RECT 56.865 117.255 57.035 117.735 ;
        RECT 57.285 117.425 57.525 117.905 ;
        RECT 57.705 117.255 57.875 117.735 ;
        RECT 56.025 117.085 57.035 117.255 ;
        RECT 57.240 117.085 57.875 117.255 ;
        RECT 59.055 117.135 62.565 117.905 ;
        RECT 56.025 116.545 56.520 117.085 ;
        RECT 57.240 116.915 57.410 117.085 ;
        RECT 56.910 116.745 57.410 116.915 ;
        RECT 54.085 115.525 54.255 116.285 ;
        RECT 54.435 115.355 54.765 116.115 ;
        RECT 54.935 115.525 55.205 116.430 ;
        RECT 55.525 115.355 55.855 116.505 ;
        RECT 56.025 116.375 57.035 116.545 ;
        RECT 56.025 115.525 56.195 116.375 ;
        RECT 56.365 115.355 56.695 116.155 ;
        RECT 56.865 115.525 57.035 116.375 ;
        RECT 57.240 116.505 57.410 116.745 ;
        RECT 57.580 116.675 57.960 116.915 ;
        RECT 57.240 116.335 57.955 116.505 ;
        RECT 57.215 115.355 57.455 116.155 ;
        RECT 57.625 115.525 57.955 116.335 ;
        RECT 59.055 116.445 60.745 116.965 ;
        RECT 60.915 116.615 62.565 117.135 ;
        RECT 62.775 117.085 63.005 117.905 ;
        RECT 63.175 117.105 63.505 117.735 ;
        RECT 62.755 116.665 63.085 116.915 ;
        RECT 63.255 116.505 63.505 117.105 ;
        RECT 63.675 117.085 63.885 117.905 ;
        RECT 64.575 117.180 64.865 117.905 ;
        RECT 65.960 117.360 71.305 117.905 ;
        RECT 59.055 115.355 62.565 116.445 ;
        RECT 62.775 115.355 63.005 116.495 ;
        RECT 63.175 115.525 63.505 116.505 ;
        RECT 63.675 115.355 63.885 116.495 ;
        RECT 64.575 115.355 64.865 116.520 ;
        RECT 67.550 115.790 67.900 117.040 ;
        RECT 69.380 116.530 69.720 117.360 ;
        RECT 71.850 117.195 72.105 117.725 ;
        RECT 72.285 117.445 72.570 117.905 ;
        RECT 71.850 116.545 72.030 117.195 ;
        RECT 72.750 116.995 73.000 117.645 ;
        RECT 72.200 116.665 73.000 116.995 ;
        RECT 71.765 116.375 72.030 116.545 ;
        RECT 71.850 116.335 72.030 116.375 ;
        RECT 65.960 115.355 71.305 115.790 ;
        RECT 71.850 115.665 72.105 116.335 ;
        RECT 72.285 115.355 72.570 116.155 ;
        RECT 72.750 116.075 73.000 116.665 ;
        RECT 73.200 117.310 73.520 117.640 ;
        RECT 73.700 117.425 74.360 117.905 ;
        RECT 74.560 117.515 75.410 117.685 ;
        RECT 73.200 116.415 73.390 117.310 ;
        RECT 73.710 116.985 74.370 117.255 ;
        RECT 74.040 116.925 74.370 116.985 ;
        RECT 73.560 116.755 73.890 116.815 ;
        RECT 74.560 116.755 74.730 117.515 ;
        RECT 75.970 117.445 76.290 117.905 ;
        RECT 76.490 117.265 76.740 117.695 ;
        RECT 77.030 117.465 77.440 117.905 ;
        RECT 77.610 117.525 78.625 117.725 ;
        RECT 74.900 117.095 76.150 117.265 ;
        RECT 74.900 116.975 75.230 117.095 ;
        RECT 73.560 116.585 75.460 116.755 ;
        RECT 73.200 116.245 75.120 116.415 ;
        RECT 73.200 116.225 73.520 116.245 ;
        RECT 72.750 115.565 73.080 116.075 ;
        RECT 73.350 115.615 73.520 116.225 ;
        RECT 75.290 116.075 75.460 116.585 ;
        RECT 75.630 116.515 75.810 116.925 ;
        RECT 75.980 116.335 76.150 117.095 ;
        RECT 73.690 115.355 74.020 116.045 ;
        RECT 74.250 115.905 75.460 116.075 ;
        RECT 75.630 116.025 76.150 116.335 ;
        RECT 76.320 116.925 76.740 117.265 ;
        RECT 77.030 116.925 77.440 117.255 ;
        RECT 76.320 116.155 76.510 116.925 ;
        RECT 77.610 116.795 77.780 117.525 ;
        RECT 78.925 117.355 79.095 117.685 ;
        RECT 79.265 117.525 79.595 117.905 ;
        RECT 77.950 116.975 78.300 117.345 ;
        RECT 77.610 116.755 78.030 116.795 ;
        RECT 76.680 116.585 78.030 116.755 ;
        RECT 76.680 116.425 76.930 116.585 ;
        RECT 77.440 116.155 77.690 116.415 ;
        RECT 76.320 115.905 77.690 116.155 ;
        RECT 74.250 115.615 74.490 115.905 ;
        RECT 75.290 115.825 75.460 115.905 ;
        RECT 74.690 115.355 75.110 115.735 ;
        RECT 75.290 115.575 75.920 115.825 ;
        RECT 76.390 115.355 76.720 115.735 ;
        RECT 76.890 115.615 77.060 115.905 ;
        RECT 77.860 115.740 78.030 116.585 ;
        RECT 78.480 116.415 78.700 117.285 ;
        RECT 78.925 117.165 79.620 117.355 ;
        RECT 78.200 116.035 78.700 116.415 ;
        RECT 78.870 116.365 79.280 116.985 ;
        RECT 79.450 116.195 79.620 117.165 ;
        RECT 78.925 116.025 79.620 116.195 ;
        RECT 77.240 115.355 77.620 115.735 ;
        RECT 77.860 115.570 78.690 115.740 ;
        RECT 78.925 115.525 79.095 116.025 ;
        RECT 79.265 115.355 79.595 115.855 ;
        RECT 79.810 115.525 80.035 117.645 ;
        RECT 80.205 117.525 80.535 117.905 ;
        RECT 80.705 117.355 80.875 117.645 ;
        RECT 80.210 117.185 80.875 117.355 ;
        RECT 80.210 116.195 80.440 117.185 ;
        RECT 81.140 117.165 81.395 117.735 ;
        RECT 81.565 117.505 81.895 117.905 ;
        RECT 82.320 117.370 82.850 117.735 ;
        RECT 83.040 117.565 83.315 117.735 ;
        RECT 83.035 117.395 83.315 117.565 ;
        RECT 82.320 117.335 82.495 117.370 ;
        RECT 81.565 117.165 82.495 117.335 ;
        RECT 80.610 116.365 80.960 117.015 ;
        RECT 81.140 116.495 81.310 117.165 ;
        RECT 81.565 116.995 81.735 117.165 ;
        RECT 81.480 116.665 81.735 116.995 ;
        RECT 81.960 116.665 82.155 116.995 ;
        RECT 80.210 116.025 80.875 116.195 ;
        RECT 80.205 115.355 80.535 115.855 ;
        RECT 80.705 115.525 80.875 116.025 ;
        RECT 81.140 115.525 81.475 116.495 ;
        RECT 81.645 115.355 81.815 116.495 ;
        RECT 81.985 115.695 82.155 116.665 ;
        RECT 82.325 116.035 82.495 117.165 ;
        RECT 82.665 116.375 82.835 117.175 ;
        RECT 83.040 116.575 83.315 117.395 ;
        RECT 83.485 116.375 83.675 117.735 ;
        RECT 83.855 117.370 84.365 117.905 ;
        RECT 84.585 117.095 84.830 117.700 ;
        RECT 86.470 117.095 86.715 117.700 ;
        RECT 86.935 117.370 87.445 117.905 ;
        RECT 83.875 116.925 85.105 117.095 ;
        RECT 82.665 116.205 83.675 116.375 ;
        RECT 83.845 116.360 84.595 116.550 ;
        RECT 82.325 115.865 83.450 116.035 ;
        RECT 83.845 115.695 84.015 116.360 ;
        RECT 84.765 116.115 85.105 116.925 ;
        RECT 81.985 115.525 84.015 115.695 ;
        RECT 84.185 115.355 84.355 116.115 ;
        RECT 84.590 115.705 85.105 116.115 ;
        RECT 86.195 116.925 87.425 117.095 ;
        RECT 86.195 116.115 86.535 116.925 ;
        RECT 86.705 116.360 87.455 116.550 ;
        RECT 86.195 115.705 86.710 116.115 ;
        RECT 86.945 115.355 87.115 116.115 ;
        RECT 87.285 115.695 87.455 116.360 ;
        RECT 87.625 116.375 87.815 117.735 ;
        RECT 87.985 117.225 88.260 117.735 ;
        RECT 88.450 117.370 88.980 117.735 ;
        RECT 89.405 117.505 89.735 117.905 ;
        RECT 88.805 117.335 88.980 117.370 ;
        RECT 87.985 117.055 88.265 117.225 ;
        RECT 87.985 116.575 88.260 117.055 ;
        RECT 88.465 116.375 88.635 117.175 ;
        RECT 87.625 116.205 88.635 116.375 ;
        RECT 88.805 117.165 89.735 117.335 ;
        RECT 89.905 117.165 90.160 117.735 ;
        RECT 90.335 117.180 90.625 117.905 ;
        RECT 92.090 117.565 92.345 117.725 ;
        RECT 92.005 117.395 92.345 117.565 ;
        RECT 92.525 117.445 92.810 117.905 ;
        RECT 92.090 117.195 92.345 117.395 ;
        RECT 88.805 116.035 88.975 117.165 ;
        RECT 89.565 116.995 89.735 117.165 ;
        RECT 87.850 115.865 88.975 116.035 ;
        RECT 89.145 116.665 89.340 116.995 ;
        RECT 89.565 116.665 89.820 116.995 ;
        RECT 89.145 115.695 89.315 116.665 ;
        RECT 89.990 116.495 90.160 117.165 ;
        RECT 87.285 115.525 89.315 115.695 ;
        RECT 89.485 115.355 89.655 116.495 ;
        RECT 89.825 115.525 90.160 116.495 ;
        RECT 90.335 115.355 90.625 116.520 ;
        RECT 92.090 116.335 92.270 117.195 ;
        RECT 92.990 116.995 93.240 117.645 ;
        RECT 92.440 116.665 93.240 116.995 ;
        RECT 92.090 115.665 92.345 116.335 ;
        RECT 92.525 115.355 92.810 116.155 ;
        RECT 92.990 116.075 93.240 116.665 ;
        RECT 93.440 117.310 93.760 117.640 ;
        RECT 93.940 117.425 94.600 117.905 ;
        RECT 94.800 117.515 95.650 117.685 ;
        RECT 93.440 116.415 93.630 117.310 ;
        RECT 93.950 116.985 94.610 117.255 ;
        RECT 94.280 116.925 94.610 116.985 ;
        RECT 93.800 116.755 94.130 116.815 ;
        RECT 94.800 116.755 94.970 117.515 ;
        RECT 96.210 117.445 96.530 117.905 ;
        RECT 96.730 117.265 96.980 117.695 ;
        RECT 97.270 117.465 97.680 117.905 ;
        RECT 97.850 117.525 98.865 117.725 ;
        RECT 95.140 117.095 96.390 117.265 ;
        RECT 95.140 116.975 95.470 117.095 ;
        RECT 93.800 116.585 95.700 116.755 ;
        RECT 93.440 116.245 95.360 116.415 ;
        RECT 93.440 116.225 93.760 116.245 ;
        RECT 92.990 115.565 93.320 116.075 ;
        RECT 93.590 115.615 93.760 116.225 ;
        RECT 95.530 116.075 95.700 116.585 ;
        RECT 95.870 116.515 96.050 116.925 ;
        RECT 96.220 116.335 96.390 117.095 ;
        RECT 93.930 115.355 94.260 116.045 ;
        RECT 94.490 115.905 95.700 116.075 ;
        RECT 95.870 116.025 96.390 116.335 ;
        RECT 96.560 116.925 96.980 117.265 ;
        RECT 97.270 116.925 97.680 117.255 ;
        RECT 96.560 116.155 96.750 116.925 ;
        RECT 97.850 116.795 98.020 117.525 ;
        RECT 99.165 117.355 99.335 117.685 ;
        RECT 99.505 117.525 99.835 117.905 ;
        RECT 98.190 116.975 98.540 117.345 ;
        RECT 97.850 116.755 98.270 116.795 ;
        RECT 96.920 116.585 98.270 116.755 ;
        RECT 96.920 116.425 97.170 116.585 ;
        RECT 97.680 116.155 97.930 116.415 ;
        RECT 96.560 115.905 97.930 116.155 ;
        RECT 94.490 115.615 94.730 115.905 ;
        RECT 95.530 115.825 95.700 115.905 ;
        RECT 94.930 115.355 95.350 115.735 ;
        RECT 95.530 115.575 96.160 115.825 ;
        RECT 96.630 115.355 96.960 115.735 ;
        RECT 97.130 115.615 97.300 115.905 ;
        RECT 98.100 115.740 98.270 116.585 ;
        RECT 98.720 116.415 98.940 117.285 ;
        RECT 99.165 117.165 99.860 117.355 ;
        RECT 98.440 116.035 98.940 116.415 ;
        RECT 99.110 116.365 99.520 116.985 ;
        RECT 99.690 116.195 99.860 117.165 ;
        RECT 99.165 116.025 99.860 116.195 ;
        RECT 97.480 115.355 97.860 115.735 ;
        RECT 98.100 115.570 98.930 115.740 ;
        RECT 99.165 115.525 99.335 116.025 ;
        RECT 99.505 115.355 99.835 115.855 ;
        RECT 100.050 115.525 100.275 117.645 ;
        RECT 100.445 117.525 100.775 117.905 ;
        RECT 100.945 117.355 101.115 117.645 ;
        RECT 100.450 117.185 101.115 117.355 ;
        RECT 101.375 117.230 101.635 117.735 ;
        RECT 101.815 117.525 102.145 117.905 ;
        RECT 102.325 117.355 102.495 117.735 ;
        RECT 100.450 116.195 100.680 117.185 ;
        RECT 100.850 116.365 101.200 117.015 ;
        RECT 101.375 116.430 101.545 117.230 ;
        RECT 101.830 117.185 102.495 117.355 ;
        RECT 101.830 116.930 102.000 117.185 ;
        RECT 103.675 117.135 107.185 117.905 ;
        RECT 101.715 116.600 102.000 116.930 ;
        RECT 102.235 116.635 102.565 117.005 ;
        RECT 101.830 116.455 102.000 116.600 ;
        RECT 100.450 116.025 101.115 116.195 ;
        RECT 100.445 115.355 100.775 115.855 ;
        RECT 100.945 115.525 101.115 116.025 ;
        RECT 101.375 115.525 101.645 116.430 ;
        RECT 101.830 116.285 102.495 116.455 ;
        RECT 101.815 115.355 102.145 116.115 ;
        RECT 102.325 115.525 102.495 116.285 ;
        RECT 103.675 116.445 105.365 116.965 ;
        RECT 105.535 116.615 107.185 117.135 ;
        RECT 107.355 117.230 107.615 117.735 ;
        RECT 107.795 117.525 108.125 117.905 ;
        RECT 108.305 117.355 108.475 117.735 ;
        RECT 103.675 115.355 107.185 116.445 ;
        RECT 107.355 116.430 107.525 117.230 ;
        RECT 107.810 117.185 108.475 117.355 ;
        RECT 108.825 117.355 108.995 117.735 ;
        RECT 109.175 117.525 109.505 117.905 ;
        RECT 108.825 117.185 109.490 117.355 ;
        RECT 109.685 117.230 109.945 117.735 ;
        RECT 110.580 117.360 115.925 117.905 ;
        RECT 107.810 116.930 107.980 117.185 ;
        RECT 107.695 116.600 107.980 116.930 ;
        RECT 108.215 116.635 108.545 117.005 ;
        RECT 108.755 116.635 109.085 117.005 ;
        RECT 109.320 116.930 109.490 117.185 ;
        RECT 107.810 116.455 107.980 116.600 ;
        RECT 109.320 116.600 109.605 116.930 ;
        RECT 109.320 116.455 109.490 116.600 ;
        RECT 107.355 115.525 107.625 116.430 ;
        RECT 107.810 116.285 108.475 116.455 ;
        RECT 107.795 115.355 108.125 116.115 ;
        RECT 108.305 115.525 108.475 116.285 ;
        RECT 108.825 116.285 109.490 116.455 ;
        RECT 109.775 116.430 109.945 117.230 ;
        RECT 108.825 115.525 108.995 116.285 ;
        RECT 109.175 115.355 109.505 116.115 ;
        RECT 109.675 115.525 109.945 116.430 ;
        RECT 112.170 115.790 112.520 117.040 ;
        RECT 114.000 116.530 114.340 117.360 ;
        RECT 116.095 117.180 116.385 117.905 ;
        RECT 116.555 117.135 118.225 117.905 ;
        RECT 110.580 115.355 115.925 115.790 ;
        RECT 116.095 115.355 116.385 116.520 ;
        RECT 116.555 116.445 117.305 116.965 ;
        RECT 117.475 116.615 118.225 117.135 ;
        RECT 118.455 117.085 118.665 117.905 ;
        RECT 118.835 117.105 119.165 117.735 ;
        RECT 118.835 116.505 119.085 117.105 ;
        RECT 119.335 117.085 119.565 117.905 ;
        RECT 119.775 117.135 122.365 117.905 ;
        RECT 122.540 117.360 127.885 117.905 ;
        RECT 119.255 116.665 119.585 116.915 ;
        RECT 116.555 115.355 118.225 116.445 ;
        RECT 118.455 115.355 118.665 116.495 ;
        RECT 118.835 115.525 119.165 116.505 ;
        RECT 119.335 115.355 119.565 116.495 ;
        RECT 119.775 116.445 120.985 116.965 ;
        RECT 121.155 116.615 122.365 117.135 ;
        RECT 119.775 115.355 122.365 116.445 ;
        RECT 124.130 115.790 124.480 117.040 ;
        RECT 125.960 116.530 126.300 117.360 ;
        RECT 128.055 117.155 129.265 117.905 ;
        RECT 128.055 116.445 128.575 116.985 ;
        RECT 128.745 116.615 129.265 117.155 ;
        RECT 122.540 115.355 127.885 115.790 ;
        RECT 128.055 115.355 129.265 116.445 ;
        RECT 9.290 115.185 129.350 115.355 ;
        RECT 9.375 114.095 10.585 115.185 ;
        RECT 12.050 114.845 12.305 114.875 ;
        RECT 11.965 114.675 12.305 114.845 ;
        RECT 9.375 113.385 9.895 113.925 ;
        RECT 10.065 113.555 10.585 114.095 ;
        RECT 12.050 114.205 12.305 114.675 ;
        RECT 12.485 114.385 12.770 115.185 ;
        RECT 12.950 114.465 13.280 114.975 ;
        RECT 9.375 112.635 10.585 113.385 ;
        RECT 12.050 113.345 12.230 114.205 ;
        RECT 12.950 113.875 13.200 114.465 ;
        RECT 13.550 114.315 13.720 114.925 ;
        RECT 13.890 114.495 14.220 115.185 ;
        RECT 14.450 114.635 14.690 114.925 ;
        RECT 14.890 114.805 15.310 115.185 ;
        RECT 15.490 114.715 16.120 114.965 ;
        RECT 16.590 114.805 16.920 115.185 ;
        RECT 15.490 114.635 15.660 114.715 ;
        RECT 17.090 114.635 17.260 114.925 ;
        RECT 17.440 114.805 17.820 115.185 ;
        RECT 18.060 114.800 18.890 114.970 ;
        RECT 14.450 114.465 15.660 114.635 ;
        RECT 12.400 113.545 13.200 113.875 ;
        RECT 12.050 112.815 12.305 113.345 ;
        RECT 12.485 112.635 12.770 113.095 ;
        RECT 12.950 112.895 13.200 113.545 ;
        RECT 13.400 114.295 13.720 114.315 ;
        RECT 13.400 114.125 15.320 114.295 ;
        RECT 13.400 113.230 13.590 114.125 ;
        RECT 15.490 113.955 15.660 114.465 ;
        RECT 15.830 114.205 16.350 114.515 ;
        RECT 13.760 113.785 15.660 113.955 ;
        RECT 13.760 113.725 14.090 113.785 ;
        RECT 14.240 113.555 14.570 113.615 ;
        RECT 13.910 113.285 14.570 113.555 ;
        RECT 13.400 112.900 13.720 113.230 ;
        RECT 13.900 112.635 14.560 113.115 ;
        RECT 14.760 113.025 14.930 113.785 ;
        RECT 15.830 113.615 16.010 114.025 ;
        RECT 15.100 113.445 15.430 113.565 ;
        RECT 16.180 113.445 16.350 114.205 ;
        RECT 15.100 113.275 16.350 113.445 ;
        RECT 16.520 114.385 17.890 114.635 ;
        RECT 16.520 113.615 16.710 114.385 ;
        RECT 17.640 114.125 17.890 114.385 ;
        RECT 16.880 113.955 17.130 114.115 ;
        RECT 18.060 113.955 18.230 114.800 ;
        RECT 19.125 114.515 19.295 115.015 ;
        RECT 19.465 114.685 19.795 115.185 ;
        RECT 18.400 114.125 18.900 114.505 ;
        RECT 19.125 114.345 19.820 114.515 ;
        RECT 16.880 113.785 18.230 113.955 ;
        RECT 17.810 113.745 18.230 113.785 ;
        RECT 16.520 113.275 16.940 113.615 ;
        RECT 17.230 113.285 17.640 113.615 ;
        RECT 14.760 112.855 15.610 113.025 ;
        RECT 16.170 112.635 16.490 113.095 ;
        RECT 16.690 112.845 16.940 113.275 ;
        RECT 17.230 112.635 17.640 113.075 ;
        RECT 17.810 113.015 17.980 113.745 ;
        RECT 18.150 113.195 18.500 113.565 ;
        RECT 18.680 113.255 18.900 114.125 ;
        RECT 19.070 113.555 19.480 114.175 ;
        RECT 19.650 113.375 19.820 114.345 ;
        RECT 19.125 113.185 19.820 113.375 ;
        RECT 17.810 112.815 18.825 113.015 ;
        RECT 19.125 112.855 19.295 113.185 ;
        RECT 19.465 112.635 19.795 113.015 ;
        RECT 20.010 112.895 20.235 115.015 ;
        RECT 20.405 114.685 20.735 115.185 ;
        RECT 20.905 114.515 21.075 115.015 ;
        RECT 20.410 114.345 21.075 114.515 ;
        RECT 20.410 113.355 20.640 114.345 ;
        RECT 20.810 113.525 21.160 114.175 ;
        RECT 21.335 114.110 21.605 115.015 ;
        RECT 21.775 114.425 22.105 115.185 ;
        RECT 22.285 114.255 22.455 115.015 ;
        RECT 20.410 113.185 21.075 113.355 ;
        RECT 20.405 112.635 20.735 113.015 ;
        RECT 20.905 112.895 21.075 113.185 ;
        RECT 21.335 113.310 21.505 114.110 ;
        RECT 21.790 114.085 22.455 114.255 ;
        RECT 23.175 114.110 23.445 115.015 ;
        RECT 23.615 114.425 23.945 115.185 ;
        RECT 24.125 114.255 24.295 115.015 ;
        RECT 21.790 113.940 21.960 114.085 ;
        RECT 21.675 113.610 21.960 113.940 ;
        RECT 21.790 113.355 21.960 113.610 ;
        RECT 22.195 113.535 22.525 113.905 ;
        RECT 21.335 112.805 21.595 113.310 ;
        RECT 21.790 113.185 22.455 113.355 ;
        RECT 21.775 112.635 22.105 113.015 ;
        RECT 22.285 112.805 22.455 113.185 ;
        RECT 23.175 113.310 23.345 114.110 ;
        RECT 23.630 114.085 24.295 114.255 ;
        RECT 24.555 114.095 25.765 115.185 ;
        RECT 23.630 113.940 23.800 114.085 ;
        RECT 23.515 113.610 23.800 113.940 ;
        RECT 23.630 113.355 23.800 113.610 ;
        RECT 24.035 113.535 24.365 113.905 ;
        RECT 24.555 113.555 25.075 114.095 ;
        RECT 25.935 114.020 26.225 115.185 ;
        RECT 26.395 114.095 28.065 115.185 ;
        RECT 25.245 113.385 25.765 113.925 ;
        RECT 26.395 113.575 27.145 114.095 ;
        RECT 28.295 114.045 28.505 115.185 ;
        RECT 28.675 114.035 29.005 115.015 ;
        RECT 29.175 114.045 29.405 115.185 ;
        RECT 30.625 114.255 30.795 115.015 ;
        RECT 30.975 114.425 31.305 115.185 ;
        RECT 30.625 114.085 31.290 114.255 ;
        RECT 31.475 114.110 31.745 115.015 ;
        RECT 27.315 113.405 28.065 113.925 ;
        RECT 23.175 112.805 23.435 113.310 ;
        RECT 23.630 113.185 24.295 113.355 ;
        RECT 23.615 112.635 23.945 113.015 ;
        RECT 24.125 112.805 24.295 113.185 ;
        RECT 24.555 112.635 25.765 113.385 ;
        RECT 25.935 112.635 26.225 113.360 ;
        RECT 26.395 112.635 28.065 113.405 ;
        RECT 28.295 112.635 28.505 113.455 ;
        RECT 28.675 113.435 28.925 114.035 ;
        RECT 31.120 113.940 31.290 114.085 ;
        RECT 29.095 113.625 29.425 113.875 ;
        RECT 30.555 113.535 30.885 113.905 ;
        RECT 31.120 113.610 31.405 113.940 ;
        RECT 28.675 112.805 29.005 113.435 ;
        RECT 29.175 112.635 29.405 113.455 ;
        RECT 31.120 113.355 31.290 113.610 ;
        RECT 30.625 113.185 31.290 113.355 ;
        RECT 31.575 113.310 31.745 114.110 ;
        RECT 30.625 112.805 30.795 113.185 ;
        RECT 30.975 112.635 31.305 113.015 ;
        RECT 31.485 112.805 31.745 113.310 ;
        RECT 32.290 114.205 32.545 114.875 ;
        RECT 32.725 114.385 33.010 115.185 ;
        RECT 33.190 114.465 33.520 114.975 ;
        RECT 32.290 113.345 32.470 114.205 ;
        RECT 33.190 113.875 33.440 114.465 ;
        RECT 33.790 114.315 33.960 114.925 ;
        RECT 34.130 114.495 34.460 115.185 ;
        RECT 34.690 114.635 34.930 114.925 ;
        RECT 35.130 114.805 35.550 115.185 ;
        RECT 35.730 114.715 36.360 114.965 ;
        RECT 36.830 114.805 37.160 115.185 ;
        RECT 35.730 114.635 35.900 114.715 ;
        RECT 37.330 114.635 37.500 114.925 ;
        RECT 37.680 114.805 38.060 115.185 ;
        RECT 38.300 114.800 39.130 114.970 ;
        RECT 34.690 114.465 35.900 114.635 ;
        RECT 32.640 113.545 33.440 113.875 ;
        RECT 32.290 113.145 32.545 113.345 ;
        RECT 32.205 112.975 32.545 113.145 ;
        RECT 32.290 112.815 32.545 112.975 ;
        RECT 32.725 112.635 33.010 113.095 ;
        RECT 33.190 112.895 33.440 113.545 ;
        RECT 33.640 114.295 33.960 114.315 ;
        RECT 33.640 114.125 35.560 114.295 ;
        RECT 33.640 113.230 33.830 114.125 ;
        RECT 35.730 113.955 35.900 114.465 ;
        RECT 36.070 114.205 36.590 114.515 ;
        RECT 34.000 113.785 35.900 113.955 ;
        RECT 34.000 113.725 34.330 113.785 ;
        RECT 34.480 113.555 34.810 113.615 ;
        RECT 34.150 113.285 34.810 113.555 ;
        RECT 33.640 112.900 33.960 113.230 ;
        RECT 34.140 112.635 34.800 113.115 ;
        RECT 35.000 113.025 35.170 113.785 ;
        RECT 36.070 113.615 36.250 114.025 ;
        RECT 35.340 113.445 35.670 113.565 ;
        RECT 36.420 113.445 36.590 114.205 ;
        RECT 35.340 113.275 36.590 113.445 ;
        RECT 36.760 114.385 38.130 114.635 ;
        RECT 36.760 113.615 36.950 114.385 ;
        RECT 37.880 114.125 38.130 114.385 ;
        RECT 37.120 113.955 37.370 114.115 ;
        RECT 38.300 113.955 38.470 114.800 ;
        RECT 39.365 114.515 39.535 115.015 ;
        RECT 39.705 114.685 40.035 115.185 ;
        RECT 38.640 114.125 39.140 114.505 ;
        RECT 39.365 114.345 40.060 114.515 ;
        RECT 37.120 113.785 38.470 113.955 ;
        RECT 38.050 113.745 38.470 113.785 ;
        RECT 36.760 113.275 37.180 113.615 ;
        RECT 37.470 113.285 37.880 113.615 ;
        RECT 35.000 112.855 35.850 113.025 ;
        RECT 36.410 112.635 36.730 113.095 ;
        RECT 36.930 112.845 37.180 113.275 ;
        RECT 37.470 112.635 37.880 113.075 ;
        RECT 38.050 113.015 38.220 113.745 ;
        RECT 38.390 113.195 38.740 113.565 ;
        RECT 38.920 113.255 39.140 114.125 ;
        RECT 39.310 113.555 39.720 114.175 ;
        RECT 39.890 113.375 40.060 114.345 ;
        RECT 39.365 113.185 40.060 113.375 ;
        RECT 38.050 112.815 39.065 113.015 ;
        RECT 39.365 112.855 39.535 113.185 ;
        RECT 39.705 112.635 40.035 113.015 ;
        RECT 40.250 112.895 40.475 115.015 ;
        RECT 40.645 114.685 40.975 115.185 ;
        RECT 41.145 114.515 41.315 115.015 ;
        RECT 40.650 114.345 41.315 114.515 ;
        RECT 40.650 113.355 40.880 114.345 ;
        RECT 41.050 113.525 41.400 114.175 ;
        RECT 41.580 114.045 41.915 115.015 ;
        RECT 42.085 114.045 42.255 115.185 ;
        RECT 42.425 114.845 44.455 115.015 ;
        RECT 41.580 113.375 41.750 114.045 ;
        RECT 42.425 113.875 42.595 114.845 ;
        RECT 41.920 113.545 42.175 113.875 ;
        RECT 42.400 113.545 42.595 113.875 ;
        RECT 42.765 114.505 43.890 114.675 ;
        RECT 42.005 113.375 42.175 113.545 ;
        RECT 42.765 113.375 42.935 114.505 ;
        RECT 40.650 113.185 41.315 113.355 ;
        RECT 40.645 112.635 40.975 113.015 ;
        RECT 41.145 112.895 41.315 113.185 ;
        RECT 41.580 112.805 41.835 113.375 ;
        RECT 42.005 113.205 42.935 113.375 ;
        RECT 43.105 114.165 44.115 114.335 ;
        RECT 43.105 113.365 43.275 114.165 ;
        RECT 42.760 113.170 42.935 113.205 ;
        RECT 42.005 112.635 42.335 113.035 ;
        RECT 42.760 112.805 43.290 113.170 ;
        RECT 43.480 113.145 43.755 113.965 ;
        RECT 43.475 112.975 43.755 113.145 ;
        RECT 43.480 112.805 43.755 112.975 ;
        RECT 43.925 112.805 44.115 114.165 ;
        RECT 44.285 114.180 44.455 114.845 ;
        RECT 44.625 114.425 44.795 115.185 ;
        RECT 45.030 114.425 45.545 114.835 ;
        RECT 44.285 113.990 45.035 114.180 ;
        RECT 45.205 113.615 45.545 114.425 ;
        RECT 46.215 114.045 46.445 115.185 ;
        RECT 46.615 114.035 46.945 115.015 ;
        RECT 47.115 114.045 47.325 115.185 ;
        RECT 47.555 114.425 48.070 114.835 ;
        RECT 48.305 114.425 48.475 115.185 ;
        RECT 48.645 114.845 50.675 115.015 ;
        RECT 46.195 113.625 46.525 113.875 ;
        RECT 44.315 113.445 45.545 113.615 ;
        RECT 44.295 112.635 44.805 113.170 ;
        RECT 45.025 112.840 45.270 113.445 ;
        RECT 46.215 112.635 46.445 113.455 ;
        RECT 46.695 113.435 46.945 114.035 ;
        RECT 47.555 113.615 47.895 114.425 ;
        RECT 48.645 114.180 48.815 114.845 ;
        RECT 49.210 114.505 50.335 114.675 ;
        RECT 48.065 113.990 48.815 114.180 ;
        RECT 48.985 114.165 49.995 114.335 ;
        RECT 46.615 112.805 46.945 113.435 ;
        RECT 47.115 112.635 47.325 113.455 ;
        RECT 47.555 113.445 48.785 113.615 ;
        RECT 47.830 112.840 48.075 113.445 ;
        RECT 48.295 112.635 48.805 113.170 ;
        RECT 48.985 112.805 49.175 114.165 ;
        RECT 49.345 113.825 49.620 113.965 ;
        RECT 49.345 113.655 49.625 113.825 ;
        RECT 49.345 112.805 49.620 113.655 ;
        RECT 49.825 113.365 49.995 114.165 ;
        RECT 50.165 113.375 50.335 114.505 ;
        RECT 50.505 113.875 50.675 114.845 ;
        RECT 50.845 114.045 51.015 115.185 ;
        RECT 51.185 114.045 51.520 115.015 ;
        RECT 50.505 113.545 50.700 113.875 ;
        RECT 50.925 113.545 51.180 113.875 ;
        RECT 50.925 113.375 51.095 113.545 ;
        RECT 51.350 113.375 51.520 114.045 ;
        RECT 51.695 114.020 51.985 115.185 ;
        RECT 52.530 114.205 52.785 114.875 ;
        RECT 52.965 114.385 53.250 115.185 ;
        RECT 53.430 114.465 53.760 114.975 ;
        RECT 52.530 114.165 52.710 114.205 ;
        RECT 52.445 113.995 52.710 114.165 ;
        RECT 50.165 113.205 51.095 113.375 ;
        RECT 50.165 113.170 50.340 113.205 ;
        RECT 49.810 112.805 50.340 113.170 ;
        RECT 50.765 112.635 51.095 113.035 ;
        RECT 51.265 112.805 51.520 113.375 ;
        RECT 51.695 112.635 51.985 113.360 ;
        RECT 52.530 113.345 52.710 113.995 ;
        RECT 53.430 113.875 53.680 114.465 ;
        RECT 54.030 114.315 54.200 114.925 ;
        RECT 54.370 114.495 54.700 115.185 ;
        RECT 54.930 114.635 55.170 114.925 ;
        RECT 55.370 114.805 55.790 115.185 ;
        RECT 55.970 114.715 56.600 114.965 ;
        RECT 57.070 114.805 57.400 115.185 ;
        RECT 55.970 114.635 56.140 114.715 ;
        RECT 57.570 114.635 57.740 114.925 ;
        RECT 57.920 114.805 58.300 115.185 ;
        RECT 58.540 114.800 59.370 114.970 ;
        RECT 54.930 114.465 56.140 114.635 ;
        RECT 52.880 113.545 53.680 113.875 ;
        RECT 52.530 112.815 52.785 113.345 ;
        RECT 52.965 112.635 53.250 113.095 ;
        RECT 53.430 112.895 53.680 113.545 ;
        RECT 53.880 114.295 54.200 114.315 ;
        RECT 53.880 114.125 55.800 114.295 ;
        RECT 53.880 113.230 54.070 114.125 ;
        RECT 55.970 113.955 56.140 114.465 ;
        RECT 56.310 114.205 56.830 114.515 ;
        RECT 54.240 113.785 56.140 113.955 ;
        RECT 54.240 113.725 54.570 113.785 ;
        RECT 54.720 113.555 55.050 113.615 ;
        RECT 54.390 113.285 55.050 113.555 ;
        RECT 53.880 112.900 54.200 113.230 ;
        RECT 54.380 112.635 55.040 113.115 ;
        RECT 55.240 113.025 55.410 113.785 ;
        RECT 56.310 113.615 56.490 114.025 ;
        RECT 55.580 113.445 55.910 113.565 ;
        RECT 56.660 113.445 56.830 114.205 ;
        RECT 55.580 113.275 56.830 113.445 ;
        RECT 57.000 114.385 58.370 114.635 ;
        RECT 57.000 113.615 57.190 114.385 ;
        RECT 58.120 114.125 58.370 114.385 ;
        RECT 57.360 113.955 57.610 114.115 ;
        RECT 58.540 113.955 58.710 114.800 ;
        RECT 59.605 114.515 59.775 115.015 ;
        RECT 59.945 114.685 60.275 115.185 ;
        RECT 58.880 114.125 59.380 114.505 ;
        RECT 59.605 114.345 60.300 114.515 ;
        RECT 57.360 113.785 58.710 113.955 ;
        RECT 58.290 113.745 58.710 113.785 ;
        RECT 57.000 113.275 57.420 113.615 ;
        RECT 57.710 113.285 58.120 113.615 ;
        RECT 55.240 112.855 56.090 113.025 ;
        RECT 56.650 112.635 56.970 113.095 ;
        RECT 57.170 112.845 57.420 113.275 ;
        RECT 57.710 112.635 58.120 113.075 ;
        RECT 58.290 113.015 58.460 113.745 ;
        RECT 58.630 113.195 58.980 113.565 ;
        RECT 59.160 113.255 59.380 114.125 ;
        RECT 59.550 113.555 59.960 114.175 ;
        RECT 60.130 113.375 60.300 114.345 ;
        RECT 59.605 113.185 60.300 113.375 ;
        RECT 58.290 112.815 59.305 113.015 ;
        RECT 59.605 112.855 59.775 113.185 ;
        RECT 59.945 112.635 60.275 113.015 ;
        RECT 60.490 112.895 60.715 115.015 ;
        RECT 60.885 114.685 61.215 115.185 ;
        RECT 61.385 114.515 61.555 115.015 ;
        RECT 62.190 114.845 62.445 114.875 ;
        RECT 62.105 114.675 62.445 114.845 ;
        RECT 60.890 114.345 61.555 114.515 ;
        RECT 60.890 113.355 61.120 114.345 ;
        RECT 62.190 114.205 62.445 114.675 ;
        RECT 62.625 114.385 62.910 115.185 ;
        RECT 63.090 114.465 63.420 114.975 ;
        RECT 61.290 113.525 61.640 114.175 ;
        RECT 60.890 113.185 61.555 113.355 ;
        RECT 60.885 112.635 61.215 113.015 ;
        RECT 61.385 112.895 61.555 113.185 ;
        RECT 62.190 113.345 62.370 114.205 ;
        RECT 63.090 113.875 63.340 114.465 ;
        RECT 63.690 114.315 63.860 114.925 ;
        RECT 64.030 114.495 64.360 115.185 ;
        RECT 64.590 114.635 64.830 114.925 ;
        RECT 65.030 114.805 65.450 115.185 ;
        RECT 65.630 114.715 66.260 114.965 ;
        RECT 66.730 114.805 67.060 115.185 ;
        RECT 65.630 114.635 65.800 114.715 ;
        RECT 67.230 114.635 67.400 114.925 ;
        RECT 67.580 114.805 67.960 115.185 ;
        RECT 68.200 114.800 69.030 114.970 ;
        RECT 64.590 114.465 65.800 114.635 ;
        RECT 62.540 113.545 63.340 113.875 ;
        RECT 62.190 112.815 62.445 113.345 ;
        RECT 62.625 112.635 62.910 113.095 ;
        RECT 63.090 112.895 63.340 113.545 ;
        RECT 63.540 114.295 63.860 114.315 ;
        RECT 63.540 114.125 65.460 114.295 ;
        RECT 63.540 113.230 63.730 114.125 ;
        RECT 65.630 113.955 65.800 114.465 ;
        RECT 65.970 114.205 66.490 114.515 ;
        RECT 63.900 113.785 65.800 113.955 ;
        RECT 63.900 113.725 64.230 113.785 ;
        RECT 64.380 113.555 64.710 113.615 ;
        RECT 64.050 113.285 64.710 113.555 ;
        RECT 63.540 112.900 63.860 113.230 ;
        RECT 64.040 112.635 64.700 113.115 ;
        RECT 64.900 113.025 65.070 113.785 ;
        RECT 65.970 113.615 66.150 114.025 ;
        RECT 65.240 113.445 65.570 113.565 ;
        RECT 66.320 113.445 66.490 114.205 ;
        RECT 65.240 113.275 66.490 113.445 ;
        RECT 66.660 114.385 68.030 114.635 ;
        RECT 66.660 113.615 66.850 114.385 ;
        RECT 67.780 114.125 68.030 114.385 ;
        RECT 67.020 113.955 67.270 114.115 ;
        RECT 68.200 113.955 68.370 114.800 ;
        RECT 69.265 114.515 69.435 115.015 ;
        RECT 69.605 114.685 69.935 115.185 ;
        RECT 68.540 114.125 69.040 114.505 ;
        RECT 69.265 114.345 69.960 114.515 ;
        RECT 67.020 113.785 68.370 113.955 ;
        RECT 67.950 113.745 68.370 113.785 ;
        RECT 66.660 113.275 67.080 113.615 ;
        RECT 67.370 113.285 67.780 113.615 ;
        RECT 64.900 112.855 65.750 113.025 ;
        RECT 66.310 112.635 66.630 113.095 ;
        RECT 66.830 112.845 67.080 113.275 ;
        RECT 67.370 112.635 67.780 113.075 ;
        RECT 67.950 113.015 68.120 113.745 ;
        RECT 68.290 113.195 68.640 113.565 ;
        RECT 68.820 113.255 69.040 114.125 ;
        RECT 69.210 113.555 69.620 114.175 ;
        RECT 69.790 113.375 69.960 114.345 ;
        RECT 69.265 113.185 69.960 113.375 ;
        RECT 67.950 112.815 68.965 113.015 ;
        RECT 69.265 112.855 69.435 113.185 ;
        RECT 69.605 112.635 69.935 113.015 ;
        RECT 70.150 112.895 70.375 115.015 ;
        RECT 70.545 114.685 70.875 115.185 ;
        RECT 71.045 114.515 71.215 115.015 ;
        RECT 70.550 114.345 71.215 114.515 ;
        RECT 70.550 113.355 70.780 114.345 ;
        RECT 70.950 113.525 71.300 114.175 ;
        RECT 71.515 114.045 71.745 115.185 ;
        RECT 71.915 114.035 72.245 115.015 ;
        RECT 72.415 114.045 72.625 115.185 ;
        RECT 72.855 114.425 73.370 114.835 ;
        RECT 73.605 114.425 73.775 115.185 ;
        RECT 73.945 114.845 75.975 115.015 ;
        RECT 71.495 113.625 71.825 113.875 ;
        RECT 70.550 113.185 71.215 113.355 ;
        RECT 70.545 112.635 70.875 113.015 ;
        RECT 71.045 112.895 71.215 113.185 ;
        RECT 71.515 112.635 71.745 113.455 ;
        RECT 71.995 113.435 72.245 114.035 ;
        RECT 72.855 113.615 73.195 114.425 ;
        RECT 73.945 114.180 74.115 114.845 ;
        RECT 74.510 114.505 75.635 114.675 ;
        RECT 73.365 113.990 74.115 114.180 ;
        RECT 74.285 114.165 75.295 114.335 ;
        RECT 71.915 112.805 72.245 113.435 ;
        RECT 72.415 112.635 72.625 113.455 ;
        RECT 72.855 113.445 74.085 113.615 ;
        RECT 73.130 112.840 73.375 113.445 ;
        RECT 73.595 112.635 74.105 113.170 ;
        RECT 74.285 112.805 74.475 114.165 ;
        RECT 74.645 113.825 74.920 113.965 ;
        RECT 74.645 113.655 74.925 113.825 ;
        RECT 74.645 112.805 74.920 113.655 ;
        RECT 75.125 113.365 75.295 114.165 ;
        RECT 75.465 113.375 75.635 114.505 ;
        RECT 75.805 113.875 75.975 114.845 ;
        RECT 76.145 114.045 76.315 115.185 ;
        RECT 76.485 114.045 76.820 115.015 ;
        RECT 75.805 113.545 76.000 113.875 ;
        RECT 76.225 113.545 76.480 113.875 ;
        RECT 76.225 113.375 76.395 113.545 ;
        RECT 76.650 113.375 76.820 114.045 ;
        RECT 77.455 114.020 77.745 115.185 ;
        RECT 77.975 114.045 78.185 115.185 ;
        RECT 78.355 114.035 78.685 115.015 ;
        RECT 78.855 114.045 79.085 115.185 ;
        RECT 79.295 114.110 79.565 115.015 ;
        RECT 79.735 114.425 80.065 115.185 ;
        RECT 80.245 114.255 80.415 115.015 ;
        RECT 75.465 113.205 76.395 113.375 ;
        RECT 75.465 113.170 75.640 113.205 ;
        RECT 75.110 112.805 75.640 113.170 ;
        RECT 76.065 112.635 76.395 113.035 ;
        RECT 76.565 112.805 76.820 113.375 ;
        RECT 77.455 112.635 77.745 113.360 ;
        RECT 77.975 112.635 78.185 113.455 ;
        RECT 78.355 113.435 78.605 114.035 ;
        RECT 78.775 113.625 79.105 113.875 ;
        RECT 78.355 112.805 78.685 113.435 ;
        RECT 78.855 112.635 79.085 113.455 ;
        RECT 79.295 113.310 79.465 114.110 ;
        RECT 79.750 114.085 80.415 114.255 ;
        RECT 80.675 114.095 81.885 115.185 ;
        RECT 82.145 114.515 82.315 115.015 ;
        RECT 82.485 114.685 82.815 115.185 ;
        RECT 82.145 114.345 82.810 114.515 ;
        RECT 79.750 113.940 79.920 114.085 ;
        RECT 79.635 113.610 79.920 113.940 ;
        RECT 79.750 113.355 79.920 113.610 ;
        RECT 80.155 113.535 80.485 113.905 ;
        RECT 80.675 113.555 81.195 114.095 ;
        RECT 81.365 113.385 81.885 113.925 ;
        RECT 82.060 113.525 82.410 114.175 ;
        RECT 79.295 112.805 79.555 113.310 ;
        RECT 79.750 113.185 80.415 113.355 ;
        RECT 79.735 112.635 80.065 113.015 ;
        RECT 80.245 112.805 80.415 113.185 ;
        RECT 80.675 112.635 81.885 113.385 ;
        RECT 82.580 113.355 82.810 114.345 ;
        RECT 82.145 113.185 82.810 113.355 ;
        RECT 82.145 112.895 82.315 113.185 ;
        RECT 82.485 112.635 82.815 113.015 ;
        RECT 82.985 112.895 83.210 115.015 ;
        RECT 83.425 114.685 83.755 115.185 ;
        RECT 83.925 114.515 84.095 115.015 ;
        RECT 84.330 114.800 85.160 114.970 ;
        RECT 85.400 114.805 85.780 115.185 ;
        RECT 83.400 114.345 84.095 114.515 ;
        RECT 83.400 113.375 83.570 114.345 ;
        RECT 83.740 113.555 84.150 114.175 ;
        RECT 84.320 114.125 84.820 114.505 ;
        RECT 83.400 113.185 84.095 113.375 ;
        RECT 84.320 113.255 84.540 114.125 ;
        RECT 84.990 113.955 85.160 114.800 ;
        RECT 85.960 114.635 86.130 114.925 ;
        RECT 86.300 114.805 86.630 115.185 ;
        RECT 87.100 114.715 87.730 114.965 ;
        RECT 87.910 114.805 88.330 115.185 ;
        RECT 87.560 114.635 87.730 114.715 ;
        RECT 88.530 114.635 88.770 114.925 ;
        RECT 85.330 114.385 86.700 114.635 ;
        RECT 85.330 114.125 85.580 114.385 ;
        RECT 86.090 113.955 86.340 114.115 ;
        RECT 84.990 113.785 86.340 113.955 ;
        RECT 84.990 113.745 85.410 113.785 ;
        RECT 84.720 113.195 85.070 113.565 ;
        RECT 83.425 112.635 83.755 113.015 ;
        RECT 83.925 112.855 84.095 113.185 ;
        RECT 85.240 113.015 85.410 113.745 ;
        RECT 86.510 113.615 86.700 114.385 ;
        RECT 85.580 113.285 85.990 113.615 ;
        RECT 86.280 113.275 86.700 113.615 ;
        RECT 86.870 114.205 87.390 114.515 ;
        RECT 87.560 114.465 88.770 114.635 ;
        RECT 89.000 114.495 89.330 115.185 ;
        RECT 86.870 113.445 87.040 114.205 ;
        RECT 87.210 113.615 87.390 114.025 ;
        RECT 87.560 113.955 87.730 114.465 ;
        RECT 89.500 114.315 89.670 114.925 ;
        RECT 89.940 114.465 90.270 114.975 ;
        RECT 89.500 114.295 89.820 114.315 ;
        RECT 87.900 114.125 89.820 114.295 ;
        RECT 87.560 113.785 89.460 113.955 ;
        RECT 87.790 113.445 88.120 113.565 ;
        RECT 86.870 113.275 88.120 113.445 ;
        RECT 84.395 112.815 85.410 113.015 ;
        RECT 85.580 112.635 85.990 113.075 ;
        RECT 86.280 112.845 86.530 113.275 ;
        RECT 86.730 112.635 87.050 113.095 ;
        RECT 88.290 113.025 88.460 113.785 ;
        RECT 89.130 113.725 89.460 113.785 ;
        RECT 88.650 113.555 88.980 113.615 ;
        RECT 88.650 113.285 89.310 113.555 ;
        RECT 89.630 113.230 89.820 114.125 ;
        RECT 87.610 112.855 88.460 113.025 ;
        RECT 88.660 112.635 89.320 113.115 ;
        RECT 89.500 112.900 89.820 113.230 ;
        RECT 90.020 113.875 90.270 114.465 ;
        RECT 90.450 114.385 90.735 115.185 ;
        RECT 90.915 114.205 91.170 114.875 ;
        RECT 90.020 113.545 90.820 113.875 ;
        RECT 90.020 112.895 90.270 113.545 ;
        RECT 90.990 113.485 91.170 114.205 ;
        RECT 91.775 114.045 91.985 115.185 ;
        RECT 92.155 114.035 92.485 115.015 ;
        RECT 92.655 114.045 92.885 115.185 ;
        RECT 93.135 114.045 93.365 115.185 ;
        RECT 93.535 114.035 93.865 115.015 ;
        RECT 94.035 114.045 94.245 115.185 ;
        RECT 94.565 114.255 94.735 115.015 ;
        RECT 94.915 114.425 95.245 115.185 ;
        RECT 94.565 114.085 95.230 114.255 ;
        RECT 95.415 114.110 95.685 115.015 ;
        RECT 90.990 113.345 91.255 113.485 ;
        RECT 90.915 113.315 91.255 113.345 ;
        RECT 90.450 112.635 90.735 113.095 ;
        RECT 90.915 112.815 91.170 113.315 ;
        RECT 91.775 112.635 91.985 113.455 ;
        RECT 92.155 113.435 92.405 114.035 ;
        RECT 92.575 113.625 92.905 113.875 ;
        RECT 93.115 113.625 93.445 113.875 ;
        RECT 92.155 112.805 92.485 113.435 ;
        RECT 92.655 112.635 92.885 113.455 ;
        RECT 93.135 112.635 93.365 113.455 ;
        RECT 93.615 113.435 93.865 114.035 ;
        RECT 95.060 113.940 95.230 114.085 ;
        RECT 94.495 113.535 94.825 113.905 ;
        RECT 95.060 113.610 95.345 113.940 ;
        RECT 93.535 112.805 93.865 113.435 ;
        RECT 94.035 112.635 94.245 113.455 ;
        RECT 95.060 113.355 95.230 113.610 ;
        RECT 94.565 113.185 95.230 113.355 ;
        RECT 95.515 113.310 95.685 114.110 ;
        RECT 95.855 114.095 97.525 115.185 ;
        RECT 97.700 114.750 103.045 115.185 ;
        RECT 95.855 113.575 96.605 114.095 ;
        RECT 96.775 113.405 97.525 113.925 ;
        RECT 99.290 113.500 99.640 114.750 ;
        RECT 103.215 114.020 103.505 115.185 ;
        RECT 104.135 114.425 104.650 114.835 ;
        RECT 104.885 114.425 105.055 115.185 ;
        RECT 105.225 114.845 107.255 115.015 ;
        RECT 94.565 112.805 94.735 113.185 ;
        RECT 94.915 112.635 95.245 113.015 ;
        RECT 95.425 112.805 95.685 113.310 ;
        RECT 95.855 112.635 97.525 113.405 ;
        RECT 101.120 113.180 101.460 114.010 ;
        RECT 104.135 113.615 104.475 114.425 ;
        RECT 105.225 114.180 105.395 114.845 ;
        RECT 105.790 114.505 106.915 114.675 ;
        RECT 104.645 113.990 105.395 114.180 ;
        RECT 105.565 114.165 106.575 114.335 ;
        RECT 104.135 113.445 105.365 113.615 ;
        RECT 97.700 112.635 103.045 113.180 ;
        RECT 103.215 112.635 103.505 113.360 ;
        RECT 104.410 112.840 104.655 113.445 ;
        RECT 104.875 112.635 105.385 113.170 ;
        RECT 105.565 112.805 105.755 114.165 ;
        RECT 105.925 113.485 106.200 113.965 ;
        RECT 105.925 113.315 106.205 113.485 ;
        RECT 106.405 113.365 106.575 114.165 ;
        RECT 106.745 113.375 106.915 114.505 ;
        RECT 107.085 113.875 107.255 114.845 ;
        RECT 107.425 114.045 107.595 115.185 ;
        RECT 107.765 114.045 108.100 115.015 ;
        RECT 108.335 114.045 108.545 115.185 ;
        RECT 107.085 113.545 107.280 113.875 ;
        RECT 107.505 113.545 107.760 113.875 ;
        RECT 107.505 113.375 107.675 113.545 ;
        RECT 107.930 113.375 108.100 114.045 ;
        RECT 108.715 114.035 109.045 115.015 ;
        RECT 109.215 114.045 109.445 115.185 ;
        RECT 110.575 114.425 111.090 114.835 ;
        RECT 111.325 114.425 111.495 115.185 ;
        RECT 111.665 114.845 113.695 115.015 ;
        RECT 105.925 112.805 106.200 113.315 ;
        RECT 106.745 113.205 107.675 113.375 ;
        RECT 106.745 113.170 106.920 113.205 ;
        RECT 106.390 112.805 106.920 113.170 ;
        RECT 107.345 112.635 107.675 113.035 ;
        RECT 107.845 112.805 108.100 113.375 ;
        RECT 108.335 112.635 108.545 113.455 ;
        RECT 108.715 113.435 108.965 114.035 ;
        RECT 109.135 113.625 109.465 113.875 ;
        RECT 110.575 113.615 110.915 114.425 ;
        RECT 111.665 114.180 111.835 114.845 ;
        RECT 112.230 114.505 113.355 114.675 ;
        RECT 111.085 113.990 111.835 114.180 ;
        RECT 112.005 114.165 113.015 114.335 ;
        RECT 108.715 112.805 109.045 113.435 ;
        RECT 109.215 112.635 109.445 113.455 ;
        RECT 110.575 113.445 111.805 113.615 ;
        RECT 110.850 112.840 111.095 113.445 ;
        RECT 111.315 112.635 111.825 113.170 ;
        RECT 112.005 112.805 112.195 114.165 ;
        RECT 112.365 113.825 112.640 113.965 ;
        RECT 112.365 113.655 112.645 113.825 ;
        RECT 112.365 112.805 112.640 113.655 ;
        RECT 112.845 113.365 113.015 114.165 ;
        RECT 113.185 113.375 113.355 114.505 ;
        RECT 113.525 113.875 113.695 114.845 ;
        RECT 113.865 114.045 114.035 115.185 ;
        RECT 114.205 114.045 114.540 115.015 ;
        RECT 115.090 114.845 115.345 114.875 ;
        RECT 115.005 114.675 115.345 114.845 ;
        RECT 113.525 113.545 113.720 113.875 ;
        RECT 113.945 113.545 114.200 113.875 ;
        RECT 113.945 113.375 114.115 113.545 ;
        RECT 114.370 113.375 114.540 114.045 ;
        RECT 113.185 113.205 114.115 113.375 ;
        RECT 113.185 113.170 113.360 113.205 ;
        RECT 112.830 112.805 113.360 113.170 ;
        RECT 113.785 112.635 114.115 113.035 ;
        RECT 114.285 112.805 114.540 113.375 ;
        RECT 115.090 114.205 115.345 114.675 ;
        RECT 115.525 114.385 115.810 115.185 ;
        RECT 115.990 114.465 116.320 114.975 ;
        RECT 115.090 113.345 115.270 114.205 ;
        RECT 115.990 113.875 116.240 114.465 ;
        RECT 116.590 114.315 116.760 114.925 ;
        RECT 116.930 114.495 117.260 115.185 ;
        RECT 117.490 114.635 117.730 114.925 ;
        RECT 117.930 114.805 118.350 115.185 ;
        RECT 118.530 114.715 119.160 114.965 ;
        RECT 119.630 114.805 119.960 115.185 ;
        RECT 118.530 114.635 118.700 114.715 ;
        RECT 120.130 114.635 120.300 114.925 ;
        RECT 120.480 114.805 120.860 115.185 ;
        RECT 121.100 114.800 121.930 114.970 ;
        RECT 117.490 114.465 118.700 114.635 ;
        RECT 115.440 113.545 116.240 113.875 ;
        RECT 115.090 112.815 115.345 113.345 ;
        RECT 115.525 112.635 115.810 113.095 ;
        RECT 115.990 112.895 116.240 113.545 ;
        RECT 116.440 114.295 116.760 114.315 ;
        RECT 116.440 114.125 118.360 114.295 ;
        RECT 116.440 113.230 116.630 114.125 ;
        RECT 118.530 113.955 118.700 114.465 ;
        RECT 118.870 114.205 119.390 114.515 ;
        RECT 116.800 113.785 118.700 113.955 ;
        RECT 116.800 113.725 117.130 113.785 ;
        RECT 117.280 113.555 117.610 113.615 ;
        RECT 116.950 113.285 117.610 113.555 ;
        RECT 116.440 112.900 116.760 113.230 ;
        RECT 116.940 112.635 117.600 113.115 ;
        RECT 117.800 113.025 117.970 113.785 ;
        RECT 118.870 113.615 119.050 114.025 ;
        RECT 118.140 113.445 118.470 113.565 ;
        RECT 119.220 113.445 119.390 114.205 ;
        RECT 118.140 113.275 119.390 113.445 ;
        RECT 119.560 114.385 120.930 114.635 ;
        RECT 119.560 113.615 119.750 114.385 ;
        RECT 120.680 114.125 120.930 114.385 ;
        RECT 119.920 113.955 120.170 114.115 ;
        RECT 121.100 113.955 121.270 114.800 ;
        RECT 122.165 114.515 122.335 115.015 ;
        RECT 122.505 114.685 122.835 115.185 ;
        RECT 121.440 114.125 121.940 114.505 ;
        RECT 122.165 114.345 122.860 114.515 ;
        RECT 119.920 113.785 121.270 113.955 ;
        RECT 120.850 113.745 121.270 113.785 ;
        RECT 119.560 113.275 119.980 113.615 ;
        RECT 120.270 113.285 120.680 113.615 ;
        RECT 117.800 112.855 118.650 113.025 ;
        RECT 119.210 112.635 119.530 113.095 ;
        RECT 119.730 112.845 119.980 113.275 ;
        RECT 120.270 112.635 120.680 113.075 ;
        RECT 120.850 113.015 121.020 113.745 ;
        RECT 121.190 113.195 121.540 113.565 ;
        RECT 121.720 113.255 121.940 114.125 ;
        RECT 122.110 113.555 122.520 114.175 ;
        RECT 122.690 113.375 122.860 114.345 ;
        RECT 122.165 113.185 122.860 113.375 ;
        RECT 120.850 112.815 121.865 113.015 ;
        RECT 122.165 112.855 122.335 113.185 ;
        RECT 122.505 112.635 122.835 113.015 ;
        RECT 123.050 112.895 123.275 115.015 ;
        RECT 123.445 114.685 123.775 115.185 ;
        RECT 123.945 114.515 124.115 115.015 ;
        RECT 123.450 114.345 124.115 114.515 ;
        RECT 123.450 113.355 123.680 114.345 ;
        RECT 123.850 113.525 124.200 114.175 ;
        RECT 124.375 114.095 127.885 115.185 ;
        RECT 128.055 114.095 129.265 115.185 ;
        RECT 124.375 113.575 126.065 114.095 ;
        RECT 126.235 113.405 127.885 113.925 ;
        RECT 128.055 113.555 128.575 114.095 ;
        RECT 123.450 113.185 124.115 113.355 ;
        RECT 123.445 112.635 123.775 113.015 ;
        RECT 123.945 112.895 124.115 113.185 ;
        RECT 124.375 112.635 127.885 113.405 ;
        RECT 128.745 113.385 129.265 113.925 ;
        RECT 128.055 112.635 129.265 113.385 ;
        RECT 9.290 112.465 129.350 112.635 ;
        RECT 9.375 111.715 10.585 112.465 ;
        RECT 9.375 111.175 9.895 111.715 ;
        RECT 11.215 111.695 12.885 112.465 ;
        RECT 13.055 111.740 13.345 112.465 ;
        RECT 13.975 111.695 15.645 112.465 ;
        RECT 10.065 111.005 10.585 111.545 ;
        RECT 9.375 109.915 10.585 111.005 ;
        RECT 11.215 111.005 11.965 111.525 ;
        RECT 12.135 111.175 12.885 111.695 ;
        RECT 11.215 109.915 12.885 111.005 ;
        RECT 13.055 109.915 13.345 111.080 ;
        RECT 13.975 111.005 14.725 111.525 ;
        RECT 14.895 111.175 15.645 111.695 ;
        RECT 15.875 111.645 16.085 112.465 ;
        RECT 16.255 111.665 16.585 112.295 ;
        RECT 16.255 111.065 16.505 111.665 ;
        RECT 16.755 111.645 16.985 112.465 ;
        RECT 17.195 111.715 18.405 112.465 ;
        RECT 16.675 111.225 17.005 111.475 ;
        RECT 13.975 109.915 15.645 111.005 ;
        RECT 15.875 109.915 16.085 111.055 ;
        RECT 16.255 110.085 16.585 111.065 ;
        RECT 16.755 109.915 16.985 111.055 ;
        RECT 17.195 111.005 17.715 111.545 ;
        RECT 17.885 111.175 18.405 111.715 ;
        RECT 18.575 111.695 22.085 112.465 ;
        RECT 22.260 111.920 27.605 112.465 ;
        RECT 27.780 111.920 33.125 112.465 ;
        RECT 33.300 111.920 38.645 112.465 ;
        RECT 18.575 111.005 20.265 111.525 ;
        RECT 20.435 111.175 22.085 111.695 ;
        RECT 17.195 109.915 18.405 111.005 ;
        RECT 18.575 109.915 22.085 111.005 ;
        RECT 23.850 110.350 24.200 111.600 ;
        RECT 25.680 111.090 26.020 111.920 ;
        RECT 29.370 110.350 29.720 111.600 ;
        RECT 31.200 111.090 31.540 111.920 ;
        RECT 34.890 110.350 35.240 111.600 ;
        RECT 36.720 111.090 37.060 111.920 ;
        RECT 38.815 111.740 39.105 112.465 ;
        RECT 40.200 111.920 45.545 112.465 ;
        RECT 46.090 112.125 46.345 112.285 ;
        RECT 46.005 111.955 46.345 112.125 ;
        RECT 46.525 112.005 46.810 112.465 ;
        RECT 22.260 109.915 27.605 110.350 ;
        RECT 27.780 109.915 33.125 110.350 ;
        RECT 33.300 109.915 38.645 110.350 ;
        RECT 38.815 109.915 39.105 111.080 ;
        RECT 41.790 110.350 42.140 111.600 ;
        RECT 43.620 111.090 43.960 111.920 ;
        RECT 46.090 111.755 46.345 111.955 ;
        RECT 46.090 110.895 46.270 111.755 ;
        RECT 46.990 111.555 47.240 112.205 ;
        RECT 46.440 111.225 47.240 111.555 ;
        RECT 40.200 109.915 45.545 110.350 ;
        RECT 46.090 110.225 46.345 110.895 ;
        RECT 46.525 109.915 46.810 110.715 ;
        RECT 46.990 110.635 47.240 111.225 ;
        RECT 47.440 111.870 47.760 112.200 ;
        RECT 47.940 111.985 48.600 112.465 ;
        RECT 48.800 112.075 49.650 112.245 ;
        RECT 47.440 110.975 47.630 111.870 ;
        RECT 47.950 111.545 48.610 111.815 ;
        RECT 48.280 111.485 48.610 111.545 ;
        RECT 47.800 111.315 48.130 111.375 ;
        RECT 48.800 111.315 48.970 112.075 ;
        RECT 50.210 112.005 50.530 112.465 ;
        RECT 50.730 111.825 50.980 112.255 ;
        RECT 51.270 112.025 51.680 112.465 ;
        RECT 51.850 112.085 52.865 112.285 ;
        RECT 49.140 111.655 50.390 111.825 ;
        RECT 49.140 111.535 49.470 111.655 ;
        RECT 47.800 111.145 49.700 111.315 ;
        RECT 47.440 110.805 49.360 110.975 ;
        RECT 47.440 110.785 47.760 110.805 ;
        RECT 46.990 110.125 47.320 110.635 ;
        RECT 47.590 110.175 47.760 110.785 ;
        RECT 49.530 110.635 49.700 111.145 ;
        RECT 49.870 111.075 50.050 111.485 ;
        RECT 50.220 110.895 50.390 111.655 ;
        RECT 47.930 109.915 48.260 110.605 ;
        RECT 48.490 110.465 49.700 110.635 ;
        RECT 49.870 110.585 50.390 110.895 ;
        RECT 50.560 111.485 50.980 111.825 ;
        RECT 51.270 111.485 51.680 111.815 ;
        RECT 50.560 110.715 50.750 111.485 ;
        RECT 51.850 111.355 52.020 112.085 ;
        RECT 53.165 111.915 53.335 112.245 ;
        RECT 53.505 112.085 53.835 112.465 ;
        RECT 52.190 111.535 52.540 111.905 ;
        RECT 51.850 111.315 52.270 111.355 ;
        RECT 50.920 111.145 52.270 111.315 ;
        RECT 50.920 110.985 51.170 111.145 ;
        RECT 51.680 110.715 51.930 110.975 ;
        RECT 50.560 110.465 51.930 110.715 ;
        RECT 48.490 110.175 48.730 110.465 ;
        RECT 49.530 110.385 49.700 110.465 ;
        RECT 48.930 109.915 49.350 110.295 ;
        RECT 49.530 110.135 50.160 110.385 ;
        RECT 50.630 109.915 50.960 110.295 ;
        RECT 51.130 110.175 51.300 110.465 ;
        RECT 52.100 110.300 52.270 111.145 ;
        RECT 52.720 110.975 52.940 111.845 ;
        RECT 53.165 111.725 53.860 111.915 ;
        RECT 52.440 110.595 52.940 110.975 ;
        RECT 53.110 110.925 53.520 111.545 ;
        RECT 53.690 110.755 53.860 111.725 ;
        RECT 53.165 110.585 53.860 110.755 ;
        RECT 51.480 109.915 51.860 110.295 ;
        RECT 52.100 110.130 52.930 110.300 ;
        RECT 53.165 110.085 53.335 110.585 ;
        RECT 53.505 109.915 53.835 110.415 ;
        RECT 54.050 110.085 54.275 112.205 ;
        RECT 54.445 112.085 54.775 112.465 ;
        RECT 54.945 111.915 55.115 112.205 ;
        RECT 54.450 111.745 55.115 111.915 ;
        RECT 54.450 110.755 54.680 111.745 ;
        RECT 55.375 111.695 58.885 112.465 ;
        RECT 59.060 111.920 64.405 112.465 ;
        RECT 54.850 110.925 55.200 111.575 ;
        RECT 55.375 111.005 57.065 111.525 ;
        RECT 57.235 111.175 58.885 111.695 ;
        RECT 54.450 110.585 55.115 110.755 ;
        RECT 54.445 109.915 54.775 110.415 ;
        RECT 54.945 110.085 55.115 110.585 ;
        RECT 55.375 109.915 58.885 111.005 ;
        RECT 60.650 110.350 61.000 111.600 ;
        RECT 62.480 111.090 62.820 111.920 ;
        RECT 64.575 111.740 64.865 112.465 ;
        RECT 65.495 111.695 68.085 112.465 ;
        RECT 68.630 112.125 68.885 112.285 ;
        RECT 68.545 111.955 68.885 112.125 ;
        RECT 69.065 112.005 69.350 112.465 ;
        RECT 59.060 109.915 64.405 110.350 ;
        RECT 64.575 109.915 64.865 111.080 ;
        RECT 65.495 111.005 66.705 111.525 ;
        RECT 66.875 111.175 68.085 111.695 ;
        RECT 68.630 111.755 68.885 111.955 ;
        RECT 65.495 109.915 68.085 111.005 ;
        RECT 68.630 110.895 68.810 111.755 ;
        RECT 69.530 111.555 69.780 112.205 ;
        RECT 68.980 111.225 69.780 111.555 ;
        RECT 68.630 110.225 68.885 110.895 ;
        RECT 69.065 109.915 69.350 110.715 ;
        RECT 69.530 110.635 69.780 111.225 ;
        RECT 69.980 111.870 70.300 112.200 ;
        RECT 70.480 111.985 71.140 112.465 ;
        RECT 71.340 112.075 72.190 112.245 ;
        RECT 69.980 110.975 70.170 111.870 ;
        RECT 70.490 111.545 71.150 111.815 ;
        RECT 70.820 111.485 71.150 111.545 ;
        RECT 70.340 111.315 70.670 111.375 ;
        RECT 71.340 111.315 71.510 112.075 ;
        RECT 72.750 112.005 73.070 112.465 ;
        RECT 73.270 111.825 73.520 112.255 ;
        RECT 73.810 112.025 74.220 112.465 ;
        RECT 74.390 112.085 75.405 112.285 ;
        RECT 71.680 111.655 72.930 111.825 ;
        RECT 71.680 111.535 72.010 111.655 ;
        RECT 70.340 111.145 72.240 111.315 ;
        RECT 69.980 110.805 71.900 110.975 ;
        RECT 69.980 110.785 70.300 110.805 ;
        RECT 69.530 110.125 69.860 110.635 ;
        RECT 70.130 110.175 70.300 110.785 ;
        RECT 72.070 110.635 72.240 111.145 ;
        RECT 72.410 111.075 72.590 111.485 ;
        RECT 72.760 110.895 72.930 111.655 ;
        RECT 70.470 109.915 70.800 110.605 ;
        RECT 71.030 110.465 72.240 110.635 ;
        RECT 72.410 110.585 72.930 110.895 ;
        RECT 73.100 111.485 73.520 111.825 ;
        RECT 73.810 111.485 74.220 111.815 ;
        RECT 73.100 110.715 73.290 111.485 ;
        RECT 74.390 111.355 74.560 112.085 ;
        RECT 75.705 111.915 75.875 112.245 ;
        RECT 76.045 112.085 76.375 112.465 ;
        RECT 74.730 111.535 75.080 111.905 ;
        RECT 74.390 111.315 74.810 111.355 ;
        RECT 73.460 111.145 74.810 111.315 ;
        RECT 73.460 110.985 73.710 111.145 ;
        RECT 74.220 110.715 74.470 110.975 ;
        RECT 73.100 110.465 74.470 110.715 ;
        RECT 71.030 110.175 71.270 110.465 ;
        RECT 72.070 110.385 72.240 110.465 ;
        RECT 71.470 109.915 71.890 110.295 ;
        RECT 72.070 110.135 72.700 110.385 ;
        RECT 73.170 109.915 73.500 110.295 ;
        RECT 73.670 110.175 73.840 110.465 ;
        RECT 74.640 110.300 74.810 111.145 ;
        RECT 75.260 110.975 75.480 111.845 ;
        RECT 75.705 111.725 76.400 111.915 ;
        RECT 74.980 110.595 75.480 110.975 ;
        RECT 75.650 110.925 76.060 111.545 ;
        RECT 76.230 110.755 76.400 111.725 ;
        RECT 75.705 110.585 76.400 110.755 ;
        RECT 74.020 109.915 74.400 110.295 ;
        RECT 74.640 110.130 75.470 110.300 ;
        RECT 75.705 110.085 75.875 110.585 ;
        RECT 76.045 109.915 76.375 110.415 ;
        RECT 76.590 110.085 76.815 112.205 ;
        RECT 76.985 112.085 77.315 112.465 ;
        RECT 77.485 111.915 77.655 112.205 ;
        RECT 78.840 111.920 84.185 112.465 ;
        RECT 76.990 111.745 77.655 111.915 ;
        RECT 76.990 110.755 77.220 111.745 ;
        RECT 77.390 110.925 77.740 111.575 ;
        RECT 76.990 110.585 77.655 110.755 ;
        RECT 76.985 109.915 77.315 110.415 ;
        RECT 77.485 110.085 77.655 110.585 ;
        RECT 80.430 110.350 80.780 111.600 ;
        RECT 82.260 111.090 82.600 111.920 ;
        RECT 84.355 111.790 84.615 112.295 ;
        RECT 84.795 112.085 85.125 112.465 ;
        RECT 85.305 111.915 85.475 112.295 ;
        RECT 84.355 110.990 84.525 111.790 ;
        RECT 84.810 111.745 85.475 111.915 ;
        RECT 84.810 111.490 84.980 111.745 ;
        RECT 85.795 111.645 86.005 112.465 ;
        RECT 86.175 111.665 86.505 112.295 ;
        RECT 84.695 111.160 84.980 111.490 ;
        RECT 85.215 111.195 85.545 111.565 ;
        RECT 84.810 111.015 84.980 111.160 ;
        RECT 86.175 111.065 86.425 111.665 ;
        RECT 86.675 111.645 86.905 112.465 ;
        RECT 87.575 111.695 90.165 112.465 ;
        RECT 90.335 111.740 90.625 112.465 ;
        RECT 90.795 111.695 92.465 112.465 ;
        RECT 92.640 111.920 97.985 112.465 ;
        RECT 98.160 111.920 103.505 112.465 ;
        RECT 86.595 111.225 86.925 111.475 ;
        RECT 78.840 109.915 84.185 110.350 ;
        RECT 84.355 110.085 84.625 110.990 ;
        RECT 84.810 110.845 85.475 111.015 ;
        RECT 84.795 109.915 85.125 110.675 ;
        RECT 85.305 110.085 85.475 110.845 ;
        RECT 85.795 109.915 86.005 111.055 ;
        RECT 86.175 110.085 86.505 111.065 ;
        RECT 86.675 109.915 86.905 111.055 ;
        RECT 87.575 111.005 88.785 111.525 ;
        RECT 88.955 111.175 90.165 111.695 ;
        RECT 87.575 109.915 90.165 111.005 ;
        RECT 90.335 109.915 90.625 111.080 ;
        RECT 90.795 111.005 91.545 111.525 ;
        RECT 91.715 111.175 92.465 111.695 ;
        RECT 90.795 109.915 92.465 111.005 ;
        RECT 94.230 110.350 94.580 111.600 ;
        RECT 96.060 111.090 96.400 111.920 ;
        RECT 99.750 110.350 100.100 111.600 ;
        RECT 101.580 111.090 101.920 111.920 ;
        RECT 103.765 111.915 103.935 112.205 ;
        RECT 104.105 112.085 104.435 112.465 ;
        RECT 103.765 111.745 104.430 111.915 ;
        RECT 103.680 110.925 104.030 111.575 ;
        RECT 104.200 110.755 104.430 111.745 ;
        RECT 103.765 110.585 104.430 110.755 ;
        RECT 92.640 109.915 97.985 110.350 ;
        RECT 98.160 109.915 103.505 110.350 ;
        RECT 103.765 110.085 103.935 110.585 ;
        RECT 104.105 109.915 104.435 110.415 ;
        RECT 104.605 110.085 104.830 112.205 ;
        RECT 105.045 112.085 105.375 112.465 ;
        RECT 105.545 111.915 105.715 112.245 ;
        RECT 106.015 112.085 107.030 112.285 ;
        RECT 105.020 111.725 105.715 111.915 ;
        RECT 105.020 110.755 105.190 111.725 ;
        RECT 105.360 110.925 105.770 111.545 ;
        RECT 105.940 110.975 106.160 111.845 ;
        RECT 106.340 111.535 106.690 111.905 ;
        RECT 106.860 111.355 107.030 112.085 ;
        RECT 107.200 112.025 107.610 112.465 ;
        RECT 107.900 111.825 108.150 112.255 ;
        RECT 108.350 112.005 108.670 112.465 ;
        RECT 109.230 112.075 110.080 112.245 ;
        RECT 107.200 111.485 107.610 111.815 ;
        RECT 107.900 111.485 108.320 111.825 ;
        RECT 106.610 111.315 107.030 111.355 ;
        RECT 106.610 111.145 107.960 111.315 ;
        RECT 105.020 110.585 105.715 110.755 ;
        RECT 105.940 110.595 106.440 110.975 ;
        RECT 105.045 109.915 105.375 110.415 ;
        RECT 105.545 110.085 105.715 110.585 ;
        RECT 106.610 110.300 106.780 111.145 ;
        RECT 107.710 110.985 107.960 111.145 ;
        RECT 106.950 110.715 107.200 110.975 ;
        RECT 108.130 110.715 108.320 111.485 ;
        RECT 106.950 110.465 108.320 110.715 ;
        RECT 108.490 111.655 109.740 111.825 ;
        RECT 108.490 110.895 108.660 111.655 ;
        RECT 109.410 111.535 109.740 111.655 ;
        RECT 108.830 111.075 109.010 111.485 ;
        RECT 109.910 111.315 110.080 112.075 ;
        RECT 110.280 111.985 110.940 112.465 ;
        RECT 111.120 111.870 111.440 112.200 ;
        RECT 110.270 111.545 110.930 111.815 ;
        RECT 110.270 111.485 110.600 111.545 ;
        RECT 110.750 111.315 111.080 111.375 ;
        RECT 109.180 111.145 111.080 111.315 ;
        RECT 108.490 110.585 109.010 110.895 ;
        RECT 109.180 110.635 109.350 111.145 ;
        RECT 111.250 110.975 111.440 111.870 ;
        RECT 109.520 110.805 111.440 110.975 ;
        RECT 111.120 110.785 111.440 110.805 ;
        RECT 111.640 111.555 111.890 112.205 ;
        RECT 112.070 112.005 112.355 112.465 ;
        RECT 112.535 112.125 112.790 112.285 ;
        RECT 112.535 111.955 112.875 112.125 ;
        RECT 112.535 111.755 112.790 111.955 ;
        RECT 111.640 111.225 112.440 111.555 ;
        RECT 109.180 110.465 110.390 110.635 ;
        RECT 105.950 110.130 106.780 110.300 ;
        RECT 107.020 109.915 107.400 110.295 ;
        RECT 107.580 110.175 107.750 110.465 ;
        RECT 109.180 110.385 109.350 110.465 ;
        RECT 107.920 109.915 108.250 110.295 ;
        RECT 108.720 110.135 109.350 110.385 ;
        RECT 109.530 109.915 109.950 110.295 ;
        RECT 110.150 110.175 110.390 110.465 ;
        RECT 110.620 109.915 110.950 110.605 ;
        RECT 111.120 110.175 111.290 110.785 ;
        RECT 111.640 110.635 111.890 111.225 ;
        RECT 112.610 110.895 112.790 111.755 ;
        RECT 113.335 111.695 115.925 112.465 ;
        RECT 116.095 111.740 116.385 112.465 ;
        RECT 116.555 111.695 119.145 112.465 ;
        RECT 119.405 111.915 119.575 112.295 ;
        RECT 119.755 112.085 120.085 112.465 ;
        RECT 119.405 111.745 120.070 111.915 ;
        RECT 120.265 111.790 120.525 112.295 ;
        RECT 111.560 110.125 111.890 110.635 ;
        RECT 112.070 109.915 112.355 110.715 ;
        RECT 112.535 110.225 112.790 110.895 ;
        RECT 113.335 111.005 114.545 111.525 ;
        RECT 114.715 111.175 115.925 111.695 ;
        RECT 113.335 109.915 115.925 111.005 ;
        RECT 116.095 109.915 116.385 111.080 ;
        RECT 116.555 111.005 117.765 111.525 ;
        RECT 117.935 111.175 119.145 111.695 ;
        RECT 119.335 111.195 119.665 111.565 ;
        RECT 119.900 111.490 120.070 111.745 ;
        RECT 119.900 111.160 120.185 111.490 ;
        RECT 119.900 111.015 120.070 111.160 ;
        RECT 116.555 109.915 119.145 111.005 ;
        RECT 119.405 110.845 120.070 111.015 ;
        RECT 120.355 110.990 120.525 111.790 ;
        RECT 120.695 111.695 122.365 112.465 ;
        RECT 122.540 111.920 127.885 112.465 ;
        RECT 119.405 110.085 119.575 110.845 ;
        RECT 119.755 109.915 120.085 110.675 ;
        RECT 120.255 110.085 120.525 110.990 ;
        RECT 120.695 111.005 121.445 111.525 ;
        RECT 121.615 111.175 122.365 111.695 ;
        RECT 120.695 109.915 122.365 111.005 ;
        RECT 124.130 110.350 124.480 111.600 ;
        RECT 125.960 111.090 126.300 111.920 ;
        RECT 128.055 111.715 129.265 112.465 ;
        RECT 128.055 111.005 128.575 111.545 ;
        RECT 128.745 111.175 129.265 111.715 ;
        RECT 122.540 109.915 127.885 110.350 ;
        RECT 128.055 109.915 129.265 111.005 ;
        RECT 9.290 109.745 129.350 109.915 ;
        RECT 9.375 108.655 10.585 109.745 ;
        RECT 9.375 107.945 9.895 108.485 ;
        RECT 10.065 108.115 10.585 108.655 ;
        RECT 10.760 108.555 11.015 109.435 ;
        RECT 11.185 108.605 11.490 109.745 ;
        RECT 11.830 109.365 12.160 109.745 ;
        RECT 12.340 109.195 12.510 109.485 ;
        RECT 12.680 109.285 12.930 109.745 ;
        RECT 11.710 109.025 12.510 109.195 ;
        RECT 13.100 109.235 13.970 109.575 ;
        RECT 9.375 107.195 10.585 107.945 ;
        RECT 10.760 107.905 10.970 108.555 ;
        RECT 11.710 108.435 11.880 109.025 ;
        RECT 13.100 108.855 13.270 109.235 ;
        RECT 14.205 109.115 14.375 109.575 ;
        RECT 14.545 109.285 14.915 109.745 ;
        RECT 15.210 109.145 15.380 109.485 ;
        RECT 15.550 109.315 15.880 109.745 ;
        RECT 16.115 109.145 16.285 109.485 ;
        RECT 12.050 108.685 13.270 108.855 ;
        RECT 13.440 108.775 13.900 109.065 ;
        RECT 14.205 108.945 14.765 109.115 ;
        RECT 15.210 108.975 16.285 109.145 ;
        RECT 16.455 109.245 17.135 109.575 ;
        RECT 17.350 109.245 17.600 109.575 ;
        RECT 17.770 109.285 18.020 109.745 ;
        RECT 14.595 108.805 14.765 108.945 ;
        RECT 13.440 108.765 14.405 108.775 ;
        RECT 13.100 108.595 13.270 108.685 ;
        RECT 13.730 108.605 14.405 108.765 ;
        RECT 11.140 108.405 11.880 108.435 ;
        RECT 11.140 108.105 12.055 108.405 ;
        RECT 11.730 107.930 12.055 108.105 ;
        RECT 10.760 107.375 11.015 107.905 ;
        RECT 11.185 107.195 11.490 107.655 ;
        RECT 11.735 107.575 12.055 107.930 ;
        RECT 12.225 108.145 12.765 108.515 ;
        RECT 13.100 108.425 13.505 108.595 ;
        RECT 12.225 107.745 12.465 108.145 ;
        RECT 12.945 107.975 13.165 108.255 ;
        RECT 12.635 107.805 13.165 107.975 ;
        RECT 12.635 107.575 12.805 107.805 ;
        RECT 13.335 107.645 13.505 108.425 ;
        RECT 13.675 107.815 14.025 108.435 ;
        RECT 14.195 107.815 14.405 108.605 ;
        RECT 14.595 108.635 16.095 108.805 ;
        RECT 14.595 107.945 14.765 108.635 ;
        RECT 16.455 108.465 16.625 109.245 ;
        RECT 17.430 109.115 17.600 109.245 ;
        RECT 14.935 108.295 16.625 108.465 ;
        RECT 16.795 108.685 17.260 109.075 ;
        RECT 17.430 108.945 17.825 109.115 ;
        RECT 14.935 108.115 15.105 108.295 ;
        RECT 11.735 107.405 12.805 107.575 ;
        RECT 12.975 107.195 13.165 107.635 ;
        RECT 13.335 107.365 14.285 107.645 ;
        RECT 14.595 107.555 14.855 107.945 ;
        RECT 15.275 107.875 16.065 108.125 ;
        RECT 14.505 107.385 14.855 107.555 ;
        RECT 15.065 107.195 15.395 107.655 ;
        RECT 16.270 107.585 16.440 108.295 ;
        RECT 16.795 108.095 16.965 108.685 ;
        RECT 16.610 107.875 16.965 108.095 ;
        RECT 17.135 107.875 17.485 108.495 ;
        RECT 17.655 107.585 17.825 108.945 ;
        RECT 18.190 108.775 18.515 109.560 ;
        RECT 17.995 107.725 18.455 108.775 ;
        RECT 16.270 107.415 17.125 107.585 ;
        RECT 17.330 107.415 17.825 107.585 ;
        RECT 17.995 107.195 18.325 107.555 ;
        RECT 18.685 107.455 18.855 109.575 ;
        RECT 19.025 109.245 19.355 109.745 ;
        RECT 19.525 109.075 19.780 109.575 ;
        RECT 19.030 108.905 19.780 109.075 ;
        RECT 19.030 107.915 19.260 108.905 ;
        RECT 19.430 108.085 19.780 108.735 ;
        RECT 19.955 108.655 21.165 109.745 ;
        RECT 21.335 108.670 21.605 109.575 ;
        RECT 21.775 108.985 22.105 109.745 ;
        RECT 22.285 108.815 22.455 109.575 ;
        RECT 19.955 108.115 20.475 108.655 ;
        RECT 20.645 107.945 21.165 108.485 ;
        RECT 19.030 107.745 19.780 107.915 ;
        RECT 19.025 107.195 19.355 107.575 ;
        RECT 19.525 107.455 19.780 107.745 ;
        RECT 19.955 107.195 21.165 107.945 ;
        RECT 21.335 107.870 21.505 108.670 ;
        RECT 21.790 108.645 22.455 108.815 ;
        RECT 23.175 108.655 25.765 109.745 ;
        RECT 21.790 108.500 21.960 108.645 ;
        RECT 21.675 108.170 21.960 108.500 ;
        RECT 21.790 107.915 21.960 108.170 ;
        RECT 22.195 108.095 22.525 108.465 ;
        RECT 23.175 108.135 24.385 108.655 ;
        RECT 25.935 108.580 26.225 109.745 ;
        RECT 27.315 108.670 27.585 109.575 ;
        RECT 27.755 108.985 28.085 109.745 ;
        RECT 28.265 108.815 28.435 109.575 ;
        RECT 29.620 109.310 34.965 109.745 ;
        RECT 35.140 109.310 40.485 109.745 ;
        RECT 40.660 109.310 46.005 109.745 ;
        RECT 46.180 109.310 51.525 109.745 ;
        RECT 24.555 107.965 25.765 108.485 ;
        RECT 21.335 107.365 21.595 107.870 ;
        RECT 21.790 107.745 22.455 107.915 ;
        RECT 21.775 107.195 22.105 107.575 ;
        RECT 22.285 107.365 22.455 107.745 ;
        RECT 23.175 107.195 25.765 107.965 ;
        RECT 25.935 107.195 26.225 107.920 ;
        RECT 27.315 107.870 27.485 108.670 ;
        RECT 27.770 108.645 28.435 108.815 ;
        RECT 27.770 108.500 27.940 108.645 ;
        RECT 27.655 108.170 27.940 108.500 ;
        RECT 27.770 107.915 27.940 108.170 ;
        RECT 28.175 108.095 28.505 108.465 ;
        RECT 31.210 108.060 31.560 109.310 ;
        RECT 27.315 107.365 27.575 107.870 ;
        RECT 27.770 107.745 28.435 107.915 ;
        RECT 27.755 107.195 28.085 107.575 ;
        RECT 28.265 107.365 28.435 107.745 ;
        RECT 33.040 107.740 33.380 108.570 ;
        RECT 36.730 108.060 37.080 109.310 ;
        RECT 38.560 107.740 38.900 108.570 ;
        RECT 42.250 108.060 42.600 109.310 ;
        RECT 44.080 107.740 44.420 108.570 ;
        RECT 47.770 108.060 48.120 109.310 ;
        RECT 51.695 108.580 51.985 109.745 ;
        RECT 52.245 108.815 52.415 109.575 ;
        RECT 52.595 108.985 52.925 109.745 ;
        RECT 52.245 108.645 52.910 108.815 ;
        RECT 53.095 108.670 53.365 109.575 ;
        RECT 49.600 107.740 49.940 108.570 ;
        RECT 52.740 108.500 52.910 108.645 ;
        RECT 52.175 108.095 52.505 108.465 ;
        RECT 52.740 108.170 53.025 108.500 ;
        RECT 29.620 107.195 34.965 107.740 ;
        RECT 35.140 107.195 40.485 107.740 ;
        RECT 40.660 107.195 46.005 107.740 ;
        RECT 46.180 107.195 51.525 107.740 ;
        RECT 51.695 107.195 51.985 107.920 ;
        RECT 52.740 107.915 52.910 108.170 ;
        RECT 52.245 107.745 52.910 107.915 ;
        RECT 53.195 107.870 53.365 108.670 ;
        RECT 53.535 108.655 55.205 109.745 ;
        RECT 55.380 109.310 60.725 109.745 ;
        RECT 60.900 109.310 66.245 109.745 ;
        RECT 66.420 109.310 71.765 109.745 ;
        RECT 71.940 109.310 77.285 109.745 ;
        RECT 53.535 108.135 54.285 108.655 ;
        RECT 54.455 107.965 55.205 108.485 ;
        RECT 56.970 108.060 57.320 109.310 ;
        RECT 52.245 107.365 52.415 107.745 ;
        RECT 52.595 107.195 52.925 107.575 ;
        RECT 53.105 107.365 53.365 107.870 ;
        RECT 53.535 107.195 55.205 107.965 ;
        RECT 58.800 107.740 59.140 108.570 ;
        RECT 62.490 108.060 62.840 109.310 ;
        RECT 64.320 107.740 64.660 108.570 ;
        RECT 68.010 108.060 68.360 109.310 ;
        RECT 69.840 107.740 70.180 108.570 ;
        RECT 73.530 108.060 73.880 109.310 ;
        RECT 77.455 108.580 77.745 109.745 ;
        RECT 78.375 108.655 80.045 109.745 ;
        RECT 80.225 108.765 80.555 109.575 ;
        RECT 80.725 108.945 80.965 109.745 ;
        RECT 75.360 107.740 75.700 108.570 ;
        RECT 78.375 108.135 79.125 108.655 ;
        RECT 80.225 108.595 80.940 108.765 ;
        RECT 79.295 107.965 80.045 108.485 ;
        RECT 80.220 108.185 80.600 108.425 ;
        RECT 80.770 108.355 80.940 108.595 ;
        RECT 81.145 108.725 81.315 109.575 ;
        RECT 81.485 108.945 81.815 109.745 ;
        RECT 81.985 108.725 82.155 109.575 ;
        RECT 81.145 108.555 82.155 108.725 ;
        RECT 82.325 108.595 82.655 109.745 ;
        RECT 83.895 108.655 87.405 109.745 ;
        RECT 87.580 109.310 92.925 109.745 ;
        RECT 93.100 109.310 98.445 109.745 ;
        RECT 80.770 108.185 81.270 108.355 ;
        RECT 80.770 108.015 80.940 108.185 ;
        RECT 81.660 108.045 82.155 108.555 ;
        RECT 83.895 108.135 85.585 108.655 ;
        RECT 81.655 108.015 82.155 108.045 ;
        RECT 55.380 107.195 60.725 107.740 ;
        RECT 60.900 107.195 66.245 107.740 ;
        RECT 66.420 107.195 71.765 107.740 ;
        RECT 71.940 107.195 77.285 107.740 ;
        RECT 77.455 107.195 77.745 107.920 ;
        RECT 78.375 107.195 80.045 107.965 ;
        RECT 80.305 107.845 80.940 108.015 ;
        RECT 81.145 107.845 82.155 108.015 ;
        RECT 80.305 107.365 80.475 107.845 ;
        RECT 80.655 107.195 80.895 107.675 ;
        RECT 81.145 107.365 81.315 107.845 ;
        RECT 81.485 107.195 81.815 107.675 ;
        RECT 81.985 107.365 82.155 107.845 ;
        RECT 82.325 107.195 82.655 107.995 ;
        RECT 85.755 107.965 87.405 108.485 ;
        RECT 89.170 108.060 89.520 109.310 ;
        RECT 83.895 107.195 87.405 107.965 ;
        RECT 91.000 107.740 91.340 108.570 ;
        RECT 94.690 108.060 95.040 109.310 ;
        RECT 98.705 108.815 98.875 109.575 ;
        RECT 99.055 108.985 99.385 109.745 ;
        RECT 98.705 108.645 99.370 108.815 ;
        RECT 99.555 108.670 99.825 109.575 ;
        RECT 96.520 107.740 96.860 108.570 ;
        RECT 99.200 108.500 99.370 108.645 ;
        RECT 98.635 108.095 98.965 108.465 ;
        RECT 99.200 108.170 99.485 108.500 ;
        RECT 99.200 107.915 99.370 108.170 ;
        RECT 98.705 107.745 99.370 107.915 ;
        RECT 99.655 107.870 99.825 108.670 ;
        RECT 100.455 108.655 103.045 109.745 ;
        RECT 100.455 108.135 101.665 108.655 ;
        RECT 103.215 108.580 103.505 109.745 ;
        RECT 103.675 108.655 104.885 109.745 ;
        RECT 105.060 109.310 110.405 109.745 ;
        RECT 110.580 109.310 115.925 109.745 ;
        RECT 116.100 109.310 121.445 109.745 ;
        RECT 101.835 107.965 103.045 108.485 ;
        RECT 103.675 108.115 104.195 108.655 ;
        RECT 87.580 107.195 92.925 107.740 ;
        RECT 93.100 107.195 98.445 107.740 ;
        RECT 98.705 107.365 98.875 107.745 ;
        RECT 99.055 107.195 99.385 107.575 ;
        RECT 99.565 107.365 99.825 107.870 ;
        RECT 100.455 107.195 103.045 107.965 ;
        RECT 104.365 107.945 104.885 108.485 ;
        RECT 106.650 108.060 107.000 109.310 ;
        RECT 103.215 107.195 103.505 107.920 ;
        RECT 103.675 107.195 104.885 107.945 ;
        RECT 108.480 107.740 108.820 108.570 ;
        RECT 112.170 108.060 112.520 109.310 ;
        RECT 114.000 107.740 114.340 108.570 ;
        RECT 117.690 108.060 118.040 109.310 ;
        RECT 121.615 108.670 121.885 109.575 ;
        RECT 122.055 108.985 122.385 109.745 ;
        RECT 122.565 108.815 122.735 109.575 ;
        RECT 119.520 107.740 119.860 108.570 ;
        RECT 121.615 107.870 121.785 108.670 ;
        RECT 122.070 108.645 122.735 108.815 ;
        RECT 122.995 108.670 123.265 109.575 ;
        RECT 123.435 108.985 123.765 109.745 ;
        RECT 123.945 108.815 124.115 109.575 ;
        RECT 122.070 108.500 122.240 108.645 ;
        RECT 121.955 108.170 122.240 108.500 ;
        RECT 122.070 107.915 122.240 108.170 ;
        RECT 122.475 108.095 122.805 108.465 ;
        RECT 105.060 107.195 110.405 107.740 ;
        RECT 110.580 107.195 115.925 107.740 ;
        RECT 116.100 107.195 121.445 107.740 ;
        RECT 121.615 107.365 121.875 107.870 ;
        RECT 122.070 107.745 122.735 107.915 ;
        RECT 122.055 107.195 122.385 107.575 ;
        RECT 122.565 107.365 122.735 107.745 ;
        RECT 122.995 107.870 123.165 108.670 ;
        RECT 123.450 108.645 124.115 108.815 ;
        RECT 124.375 108.655 127.885 109.745 ;
        RECT 128.055 108.655 129.265 109.745 ;
        RECT 123.450 108.500 123.620 108.645 ;
        RECT 123.335 108.170 123.620 108.500 ;
        RECT 123.450 107.915 123.620 108.170 ;
        RECT 123.855 108.095 124.185 108.465 ;
        RECT 124.375 108.135 126.065 108.655 ;
        RECT 126.235 107.965 127.885 108.485 ;
        RECT 128.055 108.115 128.575 108.655 ;
        RECT 122.995 107.365 123.255 107.870 ;
        RECT 123.450 107.745 124.115 107.915 ;
        RECT 123.435 107.195 123.765 107.575 ;
        RECT 123.945 107.365 124.115 107.745 ;
        RECT 124.375 107.195 127.885 107.965 ;
        RECT 128.745 107.945 129.265 108.485 ;
        RECT 128.055 107.195 129.265 107.945 ;
        RECT 9.290 107.025 129.350 107.195 ;
        RECT 9.375 106.275 10.585 107.025 ;
        RECT 9.375 105.735 9.895 106.275 ;
        RECT 11.215 106.255 12.885 107.025 ;
        RECT 13.055 106.300 13.345 107.025 ;
        RECT 10.065 105.565 10.585 106.105 ;
        RECT 9.375 104.475 10.585 105.565 ;
        RECT 11.215 105.565 11.965 106.085 ;
        RECT 12.135 105.735 12.885 106.255 ;
        RECT 14.495 106.205 14.705 107.025 ;
        RECT 14.875 106.225 15.205 106.855 ;
        RECT 11.215 104.475 12.885 105.565 ;
        RECT 13.055 104.475 13.345 105.640 ;
        RECT 14.875 105.625 15.125 106.225 ;
        RECT 15.375 106.205 15.605 107.025 ;
        RECT 15.820 106.315 16.075 106.845 ;
        RECT 16.245 106.565 16.550 107.025 ;
        RECT 16.795 106.645 17.865 106.815 ;
        RECT 15.295 105.785 15.625 106.035 ;
        RECT 15.820 105.665 16.030 106.315 ;
        RECT 16.795 106.290 17.115 106.645 ;
        RECT 16.790 106.115 17.115 106.290 ;
        RECT 16.200 105.815 17.115 106.115 ;
        RECT 17.285 106.075 17.525 106.475 ;
        RECT 17.695 106.415 17.865 106.645 ;
        RECT 18.035 106.585 18.225 107.025 ;
        RECT 18.395 106.575 19.345 106.855 ;
        RECT 19.565 106.665 19.915 106.835 ;
        RECT 17.695 106.245 18.225 106.415 ;
        RECT 16.200 105.785 16.940 105.815 ;
        RECT 14.495 104.475 14.705 105.615 ;
        RECT 14.875 104.645 15.205 105.625 ;
        RECT 15.375 104.475 15.605 105.615 ;
        RECT 15.820 104.785 16.075 105.665 ;
        RECT 16.245 104.475 16.550 105.615 ;
        RECT 16.770 105.195 16.940 105.785 ;
        RECT 17.285 105.705 17.825 106.075 ;
        RECT 18.005 105.965 18.225 106.245 ;
        RECT 18.395 105.795 18.565 106.575 ;
        RECT 18.160 105.625 18.565 105.795 ;
        RECT 18.735 105.785 19.085 106.405 ;
        RECT 18.160 105.535 18.330 105.625 ;
        RECT 19.255 105.615 19.465 106.405 ;
        RECT 17.110 105.365 18.330 105.535 ;
        RECT 18.790 105.455 19.465 105.615 ;
        RECT 16.770 105.025 17.570 105.195 ;
        RECT 16.890 104.475 17.220 104.855 ;
        RECT 17.400 104.735 17.570 105.025 ;
        RECT 18.160 104.985 18.330 105.365 ;
        RECT 18.500 105.445 19.465 105.455 ;
        RECT 19.655 106.275 19.915 106.665 ;
        RECT 20.125 106.565 20.455 107.025 ;
        RECT 21.330 106.635 22.185 106.805 ;
        RECT 22.390 106.635 22.885 106.805 ;
        RECT 23.055 106.665 23.385 107.025 ;
        RECT 19.655 105.585 19.825 106.275 ;
        RECT 19.995 105.925 20.165 106.105 ;
        RECT 20.335 106.095 21.125 106.345 ;
        RECT 21.330 105.925 21.500 106.635 ;
        RECT 21.670 106.125 22.025 106.345 ;
        RECT 19.995 105.755 21.685 105.925 ;
        RECT 18.500 105.155 18.960 105.445 ;
        RECT 19.655 105.415 21.155 105.585 ;
        RECT 19.655 105.275 19.825 105.415 ;
        RECT 19.265 105.105 19.825 105.275 ;
        RECT 17.740 104.475 17.990 104.935 ;
        RECT 18.160 104.645 19.030 104.985 ;
        RECT 19.265 104.645 19.435 105.105 ;
        RECT 20.270 105.075 21.345 105.245 ;
        RECT 19.605 104.475 19.975 104.935 ;
        RECT 20.270 104.735 20.440 105.075 ;
        RECT 20.610 104.475 20.940 104.905 ;
        RECT 21.175 104.735 21.345 105.075 ;
        RECT 21.515 104.975 21.685 105.755 ;
        RECT 21.855 105.535 22.025 106.125 ;
        RECT 22.195 105.725 22.545 106.345 ;
        RECT 21.855 105.145 22.320 105.535 ;
        RECT 22.715 105.275 22.885 106.635 ;
        RECT 23.055 105.445 23.515 106.495 ;
        RECT 22.490 105.105 22.885 105.275 ;
        RECT 22.490 104.975 22.660 105.105 ;
        RECT 21.515 104.645 22.195 104.975 ;
        RECT 22.410 104.645 22.660 104.975 ;
        RECT 22.830 104.475 23.080 104.935 ;
        RECT 23.250 104.660 23.575 105.445 ;
        RECT 23.745 104.645 23.915 106.765 ;
        RECT 24.085 106.645 24.415 107.025 ;
        RECT 24.585 106.475 24.840 106.765 ;
        RECT 24.090 106.305 24.840 106.475 ;
        RECT 24.090 105.315 24.320 106.305 ;
        RECT 25.475 106.255 27.145 107.025 ;
        RECT 24.490 105.485 24.840 106.135 ;
        RECT 25.475 105.565 26.225 106.085 ;
        RECT 26.395 105.735 27.145 106.255 ;
        RECT 27.315 106.350 27.575 106.855 ;
        RECT 27.755 106.645 28.085 107.025 ;
        RECT 28.265 106.475 28.435 106.855 ;
        RECT 24.090 105.145 24.840 105.315 ;
        RECT 24.085 104.475 24.415 104.975 ;
        RECT 24.585 104.645 24.840 105.145 ;
        RECT 25.475 104.475 27.145 105.565 ;
        RECT 27.315 105.550 27.485 106.350 ;
        RECT 27.770 106.305 28.435 106.475 ;
        RECT 27.770 106.050 27.940 106.305 ;
        RECT 28.695 106.255 31.285 107.025 ;
        RECT 27.655 105.720 27.940 106.050 ;
        RECT 28.175 105.755 28.505 106.125 ;
        RECT 27.770 105.575 27.940 105.720 ;
        RECT 27.315 104.645 27.585 105.550 ;
        RECT 27.770 105.405 28.435 105.575 ;
        RECT 27.755 104.475 28.085 105.235 ;
        RECT 28.265 104.645 28.435 105.405 ;
        RECT 28.695 105.565 29.905 106.085 ;
        RECT 30.075 105.735 31.285 106.255 ;
        RECT 31.455 106.350 31.715 106.855 ;
        RECT 31.895 106.645 32.225 107.025 ;
        RECT 32.405 106.475 32.575 106.855 ;
        RECT 28.695 104.475 31.285 105.565 ;
        RECT 31.455 105.550 31.625 106.350 ;
        RECT 31.910 106.305 32.575 106.475 ;
        RECT 31.910 106.050 32.080 106.305 ;
        RECT 33.295 106.255 36.805 107.025 ;
        RECT 31.795 105.720 32.080 106.050 ;
        RECT 32.315 105.755 32.645 106.125 ;
        RECT 31.910 105.575 32.080 105.720 ;
        RECT 31.455 104.645 31.725 105.550 ;
        RECT 31.910 105.405 32.575 105.575 ;
        RECT 31.895 104.475 32.225 105.235 ;
        RECT 32.405 104.645 32.575 105.405 ;
        RECT 33.295 105.565 34.985 106.085 ;
        RECT 35.155 105.735 36.805 106.255 ;
        RECT 36.975 106.350 37.235 106.855 ;
        RECT 37.415 106.645 37.745 107.025 ;
        RECT 37.925 106.475 38.095 106.855 ;
        RECT 33.295 104.475 36.805 105.565 ;
        RECT 36.975 105.550 37.145 106.350 ;
        RECT 37.430 106.305 38.095 106.475 ;
        RECT 37.430 106.050 37.600 106.305 ;
        RECT 38.815 106.300 39.105 107.025 ;
        RECT 40.255 106.205 40.465 107.025 ;
        RECT 40.635 106.225 40.965 106.855 ;
        RECT 37.315 105.720 37.600 106.050 ;
        RECT 37.835 105.755 38.165 106.125 ;
        RECT 37.430 105.575 37.600 105.720 ;
        RECT 36.975 104.645 37.245 105.550 ;
        RECT 37.430 105.405 38.095 105.575 ;
        RECT 37.415 104.475 37.745 105.235 ;
        RECT 37.925 104.645 38.095 105.405 ;
        RECT 38.815 104.475 39.105 105.640 ;
        RECT 40.635 105.625 40.885 106.225 ;
        RECT 41.135 106.205 41.365 107.025 ;
        RECT 41.575 106.350 41.835 106.855 ;
        RECT 42.015 106.645 42.345 107.025 ;
        RECT 42.525 106.475 42.695 106.855 ;
        RECT 41.055 105.785 41.385 106.035 ;
        RECT 40.255 104.475 40.465 105.615 ;
        RECT 40.635 104.645 40.965 105.625 ;
        RECT 41.135 104.475 41.365 105.615 ;
        RECT 41.575 105.550 41.745 106.350 ;
        RECT 42.030 106.305 42.695 106.475 ;
        RECT 42.030 106.050 42.200 106.305 ;
        RECT 43.415 106.255 45.085 107.025 ;
        RECT 45.345 106.475 45.515 106.855 ;
        RECT 45.695 106.645 46.025 107.025 ;
        RECT 45.345 106.305 46.010 106.475 ;
        RECT 46.205 106.350 46.465 106.855 ;
        RECT 41.915 105.720 42.200 106.050 ;
        RECT 42.435 105.755 42.765 106.125 ;
        RECT 42.030 105.575 42.200 105.720 ;
        RECT 41.575 104.645 41.845 105.550 ;
        RECT 42.030 105.405 42.695 105.575 ;
        RECT 42.015 104.475 42.345 105.235 ;
        RECT 42.525 104.645 42.695 105.405 ;
        RECT 43.415 105.565 44.165 106.085 ;
        RECT 44.335 105.735 45.085 106.255 ;
        RECT 45.275 105.755 45.605 106.125 ;
        RECT 45.840 106.050 46.010 106.305 ;
        RECT 45.840 105.720 46.125 106.050 ;
        RECT 45.840 105.575 46.010 105.720 ;
        RECT 43.415 104.475 45.085 105.565 ;
        RECT 45.345 105.405 46.010 105.575 ;
        RECT 46.295 105.550 46.465 106.350 ;
        RECT 47.095 106.255 48.765 107.025 ;
        RECT 48.940 106.480 54.285 107.025 ;
        RECT 45.345 104.645 45.515 105.405 ;
        RECT 45.695 104.475 46.025 105.235 ;
        RECT 46.195 104.645 46.465 105.550 ;
        RECT 47.095 105.565 47.845 106.085 ;
        RECT 48.015 105.735 48.765 106.255 ;
        RECT 47.095 104.475 48.765 105.565 ;
        RECT 50.530 104.910 50.880 106.160 ;
        RECT 52.360 105.650 52.700 106.480 ;
        RECT 54.455 106.350 54.715 106.855 ;
        RECT 54.895 106.645 55.225 107.025 ;
        RECT 55.405 106.475 55.575 106.855 ;
        RECT 54.455 105.550 54.625 106.350 ;
        RECT 54.910 106.305 55.575 106.475 ;
        RECT 54.910 106.050 55.080 106.305 ;
        RECT 55.835 106.255 57.505 107.025 ;
        RECT 57.765 106.475 57.935 106.855 ;
        RECT 58.115 106.645 58.445 107.025 ;
        RECT 57.765 106.305 58.430 106.475 ;
        RECT 58.625 106.350 58.885 106.855 ;
        RECT 54.795 105.720 55.080 106.050 ;
        RECT 55.315 105.755 55.645 106.125 ;
        RECT 54.910 105.575 55.080 105.720 ;
        RECT 48.940 104.475 54.285 104.910 ;
        RECT 54.455 104.645 54.725 105.550 ;
        RECT 54.910 105.405 55.575 105.575 ;
        RECT 54.895 104.475 55.225 105.235 ;
        RECT 55.405 104.645 55.575 105.405 ;
        RECT 55.835 105.565 56.585 106.085 ;
        RECT 56.755 105.735 57.505 106.255 ;
        RECT 57.695 105.755 58.025 106.125 ;
        RECT 58.260 106.050 58.430 106.305 ;
        RECT 58.260 105.720 58.545 106.050 ;
        RECT 58.260 105.575 58.430 105.720 ;
        RECT 55.835 104.475 57.505 105.565 ;
        RECT 57.765 105.405 58.430 105.575 ;
        RECT 58.715 105.550 58.885 106.350 ;
        RECT 59.205 106.225 59.535 107.025 ;
        RECT 59.705 106.375 59.875 106.855 ;
        RECT 60.045 106.545 60.375 107.025 ;
        RECT 60.545 106.375 60.715 106.855 ;
        RECT 60.965 106.545 61.205 107.025 ;
        RECT 61.385 106.375 61.555 106.855 ;
        RECT 59.705 106.205 60.715 106.375 ;
        RECT 60.920 106.205 61.555 106.375 ;
        RECT 61.815 106.275 63.025 107.025 ;
        RECT 59.705 105.665 60.200 106.205 ;
        RECT 60.920 106.035 61.090 106.205 ;
        RECT 60.590 105.865 61.090 106.035 ;
        RECT 57.765 104.645 57.935 105.405 ;
        RECT 58.115 104.475 58.445 105.235 ;
        RECT 58.615 104.645 58.885 105.550 ;
        RECT 59.205 104.475 59.535 105.625 ;
        RECT 59.705 105.495 60.715 105.665 ;
        RECT 59.705 104.645 59.875 105.495 ;
        RECT 60.045 104.475 60.375 105.275 ;
        RECT 60.545 104.645 60.715 105.495 ;
        RECT 60.920 105.625 61.090 105.865 ;
        RECT 61.260 105.795 61.640 106.035 ;
        RECT 60.920 105.455 61.635 105.625 ;
        RECT 60.895 104.475 61.135 105.275 ;
        RECT 61.305 104.645 61.635 105.455 ;
        RECT 61.815 105.565 62.335 106.105 ;
        RECT 62.505 105.735 63.025 106.275 ;
        RECT 63.195 106.350 63.455 106.855 ;
        RECT 63.635 106.645 63.965 107.025 ;
        RECT 64.145 106.475 64.315 106.855 ;
        RECT 61.815 104.475 63.025 105.565 ;
        RECT 63.195 105.550 63.365 106.350 ;
        RECT 63.650 106.305 64.315 106.475 ;
        RECT 63.650 106.050 63.820 106.305 ;
        RECT 64.575 106.300 64.865 107.025 ;
        RECT 65.035 106.255 67.625 107.025 ;
        RECT 67.800 106.480 73.145 107.025 ;
        RECT 63.535 105.720 63.820 106.050 ;
        RECT 64.055 105.755 64.385 106.125 ;
        RECT 63.650 105.575 63.820 105.720 ;
        RECT 63.195 104.645 63.465 105.550 ;
        RECT 63.650 105.405 64.315 105.575 ;
        RECT 63.635 104.475 63.965 105.235 ;
        RECT 64.145 104.645 64.315 105.405 ;
        RECT 64.575 104.475 64.865 105.640 ;
        RECT 65.035 105.565 66.245 106.085 ;
        RECT 66.415 105.735 67.625 106.255 ;
        RECT 65.035 104.475 67.625 105.565 ;
        RECT 69.390 104.910 69.740 106.160 ;
        RECT 71.220 105.650 71.560 106.480 ;
        RECT 73.375 106.205 73.585 107.025 ;
        RECT 73.755 106.225 74.085 106.855 ;
        RECT 73.755 105.625 74.005 106.225 ;
        RECT 74.255 106.205 74.485 107.025 ;
        RECT 74.700 106.315 74.955 106.845 ;
        RECT 75.125 106.565 75.430 107.025 ;
        RECT 75.675 106.645 76.745 106.815 ;
        RECT 74.175 105.785 74.505 106.035 ;
        RECT 74.700 105.665 74.910 106.315 ;
        RECT 75.675 106.290 75.995 106.645 ;
        RECT 75.670 106.115 75.995 106.290 ;
        RECT 75.080 105.815 75.995 106.115 ;
        RECT 76.165 106.075 76.405 106.475 ;
        RECT 76.575 106.415 76.745 106.645 ;
        RECT 76.915 106.585 77.105 107.025 ;
        RECT 77.275 106.575 78.225 106.855 ;
        RECT 78.445 106.665 78.795 106.835 ;
        RECT 76.575 106.245 77.105 106.415 ;
        RECT 75.080 105.785 75.820 105.815 ;
        RECT 67.800 104.475 73.145 104.910 ;
        RECT 73.375 104.475 73.585 105.615 ;
        RECT 73.755 104.645 74.085 105.625 ;
        RECT 74.255 104.475 74.485 105.615 ;
        RECT 74.700 104.785 74.955 105.665 ;
        RECT 75.125 104.475 75.430 105.615 ;
        RECT 75.650 105.195 75.820 105.785 ;
        RECT 76.165 105.705 76.705 106.075 ;
        RECT 76.885 105.965 77.105 106.245 ;
        RECT 77.275 105.795 77.445 106.575 ;
        RECT 77.040 105.625 77.445 105.795 ;
        RECT 77.615 105.785 77.965 106.405 ;
        RECT 77.040 105.535 77.210 105.625 ;
        RECT 78.135 105.615 78.345 106.405 ;
        RECT 75.990 105.365 77.210 105.535 ;
        RECT 77.670 105.455 78.345 105.615 ;
        RECT 75.650 105.025 76.450 105.195 ;
        RECT 75.770 104.475 76.100 104.855 ;
        RECT 76.280 104.735 76.450 105.025 ;
        RECT 77.040 104.985 77.210 105.365 ;
        RECT 77.380 105.445 78.345 105.455 ;
        RECT 78.535 106.275 78.795 106.665 ;
        RECT 79.005 106.565 79.335 107.025 ;
        RECT 80.210 106.635 81.065 106.805 ;
        RECT 81.270 106.635 81.765 106.805 ;
        RECT 81.935 106.665 82.265 107.025 ;
        RECT 78.535 105.585 78.705 106.275 ;
        RECT 78.875 105.925 79.045 106.105 ;
        RECT 79.215 106.095 80.005 106.345 ;
        RECT 80.210 105.925 80.380 106.635 ;
        RECT 80.550 106.125 80.905 106.345 ;
        RECT 78.875 105.755 80.565 105.925 ;
        RECT 77.380 105.155 77.840 105.445 ;
        RECT 78.535 105.415 80.035 105.585 ;
        RECT 78.535 105.275 78.705 105.415 ;
        RECT 78.145 105.105 78.705 105.275 ;
        RECT 76.620 104.475 76.870 104.935 ;
        RECT 77.040 104.645 77.910 104.985 ;
        RECT 78.145 104.645 78.315 105.105 ;
        RECT 79.150 105.075 80.225 105.245 ;
        RECT 78.485 104.475 78.855 104.935 ;
        RECT 79.150 104.735 79.320 105.075 ;
        RECT 79.490 104.475 79.820 104.905 ;
        RECT 80.055 104.735 80.225 105.075 ;
        RECT 80.395 104.975 80.565 105.755 ;
        RECT 80.735 105.535 80.905 106.125 ;
        RECT 81.075 105.725 81.425 106.345 ;
        RECT 80.735 105.145 81.200 105.535 ;
        RECT 81.595 105.275 81.765 106.635 ;
        RECT 81.935 105.445 82.395 106.495 ;
        RECT 81.370 105.105 81.765 105.275 ;
        RECT 81.370 104.975 81.540 105.105 ;
        RECT 80.395 104.645 81.075 104.975 ;
        RECT 81.290 104.645 81.540 104.975 ;
        RECT 81.710 104.475 81.960 104.935 ;
        RECT 82.130 104.660 82.455 105.445 ;
        RECT 82.625 104.645 82.795 106.765 ;
        RECT 82.965 106.645 83.295 107.025 ;
        RECT 83.465 106.475 83.720 106.765 ;
        RECT 84.820 106.480 90.165 107.025 ;
        RECT 82.970 106.305 83.720 106.475 ;
        RECT 82.970 105.315 83.200 106.305 ;
        RECT 83.370 105.485 83.720 106.135 ;
        RECT 82.970 105.145 83.720 105.315 ;
        RECT 82.965 104.475 83.295 104.975 ;
        RECT 83.465 104.645 83.720 105.145 ;
        RECT 86.410 104.910 86.760 106.160 ;
        RECT 88.240 105.650 88.580 106.480 ;
        RECT 90.335 106.300 90.625 107.025 ;
        RECT 91.805 106.475 91.975 106.855 ;
        RECT 92.155 106.645 92.485 107.025 ;
        RECT 91.805 106.305 92.470 106.475 ;
        RECT 92.665 106.350 92.925 106.855 ;
        RECT 91.735 105.755 92.065 106.125 ;
        RECT 92.300 106.050 92.470 106.305 ;
        RECT 92.300 105.720 92.585 106.050 ;
        RECT 84.820 104.475 90.165 104.910 ;
        RECT 90.335 104.475 90.625 105.640 ;
        RECT 92.300 105.575 92.470 105.720 ;
        RECT 91.805 105.405 92.470 105.575 ;
        RECT 92.755 105.550 92.925 106.350 ;
        RECT 91.805 104.645 91.975 105.405 ;
        RECT 92.155 104.475 92.485 105.235 ;
        RECT 92.655 104.645 92.925 105.550 ;
        RECT 93.560 106.315 93.815 106.845 ;
        RECT 93.985 106.565 94.290 107.025 ;
        RECT 94.535 106.645 95.605 106.815 ;
        RECT 93.560 105.665 93.770 106.315 ;
        RECT 94.535 106.290 94.855 106.645 ;
        RECT 94.530 106.115 94.855 106.290 ;
        RECT 93.940 105.815 94.855 106.115 ;
        RECT 95.025 106.075 95.265 106.475 ;
        RECT 95.435 106.415 95.605 106.645 ;
        RECT 95.775 106.585 95.965 107.025 ;
        RECT 96.135 106.575 97.085 106.855 ;
        RECT 97.305 106.665 97.655 106.835 ;
        RECT 95.435 106.245 95.965 106.415 ;
        RECT 93.940 105.785 94.680 105.815 ;
        RECT 93.560 104.785 93.815 105.665 ;
        RECT 93.985 104.475 94.290 105.615 ;
        RECT 94.510 105.195 94.680 105.785 ;
        RECT 95.025 105.705 95.565 106.075 ;
        RECT 95.745 105.965 95.965 106.245 ;
        RECT 96.135 105.795 96.305 106.575 ;
        RECT 95.900 105.625 96.305 105.795 ;
        RECT 96.475 105.785 96.825 106.405 ;
        RECT 95.900 105.535 96.070 105.625 ;
        RECT 96.995 105.615 97.205 106.405 ;
        RECT 94.850 105.365 96.070 105.535 ;
        RECT 96.530 105.455 97.205 105.615 ;
        RECT 94.510 105.025 95.310 105.195 ;
        RECT 94.630 104.475 94.960 104.855 ;
        RECT 95.140 104.735 95.310 105.025 ;
        RECT 95.900 104.985 96.070 105.365 ;
        RECT 96.240 105.445 97.205 105.455 ;
        RECT 97.395 106.275 97.655 106.665 ;
        RECT 97.865 106.565 98.195 107.025 ;
        RECT 99.070 106.635 99.925 106.805 ;
        RECT 100.130 106.635 100.625 106.805 ;
        RECT 100.795 106.665 101.125 107.025 ;
        RECT 97.395 105.585 97.565 106.275 ;
        RECT 97.735 105.925 97.905 106.105 ;
        RECT 98.075 106.095 98.865 106.345 ;
        RECT 99.070 105.925 99.240 106.635 ;
        RECT 99.410 106.125 99.765 106.345 ;
        RECT 97.735 105.755 99.425 105.925 ;
        RECT 96.240 105.155 96.700 105.445 ;
        RECT 97.395 105.415 98.895 105.585 ;
        RECT 97.395 105.275 97.565 105.415 ;
        RECT 97.005 105.105 97.565 105.275 ;
        RECT 95.480 104.475 95.730 104.935 ;
        RECT 95.900 104.645 96.770 104.985 ;
        RECT 97.005 104.645 97.175 105.105 ;
        RECT 98.010 105.075 99.085 105.245 ;
        RECT 97.345 104.475 97.715 104.935 ;
        RECT 98.010 104.735 98.180 105.075 ;
        RECT 98.350 104.475 98.680 104.905 ;
        RECT 98.915 104.735 99.085 105.075 ;
        RECT 99.255 104.975 99.425 105.755 ;
        RECT 99.595 105.535 99.765 106.125 ;
        RECT 99.935 105.725 100.285 106.345 ;
        RECT 99.595 105.145 100.060 105.535 ;
        RECT 100.455 105.275 100.625 106.635 ;
        RECT 100.795 105.445 101.255 106.495 ;
        RECT 100.230 105.105 100.625 105.275 ;
        RECT 100.230 104.975 100.400 105.105 ;
        RECT 99.255 104.645 99.935 104.975 ;
        RECT 100.150 104.645 100.400 104.975 ;
        RECT 100.570 104.475 100.820 104.935 ;
        RECT 100.990 104.660 101.315 105.445 ;
        RECT 101.485 104.645 101.655 106.765 ;
        RECT 101.825 106.645 102.155 107.025 ;
        RECT 102.325 106.475 102.580 106.765 ;
        RECT 101.830 106.305 102.580 106.475 ;
        RECT 101.830 105.315 102.060 106.305 ;
        RECT 103.215 106.255 104.885 107.025 ;
        RECT 105.145 106.475 105.315 106.855 ;
        RECT 105.495 106.645 105.825 107.025 ;
        RECT 105.145 106.305 105.810 106.475 ;
        RECT 106.005 106.350 106.265 106.855 ;
        RECT 102.230 105.485 102.580 106.135 ;
        RECT 103.215 105.565 103.965 106.085 ;
        RECT 104.135 105.735 104.885 106.255 ;
        RECT 105.075 105.755 105.405 106.125 ;
        RECT 105.640 106.050 105.810 106.305 ;
        RECT 105.640 105.720 105.925 106.050 ;
        RECT 105.640 105.575 105.810 105.720 ;
        RECT 101.830 105.145 102.580 105.315 ;
        RECT 101.825 104.475 102.155 104.975 ;
        RECT 102.325 104.645 102.580 105.145 ;
        RECT 103.215 104.475 104.885 105.565 ;
        RECT 105.145 105.405 105.810 105.575 ;
        RECT 106.095 105.550 106.265 106.350 ;
        RECT 107.395 106.205 107.625 107.025 ;
        RECT 107.795 106.225 108.125 106.855 ;
        RECT 107.375 105.785 107.705 106.035 ;
        RECT 107.875 105.625 108.125 106.225 ;
        RECT 108.295 106.205 108.505 107.025 ;
        RECT 108.825 106.475 108.995 106.855 ;
        RECT 109.175 106.645 109.505 107.025 ;
        RECT 108.825 106.305 109.490 106.475 ;
        RECT 109.685 106.350 109.945 106.855 ;
        RECT 108.755 105.755 109.085 106.125 ;
        RECT 109.320 106.050 109.490 106.305 ;
        RECT 105.145 104.645 105.315 105.405 ;
        RECT 105.495 104.475 105.825 105.235 ;
        RECT 105.995 104.645 106.265 105.550 ;
        RECT 107.395 104.475 107.625 105.615 ;
        RECT 107.795 104.645 108.125 105.625 ;
        RECT 109.320 105.720 109.605 106.050 ;
        RECT 108.295 104.475 108.505 105.615 ;
        RECT 109.320 105.575 109.490 105.720 ;
        RECT 108.825 105.405 109.490 105.575 ;
        RECT 109.775 105.550 109.945 106.350 ;
        RECT 110.115 106.255 113.625 107.025 ;
        RECT 113.885 106.475 114.055 106.855 ;
        RECT 114.235 106.645 114.565 107.025 ;
        RECT 113.885 106.305 114.550 106.475 ;
        RECT 114.745 106.350 115.005 106.855 ;
        RECT 108.825 104.645 108.995 105.405 ;
        RECT 109.175 104.475 109.505 105.235 ;
        RECT 109.675 104.645 109.945 105.550 ;
        RECT 110.115 105.565 111.805 106.085 ;
        RECT 111.975 105.735 113.625 106.255 ;
        RECT 113.815 105.755 114.145 106.125 ;
        RECT 114.380 106.050 114.550 106.305 ;
        RECT 114.380 105.720 114.665 106.050 ;
        RECT 114.380 105.575 114.550 105.720 ;
        RECT 110.115 104.475 113.625 105.565 ;
        RECT 113.885 105.405 114.550 105.575 ;
        RECT 114.835 105.550 115.005 106.350 ;
        RECT 116.095 106.300 116.385 107.025 ;
        RECT 117.515 106.205 117.745 107.025 ;
        RECT 117.915 106.225 118.245 106.855 ;
        RECT 117.495 105.785 117.825 106.035 ;
        RECT 113.885 104.645 114.055 105.405 ;
        RECT 114.235 104.475 114.565 105.235 ;
        RECT 114.735 104.645 115.005 105.550 ;
        RECT 116.095 104.475 116.385 105.640 ;
        RECT 117.995 105.625 118.245 106.225 ;
        RECT 118.415 106.205 118.625 107.025 ;
        RECT 118.860 106.475 119.115 106.765 ;
        RECT 119.285 106.645 119.615 107.025 ;
        RECT 118.860 106.305 119.610 106.475 ;
        RECT 117.515 104.475 117.745 105.615 ;
        RECT 117.915 104.645 118.245 105.625 ;
        RECT 118.415 104.475 118.625 105.615 ;
        RECT 118.860 105.485 119.210 106.135 ;
        RECT 119.380 105.315 119.610 106.305 ;
        RECT 118.860 105.145 119.610 105.315 ;
        RECT 118.860 104.645 119.115 105.145 ;
        RECT 119.285 104.475 119.615 104.975 ;
        RECT 119.785 104.645 119.955 106.765 ;
        RECT 120.315 106.665 120.645 107.025 ;
        RECT 120.815 106.635 121.310 106.805 ;
        RECT 121.515 106.635 122.370 106.805 ;
        RECT 120.185 105.445 120.645 106.495 ;
        RECT 120.125 104.660 120.450 105.445 ;
        RECT 120.815 105.275 120.985 106.635 ;
        RECT 121.155 105.725 121.505 106.345 ;
        RECT 121.675 106.125 122.030 106.345 ;
        RECT 121.675 105.535 121.845 106.125 ;
        RECT 122.200 105.925 122.370 106.635 ;
        RECT 123.245 106.565 123.575 107.025 ;
        RECT 123.785 106.665 124.135 106.835 ;
        RECT 122.575 106.095 123.365 106.345 ;
        RECT 123.785 106.275 124.045 106.665 ;
        RECT 124.355 106.575 125.305 106.855 ;
        RECT 125.475 106.585 125.665 107.025 ;
        RECT 125.835 106.645 126.905 106.815 ;
        RECT 123.535 105.925 123.705 106.105 ;
        RECT 120.815 105.105 121.210 105.275 ;
        RECT 121.380 105.145 121.845 105.535 ;
        RECT 122.015 105.755 123.705 105.925 ;
        RECT 121.040 104.975 121.210 105.105 ;
        RECT 122.015 104.975 122.185 105.755 ;
        RECT 123.875 105.585 124.045 106.275 ;
        RECT 122.545 105.415 124.045 105.585 ;
        RECT 124.235 105.615 124.445 106.405 ;
        RECT 124.615 105.785 124.965 106.405 ;
        RECT 125.135 105.795 125.305 106.575 ;
        RECT 125.835 106.415 126.005 106.645 ;
        RECT 125.475 106.245 126.005 106.415 ;
        RECT 125.475 105.965 125.695 106.245 ;
        RECT 126.175 106.075 126.415 106.475 ;
        RECT 125.135 105.625 125.540 105.795 ;
        RECT 125.875 105.705 126.415 106.075 ;
        RECT 126.585 106.290 126.905 106.645 ;
        RECT 127.150 106.565 127.455 107.025 ;
        RECT 127.625 106.315 127.880 106.845 ;
        RECT 126.585 106.115 126.910 106.290 ;
        RECT 126.585 105.815 127.500 106.115 ;
        RECT 126.760 105.785 127.500 105.815 ;
        RECT 124.235 105.455 124.910 105.615 ;
        RECT 125.370 105.535 125.540 105.625 ;
        RECT 124.235 105.445 125.200 105.455 ;
        RECT 123.875 105.275 124.045 105.415 ;
        RECT 120.620 104.475 120.870 104.935 ;
        RECT 121.040 104.645 121.290 104.975 ;
        RECT 121.505 104.645 122.185 104.975 ;
        RECT 122.355 105.075 123.430 105.245 ;
        RECT 123.875 105.105 124.435 105.275 ;
        RECT 124.740 105.155 125.200 105.445 ;
        RECT 125.370 105.365 126.590 105.535 ;
        RECT 122.355 104.735 122.525 105.075 ;
        RECT 122.760 104.475 123.090 104.905 ;
        RECT 123.260 104.735 123.430 105.075 ;
        RECT 123.725 104.475 124.095 104.935 ;
        RECT 124.265 104.645 124.435 105.105 ;
        RECT 125.370 104.985 125.540 105.365 ;
        RECT 126.760 105.195 126.930 105.785 ;
        RECT 127.670 105.665 127.880 106.315 ;
        RECT 128.055 106.275 129.265 107.025 ;
        RECT 124.670 104.645 125.540 104.985 ;
        RECT 126.130 105.025 126.930 105.195 ;
        RECT 125.710 104.475 125.960 104.935 ;
        RECT 126.130 104.735 126.300 105.025 ;
        RECT 126.480 104.475 126.810 104.855 ;
        RECT 127.150 104.475 127.455 105.615 ;
        RECT 127.625 104.785 127.880 105.665 ;
        RECT 128.055 105.565 128.575 106.105 ;
        RECT 128.745 105.735 129.265 106.275 ;
        RECT 128.055 104.475 129.265 105.565 ;
        RECT 9.290 104.305 129.350 104.475 ;
        RECT 9.375 103.215 10.585 104.305 ;
        RECT 9.375 102.505 9.895 103.045 ;
        RECT 10.065 102.675 10.585 103.215 ;
        RECT 11.675 103.215 15.185 104.305 ;
        RECT 11.675 102.695 13.365 103.215 ;
        RECT 15.415 103.165 15.625 104.305 ;
        RECT 15.795 103.155 16.125 104.135 ;
        RECT 16.295 103.165 16.525 104.305 ;
        RECT 13.535 102.525 15.185 103.045 ;
        RECT 9.375 101.755 10.585 102.505 ;
        RECT 11.675 101.755 15.185 102.525 ;
        RECT 15.415 101.755 15.625 102.575 ;
        RECT 15.795 102.555 16.045 103.155 ;
        RECT 16.740 103.115 16.995 103.995 ;
        RECT 17.165 103.165 17.470 104.305 ;
        RECT 17.810 103.925 18.140 104.305 ;
        RECT 18.320 103.755 18.490 104.045 ;
        RECT 18.660 103.845 18.910 104.305 ;
        RECT 17.690 103.585 18.490 103.755 ;
        RECT 19.080 103.795 19.950 104.135 ;
        RECT 16.215 102.745 16.545 102.995 ;
        RECT 15.795 101.925 16.125 102.555 ;
        RECT 16.295 101.755 16.525 102.575 ;
        RECT 16.740 102.465 16.950 103.115 ;
        RECT 17.690 102.995 17.860 103.585 ;
        RECT 19.080 103.415 19.250 103.795 ;
        RECT 20.185 103.675 20.355 104.135 ;
        RECT 20.525 103.845 20.895 104.305 ;
        RECT 21.190 103.705 21.360 104.045 ;
        RECT 21.530 103.875 21.860 104.305 ;
        RECT 22.095 103.705 22.265 104.045 ;
        RECT 18.030 103.245 19.250 103.415 ;
        RECT 19.420 103.335 19.880 103.625 ;
        RECT 20.185 103.505 20.745 103.675 ;
        RECT 21.190 103.535 22.265 103.705 ;
        RECT 22.435 103.805 23.115 104.135 ;
        RECT 23.330 103.805 23.580 104.135 ;
        RECT 23.750 103.845 24.000 104.305 ;
        RECT 20.575 103.365 20.745 103.505 ;
        RECT 19.420 103.325 20.385 103.335 ;
        RECT 19.080 103.155 19.250 103.245 ;
        RECT 19.710 103.165 20.385 103.325 ;
        RECT 17.120 102.965 17.860 102.995 ;
        RECT 17.120 102.665 18.035 102.965 ;
        RECT 17.710 102.490 18.035 102.665 ;
        RECT 16.740 101.935 16.995 102.465 ;
        RECT 17.165 101.755 17.470 102.215 ;
        RECT 17.715 102.135 18.035 102.490 ;
        RECT 18.205 102.705 18.745 103.075 ;
        RECT 19.080 102.985 19.485 103.155 ;
        RECT 18.205 102.305 18.445 102.705 ;
        RECT 18.925 102.535 19.145 102.815 ;
        RECT 18.615 102.365 19.145 102.535 ;
        RECT 18.615 102.135 18.785 102.365 ;
        RECT 19.315 102.205 19.485 102.985 ;
        RECT 19.655 102.375 20.005 102.995 ;
        RECT 20.175 102.375 20.385 103.165 ;
        RECT 20.575 103.195 22.075 103.365 ;
        RECT 20.575 102.505 20.745 103.195 ;
        RECT 22.435 103.025 22.605 103.805 ;
        RECT 23.410 103.675 23.580 103.805 ;
        RECT 20.915 102.855 22.605 103.025 ;
        RECT 22.775 103.245 23.240 103.635 ;
        RECT 23.410 103.505 23.805 103.675 ;
        RECT 20.915 102.675 21.085 102.855 ;
        RECT 17.715 101.965 18.785 102.135 ;
        RECT 18.955 101.755 19.145 102.195 ;
        RECT 19.315 101.925 20.265 102.205 ;
        RECT 20.575 102.115 20.835 102.505 ;
        RECT 21.255 102.435 22.045 102.685 ;
        RECT 20.485 101.945 20.835 102.115 ;
        RECT 21.045 101.755 21.375 102.215 ;
        RECT 22.250 102.145 22.420 102.855 ;
        RECT 22.775 102.655 22.945 103.245 ;
        RECT 22.590 102.435 22.945 102.655 ;
        RECT 23.115 102.435 23.465 103.055 ;
        RECT 23.635 102.145 23.805 103.505 ;
        RECT 24.170 103.335 24.495 104.120 ;
        RECT 23.975 102.285 24.435 103.335 ;
        RECT 22.250 101.975 23.105 102.145 ;
        RECT 23.310 101.975 23.805 102.145 ;
        RECT 23.975 101.755 24.305 102.115 ;
        RECT 24.665 102.015 24.835 104.135 ;
        RECT 25.005 103.805 25.335 104.305 ;
        RECT 25.505 103.635 25.760 104.135 ;
        RECT 25.010 103.465 25.760 103.635 ;
        RECT 25.010 102.475 25.240 103.465 ;
        RECT 25.410 102.645 25.760 103.295 ;
        RECT 25.935 103.140 26.225 104.305 ;
        RECT 26.915 103.165 27.125 104.305 ;
        RECT 27.295 103.155 27.625 104.135 ;
        RECT 27.795 103.165 28.025 104.305 ;
        RECT 28.235 103.215 31.745 104.305 ;
        RECT 25.010 102.305 25.760 102.475 ;
        RECT 25.005 101.755 25.335 102.135 ;
        RECT 25.505 102.015 25.760 102.305 ;
        RECT 25.935 101.755 26.225 102.480 ;
        RECT 26.915 101.755 27.125 102.575 ;
        RECT 27.295 102.555 27.545 103.155 ;
        RECT 27.715 102.745 28.045 102.995 ;
        RECT 28.235 102.695 29.925 103.215 ;
        RECT 31.955 103.165 32.185 104.305 ;
        RECT 32.355 103.155 32.685 104.135 ;
        RECT 32.855 103.165 33.065 104.305 ;
        RECT 33.300 103.635 33.555 104.135 ;
        RECT 33.725 103.805 34.055 104.305 ;
        RECT 33.300 103.465 34.050 103.635 ;
        RECT 27.295 101.925 27.625 102.555 ;
        RECT 27.795 101.755 28.025 102.575 ;
        RECT 30.095 102.525 31.745 103.045 ;
        RECT 31.935 102.745 32.265 102.995 ;
        RECT 28.235 101.755 31.745 102.525 ;
        RECT 31.955 101.755 32.185 102.575 ;
        RECT 32.435 102.555 32.685 103.155 ;
        RECT 33.300 102.645 33.650 103.295 ;
        RECT 32.355 101.925 32.685 102.555 ;
        RECT 32.855 101.755 33.065 102.575 ;
        RECT 33.820 102.475 34.050 103.465 ;
        RECT 33.300 102.305 34.050 102.475 ;
        RECT 33.300 102.015 33.555 102.305 ;
        RECT 33.725 101.755 34.055 102.135 ;
        RECT 34.225 102.015 34.395 104.135 ;
        RECT 34.565 103.335 34.890 104.120 ;
        RECT 35.060 103.845 35.310 104.305 ;
        RECT 35.480 103.805 35.730 104.135 ;
        RECT 35.945 103.805 36.625 104.135 ;
        RECT 35.480 103.675 35.650 103.805 ;
        RECT 35.255 103.505 35.650 103.675 ;
        RECT 34.625 102.285 35.085 103.335 ;
        RECT 35.255 102.145 35.425 103.505 ;
        RECT 35.820 103.245 36.285 103.635 ;
        RECT 35.595 102.435 35.945 103.055 ;
        RECT 36.115 102.655 36.285 103.245 ;
        RECT 36.455 103.025 36.625 103.805 ;
        RECT 36.795 103.705 36.965 104.045 ;
        RECT 37.200 103.875 37.530 104.305 ;
        RECT 37.700 103.705 37.870 104.045 ;
        RECT 38.165 103.845 38.535 104.305 ;
        RECT 36.795 103.535 37.870 103.705 ;
        RECT 38.705 103.675 38.875 104.135 ;
        RECT 39.110 103.795 39.980 104.135 ;
        RECT 40.150 103.845 40.400 104.305 ;
        RECT 38.315 103.505 38.875 103.675 ;
        RECT 38.315 103.365 38.485 103.505 ;
        RECT 36.985 103.195 38.485 103.365 ;
        RECT 39.180 103.335 39.640 103.625 ;
        RECT 36.455 102.855 38.145 103.025 ;
        RECT 36.115 102.435 36.470 102.655 ;
        RECT 36.640 102.145 36.810 102.855 ;
        RECT 37.015 102.435 37.805 102.685 ;
        RECT 37.975 102.675 38.145 102.855 ;
        RECT 38.315 102.505 38.485 103.195 ;
        RECT 34.755 101.755 35.085 102.115 ;
        RECT 35.255 101.975 35.750 102.145 ;
        RECT 35.955 101.975 36.810 102.145 ;
        RECT 37.685 101.755 38.015 102.215 ;
        RECT 38.225 102.115 38.485 102.505 ;
        RECT 38.675 103.325 39.640 103.335 ;
        RECT 39.810 103.415 39.980 103.795 ;
        RECT 40.570 103.755 40.740 104.045 ;
        RECT 40.920 103.925 41.250 104.305 ;
        RECT 40.570 103.585 41.370 103.755 ;
        RECT 38.675 103.165 39.350 103.325 ;
        RECT 39.810 103.245 41.030 103.415 ;
        RECT 38.675 102.375 38.885 103.165 ;
        RECT 39.810 103.155 39.980 103.245 ;
        RECT 39.055 102.375 39.405 102.995 ;
        RECT 39.575 102.985 39.980 103.155 ;
        RECT 39.575 102.205 39.745 102.985 ;
        RECT 39.915 102.535 40.135 102.815 ;
        RECT 40.315 102.705 40.855 103.075 ;
        RECT 41.200 102.995 41.370 103.585 ;
        RECT 41.590 103.165 41.895 104.305 ;
        RECT 42.065 103.115 42.320 103.995 ;
        RECT 41.200 102.965 41.940 102.995 ;
        RECT 39.915 102.365 40.445 102.535 ;
        RECT 38.225 101.945 38.575 102.115 ;
        RECT 38.795 101.925 39.745 102.205 ;
        RECT 39.915 101.755 40.105 102.195 ;
        RECT 40.275 102.135 40.445 102.365 ;
        RECT 40.615 102.305 40.855 102.705 ;
        RECT 41.025 102.665 41.940 102.965 ;
        RECT 41.025 102.490 41.350 102.665 ;
        RECT 41.025 102.135 41.345 102.490 ;
        RECT 42.110 102.465 42.320 103.115 ;
        RECT 40.275 101.965 41.345 102.135 ;
        RECT 41.590 101.755 41.895 102.215 ;
        RECT 42.065 101.935 42.320 102.465 ;
        RECT 42.500 103.115 42.755 103.995 ;
        RECT 42.925 103.165 43.230 104.305 ;
        RECT 43.570 103.925 43.900 104.305 ;
        RECT 44.080 103.755 44.250 104.045 ;
        RECT 44.420 103.845 44.670 104.305 ;
        RECT 43.450 103.585 44.250 103.755 ;
        RECT 44.840 103.795 45.710 104.135 ;
        RECT 42.500 102.465 42.710 103.115 ;
        RECT 43.450 102.995 43.620 103.585 ;
        RECT 44.840 103.415 45.010 103.795 ;
        RECT 45.945 103.675 46.115 104.135 ;
        RECT 46.285 103.845 46.655 104.305 ;
        RECT 46.950 103.705 47.120 104.045 ;
        RECT 47.290 103.875 47.620 104.305 ;
        RECT 47.855 103.705 48.025 104.045 ;
        RECT 43.790 103.245 45.010 103.415 ;
        RECT 45.180 103.335 45.640 103.625 ;
        RECT 45.945 103.505 46.505 103.675 ;
        RECT 46.950 103.535 48.025 103.705 ;
        RECT 48.195 103.805 48.875 104.135 ;
        RECT 49.090 103.805 49.340 104.135 ;
        RECT 49.510 103.845 49.760 104.305 ;
        RECT 46.335 103.365 46.505 103.505 ;
        RECT 45.180 103.325 46.145 103.335 ;
        RECT 44.840 103.155 45.010 103.245 ;
        RECT 45.470 103.165 46.145 103.325 ;
        RECT 42.880 102.965 43.620 102.995 ;
        RECT 42.880 102.665 43.795 102.965 ;
        RECT 43.470 102.490 43.795 102.665 ;
        RECT 42.500 101.935 42.755 102.465 ;
        RECT 42.925 101.755 43.230 102.215 ;
        RECT 43.475 102.135 43.795 102.490 ;
        RECT 43.965 102.705 44.505 103.075 ;
        RECT 44.840 102.985 45.245 103.155 ;
        RECT 43.965 102.305 44.205 102.705 ;
        RECT 44.685 102.535 44.905 102.815 ;
        RECT 44.375 102.365 44.905 102.535 ;
        RECT 44.375 102.135 44.545 102.365 ;
        RECT 45.075 102.205 45.245 102.985 ;
        RECT 45.415 102.375 45.765 102.995 ;
        RECT 45.935 102.375 46.145 103.165 ;
        RECT 46.335 103.195 47.835 103.365 ;
        RECT 46.335 102.505 46.505 103.195 ;
        RECT 48.195 103.025 48.365 103.805 ;
        RECT 49.170 103.675 49.340 103.805 ;
        RECT 46.675 102.855 48.365 103.025 ;
        RECT 48.535 103.245 49.000 103.635 ;
        RECT 49.170 103.505 49.565 103.675 ;
        RECT 46.675 102.675 46.845 102.855 ;
        RECT 43.475 101.965 44.545 102.135 ;
        RECT 44.715 101.755 44.905 102.195 ;
        RECT 45.075 101.925 46.025 102.205 ;
        RECT 46.335 102.115 46.595 102.505 ;
        RECT 47.015 102.435 47.805 102.685 ;
        RECT 46.245 101.945 46.595 102.115 ;
        RECT 46.805 101.755 47.135 102.215 ;
        RECT 48.010 102.145 48.180 102.855 ;
        RECT 48.535 102.655 48.705 103.245 ;
        RECT 48.350 102.435 48.705 102.655 ;
        RECT 48.875 102.435 49.225 103.055 ;
        RECT 49.395 102.145 49.565 103.505 ;
        RECT 49.930 103.335 50.255 104.120 ;
        RECT 49.735 102.285 50.195 103.335 ;
        RECT 48.010 101.975 48.865 102.145 ;
        RECT 49.070 101.975 49.565 102.145 ;
        RECT 49.735 101.755 50.065 102.115 ;
        RECT 50.425 102.015 50.595 104.135 ;
        RECT 50.765 103.805 51.095 104.305 ;
        RECT 51.265 103.635 51.520 104.135 ;
        RECT 50.770 103.465 51.520 103.635 ;
        RECT 50.770 102.475 51.000 103.465 ;
        RECT 51.170 102.645 51.520 103.295 ;
        RECT 51.695 103.140 51.985 104.305 ;
        RECT 52.155 103.215 53.825 104.305 ;
        RECT 52.155 102.695 52.905 103.215 ;
        RECT 54.055 103.165 54.265 104.305 ;
        RECT 54.435 103.155 54.765 104.135 ;
        RECT 54.935 103.165 55.165 104.305 ;
        RECT 55.835 103.215 57.505 104.305 ;
        RECT 53.075 102.525 53.825 103.045 ;
        RECT 50.770 102.305 51.520 102.475 ;
        RECT 50.765 101.755 51.095 102.135 ;
        RECT 51.265 102.015 51.520 102.305 ;
        RECT 51.695 101.755 51.985 102.480 ;
        RECT 52.155 101.755 53.825 102.525 ;
        RECT 54.055 101.755 54.265 102.575 ;
        RECT 54.435 102.555 54.685 103.155 ;
        RECT 54.855 102.745 55.185 102.995 ;
        RECT 55.835 102.695 56.585 103.215 ;
        RECT 57.715 103.165 57.945 104.305 ;
        RECT 58.115 103.155 58.445 104.135 ;
        RECT 58.615 103.165 58.825 104.305 ;
        RECT 59.095 103.165 59.325 104.305 ;
        RECT 59.495 103.155 59.825 104.135 ;
        RECT 59.995 103.165 60.205 104.305 ;
        RECT 60.440 103.635 60.695 104.135 ;
        RECT 60.865 103.805 61.195 104.305 ;
        RECT 60.440 103.465 61.190 103.635 ;
        RECT 54.435 101.925 54.765 102.555 ;
        RECT 54.935 101.755 55.165 102.575 ;
        RECT 56.755 102.525 57.505 103.045 ;
        RECT 57.695 102.745 58.025 102.995 ;
        RECT 55.835 101.755 57.505 102.525 ;
        RECT 57.715 101.755 57.945 102.575 ;
        RECT 58.195 102.555 58.445 103.155 ;
        RECT 59.075 102.745 59.405 102.995 ;
        RECT 58.115 101.925 58.445 102.555 ;
        RECT 58.615 101.755 58.825 102.575 ;
        RECT 59.095 101.755 59.325 102.575 ;
        RECT 59.575 102.555 59.825 103.155 ;
        RECT 60.440 102.645 60.790 103.295 ;
        RECT 59.495 101.925 59.825 102.555 ;
        RECT 59.995 101.755 60.205 102.575 ;
        RECT 60.960 102.475 61.190 103.465 ;
        RECT 60.440 102.305 61.190 102.475 ;
        RECT 60.440 102.015 60.695 102.305 ;
        RECT 60.865 101.755 61.195 102.135 ;
        RECT 61.365 102.015 61.535 104.135 ;
        RECT 61.705 103.335 62.030 104.120 ;
        RECT 62.200 103.845 62.450 104.305 ;
        RECT 62.620 103.805 62.870 104.135 ;
        RECT 63.085 103.805 63.765 104.135 ;
        RECT 62.620 103.675 62.790 103.805 ;
        RECT 62.395 103.505 62.790 103.675 ;
        RECT 61.765 102.285 62.225 103.335 ;
        RECT 62.395 102.145 62.565 103.505 ;
        RECT 62.960 103.245 63.425 103.635 ;
        RECT 62.735 102.435 63.085 103.055 ;
        RECT 63.255 102.655 63.425 103.245 ;
        RECT 63.595 103.025 63.765 103.805 ;
        RECT 63.935 103.705 64.105 104.045 ;
        RECT 64.340 103.875 64.670 104.305 ;
        RECT 64.840 103.705 65.010 104.045 ;
        RECT 65.305 103.845 65.675 104.305 ;
        RECT 63.935 103.535 65.010 103.705 ;
        RECT 65.845 103.675 66.015 104.135 ;
        RECT 66.250 103.795 67.120 104.135 ;
        RECT 67.290 103.845 67.540 104.305 ;
        RECT 65.455 103.505 66.015 103.675 ;
        RECT 65.455 103.365 65.625 103.505 ;
        RECT 64.125 103.195 65.625 103.365 ;
        RECT 66.320 103.335 66.780 103.625 ;
        RECT 63.595 102.855 65.285 103.025 ;
        RECT 63.255 102.435 63.610 102.655 ;
        RECT 63.780 102.145 63.950 102.855 ;
        RECT 64.155 102.435 64.945 102.685 ;
        RECT 65.115 102.675 65.285 102.855 ;
        RECT 65.455 102.505 65.625 103.195 ;
        RECT 61.895 101.755 62.225 102.115 ;
        RECT 62.395 101.975 62.890 102.145 ;
        RECT 63.095 101.975 63.950 102.145 ;
        RECT 64.825 101.755 65.155 102.215 ;
        RECT 65.365 102.115 65.625 102.505 ;
        RECT 65.815 103.325 66.780 103.335 ;
        RECT 66.950 103.415 67.120 103.795 ;
        RECT 67.710 103.755 67.880 104.045 ;
        RECT 68.060 103.925 68.390 104.305 ;
        RECT 67.710 103.585 68.510 103.755 ;
        RECT 65.815 103.165 66.490 103.325 ;
        RECT 66.950 103.245 68.170 103.415 ;
        RECT 65.815 102.375 66.025 103.165 ;
        RECT 66.950 103.155 67.120 103.245 ;
        RECT 66.195 102.375 66.545 102.995 ;
        RECT 66.715 102.985 67.120 103.155 ;
        RECT 66.715 102.205 66.885 102.985 ;
        RECT 67.055 102.535 67.275 102.815 ;
        RECT 67.455 102.705 67.995 103.075 ;
        RECT 68.340 102.995 68.510 103.585 ;
        RECT 68.730 103.165 69.035 104.305 ;
        RECT 69.205 103.115 69.460 103.995 ;
        RECT 68.340 102.965 69.080 102.995 ;
        RECT 67.055 102.365 67.585 102.535 ;
        RECT 65.365 101.945 65.715 102.115 ;
        RECT 65.935 101.925 66.885 102.205 ;
        RECT 67.055 101.755 67.245 102.195 ;
        RECT 67.415 102.135 67.585 102.365 ;
        RECT 67.755 102.305 67.995 102.705 ;
        RECT 68.165 102.665 69.080 102.965 ;
        RECT 68.165 102.490 68.490 102.665 ;
        RECT 68.165 102.135 68.485 102.490 ;
        RECT 69.250 102.465 69.460 103.115 ;
        RECT 69.635 103.215 70.845 104.305 ;
        RECT 71.015 103.215 74.525 104.305 ;
        RECT 69.635 102.675 70.155 103.215 ;
        RECT 70.325 102.505 70.845 103.045 ;
        RECT 71.015 102.695 72.705 103.215 ;
        RECT 74.755 103.165 74.965 104.305 ;
        RECT 75.135 103.155 75.465 104.135 ;
        RECT 75.635 103.165 75.865 104.305 ;
        RECT 76.135 103.165 76.345 104.305 ;
        RECT 76.515 103.155 76.845 104.135 ;
        RECT 77.015 103.165 77.245 104.305 ;
        RECT 72.875 102.525 74.525 103.045 ;
        RECT 67.415 101.965 68.485 102.135 ;
        RECT 68.730 101.755 69.035 102.215 ;
        RECT 69.205 101.935 69.460 102.465 ;
        RECT 69.635 101.755 70.845 102.505 ;
        RECT 71.015 101.755 74.525 102.525 ;
        RECT 74.755 101.755 74.965 102.575 ;
        RECT 75.135 102.555 75.385 103.155 ;
        RECT 75.555 102.745 75.885 102.995 ;
        RECT 75.135 101.925 75.465 102.555 ;
        RECT 75.635 101.755 75.865 102.575 ;
        RECT 76.135 101.755 76.345 102.575 ;
        RECT 76.515 102.555 76.765 103.155 ;
        RECT 77.455 103.140 77.745 104.305 ;
        RECT 78.005 103.375 78.175 104.135 ;
        RECT 78.355 103.545 78.685 104.305 ;
        RECT 78.005 103.205 78.670 103.375 ;
        RECT 78.855 103.230 79.125 104.135 ;
        RECT 78.500 103.060 78.670 103.205 ;
        RECT 76.935 102.745 77.265 102.995 ;
        RECT 77.935 102.655 78.265 103.025 ;
        RECT 78.500 102.730 78.785 103.060 ;
        RECT 76.515 101.925 76.845 102.555 ;
        RECT 77.015 101.755 77.245 102.575 ;
        RECT 77.455 101.755 77.745 102.480 ;
        RECT 78.500 102.475 78.670 102.730 ;
        RECT 78.005 102.305 78.670 102.475 ;
        RECT 78.955 102.430 79.125 103.230 ;
        RECT 79.385 103.375 79.555 104.135 ;
        RECT 79.735 103.545 80.065 104.305 ;
        RECT 79.385 103.205 80.050 103.375 ;
        RECT 80.235 103.230 80.505 104.135 ;
        RECT 79.880 103.060 80.050 103.205 ;
        RECT 79.315 102.655 79.645 103.025 ;
        RECT 79.880 102.730 80.165 103.060 ;
        RECT 79.880 102.475 80.050 102.730 ;
        RECT 78.005 101.925 78.175 102.305 ;
        RECT 78.355 101.755 78.685 102.135 ;
        RECT 78.865 101.925 79.125 102.430 ;
        RECT 79.385 102.305 80.050 102.475 ;
        RECT 80.335 102.430 80.505 103.230 ;
        RECT 80.675 103.215 84.185 104.305 ;
        RECT 80.675 102.695 82.365 103.215 ;
        RECT 84.415 103.165 84.625 104.305 ;
        RECT 84.795 103.155 85.125 104.135 ;
        RECT 85.295 103.165 85.525 104.305 ;
        RECT 85.825 103.375 85.995 104.135 ;
        RECT 86.175 103.545 86.505 104.305 ;
        RECT 85.825 103.205 86.490 103.375 ;
        RECT 86.675 103.230 86.945 104.135 ;
        RECT 82.535 102.525 84.185 103.045 ;
        RECT 79.385 101.925 79.555 102.305 ;
        RECT 79.735 101.755 80.065 102.135 ;
        RECT 80.245 101.925 80.505 102.430 ;
        RECT 80.675 101.755 84.185 102.525 ;
        RECT 84.415 101.755 84.625 102.575 ;
        RECT 84.795 102.555 85.045 103.155 ;
        RECT 86.320 103.060 86.490 103.205 ;
        RECT 85.215 102.745 85.545 102.995 ;
        RECT 85.755 102.655 86.085 103.025 ;
        RECT 86.320 102.730 86.605 103.060 ;
        RECT 84.795 101.925 85.125 102.555 ;
        RECT 85.295 101.755 85.525 102.575 ;
        RECT 86.320 102.475 86.490 102.730 ;
        RECT 85.825 102.305 86.490 102.475 ;
        RECT 86.775 102.430 86.945 103.230 ;
        RECT 87.155 103.165 87.385 104.305 ;
        RECT 87.555 103.155 87.885 104.135 ;
        RECT 88.055 103.165 88.265 104.305 ;
        RECT 87.135 102.745 87.465 102.995 ;
        RECT 85.825 101.925 85.995 102.305 ;
        RECT 86.175 101.755 86.505 102.135 ;
        RECT 86.685 101.925 86.945 102.430 ;
        RECT 87.155 101.755 87.385 102.575 ;
        RECT 87.635 102.555 87.885 103.155 ;
        RECT 88.500 103.115 88.755 103.995 ;
        RECT 88.925 103.165 89.230 104.305 ;
        RECT 89.570 103.925 89.900 104.305 ;
        RECT 90.080 103.755 90.250 104.045 ;
        RECT 90.420 103.845 90.670 104.305 ;
        RECT 89.450 103.585 90.250 103.755 ;
        RECT 90.840 103.795 91.710 104.135 ;
        RECT 87.555 101.925 87.885 102.555 ;
        RECT 88.055 101.755 88.265 102.575 ;
        RECT 88.500 102.465 88.710 103.115 ;
        RECT 89.450 102.995 89.620 103.585 ;
        RECT 90.840 103.415 91.010 103.795 ;
        RECT 91.945 103.675 92.115 104.135 ;
        RECT 92.285 103.845 92.655 104.305 ;
        RECT 92.950 103.705 93.120 104.045 ;
        RECT 93.290 103.875 93.620 104.305 ;
        RECT 93.855 103.705 94.025 104.045 ;
        RECT 89.790 103.245 91.010 103.415 ;
        RECT 91.180 103.335 91.640 103.625 ;
        RECT 91.945 103.505 92.505 103.675 ;
        RECT 92.950 103.535 94.025 103.705 ;
        RECT 94.195 103.805 94.875 104.135 ;
        RECT 95.090 103.805 95.340 104.135 ;
        RECT 95.510 103.845 95.760 104.305 ;
        RECT 92.335 103.365 92.505 103.505 ;
        RECT 91.180 103.325 92.145 103.335 ;
        RECT 90.840 103.155 91.010 103.245 ;
        RECT 91.470 103.165 92.145 103.325 ;
        RECT 88.880 102.965 89.620 102.995 ;
        RECT 88.880 102.665 89.795 102.965 ;
        RECT 89.470 102.490 89.795 102.665 ;
        RECT 88.500 101.935 88.755 102.465 ;
        RECT 88.925 101.755 89.230 102.215 ;
        RECT 89.475 102.135 89.795 102.490 ;
        RECT 89.965 102.705 90.505 103.075 ;
        RECT 90.840 102.985 91.245 103.155 ;
        RECT 89.965 102.305 90.205 102.705 ;
        RECT 90.685 102.535 90.905 102.815 ;
        RECT 90.375 102.365 90.905 102.535 ;
        RECT 90.375 102.135 90.545 102.365 ;
        RECT 91.075 102.205 91.245 102.985 ;
        RECT 91.415 102.375 91.765 102.995 ;
        RECT 91.935 102.375 92.145 103.165 ;
        RECT 92.335 103.195 93.835 103.365 ;
        RECT 92.335 102.505 92.505 103.195 ;
        RECT 94.195 103.025 94.365 103.805 ;
        RECT 95.170 103.675 95.340 103.805 ;
        RECT 92.675 102.855 94.365 103.025 ;
        RECT 94.535 103.245 95.000 103.635 ;
        RECT 95.170 103.505 95.565 103.675 ;
        RECT 92.675 102.675 92.845 102.855 ;
        RECT 89.475 101.965 90.545 102.135 ;
        RECT 90.715 101.755 90.905 102.195 ;
        RECT 91.075 101.925 92.025 102.205 ;
        RECT 92.335 102.115 92.595 102.505 ;
        RECT 93.015 102.435 93.805 102.685 ;
        RECT 92.245 101.945 92.595 102.115 ;
        RECT 92.805 101.755 93.135 102.215 ;
        RECT 94.010 102.145 94.180 102.855 ;
        RECT 94.535 102.655 94.705 103.245 ;
        RECT 94.350 102.435 94.705 102.655 ;
        RECT 94.875 102.435 95.225 103.055 ;
        RECT 95.395 102.145 95.565 103.505 ;
        RECT 95.930 103.335 96.255 104.120 ;
        RECT 95.735 102.285 96.195 103.335 ;
        RECT 94.010 101.975 94.865 102.145 ;
        RECT 95.070 101.975 95.565 102.145 ;
        RECT 95.735 101.755 96.065 102.115 ;
        RECT 96.425 102.015 96.595 104.135 ;
        RECT 96.765 103.805 97.095 104.305 ;
        RECT 97.265 103.635 97.520 104.135 ;
        RECT 96.770 103.465 97.520 103.635 ;
        RECT 96.770 102.475 97.000 103.465 ;
        RECT 97.170 102.645 97.520 103.295 ;
        RECT 97.755 103.165 97.965 104.305 ;
        RECT 98.135 103.155 98.465 104.135 ;
        RECT 98.635 103.165 98.865 104.305 ;
        RECT 99.075 103.215 101.665 104.305 ;
        RECT 96.770 102.305 97.520 102.475 ;
        RECT 96.765 101.755 97.095 102.135 ;
        RECT 97.265 102.015 97.520 102.305 ;
        RECT 97.755 101.755 97.965 102.575 ;
        RECT 98.135 102.555 98.385 103.155 ;
        RECT 98.555 102.745 98.885 102.995 ;
        RECT 99.075 102.695 100.285 103.215 ;
        RECT 101.875 103.165 102.105 104.305 ;
        RECT 102.275 103.155 102.605 104.135 ;
        RECT 102.775 103.165 102.985 104.305 ;
        RECT 98.135 101.925 98.465 102.555 ;
        RECT 98.635 101.755 98.865 102.575 ;
        RECT 100.455 102.525 101.665 103.045 ;
        RECT 101.855 102.745 102.185 102.995 ;
        RECT 99.075 101.755 101.665 102.525 ;
        RECT 101.875 101.755 102.105 102.575 ;
        RECT 102.355 102.555 102.605 103.155 ;
        RECT 103.215 103.140 103.505 104.305 ;
        RECT 104.600 103.635 104.855 104.135 ;
        RECT 105.025 103.805 105.355 104.305 ;
        RECT 104.600 103.465 105.350 103.635 ;
        RECT 104.600 102.645 104.950 103.295 ;
        RECT 102.275 101.925 102.605 102.555 ;
        RECT 102.775 101.755 102.985 102.575 ;
        RECT 103.215 101.755 103.505 102.480 ;
        RECT 105.120 102.475 105.350 103.465 ;
        RECT 104.600 102.305 105.350 102.475 ;
        RECT 104.600 102.015 104.855 102.305 ;
        RECT 105.025 101.755 105.355 102.135 ;
        RECT 105.525 102.015 105.695 104.135 ;
        RECT 105.865 103.335 106.190 104.120 ;
        RECT 106.360 103.845 106.610 104.305 ;
        RECT 106.780 103.805 107.030 104.135 ;
        RECT 107.245 103.805 107.925 104.135 ;
        RECT 106.780 103.675 106.950 103.805 ;
        RECT 106.555 103.505 106.950 103.675 ;
        RECT 105.925 102.285 106.385 103.335 ;
        RECT 106.555 102.145 106.725 103.505 ;
        RECT 107.120 103.245 107.585 103.635 ;
        RECT 106.895 102.435 107.245 103.055 ;
        RECT 107.415 102.655 107.585 103.245 ;
        RECT 107.755 103.025 107.925 103.805 ;
        RECT 108.095 103.705 108.265 104.045 ;
        RECT 108.500 103.875 108.830 104.305 ;
        RECT 109.000 103.705 109.170 104.045 ;
        RECT 109.465 103.845 109.835 104.305 ;
        RECT 108.095 103.535 109.170 103.705 ;
        RECT 110.005 103.675 110.175 104.135 ;
        RECT 110.410 103.795 111.280 104.135 ;
        RECT 111.450 103.845 111.700 104.305 ;
        RECT 109.615 103.505 110.175 103.675 ;
        RECT 109.615 103.365 109.785 103.505 ;
        RECT 108.285 103.195 109.785 103.365 ;
        RECT 110.480 103.335 110.940 103.625 ;
        RECT 107.755 102.855 109.445 103.025 ;
        RECT 107.415 102.435 107.770 102.655 ;
        RECT 107.940 102.145 108.110 102.855 ;
        RECT 108.315 102.435 109.105 102.685 ;
        RECT 109.275 102.675 109.445 102.855 ;
        RECT 109.615 102.505 109.785 103.195 ;
        RECT 106.055 101.755 106.385 102.115 ;
        RECT 106.555 101.975 107.050 102.145 ;
        RECT 107.255 101.975 108.110 102.145 ;
        RECT 108.985 101.755 109.315 102.215 ;
        RECT 109.525 102.115 109.785 102.505 ;
        RECT 109.975 103.325 110.940 103.335 ;
        RECT 111.110 103.415 111.280 103.795 ;
        RECT 111.870 103.755 112.040 104.045 ;
        RECT 112.220 103.925 112.550 104.305 ;
        RECT 111.870 103.585 112.670 103.755 ;
        RECT 109.975 103.165 110.650 103.325 ;
        RECT 111.110 103.245 112.330 103.415 ;
        RECT 109.975 102.375 110.185 103.165 ;
        RECT 111.110 103.155 111.280 103.245 ;
        RECT 110.355 102.375 110.705 102.995 ;
        RECT 110.875 102.985 111.280 103.155 ;
        RECT 110.875 102.205 111.045 102.985 ;
        RECT 111.215 102.535 111.435 102.815 ;
        RECT 111.615 102.705 112.155 103.075 ;
        RECT 112.500 102.995 112.670 103.585 ;
        RECT 112.890 103.165 113.195 104.305 ;
        RECT 113.365 103.115 113.620 103.995 ;
        RECT 112.500 102.965 113.240 102.995 ;
        RECT 111.215 102.365 111.745 102.535 ;
        RECT 109.525 101.945 109.875 102.115 ;
        RECT 110.095 101.925 111.045 102.205 ;
        RECT 111.215 101.755 111.405 102.195 ;
        RECT 111.575 102.135 111.745 102.365 ;
        RECT 111.915 102.305 112.155 102.705 ;
        RECT 112.325 102.665 113.240 102.965 ;
        RECT 112.325 102.490 112.650 102.665 ;
        RECT 112.325 102.135 112.645 102.490 ;
        RECT 113.410 102.465 113.620 103.115 ;
        RECT 113.795 103.215 115.465 104.305 ;
        RECT 113.795 102.695 114.545 103.215 ;
        RECT 115.675 103.165 115.905 104.305 ;
        RECT 116.075 103.155 116.405 104.135 ;
        RECT 116.575 103.165 116.785 104.305 ;
        RECT 117.515 103.165 117.745 104.305 ;
        RECT 117.915 103.155 118.245 104.135 ;
        RECT 118.415 103.165 118.625 104.305 ;
        RECT 118.860 103.635 119.115 104.135 ;
        RECT 119.285 103.805 119.615 104.305 ;
        RECT 118.860 103.465 119.610 103.635 ;
        RECT 114.715 102.525 115.465 103.045 ;
        RECT 115.655 102.745 115.985 102.995 ;
        RECT 111.575 101.965 112.645 102.135 ;
        RECT 112.890 101.755 113.195 102.215 ;
        RECT 113.365 101.935 113.620 102.465 ;
        RECT 113.795 101.755 115.465 102.525 ;
        RECT 115.675 101.755 115.905 102.575 ;
        RECT 116.155 102.555 116.405 103.155 ;
        RECT 117.495 102.745 117.825 102.995 ;
        RECT 116.075 101.925 116.405 102.555 ;
        RECT 116.575 101.755 116.785 102.575 ;
        RECT 117.515 101.755 117.745 102.575 ;
        RECT 117.995 102.555 118.245 103.155 ;
        RECT 118.860 102.645 119.210 103.295 ;
        RECT 117.915 101.925 118.245 102.555 ;
        RECT 118.415 101.755 118.625 102.575 ;
        RECT 119.380 102.475 119.610 103.465 ;
        RECT 118.860 102.305 119.610 102.475 ;
        RECT 118.860 102.015 119.115 102.305 ;
        RECT 119.285 101.755 119.615 102.135 ;
        RECT 119.785 102.015 119.955 104.135 ;
        RECT 120.125 103.335 120.450 104.120 ;
        RECT 120.620 103.845 120.870 104.305 ;
        RECT 121.040 103.805 121.290 104.135 ;
        RECT 121.505 103.805 122.185 104.135 ;
        RECT 121.040 103.675 121.210 103.805 ;
        RECT 120.815 103.505 121.210 103.675 ;
        RECT 120.185 102.285 120.645 103.335 ;
        RECT 120.815 102.145 120.985 103.505 ;
        RECT 121.380 103.245 121.845 103.635 ;
        RECT 121.155 102.435 121.505 103.055 ;
        RECT 121.675 102.655 121.845 103.245 ;
        RECT 122.015 103.025 122.185 103.805 ;
        RECT 122.355 103.705 122.525 104.045 ;
        RECT 122.760 103.875 123.090 104.305 ;
        RECT 123.260 103.705 123.430 104.045 ;
        RECT 123.725 103.845 124.095 104.305 ;
        RECT 122.355 103.535 123.430 103.705 ;
        RECT 124.265 103.675 124.435 104.135 ;
        RECT 124.670 103.795 125.540 104.135 ;
        RECT 125.710 103.845 125.960 104.305 ;
        RECT 123.875 103.505 124.435 103.675 ;
        RECT 123.875 103.365 124.045 103.505 ;
        RECT 122.545 103.195 124.045 103.365 ;
        RECT 124.740 103.335 125.200 103.625 ;
        RECT 122.015 102.855 123.705 103.025 ;
        RECT 121.675 102.435 122.030 102.655 ;
        RECT 122.200 102.145 122.370 102.855 ;
        RECT 122.575 102.435 123.365 102.685 ;
        RECT 123.535 102.675 123.705 102.855 ;
        RECT 123.875 102.505 124.045 103.195 ;
        RECT 120.315 101.755 120.645 102.115 ;
        RECT 120.815 101.975 121.310 102.145 ;
        RECT 121.515 101.975 122.370 102.145 ;
        RECT 123.245 101.755 123.575 102.215 ;
        RECT 123.785 102.115 124.045 102.505 ;
        RECT 124.235 103.325 125.200 103.335 ;
        RECT 125.370 103.415 125.540 103.795 ;
        RECT 126.130 103.755 126.300 104.045 ;
        RECT 126.480 103.925 126.810 104.305 ;
        RECT 126.130 103.585 126.930 103.755 ;
        RECT 124.235 103.165 124.910 103.325 ;
        RECT 125.370 103.245 126.590 103.415 ;
        RECT 124.235 102.375 124.445 103.165 ;
        RECT 125.370 103.155 125.540 103.245 ;
        RECT 124.615 102.375 124.965 102.995 ;
        RECT 125.135 102.985 125.540 103.155 ;
        RECT 125.135 102.205 125.305 102.985 ;
        RECT 125.475 102.535 125.695 102.815 ;
        RECT 125.875 102.705 126.415 103.075 ;
        RECT 126.760 102.995 126.930 103.585 ;
        RECT 127.150 103.165 127.455 104.305 ;
        RECT 127.625 103.115 127.880 103.995 ;
        RECT 126.760 102.965 127.500 102.995 ;
        RECT 125.475 102.365 126.005 102.535 ;
        RECT 123.785 101.945 124.135 102.115 ;
        RECT 124.355 101.925 125.305 102.205 ;
        RECT 125.475 101.755 125.665 102.195 ;
        RECT 125.835 102.135 126.005 102.365 ;
        RECT 126.175 102.305 126.415 102.705 ;
        RECT 126.585 102.665 127.500 102.965 ;
        RECT 126.585 102.490 126.910 102.665 ;
        RECT 126.585 102.135 126.905 102.490 ;
        RECT 127.670 102.465 127.880 103.115 ;
        RECT 128.055 103.215 129.265 104.305 ;
        RECT 128.055 102.675 128.575 103.215 ;
        RECT 128.745 102.505 129.265 103.045 ;
        RECT 125.835 101.965 126.905 102.135 ;
        RECT 127.150 101.755 127.455 102.215 ;
        RECT 127.625 101.935 127.880 102.465 ;
        RECT 128.055 101.755 129.265 102.505 ;
        RECT 9.290 101.585 129.350 101.755 ;
        RECT 9.375 100.835 10.585 101.585 ;
        RECT 9.375 100.295 9.895 100.835 ;
        RECT 11.215 100.815 12.885 101.585 ;
        RECT 13.055 100.860 13.345 101.585 ;
        RECT 13.520 101.040 18.865 101.585 ;
        RECT 10.065 100.125 10.585 100.665 ;
        RECT 9.375 99.035 10.585 100.125 ;
        RECT 11.215 100.125 11.965 100.645 ;
        RECT 12.135 100.295 12.885 100.815 ;
        RECT 11.215 99.035 12.885 100.125 ;
        RECT 13.055 99.035 13.345 100.200 ;
        RECT 15.110 99.470 15.460 100.720 ;
        RECT 16.940 100.210 17.280 101.040 ;
        RECT 19.075 100.765 19.305 101.585 ;
        RECT 19.475 100.785 19.805 101.415 ;
        RECT 19.055 100.345 19.385 100.595 ;
        RECT 19.555 100.185 19.805 100.785 ;
        RECT 19.975 100.765 20.185 101.585 ;
        RECT 20.420 101.035 20.675 101.325 ;
        RECT 20.845 101.205 21.175 101.585 ;
        RECT 20.420 100.865 21.170 101.035 ;
        RECT 13.520 99.035 18.865 99.470 ;
        RECT 19.075 99.035 19.305 100.175 ;
        RECT 19.475 99.205 19.805 100.185 ;
        RECT 19.975 99.035 20.185 100.175 ;
        RECT 20.420 100.045 20.770 100.695 ;
        RECT 20.940 99.875 21.170 100.865 ;
        RECT 20.420 99.705 21.170 99.875 ;
        RECT 20.420 99.205 20.675 99.705 ;
        RECT 20.845 99.035 21.175 99.535 ;
        RECT 21.345 99.205 21.515 101.325 ;
        RECT 21.875 101.225 22.205 101.585 ;
        RECT 22.375 101.195 22.870 101.365 ;
        RECT 23.075 101.195 23.930 101.365 ;
        RECT 21.745 100.005 22.205 101.055 ;
        RECT 21.685 99.220 22.010 100.005 ;
        RECT 22.375 99.835 22.545 101.195 ;
        RECT 22.715 100.285 23.065 100.905 ;
        RECT 23.235 100.685 23.590 100.905 ;
        RECT 23.235 100.095 23.405 100.685 ;
        RECT 23.760 100.485 23.930 101.195 ;
        RECT 24.805 101.125 25.135 101.585 ;
        RECT 25.345 101.225 25.695 101.395 ;
        RECT 24.135 100.655 24.925 100.905 ;
        RECT 25.345 100.835 25.605 101.225 ;
        RECT 25.915 101.135 26.865 101.415 ;
        RECT 27.035 101.145 27.225 101.585 ;
        RECT 27.395 101.205 28.465 101.375 ;
        RECT 25.095 100.485 25.265 100.665 ;
        RECT 22.375 99.665 22.770 99.835 ;
        RECT 22.940 99.705 23.405 100.095 ;
        RECT 23.575 100.315 25.265 100.485 ;
        RECT 22.600 99.535 22.770 99.665 ;
        RECT 23.575 99.535 23.745 100.315 ;
        RECT 25.435 100.145 25.605 100.835 ;
        RECT 24.105 99.975 25.605 100.145 ;
        RECT 25.795 100.175 26.005 100.965 ;
        RECT 26.175 100.345 26.525 100.965 ;
        RECT 26.695 100.355 26.865 101.135 ;
        RECT 27.395 100.975 27.565 101.205 ;
        RECT 27.035 100.805 27.565 100.975 ;
        RECT 27.035 100.525 27.255 100.805 ;
        RECT 27.735 100.635 27.975 101.035 ;
        RECT 26.695 100.185 27.100 100.355 ;
        RECT 27.435 100.265 27.975 100.635 ;
        RECT 28.145 100.850 28.465 101.205 ;
        RECT 28.710 101.125 29.015 101.585 ;
        RECT 29.185 100.875 29.440 101.405 ;
        RECT 28.145 100.675 28.470 100.850 ;
        RECT 28.145 100.375 29.060 100.675 ;
        RECT 28.320 100.345 29.060 100.375 ;
        RECT 25.795 100.015 26.470 100.175 ;
        RECT 26.930 100.095 27.100 100.185 ;
        RECT 25.795 100.005 26.760 100.015 ;
        RECT 25.435 99.835 25.605 99.975 ;
        RECT 22.180 99.035 22.430 99.495 ;
        RECT 22.600 99.205 22.850 99.535 ;
        RECT 23.065 99.205 23.745 99.535 ;
        RECT 23.915 99.635 24.990 99.805 ;
        RECT 25.435 99.665 25.995 99.835 ;
        RECT 26.300 99.715 26.760 100.005 ;
        RECT 26.930 99.925 28.150 100.095 ;
        RECT 23.915 99.295 24.085 99.635 ;
        RECT 24.320 99.035 24.650 99.465 ;
        RECT 24.820 99.295 24.990 99.635 ;
        RECT 25.285 99.035 25.655 99.495 ;
        RECT 25.825 99.205 25.995 99.665 ;
        RECT 26.930 99.545 27.100 99.925 ;
        RECT 28.320 99.755 28.490 100.345 ;
        RECT 29.230 100.225 29.440 100.875 ;
        RECT 26.230 99.205 27.100 99.545 ;
        RECT 27.690 99.585 28.490 99.755 ;
        RECT 27.270 99.035 27.520 99.495 ;
        RECT 27.690 99.295 27.860 99.585 ;
        RECT 28.040 99.035 28.370 99.415 ;
        RECT 28.710 99.035 29.015 100.175 ;
        RECT 29.185 99.345 29.440 100.225 ;
        RECT 29.620 100.875 29.875 101.405 ;
        RECT 30.045 101.125 30.350 101.585 ;
        RECT 30.595 101.205 31.665 101.375 ;
        RECT 29.620 100.225 29.830 100.875 ;
        RECT 30.595 100.850 30.915 101.205 ;
        RECT 30.590 100.675 30.915 100.850 ;
        RECT 30.000 100.375 30.915 100.675 ;
        RECT 31.085 100.635 31.325 101.035 ;
        RECT 31.495 100.975 31.665 101.205 ;
        RECT 31.835 101.145 32.025 101.585 ;
        RECT 32.195 101.135 33.145 101.415 ;
        RECT 33.365 101.225 33.715 101.395 ;
        RECT 31.495 100.805 32.025 100.975 ;
        RECT 30.000 100.345 30.740 100.375 ;
        RECT 29.620 99.345 29.875 100.225 ;
        RECT 30.045 99.035 30.350 100.175 ;
        RECT 30.570 99.755 30.740 100.345 ;
        RECT 31.085 100.265 31.625 100.635 ;
        RECT 31.805 100.525 32.025 100.805 ;
        RECT 32.195 100.355 32.365 101.135 ;
        RECT 31.960 100.185 32.365 100.355 ;
        RECT 32.535 100.345 32.885 100.965 ;
        RECT 31.960 100.095 32.130 100.185 ;
        RECT 33.055 100.175 33.265 100.965 ;
        RECT 30.910 99.925 32.130 100.095 ;
        RECT 32.590 100.015 33.265 100.175 ;
        RECT 30.570 99.585 31.370 99.755 ;
        RECT 30.690 99.035 31.020 99.415 ;
        RECT 31.200 99.295 31.370 99.585 ;
        RECT 31.960 99.545 32.130 99.925 ;
        RECT 32.300 100.005 33.265 100.015 ;
        RECT 33.455 100.835 33.715 101.225 ;
        RECT 33.925 101.125 34.255 101.585 ;
        RECT 35.130 101.195 35.985 101.365 ;
        RECT 36.190 101.195 36.685 101.365 ;
        RECT 36.855 101.225 37.185 101.585 ;
        RECT 33.455 100.145 33.625 100.835 ;
        RECT 33.795 100.485 33.965 100.665 ;
        RECT 34.135 100.655 34.925 100.905 ;
        RECT 35.130 100.485 35.300 101.195 ;
        RECT 35.470 100.685 35.825 100.905 ;
        RECT 33.795 100.315 35.485 100.485 ;
        RECT 32.300 99.715 32.760 100.005 ;
        RECT 33.455 99.975 34.955 100.145 ;
        RECT 33.455 99.835 33.625 99.975 ;
        RECT 33.065 99.665 33.625 99.835 ;
        RECT 31.540 99.035 31.790 99.495 ;
        RECT 31.960 99.205 32.830 99.545 ;
        RECT 33.065 99.205 33.235 99.665 ;
        RECT 34.070 99.635 35.145 99.805 ;
        RECT 33.405 99.035 33.775 99.495 ;
        RECT 34.070 99.295 34.240 99.635 ;
        RECT 34.410 99.035 34.740 99.465 ;
        RECT 34.975 99.295 35.145 99.635 ;
        RECT 35.315 99.535 35.485 100.315 ;
        RECT 35.655 100.095 35.825 100.685 ;
        RECT 35.995 100.285 36.345 100.905 ;
        RECT 35.655 99.705 36.120 100.095 ;
        RECT 36.515 99.835 36.685 101.195 ;
        RECT 36.855 100.005 37.315 101.055 ;
        RECT 36.290 99.665 36.685 99.835 ;
        RECT 36.290 99.535 36.460 99.665 ;
        RECT 35.315 99.205 35.995 99.535 ;
        RECT 36.210 99.205 36.460 99.535 ;
        RECT 36.630 99.035 36.880 99.495 ;
        RECT 37.050 99.220 37.375 100.005 ;
        RECT 37.545 99.205 37.715 101.325 ;
        RECT 37.885 101.205 38.215 101.585 ;
        RECT 38.385 101.035 38.640 101.325 ;
        RECT 37.890 100.865 38.640 101.035 ;
        RECT 37.890 99.875 38.120 100.865 ;
        RECT 38.815 100.860 39.105 101.585 ;
        RECT 39.280 101.040 44.625 101.585 ;
        RECT 38.290 100.045 38.640 100.695 ;
        RECT 37.890 99.705 38.640 99.875 ;
        RECT 37.885 99.035 38.215 99.535 ;
        RECT 38.385 99.205 38.640 99.705 ;
        RECT 38.815 99.035 39.105 100.200 ;
        RECT 40.870 99.470 41.220 100.720 ;
        RECT 42.700 100.210 43.040 101.040 ;
        RECT 44.835 100.765 45.065 101.585 ;
        RECT 45.235 100.785 45.565 101.415 ;
        RECT 44.815 100.345 45.145 100.595 ;
        RECT 45.315 100.185 45.565 100.785 ;
        RECT 45.735 100.765 45.945 101.585 ;
        RECT 46.180 101.035 46.435 101.325 ;
        RECT 46.605 101.205 46.935 101.585 ;
        RECT 46.180 100.865 46.930 101.035 ;
        RECT 39.280 99.035 44.625 99.470 ;
        RECT 44.835 99.035 45.065 100.175 ;
        RECT 45.235 99.205 45.565 100.185 ;
        RECT 45.735 99.035 45.945 100.175 ;
        RECT 46.180 100.045 46.530 100.695 ;
        RECT 46.700 99.875 46.930 100.865 ;
        RECT 46.180 99.705 46.930 99.875 ;
        RECT 46.180 99.205 46.435 99.705 ;
        RECT 46.605 99.035 46.935 99.535 ;
        RECT 47.105 99.205 47.275 101.325 ;
        RECT 47.635 101.225 47.965 101.585 ;
        RECT 48.135 101.195 48.630 101.365 ;
        RECT 48.835 101.195 49.690 101.365 ;
        RECT 47.505 100.005 47.965 101.055 ;
        RECT 47.445 99.220 47.770 100.005 ;
        RECT 48.135 99.835 48.305 101.195 ;
        RECT 48.475 100.285 48.825 100.905 ;
        RECT 48.995 100.685 49.350 100.905 ;
        RECT 48.995 100.095 49.165 100.685 ;
        RECT 49.520 100.485 49.690 101.195 ;
        RECT 50.565 101.125 50.895 101.585 ;
        RECT 51.105 101.225 51.455 101.395 ;
        RECT 49.895 100.655 50.685 100.905 ;
        RECT 51.105 100.835 51.365 101.225 ;
        RECT 51.675 101.135 52.625 101.415 ;
        RECT 52.795 101.145 52.985 101.585 ;
        RECT 53.155 101.205 54.225 101.375 ;
        RECT 50.855 100.485 51.025 100.665 ;
        RECT 48.135 99.665 48.530 99.835 ;
        RECT 48.700 99.705 49.165 100.095 ;
        RECT 49.335 100.315 51.025 100.485 ;
        RECT 48.360 99.535 48.530 99.665 ;
        RECT 49.335 99.535 49.505 100.315 ;
        RECT 51.195 100.145 51.365 100.835 ;
        RECT 49.865 99.975 51.365 100.145 ;
        RECT 51.555 100.175 51.765 100.965 ;
        RECT 51.935 100.345 52.285 100.965 ;
        RECT 52.455 100.355 52.625 101.135 ;
        RECT 53.155 100.975 53.325 101.205 ;
        RECT 52.795 100.805 53.325 100.975 ;
        RECT 52.795 100.525 53.015 100.805 ;
        RECT 53.495 100.635 53.735 101.035 ;
        RECT 52.455 100.185 52.860 100.355 ;
        RECT 53.195 100.265 53.735 100.635 ;
        RECT 53.905 100.850 54.225 101.205 ;
        RECT 54.470 101.125 54.775 101.585 ;
        RECT 54.945 100.875 55.200 101.405 ;
        RECT 53.905 100.675 54.230 100.850 ;
        RECT 53.905 100.375 54.820 100.675 ;
        RECT 54.080 100.345 54.820 100.375 ;
        RECT 51.555 100.015 52.230 100.175 ;
        RECT 52.690 100.095 52.860 100.185 ;
        RECT 51.555 100.005 52.520 100.015 ;
        RECT 51.195 99.835 51.365 99.975 ;
        RECT 47.940 99.035 48.190 99.495 ;
        RECT 48.360 99.205 48.610 99.535 ;
        RECT 48.825 99.205 49.505 99.535 ;
        RECT 49.675 99.635 50.750 99.805 ;
        RECT 51.195 99.665 51.755 99.835 ;
        RECT 52.060 99.715 52.520 100.005 ;
        RECT 52.690 99.925 53.910 100.095 ;
        RECT 49.675 99.295 49.845 99.635 ;
        RECT 50.080 99.035 50.410 99.465 ;
        RECT 50.580 99.295 50.750 99.635 ;
        RECT 51.045 99.035 51.415 99.495 ;
        RECT 51.585 99.205 51.755 99.665 ;
        RECT 52.690 99.545 52.860 99.925 ;
        RECT 54.080 99.755 54.250 100.345 ;
        RECT 54.990 100.225 55.200 100.875 ;
        RECT 51.990 99.205 52.860 99.545 ;
        RECT 53.450 99.585 54.250 99.755 ;
        RECT 53.030 99.035 53.280 99.495 ;
        RECT 53.450 99.295 53.620 99.585 ;
        RECT 53.800 99.035 54.130 99.415 ;
        RECT 54.470 99.035 54.775 100.175 ;
        RECT 54.945 99.345 55.200 100.225 ;
        RECT 55.380 100.875 55.635 101.405 ;
        RECT 55.805 101.125 56.110 101.585 ;
        RECT 56.355 101.205 57.425 101.375 ;
        RECT 55.380 100.225 55.590 100.875 ;
        RECT 56.355 100.850 56.675 101.205 ;
        RECT 56.350 100.675 56.675 100.850 ;
        RECT 55.760 100.375 56.675 100.675 ;
        RECT 56.845 100.635 57.085 101.035 ;
        RECT 57.255 100.975 57.425 101.205 ;
        RECT 57.595 101.145 57.785 101.585 ;
        RECT 57.955 101.135 58.905 101.415 ;
        RECT 59.125 101.225 59.475 101.395 ;
        RECT 57.255 100.805 57.785 100.975 ;
        RECT 55.760 100.345 56.500 100.375 ;
        RECT 55.380 99.345 55.635 100.225 ;
        RECT 55.805 99.035 56.110 100.175 ;
        RECT 56.330 99.755 56.500 100.345 ;
        RECT 56.845 100.265 57.385 100.635 ;
        RECT 57.565 100.525 57.785 100.805 ;
        RECT 57.955 100.355 58.125 101.135 ;
        RECT 57.720 100.185 58.125 100.355 ;
        RECT 58.295 100.345 58.645 100.965 ;
        RECT 57.720 100.095 57.890 100.185 ;
        RECT 58.815 100.175 59.025 100.965 ;
        RECT 56.670 99.925 57.890 100.095 ;
        RECT 58.350 100.015 59.025 100.175 ;
        RECT 56.330 99.585 57.130 99.755 ;
        RECT 56.450 99.035 56.780 99.415 ;
        RECT 56.960 99.295 57.130 99.585 ;
        RECT 57.720 99.545 57.890 99.925 ;
        RECT 58.060 100.005 59.025 100.015 ;
        RECT 59.215 100.835 59.475 101.225 ;
        RECT 59.685 101.125 60.015 101.585 ;
        RECT 60.890 101.195 61.745 101.365 ;
        RECT 61.950 101.195 62.445 101.365 ;
        RECT 62.615 101.225 62.945 101.585 ;
        RECT 59.215 100.145 59.385 100.835 ;
        RECT 59.555 100.485 59.725 100.665 ;
        RECT 59.895 100.655 60.685 100.905 ;
        RECT 60.890 100.485 61.060 101.195 ;
        RECT 61.230 100.685 61.585 100.905 ;
        RECT 59.555 100.315 61.245 100.485 ;
        RECT 58.060 99.715 58.520 100.005 ;
        RECT 59.215 99.975 60.715 100.145 ;
        RECT 59.215 99.835 59.385 99.975 ;
        RECT 58.825 99.665 59.385 99.835 ;
        RECT 57.300 99.035 57.550 99.495 ;
        RECT 57.720 99.205 58.590 99.545 ;
        RECT 58.825 99.205 58.995 99.665 ;
        RECT 59.830 99.635 60.905 99.805 ;
        RECT 59.165 99.035 59.535 99.495 ;
        RECT 59.830 99.295 60.000 99.635 ;
        RECT 60.170 99.035 60.500 99.465 ;
        RECT 60.735 99.295 60.905 99.635 ;
        RECT 61.075 99.535 61.245 100.315 ;
        RECT 61.415 100.095 61.585 100.685 ;
        RECT 61.755 100.285 62.105 100.905 ;
        RECT 61.415 99.705 61.880 100.095 ;
        RECT 62.275 99.835 62.445 101.195 ;
        RECT 62.615 100.005 63.075 101.055 ;
        RECT 62.050 99.665 62.445 99.835 ;
        RECT 62.050 99.535 62.220 99.665 ;
        RECT 61.075 99.205 61.755 99.535 ;
        RECT 61.970 99.205 62.220 99.535 ;
        RECT 62.390 99.035 62.640 99.495 ;
        RECT 62.810 99.220 63.135 100.005 ;
        RECT 63.305 99.205 63.475 101.325 ;
        RECT 63.645 101.205 63.975 101.585 ;
        RECT 64.145 101.035 64.400 101.325 ;
        RECT 63.650 100.865 64.400 101.035 ;
        RECT 63.650 99.875 63.880 100.865 ;
        RECT 64.575 100.860 64.865 101.585 ;
        RECT 65.960 101.040 71.305 101.585 ;
        RECT 64.050 100.045 64.400 100.695 ;
        RECT 63.650 99.705 64.400 99.875 ;
        RECT 63.645 99.035 63.975 99.535 ;
        RECT 64.145 99.205 64.400 99.705 ;
        RECT 64.575 99.035 64.865 100.200 ;
        RECT 67.550 99.470 67.900 100.720 ;
        RECT 69.380 100.210 69.720 101.040 ;
        RECT 71.480 100.875 71.735 101.405 ;
        RECT 71.905 101.125 72.210 101.585 ;
        RECT 72.455 101.205 73.525 101.375 ;
        RECT 71.480 100.225 71.690 100.875 ;
        RECT 72.455 100.850 72.775 101.205 ;
        RECT 72.450 100.675 72.775 100.850 ;
        RECT 71.860 100.375 72.775 100.675 ;
        RECT 72.945 100.635 73.185 101.035 ;
        RECT 73.355 100.975 73.525 101.205 ;
        RECT 73.695 101.145 73.885 101.585 ;
        RECT 74.055 101.135 75.005 101.415 ;
        RECT 75.225 101.225 75.575 101.395 ;
        RECT 73.355 100.805 73.885 100.975 ;
        RECT 71.860 100.345 72.600 100.375 ;
        RECT 65.960 99.035 71.305 99.470 ;
        RECT 71.480 99.345 71.735 100.225 ;
        RECT 71.905 99.035 72.210 100.175 ;
        RECT 72.430 99.755 72.600 100.345 ;
        RECT 72.945 100.265 73.485 100.635 ;
        RECT 73.665 100.525 73.885 100.805 ;
        RECT 74.055 100.355 74.225 101.135 ;
        RECT 73.820 100.185 74.225 100.355 ;
        RECT 74.395 100.345 74.745 100.965 ;
        RECT 73.820 100.095 73.990 100.185 ;
        RECT 74.915 100.175 75.125 100.965 ;
        RECT 72.770 99.925 73.990 100.095 ;
        RECT 74.450 100.015 75.125 100.175 ;
        RECT 72.430 99.585 73.230 99.755 ;
        RECT 72.550 99.035 72.880 99.415 ;
        RECT 73.060 99.295 73.230 99.585 ;
        RECT 73.820 99.545 73.990 99.925 ;
        RECT 74.160 100.005 75.125 100.015 ;
        RECT 75.315 100.835 75.575 101.225 ;
        RECT 75.785 101.125 76.115 101.585 ;
        RECT 76.990 101.195 77.845 101.365 ;
        RECT 78.050 101.195 78.545 101.365 ;
        RECT 78.715 101.225 79.045 101.585 ;
        RECT 75.315 100.145 75.485 100.835 ;
        RECT 75.655 100.485 75.825 100.665 ;
        RECT 75.995 100.655 76.785 100.905 ;
        RECT 76.990 100.485 77.160 101.195 ;
        RECT 77.330 100.685 77.685 100.905 ;
        RECT 75.655 100.315 77.345 100.485 ;
        RECT 74.160 99.715 74.620 100.005 ;
        RECT 75.315 99.975 76.815 100.145 ;
        RECT 75.315 99.835 75.485 99.975 ;
        RECT 74.925 99.665 75.485 99.835 ;
        RECT 73.400 99.035 73.650 99.495 ;
        RECT 73.820 99.205 74.690 99.545 ;
        RECT 74.925 99.205 75.095 99.665 ;
        RECT 75.930 99.635 77.005 99.805 ;
        RECT 75.265 99.035 75.635 99.495 ;
        RECT 75.930 99.295 76.100 99.635 ;
        RECT 76.270 99.035 76.600 99.465 ;
        RECT 76.835 99.295 77.005 99.635 ;
        RECT 77.175 99.535 77.345 100.315 ;
        RECT 77.515 100.095 77.685 100.685 ;
        RECT 77.855 100.285 78.205 100.905 ;
        RECT 77.515 99.705 77.980 100.095 ;
        RECT 78.375 99.835 78.545 101.195 ;
        RECT 78.715 100.005 79.175 101.055 ;
        RECT 78.150 99.665 78.545 99.835 ;
        RECT 78.150 99.535 78.320 99.665 ;
        RECT 77.175 99.205 77.855 99.535 ;
        RECT 78.070 99.205 78.320 99.535 ;
        RECT 78.490 99.035 78.740 99.495 ;
        RECT 78.910 99.220 79.235 100.005 ;
        RECT 79.405 99.205 79.575 101.325 ;
        RECT 79.745 101.205 80.075 101.585 ;
        RECT 80.245 101.035 80.500 101.325 ;
        RECT 79.750 100.865 80.500 101.035 ;
        RECT 81.140 100.875 81.395 101.405 ;
        RECT 81.565 101.125 81.870 101.585 ;
        RECT 82.115 101.205 83.185 101.375 ;
        RECT 79.750 99.875 79.980 100.865 ;
        RECT 80.150 100.045 80.500 100.695 ;
        RECT 81.140 100.225 81.350 100.875 ;
        RECT 82.115 100.850 82.435 101.205 ;
        RECT 82.110 100.675 82.435 100.850 ;
        RECT 81.520 100.375 82.435 100.675 ;
        RECT 82.605 100.635 82.845 101.035 ;
        RECT 83.015 100.975 83.185 101.205 ;
        RECT 83.355 101.145 83.545 101.585 ;
        RECT 83.715 101.135 84.665 101.415 ;
        RECT 84.885 101.225 85.235 101.395 ;
        RECT 83.015 100.805 83.545 100.975 ;
        RECT 81.520 100.345 82.260 100.375 ;
        RECT 79.750 99.705 80.500 99.875 ;
        RECT 79.745 99.035 80.075 99.535 ;
        RECT 80.245 99.205 80.500 99.705 ;
        RECT 81.140 99.345 81.395 100.225 ;
        RECT 81.565 99.035 81.870 100.175 ;
        RECT 82.090 99.755 82.260 100.345 ;
        RECT 82.605 100.265 83.145 100.635 ;
        RECT 83.325 100.525 83.545 100.805 ;
        RECT 83.715 100.355 83.885 101.135 ;
        RECT 83.480 100.185 83.885 100.355 ;
        RECT 84.055 100.345 84.405 100.965 ;
        RECT 83.480 100.095 83.650 100.185 ;
        RECT 84.575 100.175 84.785 100.965 ;
        RECT 82.430 99.925 83.650 100.095 ;
        RECT 84.110 100.015 84.785 100.175 ;
        RECT 82.090 99.585 82.890 99.755 ;
        RECT 82.210 99.035 82.540 99.415 ;
        RECT 82.720 99.295 82.890 99.585 ;
        RECT 83.480 99.545 83.650 99.925 ;
        RECT 83.820 100.005 84.785 100.015 ;
        RECT 84.975 100.835 85.235 101.225 ;
        RECT 85.445 101.125 85.775 101.585 ;
        RECT 86.650 101.195 87.505 101.365 ;
        RECT 87.710 101.195 88.205 101.365 ;
        RECT 88.375 101.225 88.705 101.585 ;
        RECT 84.975 100.145 85.145 100.835 ;
        RECT 85.315 100.485 85.485 100.665 ;
        RECT 85.655 100.655 86.445 100.905 ;
        RECT 86.650 100.485 86.820 101.195 ;
        RECT 86.990 100.685 87.345 100.905 ;
        RECT 85.315 100.315 87.005 100.485 ;
        RECT 83.820 99.715 84.280 100.005 ;
        RECT 84.975 99.975 86.475 100.145 ;
        RECT 84.975 99.835 85.145 99.975 ;
        RECT 84.585 99.665 85.145 99.835 ;
        RECT 83.060 99.035 83.310 99.495 ;
        RECT 83.480 99.205 84.350 99.545 ;
        RECT 84.585 99.205 84.755 99.665 ;
        RECT 85.590 99.635 86.665 99.805 ;
        RECT 84.925 99.035 85.295 99.495 ;
        RECT 85.590 99.295 85.760 99.635 ;
        RECT 85.930 99.035 86.260 99.465 ;
        RECT 86.495 99.295 86.665 99.635 ;
        RECT 86.835 99.535 87.005 100.315 ;
        RECT 87.175 100.095 87.345 100.685 ;
        RECT 87.515 100.285 87.865 100.905 ;
        RECT 87.175 99.705 87.640 100.095 ;
        RECT 88.035 99.835 88.205 101.195 ;
        RECT 88.375 100.005 88.835 101.055 ;
        RECT 87.810 99.665 88.205 99.835 ;
        RECT 87.810 99.535 87.980 99.665 ;
        RECT 86.835 99.205 87.515 99.535 ;
        RECT 87.730 99.205 87.980 99.535 ;
        RECT 88.150 99.035 88.400 99.495 ;
        RECT 88.570 99.220 88.895 100.005 ;
        RECT 89.065 99.205 89.235 101.325 ;
        RECT 89.405 101.205 89.735 101.585 ;
        RECT 89.905 101.035 90.160 101.325 ;
        RECT 89.410 100.865 90.160 101.035 ;
        RECT 89.410 99.875 89.640 100.865 ;
        RECT 90.335 100.860 90.625 101.585 ;
        RECT 90.795 100.815 94.305 101.585 ;
        RECT 94.480 101.040 99.825 101.585 ;
        RECT 89.810 100.045 90.160 100.695 ;
        RECT 89.410 99.705 90.160 99.875 ;
        RECT 89.405 99.035 89.735 99.535 ;
        RECT 89.905 99.205 90.160 99.705 ;
        RECT 90.335 99.035 90.625 100.200 ;
        RECT 90.795 100.125 92.485 100.645 ;
        RECT 92.655 100.295 94.305 100.815 ;
        RECT 90.795 99.035 94.305 100.125 ;
        RECT 96.070 99.470 96.420 100.720 ;
        RECT 97.900 100.210 98.240 101.040 ;
        RECT 100.000 100.875 100.255 101.405 ;
        RECT 100.425 101.125 100.730 101.585 ;
        RECT 100.975 101.205 102.045 101.375 ;
        RECT 100.000 100.225 100.210 100.875 ;
        RECT 100.975 100.850 101.295 101.205 ;
        RECT 100.970 100.675 101.295 100.850 ;
        RECT 100.380 100.375 101.295 100.675 ;
        RECT 101.465 100.635 101.705 101.035 ;
        RECT 101.875 100.975 102.045 101.205 ;
        RECT 102.215 101.145 102.405 101.585 ;
        RECT 102.575 101.135 103.525 101.415 ;
        RECT 103.745 101.225 104.095 101.395 ;
        RECT 101.875 100.805 102.405 100.975 ;
        RECT 100.380 100.345 101.120 100.375 ;
        RECT 94.480 99.035 99.825 99.470 ;
        RECT 100.000 99.345 100.255 100.225 ;
        RECT 100.425 99.035 100.730 100.175 ;
        RECT 100.950 99.755 101.120 100.345 ;
        RECT 101.465 100.265 102.005 100.635 ;
        RECT 102.185 100.525 102.405 100.805 ;
        RECT 102.575 100.355 102.745 101.135 ;
        RECT 102.340 100.185 102.745 100.355 ;
        RECT 102.915 100.345 103.265 100.965 ;
        RECT 102.340 100.095 102.510 100.185 ;
        RECT 103.435 100.175 103.645 100.965 ;
        RECT 101.290 99.925 102.510 100.095 ;
        RECT 102.970 100.015 103.645 100.175 ;
        RECT 100.950 99.585 101.750 99.755 ;
        RECT 101.070 99.035 101.400 99.415 ;
        RECT 101.580 99.295 101.750 99.585 ;
        RECT 102.340 99.545 102.510 99.925 ;
        RECT 102.680 100.005 103.645 100.015 ;
        RECT 103.835 100.835 104.095 101.225 ;
        RECT 104.305 101.125 104.635 101.585 ;
        RECT 105.510 101.195 106.365 101.365 ;
        RECT 106.570 101.195 107.065 101.365 ;
        RECT 107.235 101.225 107.565 101.585 ;
        RECT 103.835 100.145 104.005 100.835 ;
        RECT 104.175 100.485 104.345 100.665 ;
        RECT 104.515 100.655 105.305 100.905 ;
        RECT 105.510 100.485 105.680 101.195 ;
        RECT 105.850 100.685 106.205 100.905 ;
        RECT 104.175 100.315 105.865 100.485 ;
        RECT 102.680 99.715 103.140 100.005 ;
        RECT 103.835 99.975 105.335 100.145 ;
        RECT 103.835 99.835 104.005 99.975 ;
        RECT 103.445 99.665 104.005 99.835 ;
        RECT 101.920 99.035 102.170 99.495 ;
        RECT 102.340 99.205 103.210 99.545 ;
        RECT 103.445 99.205 103.615 99.665 ;
        RECT 104.450 99.635 105.525 99.805 ;
        RECT 103.785 99.035 104.155 99.495 ;
        RECT 104.450 99.295 104.620 99.635 ;
        RECT 104.790 99.035 105.120 99.465 ;
        RECT 105.355 99.295 105.525 99.635 ;
        RECT 105.695 99.535 105.865 100.315 ;
        RECT 106.035 100.095 106.205 100.685 ;
        RECT 106.375 100.285 106.725 100.905 ;
        RECT 106.035 99.705 106.500 100.095 ;
        RECT 106.895 99.835 107.065 101.195 ;
        RECT 107.235 100.005 107.695 101.055 ;
        RECT 106.670 99.665 107.065 99.835 ;
        RECT 106.670 99.535 106.840 99.665 ;
        RECT 105.695 99.205 106.375 99.535 ;
        RECT 106.590 99.205 106.840 99.535 ;
        RECT 107.010 99.035 107.260 99.495 ;
        RECT 107.430 99.220 107.755 100.005 ;
        RECT 107.925 99.205 108.095 101.325 ;
        RECT 108.265 101.205 108.595 101.585 ;
        RECT 108.765 101.035 109.020 101.325 ;
        RECT 108.270 100.865 109.020 101.035 ;
        RECT 108.270 99.875 108.500 100.865 ;
        RECT 109.195 100.835 110.405 101.585 ;
        RECT 110.580 101.040 115.925 101.585 ;
        RECT 108.670 100.045 109.020 100.695 ;
        RECT 109.195 100.125 109.715 100.665 ;
        RECT 109.885 100.295 110.405 100.835 ;
        RECT 108.270 99.705 109.020 99.875 ;
        RECT 108.265 99.035 108.595 99.535 ;
        RECT 108.765 99.205 109.020 99.705 ;
        RECT 109.195 99.035 110.405 100.125 ;
        RECT 112.170 99.470 112.520 100.720 ;
        RECT 114.000 100.210 114.340 101.040 ;
        RECT 116.095 100.860 116.385 101.585 ;
        RECT 116.560 100.875 116.815 101.405 ;
        RECT 116.985 101.125 117.290 101.585 ;
        RECT 117.535 101.205 118.605 101.375 ;
        RECT 116.560 100.225 116.770 100.875 ;
        RECT 117.535 100.850 117.855 101.205 ;
        RECT 117.530 100.675 117.855 100.850 ;
        RECT 116.940 100.375 117.855 100.675 ;
        RECT 118.025 100.635 118.265 101.035 ;
        RECT 118.435 100.975 118.605 101.205 ;
        RECT 118.775 101.145 118.965 101.585 ;
        RECT 119.135 101.135 120.085 101.415 ;
        RECT 120.305 101.225 120.655 101.395 ;
        RECT 118.435 100.805 118.965 100.975 ;
        RECT 116.940 100.345 117.680 100.375 ;
        RECT 110.580 99.035 115.925 99.470 ;
        RECT 116.095 99.035 116.385 100.200 ;
        RECT 116.560 99.345 116.815 100.225 ;
        RECT 116.985 99.035 117.290 100.175 ;
        RECT 117.510 99.755 117.680 100.345 ;
        RECT 118.025 100.265 118.565 100.635 ;
        RECT 118.745 100.525 118.965 100.805 ;
        RECT 119.135 100.355 119.305 101.135 ;
        RECT 118.900 100.185 119.305 100.355 ;
        RECT 119.475 100.345 119.825 100.965 ;
        RECT 118.900 100.095 119.070 100.185 ;
        RECT 119.995 100.175 120.205 100.965 ;
        RECT 117.850 99.925 119.070 100.095 ;
        RECT 119.530 100.015 120.205 100.175 ;
        RECT 117.510 99.585 118.310 99.755 ;
        RECT 117.630 99.035 117.960 99.415 ;
        RECT 118.140 99.295 118.310 99.585 ;
        RECT 118.900 99.545 119.070 99.925 ;
        RECT 119.240 100.005 120.205 100.015 ;
        RECT 120.395 100.835 120.655 101.225 ;
        RECT 120.865 101.125 121.195 101.585 ;
        RECT 122.070 101.195 122.925 101.365 ;
        RECT 123.130 101.195 123.625 101.365 ;
        RECT 123.795 101.225 124.125 101.585 ;
        RECT 120.395 100.145 120.565 100.835 ;
        RECT 120.735 100.485 120.905 100.665 ;
        RECT 121.075 100.655 121.865 100.905 ;
        RECT 122.070 100.485 122.240 101.195 ;
        RECT 122.410 100.685 122.765 100.905 ;
        RECT 120.735 100.315 122.425 100.485 ;
        RECT 119.240 99.715 119.700 100.005 ;
        RECT 120.395 99.975 121.895 100.145 ;
        RECT 120.395 99.835 120.565 99.975 ;
        RECT 120.005 99.665 120.565 99.835 ;
        RECT 118.480 99.035 118.730 99.495 ;
        RECT 118.900 99.205 119.770 99.545 ;
        RECT 120.005 99.205 120.175 99.665 ;
        RECT 121.010 99.635 122.085 99.805 ;
        RECT 120.345 99.035 120.715 99.495 ;
        RECT 121.010 99.295 121.180 99.635 ;
        RECT 121.350 99.035 121.680 99.465 ;
        RECT 121.915 99.295 122.085 99.635 ;
        RECT 122.255 99.535 122.425 100.315 ;
        RECT 122.595 100.095 122.765 100.685 ;
        RECT 122.935 100.285 123.285 100.905 ;
        RECT 122.595 99.705 123.060 100.095 ;
        RECT 123.455 99.835 123.625 101.195 ;
        RECT 123.795 100.005 124.255 101.055 ;
        RECT 123.230 99.665 123.625 99.835 ;
        RECT 123.230 99.535 123.400 99.665 ;
        RECT 122.255 99.205 122.935 99.535 ;
        RECT 123.150 99.205 123.400 99.535 ;
        RECT 123.570 99.035 123.820 99.495 ;
        RECT 123.990 99.220 124.315 100.005 ;
        RECT 124.485 99.205 124.655 101.325 ;
        RECT 124.825 101.205 125.155 101.585 ;
        RECT 125.325 101.035 125.580 101.325 ;
        RECT 124.830 100.865 125.580 101.035 ;
        RECT 126.675 100.910 126.935 101.415 ;
        RECT 127.115 101.205 127.445 101.585 ;
        RECT 127.625 101.035 127.795 101.415 ;
        RECT 124.830 99.875 125.060 100.865 ;
        RECT 125.230 100.045 125.580 100.695 ;
        RECT 126.675 100.110 126.855 100.910 ;
        RECT 127.130 100.865 127.795 101.035 ;
        RECT 127.130 100.610 127.300 100.865 ;
        RECT 128.055 100.835 129.265 101.585 ;
        RECT 127.025 100.280 127.300 100.610 ;
        RECT 127.525 100.315 127.865 100.685 ;
        RECT 127.130 100.135 127.300 100.280 ;
        RECT 124.830 99.705 125.580 99.875 ;
        RECT 124.825 99.035 125.155 99.535 ;
        RECT 125.325 99.205 125.580 99.705 ;
        RECT 126.675 99.205 126.945 100.110 ;
        RECT 127.130 99.965 127.805 100.135 ;
        RECT 127.115 99.035 127.445 99.795 ;
        RECT 127.625 99.205 127.805 99.965 ;
        RECT 128.055 100.125 128.575 100.665 ;
        RECT 128.745 100.295 129.265 100.835 ;
        RECT 128.055 99.035 129.265 100.125 ;
        RECT 9.290 98.865 129.350 99.035 ;
        RECT 9.375 97.775 10.585 98.865 ;
        RECT 9.375 97.065 9.895 97.605 ;
        RECT 10.065 97.235 10.585 97.775 ;
        RECT 11.215 97.775 12.885 98.865 ;
        RECT 11.215 97.255 11.965 97.775 ;
        RECT 13.055 97.700 13.345 98.865 ;
        RECT 13.515 97.775 14.725 98.865 ;
        RECT 14.900 98.430 20.245 98.865 ;
        RECT 20.420 98.430 25.765 98.865 ;
        RECT 12.135 97.085 12.885 97.605 ;
        RECT 13.515 97.235 14.035 97.775 ;
        RECT 9.375 96.315 10.585 97.065 ;
        RECT 11.215 96.315 12.885 97.085 ;
        RECT 14.205 97.065 14.725 97.605 ;
        RECT 16.490 97.180 16.840 98.430 ;
        RECT 13.055 96.315 13.345 97.040 ;
        RECT 13.515 96.315 14.725 97.065 ;
        RECT 18.320 96.860 18.660 97.690 ;
        RECT 22.010 97.180 22.360 98.430 ;
        RECT 25.935 97.700 26.225 98.865 ;
        RECT 26.395 97.775 27.605 98.865 ;
        RECT 27.780 98.430 33.125 98.865 ;
        RECT 33.300 98.430 38.645 98.865 ;
        RECT 23.840 96.860 24.180 97.690 ;
        RECT 26.395 97.235 26.915 97.775 ;
        RECT 27.085 97.065 27.605 97.605 ;
        RECT 29.370 97.180 29.720 98.430 ;
        RECT 14.900 96.315 20.245 96.860 ;
        RECT 20.420 96.315 25.765 96.860 ;
        RECT 25.935 96.315 26.225 97.040 ;
        RECT 26.395 96.315 27.605 97.065 ;
        RECT 31.200 96.860 31.540 97.690 ;
        RECT 34.890 97.180 35.240 98.430 ;
        RECT 38.815 97.700 39.105 98.865 ;
        RECT 39.275 97.775 40.485 98.865 ;
        RECT 40.660 98.430 46.005 98.865 ;
        RECT 46.180 98.430 51.525 98.865 ;
        RECT 36.720 96.860 37.060 97.690 ;
        RECT 39.275 97.235 39.795 97.775 ;
        RECT 39.965 97.065 40.485 97.605 ;
        RECT 42.250 97.180 42.600 98.430 ;
        RECT 27.780 96.315 33.125 96.860 ;
        RECT 33.300 96.315 38.645 96.860 ;
        RECT 38.815 96.315 39.105 97.040 ;
        RECT 39.275 96.315 40.485 97.065 ;
        RECT 44.080 96.860 44.420 97.690 ;
        RECT 47.770 97.180 48.120 98.430 ;
        RECT 51.695 97.700 51.985 98.865 ;
        RECT 52.155 97.775 53.365 98.865 ;
        RECT 53.540 98.430 58.885 98.865 ;
        RECT 59.060 98.430 64.405 98.865 ;
        RECT 49.600 96.860 49.940 97.690 ;
        RECT 52.155 97.235 52.675 97.775 ;
        RECT 52.845 97.065 53.365 97.605 ;
        RECT 55.130 97.180 55.480 98.430 ;
        RECT 40.660 96.315 46.005 96.860 ;
        RECT 46.180 96.315 51.525 96.860 ;
        RECT 51.695 96.315 51.985 97.040 ;
        RECT 52.155 96.315 53.365 97.065 ;
        RECT 56.960 96.860 57.300 97.690 ;
        RECT 60.650 97.180 61.000 98.430 ;
        RECT 64.575 97.700 64.865 98.865 ;
        RECT 65.035 97.775 66.245 98.865 ;
        RECT 66.420 98.430 71.765 98.865 ;
        RECT 71.940 98.430 77.285 98.865 ;
        RECT 62.480 96.860 62.820 97.690 ;
        RECT 65.035 97.235 65.555 97.775 ;
        RECT 65.725 97.065 66.245 97.605 ;
        RECT 68.010 97.180 68.360 98.430 ;
        RECT 53.540 96.315 58.885 96.860 ;
        RECT 59.060 96.315 64.405 96.860 ;
        RECT 64.575 96.315 64.865 97.040 ;
        RECT 65.035 96.315 66.245 97.065 ;
        RECT 69.840 96.860 70.180 97.690 ;
        RECT 73.530 97.180 73.880 98.430 ;
        RECT 77.455 97.700 77.745 98.865 ;
        RECT 77.915 97.775 79.125 98.865 ;
        RECT 79.300 98.430 84.645 98.865 ;
        RECT 84.820 98.430 90.165 98.865 ;
        RECT 75.360 96.860 75.700 97.690 ;
        RECT 77.915 97.235 78.435 97.775 ;
        RECT 78.605 97.065 79.125 97.605 ;
        RECT 80.890 97.180 81.240 98.430 ;
        RECT 66.420 96.315 71.765 96.860 ;
        RECT 71.940 96.315 77.285 96.860 ;
        RECT 77.455 96.315 77.745 97.040 ;
        RECT 77.915 96.315 79.125 97.065 ;
        RECT 82.720 96.860 83.060 97.690 ;
        RECT 86.410 97.180 86.760 98.430 ;
        RECT 90.335 97.700 90.625 98.865 ;
        RECT 90.795 97.775 92.005 98.865 ;
        RECT 92.180 98.430 97.525 98.865 ;
        RECT 97.700 98.430 103.045 98.865 ;
        RECT 88.240 96.860 88.580 97.690 ;
        RECT 90.795 97.235 91.315 97.775 ;
        RECT 91.485 97.065 92.005 97.605 ;
        RECT 93.770 97.180 94.120 98.430 ;
        RECT 79.300 96.315 84.645 96.860 ;
        RECT 84.820 96.315 90.165 96.860 ;
        RECT 90.335 96.315 90.625 97.040 ;
        RECT 90.795 96.315 92.005 97.065 ;
        RECT 95.600 96.860 95.940 97.690 ;
        RECT 99.290 97.180 99.640 98.430 ;
        RECT 103.215 97.700 103.505 98.865 ;
        RECT 103.675 97.775 104.885 98.865 ;
        RECT 105.060 98.430 110.405 98.865 ;
        RECT 110.580 98.430 115.925 98.865 ;
        RECT 101.120 96.860 101.460 97.690 ;
        RECT 103.675 97.235 104.195 97.775 ;
        RECT 104.365 97.065 104.885 97.605 ;
        RECT 106.650 97.180 107.000 98.430 ;
        RECT 92.180 96.315 97.525 96.860 ;
        RECT 97.700 96.315 103.045 96.860 ;
        RECT 103.215 96.315 103.505 97.040 ;
        RECT 103.675 96.315 104.885 97.065 ;
        RECT 108.480 96.860 108.820 97.690 ;
        RECT 112.170 97.180 112.520 98.430 ;
        RECT 116.095 97.700 116.385 98.865 ;
        RECT 117.020 98.430 122.365 98.865 ;
        RECT 122.540 98.430 127.885 98.865 ;
        RECT 114.000 96.860 114.340 97.690 ;
        RECT 118.610 97.180 118.960 98.430 ;
        RECT 105.060 96.315 110.405 96.860 ;
        RECT 110.580 96.315 115.925 96.860 ;
        RECT 116.095 96.315 116.385 97.040 ;
        RECT 120.440 96.860 120.780 97.690 ;
        RECT 124.130 97.180 124.480 98.430 ;
        RECT 128.055 97.775 129.265 98.865 ;
        RECT 125.960 96.860 126.300 97.690 ;
        RECT 128.055 97.235 128.575 97.775 ;
        RECT 128.745 97.065 129.265 97.605 ;
        RECT 117.020 96.315 122.365 96.860 ;
        RECT 122.540 96.315 127.885 96.860 ;
        RECT 128.055 96.315 129.265 97.065 ;
        RECT 9.290 96.145 129.350 96.315 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 9.290 215.670 129.350 216.150 ;
        RECT 9.290 212.950 129.350 213.430 ;
        RECT 9.290 210.230 129.350 210.710 ;
        RECT 9.290 207.510 129.350 207.990 ;
        RECT 9.290 204.790 129.350 205.270 ;
        RECT 9.290 202.070 129.350 202.550 ;
        RECT 9.290 199.350 129.350 199.830 ;
        RECT 58.575 198.810 59.225 198.855 ;
        RECT 62.175 198.810 62.465 198.855 ;
        RECT 65.495 198.810 65.785 198.855 ;
        RECT 58.575 198.670 65.785 198.810 ;
        RECT 58.575 198.625 59.225 198.670 ;
        RECT 61.875 198.625 62.465 198.670 ;
        RECT 65.495 198.625 65.785 198.670 ;
        RECT 66.030 198.670 73.070 198.810 ;
        RECT 55.380 198.470 55.670 198.515 ;
        RECT 57.215 198.470 57.505 198.515 ;
        RECT 60.795 198.470 61.085 198.515 ;
        RECT 55.380 198.330 61.085 198.470 ;
        RECT 55.380 198.285 55.670 198.330 ;
        RECT 57.215 198.285 57.505 198.330 ;
        RECT 60.795 198.285 61.085 198.330 ;
        RECT 61.875 198.310 62.165 198.625 ;
        RECT 62.720 198.470 63.040 198.530 ;
        RECT 66.030 198.515 66.170 198.670 ;
        RECT 65.955 198.470 66.245 198.515 ;
        RECT 62.720 198.330 66.245 198.470 ;
        RECT 62.720 198.270 63.040 198.330 ;
        RECT 65.955 198.285 66.245 198.330 ;
        RECT 66.400 198.470 66.720 198.530 ;
        RECT 68.715 198.470 69.005 198.515 ;
        RECT 66.400 198.330 69.005 198.470 ;
        RECT 66.400 198.270 66.720 198.330 ;
        RECT 68.715 198.285 69.005 198.330 ;
        RECT 72.930 198.190 73.070 198.670 ;
        RECT 99.075 198.285 99.365 198.515 ;
        RECT 54.900 197.930 55.220 198.190 ;
        RECT 56.295 198.130 56.585 198.175 ;
        RECT 56.295 197.990 67.090 198.130 ;
        RECT 56.295 197.945 56.585 197.990 ;
        RECT 66.950 197.835 67.090 197.990 ;
        RECT 68.240 197.930 68.560 198.190 ;
        RECT 72.840 198.130 73.160 198.190 ;
        RECT 99.150 198.130 99.290 198.285 ;
        RECT 100.440 198.270 100.760 198.530 ;
        RECT 115.175 198.470 115.465 198.515 ;
        RECT 116.080 198.470 116.400 198.530 ;
        RECT 111.110 198.330 116.400 198.470 ;
        RECT 111.110 198.190 111.250 198.330 ;
        RECT 115.175 198.285 115.465 198.330 ;
        RECT 116.080 198.270 116.400 198.330 ;
        RECT 111.020 198.130 111.340 198.190 ;
        RECT 72.840 197.990 111.340 198.130 ;
        RECT 72.840 197.930 73.160 197.990 ;
        RECT 111.020 197.930 111.340 197.990 ;
        RECT 55.785 197.790 56.075 197.835 ;
        RECT 57.675 197.790 57.965 197.835 ;
        RECT 60.795 197.790 61.085 197.835 ;
        RECT 55.785 197.650 61.085 197.790 ;
        RECT 55.785 197.605 56.075 197.650 ;
        RECT 57.675 197.605 57.965 197.650 ;
        RECT 60.795 197.605 61.085 197.650 ;
        RECT 66.875 197.605 67.165 197.835 ;
        RECT 63.655 197.450 63.945 197.495 ;
        RECT 66.400 197.450 66.720 197.510 ;
        RECT 63.655 197.310 66.720 197.450 ;
        RECT 63.655 197.265 63.945 197.310 ;
        RECT 66.400 197.250 66.720 197.310 ;
        RECT 98.600 197.250 98.920 197.510 ;
        RECT 101.360 197.250 101.680 197.510 ;
        RECT 114.715 197.450 115.005 197.495 ;
        RECT 115.160 197.450 115.480 197.510 ;
        RECT 114.715 197.310 115.480 197.450 ;
        RECT 114.715 197.265 115.005 197.310 ;
        RECT 115.160 197.250 115.480 197.310 ;
        RECT 9.290 196.630 129.350 197.110 ;
        RECT 83.420 196.430 83.740 196.490 ;
        RECT 84.125 196.430 84.415 196.475 ;
        RECT 91.240 196.430 91.560 196.490 ;
        RECT 83.420 196.290 91.560 196.430 ;
        RECT 83.420 196.230 83.740 196.290 ;
        RECT 84.125 196.245 84.415 196.290 ;
        RECT 91.240 196.230 91.560 196.290 ;
        RECT 57.625 196.090 57.915 196.135 ;
        RECT 59.515 196.090 59.805 196.135 ;
        RECT 62.635 196.090 62.925 196.135 ;
        RECT 57.625 195.950 62.925 196.090 ;
        RECT 57.625 195.905 57.915 195.950 ;
        RECT 59.515 195.905 59.805 195.950 ;
        RECT 62.635 195.905 62.925 195.950 ;
        RECT 87.990 196.090 88.280 196.135 ;
        RECT 90.770 196.090 91.060 196.135 ;
        RECT 92.630 196.090 92.920 196.135 ;
        RECT 87.990 195.950 92.920 196.090 ;
        RECT 87.990 195.905 88.280 195.950 ;
        RECT 90.770 195.905 91.060 195.950 ;
        RECT 92.630 195.905 92.920 195.950 ;
        RECT 96.875 196.090 97.165 196.135 ;
        RECT 99.995 196.090 100.285 196.135 ;
        RECT 101.885 196.090 102.175 196.135 ;
        RECT 96.875 195.950 102.175 196.090 ;
        RECT 96.875 195.905 97.165 195.950 ;
        RECT 99.995 195.905 100.285 195.950 ;
        RECT 101.885 195.905 102.175 195.950 ;
        RECT 114.355 196.090 114.645 196.135 ;
        RECT 117.475 196.090 117.765 196.135 ;
        RECT 119.365 196.090 119.655 196.135 ;
        RECT 114.355 195.950 119.655 196.090 ;
        RECT 114.355 195.905 114.645 195.950 ;
        RECT 117.475 195.905 117.765 195.950 ;
        RECT 119.365 195.905 119.655 195.950 ;
        RECT 54.900 195.750 55.220 195.810 ;
        RECT 56.740 195.750 57.060 195.810 ;
        RECT 54.900 195.610 57.060 195.750 ;
        RECT 54.900 195.550 55.220 195.610 ;
        RECT 56.740 195.550 57.060 195.610 ;
        RECT 74.680 195.550 75.000 195.810 ;
        RECT 91.255 195.750 91.545 195.795 ;
        RECT 93.540 195.750 93.860 195.810 ;
        RECT 91.255 195.610 93.860 195.750 ;
        RECT 91.255 195.565 91.545 195.610 ;
        RECT 93.540 195.550 93.860 195.610 ;
        RECT 101.360 195.550 101.680 195.810 ;
        RECT 38.340 195.410 38.660 195.470 ;
        RECT 44.335 195.410 44.625 195.455 ;
        RECT 38.340 195.270 44.625 195.410 ;
        RECT 38.340 195.210 38.660 195.270 ;
        RECT 44.335 195.225 44.625 195.270 ;
        RECT 46.635 195.410 46.925 195.455 ;
        RECT 50.315 195.410 50.605 195.455 ;
        RECT 51.680 195.410 52.000 195.470 ;
        RECT 46.635 195.270 52.000 195.410 ;
        RECT 46.635 195.225 46.925 195.270 ;
        RECT 50.315 195.225 50.605 195.270 ;
        RECT 51.680 195.210 52.000 195.270 ;
        RECT 53.980 195.210 54.300 195.470 ;
        RECT 57.220 195.410 57.510 195.455 ;
        RECT 59.055 195.410 59.345 195.455 ;
        RECT 62.635 195.410 62.925 195.455 ;
        RECT 57.220 195.270 62.925 195.410 ;
        RECT 57.220 195.225 57.510 195.270 ;
        RECT 59.055 195.225 59.345 195.270 ;
        RECT 62.635 195.225 62.925 195.270 ;
        RECT 58.135 194.885 58.425 195.115 ;
        RECT 60.415 195.070 61.065 195.115 ;
        RECT 63.180 195.070 63.500 195.130 ;
        RECT 63.715 195.115 64.005 195.430 ;
        RECT 65.480 195.410 65.800 195.470 ;
        RECT 68.255 195.410 68.545 195.455 ;
        RECT 65.480 195.270 68.545 195.410 ;
        RECT 65.480 195.210 65.800 195.270 ;
        RECT 68.255 195.225 68.545 195.270 ;
        RECT 72.840 195.210 73.160 195.470 ;
        RECT 75.155 195.225 75.445 195.455 ;
        RECT 87.990 195.410 88.280 195.455 ;
        RECT 90.780 195.410 91.100 195.470 ;
        RECT 92.620 195.410 92.940 195.470 ;
        RECT 93.095 195.410 93.385 195.455 ;
        RECT 87.990 195.270 90.525 195.410 ;
        RECT 87.990 195.225 88.280 195.270 ;
        RECT 63.715 195.070 64.305 195.115 ;
        RECT 60.415 194.930 64.305 195.070 ;
        RECT 60.415 194.885 61.065 194.930 ;
        RECT 40.640 194.730 40.960 194.790 ;
        RECT 43.415 194.730 43.705 194.775 ;
        RECT 40.640 194.590 43.705 194.730 ;
        RECT 40.640 194.530 40.960 194.590 ;
        RECT 43.415 194.545 43.705 194.590 ;
        RECT 46.160 194.530 46.480 194.790 ;
        RECT 50.760 194.530 51.080 194.790 ;
        RECT 54.915 194.730 55.205 194.775 ;
        RECT 56.280 194.730 56.600 194.790 ;
        RECT 54.915 194.590 56.600 194.730 ;
        RECT 58.210 194.730 58.350 194.885 ;
        RECT 63.180 194.870 63.500 194.930 ;
        RECT 64.015 194.885 64.305 194.930 ;
        RECT 66.860 194.870 67.180 195.130 ;
        RECT 69.160 195.070 69.480 195.130 ;
        RECT 71.460 195.070 71.780 195.130 ;
        RECT 75.230 195.070 75.370 195.225 ;
        RECT 90.310 195.115 90.525 195.270 ;
        RECT 90.780 195.270 93.385 195.410 ;
        RECT 90.780 195.210 91.100 195.270 ;
        RECT 92.620 195.210 92.940 195.270 ;
        RECT 93.095 195.225 93.385 195.270 ;
        RECT 95.795 195.115 96.085 195.430 ;
        RECT 96.875 195.410 97.165 195.455 ;
        RECT 100.455 195.410 100.745 195.455 ;
        RECT 102.290 195.410 102.580 195.455 ;
        RECT 96.875 195.270 102.580 195.410 ;
        RECT 96.875 195.225 97.165 195.270 ;
        RECT 100.455 195.225 100.745 195.270 ;
        RECT 102.290 195.225 102.580 195.270 ;
        RECT 102.740 195.210 103.060 195.470 ;
        RECT 111.020 195.210 111.340 195.470 ;
        RECT 69.160 194.930 75.370 195.070 ;
        RECT 86.130 195.070 86.420 195.115 ;
        RECT 89.390 195.070 89.680 195.115 ;
        RECT 90.310 195.070 90.600 195.115 ;
        RECT 92.170 195.070 92.460 195.115 ;
        RECT 86.130 194.930 90.090 195.070 ;
        RECT 69.160 194.870 69.480 194.930 ;
        RECT 71.460 194.870 71.780 194.930 ;
        RECT 86.130 194.885 86.420 194.930 ;
        RECT 89.390 194.885 89.680 194.930 ;
        RECT 67.335 194.730 67.625 194.775 ;
        RECT 58.210 194.590 67.625 194.730 ;
        RECT 54.915 194.545 55.205 194.590 ;
        RECT 56.280 194.530 56.600 194.590 ;
        RECT 67.335 194.545 67.625 194.590 ;
        RECT 73.300 194.530 73.620 194.790 ;
        RECT 76.995 194.730 77.285 194.775 ;
        RECT 77.440 194.730 77.760 194.790 ;
        RECT 76.995 194.590 77.760 194.730 ;
        RECT 89.950 194.730 90.090 194.930 ;
        RECT 90.310 194.930 92.460 195.070 ;
        RECT 90.310 194.885 90.600 194.930 ;
        RECT 92.170 194.885 92.460 194.930 ;
        RECT 95.495 195.070 96.085 195.115 ;
        RECT 98.600 195.115 98.920 195.130 ;
        RECT 113.275 195.115 113.565 195.430 ;
        RECT 114.355 195.410 114.645 195.455 ;
        RECT 117.935 195.410 118.225 195.455 ;
        RECT 119.770 195.410 120.060 195.455 ;
        RECT 114.355 195.270 120.060 195.410 ;
        RECT 114.355 195.225 114.645 195.270 ;
        RECT 117.935 195.225 118.225 195.270 ;
        RECT 119.770 195.225 120.060 195.270 ;
        RECT 120.220 195.210 120.540 195.470 ;
        RECT 98.600 195.070 99.385 195.115 ;
        RECT 95.495 194.930 99.385 195.070 ;
        RECT 95.495 194.885 95.785 194.930 ;
        RECT 98.600 194.885 99.385 194.930 ;
        RECT 112.975 195.070 113.565 195.115 ;
        RECT 115.160 195.070 115.480 195.130 ;
        RECT 116.215 195.070 116.865 195.115 ;
        RECT 112.975 194.930 116.865 195.070 ;
        RECT 112.975 194.885 113.265 194.930 ;
        RECT 98.600 194.870 98.920 194.885 ;
        RECT 115.160 194.870 115.480 194.930 ;
        RECT 116.215 194.885 116.865 194.930 ;
        RECT 117.460 195.070 117.780 195.130 ;
        RECT 118.855 195.070 119.145 195.115 ;
        RECT 117.460 194.930 119.145 195.070 ;
        RECT 117.460 194.870 117.780 194.930 ;
        RECT 118.855 194.885 119.145 194.930 ;
        RECT 91.700 194.730 92.020 194.790 ;
        RECT 89.950 194.590 92.020 194.730 ;
        RECT 76.995 194.545 77.285 194.590 ;
        RECT 77.440 194.530 77.760 194.590 ;
        RECT 91.700 194.530 92.020 194.590 ;
        RECT 94.015 194.730 94.305 194.775 ;
        RECT 96.760 194.730 97.080 194.790 ;
        RECT 94.015 194.590 97.080 194.730 ;
        RECT 94.015 194.545 94.305 194.590 ;
        RECT 96.760 194.530 97.080 194.590 ;
        RECT 110.560 194.530 110.880 194.790 ;
        RECT 111.480 194.530 111.800 194.790 ;
        RECT 9.290 193.910 129.350 194.390 ;
        RECT 36.055 193.710 36.345 193.755 ;
        RECT 62.735 193.710 63.025 193.755 ;
        RECT 63.180 193.710 63.500 193.770 ;
        RECT 36.055 193.570 48.230 193.710 ;
        RECT 36.055 193.525 36.345 193.570 ;
        RECT 40.640 193.170 40.960 193.430 ;
        RECT 42.935 193.370 43.585 193.415 ;
        RECT 46.535 193.370 46.825 193.415 ;
        RECT 42.935 193.230 46.825 193.370 ;
        RECT 42.935 193.185 43.585 193.230 ;
        RECT 46.235 193.185 46.825 193.230 ;
        RECT 46.235 193.090 46.525 193.185 ;
        RECT 36.040 193.030 36.360 193.090 ;
        RECT 36.515 193.030 36.805 193.075 ;
        RECT 36.040 192.890 36.805 193.030 ;
        RECT 36.040 192.830 36.360 192.890 ;
        RECT 36.515 192.845 36.805 192.890 ;
        RECT 39.740 193.030 40.030 193.075 ;
        RECT 41.575 193.030 41.865 193.075 ;
        RECT 45.155 193.030 45.445 193.075 ;
        RECT 39.740 192.890 45.445 193.030 ;
        RECT 39.740 192.845 40.030 192.890 ;
        RECT 41.575 192.845 41.865 192.890 ;
        RECT 45.155 192.845 45.445 192.890 ;
        RECT 46.160 192.870 46.525 193.090 ;
        RECT 46.160 192.830 46.480 192.870 ;
        RECT 35.580 192.490 35.900 192.750 ;
        RECT 38.800 192.690 39.120 192.750 ;
        RECT 39.275 192.690 39.565 192.735 ;
        RECT 38.800 192.550 39.565 192.690 ;
        RECT 38.800 192.490 39.120 192.550 ;
        RECT 39.275 192.505 39.565 192.550 ;
        RECT 38.340 192.150 38.660 192.410 ;
        RECT 40.145 192.350 40.435 192.395 ;
        RECT 42.035 192.350 42.325 192.395 ;
        RECT 45.155 192.350 45.445 192.395 ;
        RECT 40.145 192.210 45.445 192.350 ;
        RECT 40.145 192.165 40.435 192.210 ;
        RECT 42.035 192.165 42.325 192.210 ;
        RECT 45.155 192.165 45.445 192.210 ;
        RECT 46.620 192.010 46.940 192.070 ;
        RECT 48.090 192.055 48.230 193.570 ;
        RECT 62.735 193.570 63.500 193.710 ;
        RECT 62.735 193.525 63.025 193.570 ;
        RECT 63.180 193.510 63.500 193.570 ;
        RECT 65.480 193.510 65.800 193.770 ;
        RECT 68.240 193.510 68.560 193.770 ;
        RECT 68.715 193.525 69.005 193.755 ;
        RECT 50.415 193.370 50.705 193.415 ;
        RECT 53.655 193.370 54.305 193.415 ;
        RECT 50.415 193.230 54.305 193.370 ;
        RECT 50.415 193.185 51.005 193.230 ;
        RECT 53.655 193.185 54.305 193.230 ;
        RECT 50.715 193.090 51.005 193.185 ;
        RECT 56.280 193.170 56.600 193.430 ;
        RECT 56.740 193.370 57.060 193.430 ;
        RECT 66.255 193.370 66.545 193.415 ;
        RECT 56.740 193.230 57.890 193.370 ;
        RECT 56.740 193.170 57.060 193.230 ;
        RECT 50.715 192.870 51.080 193.090 ;
        RECT 57.750 193.075 57.890 193.230 ;
        RECT 65.570 193.230 66.545 193.370 ;
        RECT 65.570 193.090 65.710 193.230 ;
        RECT 66.255 193.185 66.545 193.230 ;
        RECT 67.320 193.170 67.640 193.430 ;
        RECT 68.790 193.370 68.930 193.525 ;
        RECT 69.160 193.510 69.480 193.770 ;
        RECT 71.015 193.710 71.305 193.755 ;
        RECT 74.680 193.710 75.000 193.770 ;
        RECT 91.255 193.710 91.545 193.755 ;
        RECT 71.015 193.570 75.000 193.710 ;
        RECT 71.015 193.525 71.305 193.570 ;
        RECT 74.680 193.510 75.000 193.570 ;
        RECT 86.730 193.570 91.545 193.710 ;
        RECT 71.920 193.370 72.240 193.430 ;
        RECT 68.790 193.230 72.240 193.370 ;
        RECT 50.760 192.830 51.080 192.870 ;
        RECT 51.795 193.030 52.085 193.075 ;
        RECT 55.375 193.030 55.665 193.075 ;
        RECT 57.210 193.030 57.500 193.075 ;
        RECT 51.795 192.890 57.500 193.030 ;
        RECT 51.795 192.845 52.085 192.890 ;
        RECT 55.375 192.845 55.665 192.890 ;
        RECT 57.210 192.845 57.500 192.890 ;
        RECT 57.675 193.030 57.965 193.075 ;
        RECT 58.120 193.030 58.440 193.090 ;
        RECT 57.675 192.890 58.440 193.030 ;
        RECT 57.675 192.845 57.965 192.890 ;
        RECT 58.120 192.830 58.440 192.890 ;
        RECT 62.720 193.030 63.040 193.090 ;
        RECT 63.195 193.030 63.485 193.075 ;
        RECT 62.720 192.890 63.485 193.030 ;
        RECT 62.720 192.830 63.040 192.890 ;
        RECT 63.195 192.845 63.485 192.890 ;
        RECT 65.480 192.830 65.800 193.090 ;
        RECT 66.860 193.030 67.180 193.090 ;
        RECT 69.620 193.030 69.940 193.090 ;
        RECT 70.170 193.075 70.310 193.230 ;
        RECT 71.920 193.170 72.240 193.230 ;
        RECT 72.955 193.370 73.245 193.415 ;
        RECT 76.195 193.370 76.845 193.415 ;
        RECT 72.955 193.230 76.845 193.370 ;
        RECT 72.955 193.185 73.545 193.230 ;
        RECT 76.195 193.185 76.845 193.230 ;
        RECT 77.440 193.370 77.760 193.430 ;
        RECT 78.835 193.370 79.125 193.415 ;
        RECT 77.440 193.230 79.125 193.370 ;
        RECT 73.255 193.090 73.545 193.185 ;
        RECT 77.440 193.170 77.760 193.230 ;
        RECT 78.835 193.185 79.125 193.230 ;
        RECT 82.910 193.370 83.200 193.415 ;
        RECT 86.170 193.370 86.460 193.415 ;
        RECT 86.730 193.370 86.870 193.570 ;
        RECT 91.255 193.525 91.545 193.570 ;
        RECT 91.700 193.710 92.020 193.770 ;
        RECT 92.635 193.710 92.925 193.755 ;
        RECT 91.700 193.570 92.925 193.710 ;
        RECT 91.700 193.510 92.020 193.570 ;
        RECT 92.635 193.525 92.925 193.570 ;
        RECT 93.540 193.510 93.860 193.770 ;
        RECT 99.075 193.710 99.365 193.755 ;
        RECT 100.440 193.710 100.760 193.770 ;
        RECT 99.075 193.570 100.760 193.710 ;
        RECT 99.075 193.525 99.365 193.570 ;
        RECT 100.440 193.510 100.760 193.570 ;
        RECT 117.460 193.510 117.780 193.770 ;
        RECT 82.910 193.230 86.870 193.370 ;
        RECT 87.090 193.370 87.380 193.415 ;
        RECT 88.950 193.370 89.240 193.415 ;
        RECT 90.320 193.370 90.640 193.430 ;
        RECT 95.840 193.370 96.160 193.430 ;
        RECT 108.375 193.370 108.665 193.415 ;
        RECT 110.560 193.370 110.880 193.430 ;
        RECT 111.615 193.370 112.265 193.415 ;
        RECT 87.090 193.230 89.240 193.370 ;
        RECT 82.910 193.185 83.200 193.230 ;
        RECT 86.170 193.185 86.460 193.230 ;
        RECT 87.090 193.185 87.380 193.230 ;
        RECT 88.950 193.185 89.240 193.230 ;
        RECT 89.490 193.230 90.640 193.370 ;
        RECT 66.860 192.890 69.940 193.030 ;
        RECT 66.860 192.830 67.180 192.890 ;
        RECT 69.620 192.830 69.940 192.890 ;
        RECT 70.095 192.845 70.385 193.075 ;
        RECT 71.015 192.845 71.305 193.075 ;
        RECT 73.255 192.870 73.620 193.090 ;
        RECT 67.780 192.690 68.100 192.750 ;
        RECT 71.090 192.690 71.230 192.845 ;
        RECT 73.300 192.830 73.620 192.870 ;
        RECT 74.335 193.030 74.625 193.075 ;
        RECT 77.915 193.030 78.205 193.075 ;
        RECT 79.750 193.030 80.040 193.075 ;
        RECT 74.335 192.890 80.040 193.030 ;
        RECT 74.335 192.845 74.625 192.890 ;
        RECT 77.915 192.845 78.205 192.890 ;
        RECT 79.750 192.845 80.040 192.890 ;
        RECT 84.770 193.030 85.060 193.075 ;
        RECT 87.090 193.030 87.305 193.185 ;
        RECT 84.770 192.890 87.305 193.030 ;
        RECT 88.035 193.030 88.325 193.075 ;
        RECT 89.490 193.030 89.630 193.230 ;
        RECT 90.320 193.170 90.640 193.230 ;
        RECT 93.170 193.230 100.440 193.370 ;
        RECT 88.035 192.890 89.630 193.030 ;
        RECT 89.875 193.030 90.165 193.075 ;
        RECT 90.780 193.030 91.100 193.090 ;
        RECT 93.170 193.075 93.310 193.230 ;
        RECT 95.840 193.170 96.160 193.230 ;
        RECT 89.875 192.890 91.100 193.030 ;
        RECT 84.770 192.845 85.060 192.890 ;
        RECT 88.035 192.845 88.325 192.890 ;
        RECT 89.875 192.845 90.165 192.890 ;
        RECT 67.780 192.550 71.230 192.690 ;
        RECT 80.215 192.690 80.505 192.735 ;
        RECT 80.660 192.690 80.980 192.750 ;
        RECT 86.640 192.690 86.960 192.750 ;
        RECT 89.950 192.690 90.090 192.845 ;
        RECT 90.780 192.830 91.100 192.890 ;
        RECT 91.715 193.030 92.005 193.075 ;
        RECT 93.095 193.030 93.385 193.075 ;
        RECT 91.715 192.890 93.385 193.030 ;
        RECT 91.715 192.845 92.005 192.890 ;
        RECT 93.095 192.845 93.385 192.890 ;
        RECT 94.475 192.845 94.765 193.075 ;
        RECT 97.235 193.030 97.525 193.075 ;
        RECT 95.010 192.890 97.525 193.030 ;
        RECT 100.300 193.030 100.440 193.230 ;
        RECT 108.375 193.230 112.265 193.370 ;
        RECT 108.375 193.185 108.965 193.230 ;
        RECT 101.835 193.030 102.125 193.075 ;
        RECT 107.800 193.030 108.120 193.090 ;
        RECT 100.300 192.890 102.125 193.030 ;
        RECT 80.215 192.550 90.090 192.690 ;
        RECT 92.160 192.690 92.480 192.750 ;
        RECT 94.550 192.690 94.690 192.845 ;
        RECT 92.160 192.550 94.690 192.690 ;
        RECT 67.780 192.490 68.100 192.550 ;
        RECT 80.215 192.505 80.505 192.550 ;
        RECT 80.660 192.490 80.980 192.550 ;
        RECT 86.640 192.490 86.960 192.550 ;
        RECT 92.160 192.490 92.480 192.550 ;
        RECT 51.795 192.350 52.085 192.395 ;
        RECT 54.915 192.350 55.205 192.395 ;
        RECT 56.805 192.350 57.095 192.395 ;
        RECT 51.795 192.210 57.095 192.350 ;
        RECT 51.795 192.165 52.085 192.210 ;
        RECT 54.915 192.165 55.205 192.210 ;
        RECT 56.805 192.165 57.095 192.210 ;
        RECT 74.335 192.350 74.625 192.395 ;
        RECT 77.455 192.350 77.745 192.395 ;
        RECT 79.345 192.350 79.635 192.395 ;
        RECT 74.335 192.210 79.635 192.350 ;
        RECT 74.335 192.165 74.625 192.210 ;
        RECT 77.455 192.165 77.745 192.210 ;
        RECT 79.345 192.165 79.635 192.210 ;
        RECT 84.770 192.350 85.060 192.395 ;
        RECT 87.550 192.350 87.840 192.395 ;
        RECT 89.410 192.350 89.700 192.395 ;
        RECT 84.770 192.210 89.700 192.350 ;
        RECT 84.770 192.165 85.060 192.210 ;
        RECT 87.550 192.165 87.840 192.210 ;
        RECT 89.410 192.165 89.700 192.210 ;
        RECT 91.240 192.350 91.560 192.410 ;
        RECT 95.010 192.350 95.150 192.890 ;
        RECT 97.235 192.845 97.525 192.890 ;
        RECT 101.835 192.845 102.125 192.890 ;
        RECT 102.370 192.890 108.120 193.030 ;
        RECT 96.300 192.490 96.620 192.750 ;
        RECT 96.760 192.690 97.080 192.750 ;
        RECT 100.900 192.690 101.220 192.750 ;
        RECT 101.375 192.690 101.665 192.735 ;
        RECT 102.370 192.690 102.510 192.890 ;
        RECT 107.800 192.830 108.120 192.890 ;
        RECT 108.675 192.870 108.965 193.185 ;
        RECT 110.560 193.170 110.880 193.230 ;
        RECT 111.615 193.185 112.265 193.230 ;
        RECT 109.755 193.030 110.045 193.075 ;
        RECT 113.335 193.030 113.625 193.075 ;
        RECT 115.170 193.030 115.460 193.075 ;
        RECT 109.755 192.890 115.460 193.030 ;
        RECT 109.755 192.845 110.045 192.890 ;
        RECT 113.335 192.845 113.625 192.890 ;
        RECT 115.170 192.845 115.460 192.890 ;
        RECT 116.540 192.830 116.860 193.090 ;
        RECT 96.760 192.550 100.670 192.690 ;
        RECT 96.760 192.490 97.080 192.550 ;
        RECT 91.240 192.210 95.150 192.350 ;
        RECT 100.530 192.350 100.670 192.550 ;
        RECT 100.900 192.550 101.665 192.690 ;
        RECT 100.900 192.490 101.220 192.550 ;
        RECT 101.375 192.505 101.665 192.550 ;
        RECT 101.910 192.550 102.510 192.690 ;
        RECT 102.740 192.690 103.060 192.750 ;
        RECT 115.635 192.690 115.925 192.735 ;
        RECT 120.220 192.690 120.540 192.750 ;
        RECT 102.740 192.550 120.540 192.690 ;
        RECT 101.910 192.350 102.050 192.550 ;
        RECT 102.740 192.490 103.060 192.550 ;
        RECT 115.635 192.505 115.925 192.550 ;
        RECT 120.220 192.490 120.540 192.550 ;
        RECT 100.530 192.210 102.050 192.350 ;
        RECT 109.755 192.350 110.045 192.395 ;
        RECT 112.875 192.350 113.165 192.395 ;
        RECT 114.765 192.350 115.055 192.395 ;
        RECT 109.755 192.210 115.055 192.350 ;
        RECT 91.240 192.150 91.560 192.210 ;
        RECT 109.755 192.165 110.045 192.210 ;
        RECT 112.875 192.165 113.165 192.210 ;
        RECT 114.765 192.165 115.055 192.210 ;
        RECT 48.015 192.010 48.305 192.055 ;
        RECT 46.620 191.870 48.305 192.010 ;
        RECT 46.620 191.810 46.940 191.870 ;
        RECT 48.015 191.825 48.305 191.870 ;
        RECT 48.935 192.010 49.225 192.055 ;
        RECT 50.760 192.010 51.080 192.070 ;
        RECT 48.935 191.870 51.080 192.010 ;
        RECT 48.935 191.825 49.225 191.870 ;
        RECT 50.760 191.810 51.080 191.870 ;
        RECT 66.415 192.010 66.705 192.055 ;
        RECT 68.240 192.010 68.560 192.070 ;
        RECT 66.415 191.870 68.560 192.010 ;
        RECT 66.415 191.825 66.705 191.870 ;
        RECT 68.240 191.810 68.560 191.870 ;
        RECT 70.080 192.010 70.400 192.070 ;
        RECT 71.475 192.010 71.765 192.055 ;
        RECT 70.080 191.870 71.765 192.010 ;
        RECT 70.080 191.810 70.400 191.870 ;
        RECT 71.475 191.825 71.765 191.870 ;
        RECT 80.905 192.010 81.195 192.055 ;
        RECT 84.340 192.010 84.660 192.070 ;
        RECT 80.905 191.870 84.660 192.010 ;
        RECT 80.905 191.825 81.195 191.870 ;
        RECT 84.340 191.810 84.660 191.870 ;
        RECT 106.880 191.810 107.200 192.070 ;
        RECT 114.350 192.010 114.640 192.055 ;
        RECT 115.160 192.010 115.480 192.070 ;
        RECT 114.350 191.870 115.480 192.010 ;
        RECT 114.350 191.825 114.640 191.870 ;
        RECT 115.160 191.810 115.480 191.870 ;
        RECT 9.290 191.190 129.350 191.670 ;
        RECT 52.615 190.990 52.905 191.035 ;
        RECT 44.410 190.850 52.905 190.990 ;
        RECT 35.090 190.650 35.380 190.695 ;
        RECT 37.870 190.650 38.160 190.695 ;
        RECT 39.730 190.650 40.020 190.695 ;
        RECT 35.090 190.510 40.020 190.650 ;
        RECT 35.090 190.465 35.380 190.510 ;
        RECT 37.870 190.465 38.160 190.510 ;
        RECT 39.730 190.465 40.020 190.510 ;
        RECT 31.440 190.310 31.760 190.370 ;
        RECT 38.800 190.310 39.120 190.370 ;
        RECT 40.195 190.310 40.485 190.355 ;
        RECT 31.440 190.170 40.485 190.310 ;
        RECT 31.440 190.110 31.760 190.170 ;
        RECT 38.800 190.110 39.120 190.170 ;
        RECT 40.195 190.125 40.485 190.170 ;
        RECT 22.700 189.970 23.020 190.030 ;
        RECT 29.615 189.970 29.905 190.015 ;
        RECT 22.700 189.830 29.905 189.970 ;
        RECT 22.700 189.770 23.020 189.830 ;
        RECT 29.615 189.785 29.905 189.830 ;
        RECT 35.090 189.970 35.380 190.015 ;
        RECT 38.355 189.970 38.645 190.015 ;
        RECT 35.090 189.830 37.625 189.970 ;
        RECT 35.090 189.785 35.380 189.830 ;
        RECT 37.410 189.675 37.625 189.830 ;
        RECT 38.355 189.830 40.870 189.970 ;
        RECT 38.355 189.785 38.645 189.830 ;
        RECT 30.075 189.630 30.365 189.675 ;
        RECT 33.230 189.630 33.520 189.675 ;
        RECT 36.490 189.630 36.780 189.675 ;
        RECT 30.075 189.490 36.780 189.630 ;
        RECT 30.075 189.445 30.365 189.490 ;
        RECT 33.230 189.445 33.520 189.490 ;
        RECT 36.490 189.445 36.780 189.490 ;
        RECT 37.410 189.630 37.700 189.675 ;
        RECT 39.270 189.630 39.560 189.675 ;
        RECT 37.410 189.490 39.560 189.630 ;
        RECT 37.410 189.445 37.700 189.490 ;
        RECT 39.270 189.445 39.560 189.490 ;
        RECT 31.225 189.290 31.515 189.335 ;
        RECT 36.040 189.290 36.360 189.350 ;
        RECT 40.730 189.335 40.870 189.830 ;
        RECT 41.560 189.770 41.880 190.030 ;
        RECT 44.410 189.990 44.550 190.850 ;
        RECT 52.615 190.805 52.905 190.850 ;
        RECT 64.575 190.990 64.865 191.035 ;
        RECT 65.480 190.990 65.800 191.050 ;
        RECT 64.575 190.850 65.800 190.990 ;
        RECT 64.575 190.805 64.865 190.850 ;
        RECT 65.480 190.790 65.800 190.850 ;
        RECT 66.860 190.790 67.180 191.050 ;
        RECT 70.555 190.990 70.845 191.035 ;
        RECT 71.460 190.990 71.780 191.050 ;
        RECT 67.410 190.850 71.780 190.990 ;
        RECT 45.355 190.650 45.645 190.695 ;
        RECT 48.475 190.650 48.765 190.695 ;
        RECT 50.365 190.650 50.655 190.695 ;
        RECT 67.410 190.650 67.550 190.850 ;
        RECT 70.555 190.805 70.845 190.850 ;
        RECT 71.460 190.790 71.780 190.850 ;
        RECT 73.315 190.990 73.605 191.035 ;
        RECT 74.695 190.990 74.985 191.035 ;
        RECT 73.315 190.850 74.985 190.990 ;
        RECT 73.315 190.805 73.605 190.850 ;
        RECT 74.695 190.805 74.985 190.850 ;
        RECT 90.320 190.790 90.640 191.050 ;
        RECT 114.715 190.990 115.005 191.035 ;
        RECT 115.160 190.990 115.480 191.050 ;
        RECT 114.715 190.850 115.480 190.990 ;
        RECT 114.715 190.805 115.005 190.850 ;
        RECT 115.160 190.790 115.480 190.850 ;
        RECT 45.355 190.510 50.655 190.650 ;
        RECT 45.355 190.465 45.645 190.510 ;
        RECT 48.475 190.465 48.765 190.510 ;
        RECT 50.365 190.465 50.655 190.510 ;
        RECT 66.030 190.510 67.550 190.650 ;
        RECT 67.795 190.650 68.085 190.695 ;
        RECT 89.875 190.650 90.165 190.695 ;
        RECT 92.160 190.650 92.480 190.710 ;
        RECT 67.795 190.510 69.850 190.650 ;
        RECT 62.735 190.310 63.025 190.355 ;
        RECT 61.890 190.170 63.025 190.310 ;
        RECT 44.275 189.675 44.565 189.990 ;
        RECT 45.355 189.970 45.645 190.015 ;
        RECT 48.935 189.970 49.225 190.015 ;
        RECT 50.770 189.970 51.060 190.015 ;
        RECT 45.355 189.830 51.060 189.970 ;
        RECT 45.355 189.785 45.645 189.830 ;
        RECT 48.935 189.785 49.225 189.830 ;
        RECT 50.770 189.785 51.060 189.830 ;
        RECT 51.220 189.770 51.540 190.030 ;
        RECT 51.680 189.970 52.000 190.030 ;
        RECT 53.075 189.970 53.365 190.015 ;
        RECT 53.520 189.970 53.840 190.030 ;
        RECT 51.680 189.830 53.840 189.970 ;
        RECT 51.680 189.770 52.000 189.830 ;
        RECT 53.075 189.785 53.365 189.830 ;
        RECT 53.520 189.770 53.840 189.830 ;
        RECT 43.975 189.630 44.565 189.675 ;
        RECT 47.215 189.630 47.865 189.675 ;
        RECT 49.855 189.630 50.145 189.675 ;
        RECT 43.975 189.490 47.865 189.630 ;
        RECT 43.975 189.445 44.265 189.490 ;
        RECT 47.215 189.445 47.865 189.490 ;
        RECT 48.090 189.490 50.145 189.630 ;
        RECT 48.090 189.350 48.230 189.490 ;
        RECT 49.855 189.445 50.145 189.490 ;
        RECT 31.225 189.150 36.360 189.290 ;
        RECT 31.225 189.105 31.515 189.150 ;
        RECT 36.040 189.090 36.360 189.150 ;
        RECT 40.655 189.105 40.945 189.335 ;
        RECT 41.100 189.290 41.420 189.350 ;
        RECT 42.495 189.290 42.785 189.335 ;
        RECT 41.100 189.150 42.785 189.290 ;
        RECT 41.100 189.090 41.420 189.150 ;
        RECT 42.495 189.105 42.785 189.150 ;
        RECT 48.000 189.090 48.320 189.350 ;
        RECT 61.890 189.290 62.030 190.170 ;
        RECT 62.735 190.125 63.025 190.170 ;
        RECT 63.655 190.310 63.945 190.355 ;
        RECT 66.030 190.310 66.170 190.510 ;
        RECT 67.795 190.465 68.085 190.510 ;
        RECT 63.655 190.170 66.170 190.310 ;
        RECT 66.400 190.310 66.720 190.370 ;
        RECT 68.240 190.310 68.560 190.370 ;
        RECT 69.710 190.355 69.850 190.510 ;
        RECT 89.875 190.510 92.480 190.650 ;
        RECT 89.875 190.465 90.165 190.510 ;
        RECT 92.160 190.450 92.480 190.510 ;
        RECT 94.885 190.650 95.175 190.695 ;
        RECT 96.775 190.650 97.065 190.695 ;
        RECT 99.895 190.650 100.185 190.695 ;
        RECT 94.885 190.510 100.185 190.650 ;
        RECT 94.885 190.465 95.175 190.510 ;
        RECT 96.775 190.465 97.065 190.510 ;
        RECT 99.895 190.465 100.185 190.510 ;
        RECT 114.255 190.650 114.545 190.695 ;
        RECT 116.540 190.650 116.860 190.710 ;
        RECT 114.255 190.510 116.860 190.650 ;
        RECT 114.255 190.465 114.545 190.510 ;
        RECT 116.540 190.450 116.860 190.510 ;
        RECT 66.400 190.170 68.560 190.310 ;
        RECT 63.655 190.125 63.945 190.170 ;
        RECT 66.400 190.110 66.720 190.170 ;
        RECT 68.240 190.110 68.560 190.170 ;
        RECT 69.635 190.125 69.925 190.355 ;
        RECT 70.170 190.170 71.690 190.310 ;
        RECT 62.275 189.785 62.565 190.015 ;
        RECT 63.195 189.970 63.485 190.015 ;
        RECT 65.035 189.970 65.325 190.015 ;
        RECT 65.940 189.970 66.260 190.030 ;
        RECT 70.170 189.970 70.310 190.170 ;
        RECT 63.195 189.830 70.310 189.970 ;
        RECT 63.195 189.785 63.485 189.830 ;
        RECT 65.035 189.785 65.325 189.830 ;
        RECT 62.350 189.630 62.490 189.785 ;
        RECT 65.940 189.770 66.260 189.830 ;
        RECT 71.000 189.770 71.320 190.030 ;
        RECT 71.550 190.015 71.690 190.170 ;
        RECT 87.100 190.110 87.420 190.370 ;
        RECT 87.575 190.310 87.865 190.355 ;
        RECT 90.780 190.310 91.100 190.370 ;
        RECT 87.575 190.170 91.100 190.310 ;
        RECT 87.575 190.125 87.865 190.170 ;
        RECT 90.780 190.110 91.100 190.170 ;
        RECT 92.620 190.310 92.940 190.370 ;
        RECT 94.015 190.310 94.305 190.355 ;
        RECT 92.620 190.170 94.305 190.310 ;
        RECT 92.620 190.110 92.940 190.170 ;
        RECT 94.015 190.125 94.305 190.170 ;
        RECT 110.560 190.310 110.880 190.370 ;
        RECT 111.035 190.310 111.325 190.355 ;
        RECT 110.560 190.170 111.325 190.310 ;
        RECT 110.560 190.110 110.880 190.170 ;
        RECT 111.035 190.125 111.325 190.170 ;
        RECT 71.475 189.970 71.765 190.015 ;
        RECT 71.920 189.970 72.240 190.030 ;
        RECT 71.475 189.830 72.240 189.970 ;
        RECT 71.475 189.785 71.765 189.830 ;
        RECT 71.920 189.770 72.240 189.830 ;
        RECT 72.380 189.770 72.700 190.030 ;
        RECT 91.240 189.770 91.560 190.030 ;
        RECT 94.480 189.970 94.770 190.015 ;
        RECT 96.315 189.970 96.605 190.015 ;
        RECT 99.895 189.970 100.185 190.015 ;
        RECT 94.480 189.830 100.185 189.970 ;
        RECT 94.480 189.785 94.770 189.830 ;
        RECT 96.315 189.785 96.605 189.830 ;
        RECT 99.895 189.785 100.185 189.830 ;
        RECT 100.900 189.990 101.220 190.030 ;
        RECT 100.900 189.770 101.265 189.990 ;
        RECT 115.620 189.770 115.940 190.030 ;
        RECT 69.620 189.630 69.940 189.690 ;
        RECT 74.535 189.630 74.825 189.675 ;
        RECT 62.350 189.490 69.940 189.630 ;
        RECT 69.620 189.430 69.940 189.490 ;
        RECT 70.170 189.490 74.825 189.630 ;
        RECT 66.400 189.290 66.720 189.350 ;
        RECT 61.890 189.150 66.720 189.290 ;
        RECT 66.400 189.090 66.720 189.150 ;
        RECT 67.320 189.290 67.640 189.350 ;
        RECT 68.255 189.290 68.545 189.335 ;
        RECT 70.170 189.290 70.310 189.490 ;
        RECT 74.535 189.445 74.825 189.490 ;
        RECT 75.140 189.630 75.460 189.690 ;
        RECT 75.615 189.630 75.905 189.675 ;
        RECT 75.140 189.490 75.905 189.630 ;
        RECT 75.140 189.430 75.460 189.490 ;
        RECT 75.615 189.445 75.905 189.490 ;
        RECT 95.380 189.430 95.700 189.690 ;
        RECT 100.975 189.675 101.265 189.770 ;
        RECT 97.675 189.630 98.325 189.675 ;
        RECT 100.975 189.630 101.565 189.675 ;
        RECT 97.675 189.490 101.565 189.630 ;
        RECT 97.675 189.445 98.325 189.490 ;
        RECT 101.275 189.445 101.565 189.490 ;
        RECT 111.480 189.630 111.800 189.690 ;
        RECT 111.955 189.630 112.245 189.675 ;
        RECT 113.780 189.630 114.100 189.690 ;
        RECT 111.480 189.490 114.100 189.630 ;
        RECT 111.480 189.430 111.800 189.490 ;
        RECT 111.955 189.445 112.245 189.490 ;
        RECT 113.780 189.430 114.100 189.490 ;
        RECT 67.320 189.150 70.310 189.290 ;
        RECT 67.320 189.090 67.640 189.150 ;
        RECT 68.255 189.105 68.545 189.150 ;
        RECT 73.760 189.090 74.080 189.350 ;
        RECT 84.800 189.290 85.120 189.350 ;
        RECT 88.035 189.290 88.325 189.335 ;
        RECT 84.800 189.150 88.325 189.290 ;
        RECT 84.800 189.090 85.120 189.150 ;
        RECT 88.035 189.105 88.325 189.150 ;
        RECT 102.280 189.290 102.600 189.350 ;
        RECT 102.755 189.290 103.045 189.335 ;
        RECT 102.280 189.150 103.045 189.290 ;
        RECT 102.280 189.090 102.600 189.150 ;
        RECT 102.755 189.105 103.045 189.150 ;
        RECT 107.800 189.290 108.120 189.350 ;
        RECT 112.415 189.290 112.705 189.335 ;
        RECT 107.800 189.150 112.705 189.290 ;
        RECT 107.800 189.090 108.120 189.150 ;
        RECT 112.415 189.105 112.705 189.150 ;
        RECT 9.290 188.470 129.350 188.950 ;
        RECT 30.995 188.270 31.285 188.315 ;
        RECT 36.055 188.270 36.345 188.315 ;
        RECT 29.230 188.130 31.285 188.270 ;
        RECT 29.230 187.975 29.370 188.130 ;
        RECT 30.995 188.085 31.285 188.130 ;
        RECT 32.450 188.130 36.345 188.270 ;
        RECT 20.875 187.930 21.165 187.975 ;
        RECT 23.275 187.930 23.565 187.975 ;
        RECT 26.515 187.930 27.165 187.975 ;
        RECT 20.875 187.790 27.165 187.930 ;
        RECT 20.875 187.745 21.165 187.790 ;
        RECT 23.275 187.745 23.865 187.790 ;
        RECT 26.515 187.745 27.165 187.790 ;
        RECT 29.155 187.745 29.445 187.975 ;
        RECT 31.440 187.930 31.760 187.990 ;
        RECT 30.610 187.790 31.760 187.930 ;
        RECT 20.415 187.590 20.705 187.635 ;
        RECT 22.700 187.590 23.020 187.650 ;
        RECT 20.415 187.450 23.020 187.590 ;
        RECT 20.415 187.405 20.705 187.450 ;
        RECT 22.700 187.390 23.020 187.450 ;
        RECT 23.575 187.430 23.865 187.745 ;
        RECT 30.610 187.635 30.750 187.790 ;
        RECT 31.440 187.730 31.760 187.790 ;
        RECT 24.655 187.590 24.945 187.635 ;
        RECT 28.235 187.590 28.525 187.635 ;
        RECT 30.070 187.590 30.360 187.635 ;
        RECT 24.655 187.450 30.360 187.590 ;
        RECT 24.655 187.405 24.945 187.450 ;
        RECT 28.235 187.405 28.525 187.450 ;
        RECT 30.070 187.405 30.360 187.450 ;
        RECT 30.535 187.405 30.825 187.635 ;
        RECT 30.980 187.590 31.300 187.650 ;
        RECT 31.915 187.590 32.205 187.635 ;
        RECT 30.980 187.450 32.205 187.590 ;
        RECT 30.980 187.390 31.300 187.450 ;
        RECT 31.915 187.405 32.205 187.450 ;
        RECT 21.795 187.250 22.085 187.295 ;
        RECT 27.300 187.250 27.620 187.310 ;
        RECT 32.450 187.250 32.590 188.130 ;
        RECT 36.055 188.085 36.345 188.130 ;
        RECT 37.895 188.270 38.185 188.315 ;
        RECT 41.560 188.270 41.880 188.330 ;
        RECT 37.895 188.130 41.880 188.270 ;
        RECT 37.895 188.085 38.185 188.130 ;
        RECT 41.560 188.070 41.880 188.130 ;
        RECT 48.000 188.270 48.320 188.330 ;
        RECT 48.935 188.270 49.225 188.315 ;
        RECT 48.000 188.130 49.225 188.270 ;
        RECT 48.000 188.070 48.320 188.130 ;
        RECT 48.935 188.085 49.225 188.130 ;
        RECT 53.075 188.270 53.365 188.315 ;
        RECT 53.980 188.270 54.300 188.330 ;
        RECT 53.075 188.130 54.300 188.270 ;
        RECT 53.075 188.085 53.365 188.130 ;
        RECT 53.980 188.070 54.300 188.130 ;
        RECT 70.095 188.270 70.385 188.315 ;
        RECT 71.460 188.270 71.780 188.330 ;
        RECT 70.095 188.130 71.780 188.270 ;
        RECT 70.095 188.085 70.385 188.130 ;
        RECT 71.460 188.070 71.780 188.130 ;
        RECT 89.415 188.270 89.705 188.315 ;
        RECT 91.240 188.270 91.560 188.330 ;
        RECT 89.415 188.130 91.560 188.270 ;
        RECT 89.415 188.085 89.705 188.130 ;
        RECT 91.240 188.070 91.560 188.130 ;
        RECT 95.380 188.270 95.700 188.330 ;
        RECT 101.375 188.270 101.665 188.315 ;
        RECT 95.380 188.130 101.665 188.270 ;
        RECT 95.380 188.070 95.700 188.130 ;
        RECT 101.375 188.085 101.665 188.130 ;
        RECT 102.280 188.070 102.600 188.330 ;
        RECT 111.020 188.270 111.340 188.330 ;
        RECT 111.495 188.270 111.785 188.315 ;
        RECT 111.020 188.130 111.785 188.270 ;
        RECT 111.020 188.070 111.340 188.130 ;
        RECT 111.495 188.085 111.785 188.130 ;
        RECT 113.335 188.270 113.625 188.315 ;
        RECT 115.620 188.270 115.940 188.330 ;
        RECT 113.335 188.130 115.940 188.270 ;
        RECT 113.335 188.085 113.625 188.130 ;
        RECT 115.620 188.070 115.940 188.130 ;
        RECT 46.620 187.930 46.940 187.990 ;
        RECT 51.235 187.930 51.525 187.975 ;
        RECT 46.620 187.790 51.525 187.930 ;
        RECT 46.620 187.730 46.940 187.790 ;
        RECT 51.235 187.745 51.525 187.790 ;
        RECT 72.955 187.930 73.245 187.975 ;
        RECT 75.600 187.930 75.920 187.990 ;
        RECT 76.195 187.930 76.845 187.975 ;
        RECT 72.955 187.790 76.845 187.930 ;
        RECT 102.370 187.930 102.510 188.070 ;
        RECT 105.055 187.930 105.345 187.975 ;
        RECT 102.370 187.790 105.345 187.930 ;
        RECT 72.955 187.745 73.545 187.790 ;
        RECT 48.000 187.390 48.320 187.650 ;
        RECT 70.080 187.590 70.400 187.650 ;
        RECT 71.015 187.590 71.305 187.635 ;
        RECT 70.080 187.450 71.305 187.590 ;
        RECT 70.080 187.390 70.400 187.450 ;
        RECT 71.015 187.405 71.305 187.450 ;
        RECT 73.255 187.430 73.545 187.745 ;
        RECT 75.600 187.730 75.920 187.790 ;
        RECT 76.195 187.745 76.845 187.790 ;
        RECT 105.055 187.745 105.345 187.790 ;
        RECT 74.335 187.590 74.625 187.635 ;
        RECT 77.915 187.590 78.205 187.635 ;
        RECT 79.750 187.590 80.040 187.635 ;
        RECT 74.335 187.450 80.040 187.590 ;
        RECT 74.335 187.405 74.625 187.450 ;
        RECT 77.915 187.405 78.205 187.450 ;
        RECT 79.750 187.405 80.040 187.450 ;
        RECT 84.800 187.590 85.120 187.650 ;
        RECT 87.115 187.590 87.405 187.635 ;
        RECT 84.800 187.450 87.405 187.590 ;
        RECT 84.800 187.390 85.120 187.450 ;
        RECT 87.115 187.405 87.405 187.450 ;
        RECT 87.560 187.390 87.880 187.650 ;
        RECT 102.295 187.590 102.585 187.635 ;
        RECT 104.595 187.590 104.885 187.635 ;
        RECT 106.880 187.590 107.200 187.650 ;
        RECT 111.035 187.590 111.325 187.635 ;
        RECT 102.295 187.450 102.970 187.590 ;
        RECT 102.295 187.405 102.585 187.450 ;
        RECT 21.795 187.110 32.590 187.250 ;
        RECT 21.795 187.065 22.085 187.110 ;
        RECT 27.300 187.050 27.620 187.110 ;
        RECT 35.120 187.050 35.440 187.310 ;
        RECT 35.595 187.250 35.885 187.295 ;
        RECT 36.040 187.250 36.360 187.310 ;
        RECT 35.595 187.110 36.360 187.250 ;
        RECT 35.595 187.065 35.885 187.110 ;
        RECT 36.040 187.050 36.360 187.110 ;
        RECT 49.840 187.050 50.160 187.310 ;
        RECT 50.760 187.050 51.080 187.310 ;
        RECT 78.820 187.050 79.140 187.310 ;
        RECT 80.215 187.250 80.505 187.295 ;
        RECT 80.660 187.250 80.980 187.310 ;
        RECT 80.215 187.110 80.980 187.250 ;
        RECT 80.215 187.065 80.505 187.110 ;
        RECT 80.660 187.050 80.980 187.110 ;
        RECT 86.655 187.065 86.945 187.295 ;
        RECT 24.655 186.910 24.945 186.955 ;
        RECT 27.775 186.910 28.065 186.955 ;
        RECT 29.665 186.910 29.955 186.955 ;
        RECT 24.655 186.770 29.955 186.910 ;
        RECT 24.655 186.725 24.945 186.770 ;
        RECT 27.775 186.725 28.065 186.770 ;
        RECT 29.665 186.725 29.955 186.770 ;
        RECT 74.335 186.910 74.625 186.955 ;
        RECT 77.455 186.910 77.745 186.955 ;
        RECT 79.345 186.910 79.635 186.955 ;
        RECT 74.335 186.770 79.635 186.910 ;
        RECT 86.730 186.910 86.870 187.065 ;
        RECT 87.100 186.910 87.420 186.970 ;
        RECT 102.830 186.955 102.970 187.450 ;
        RECT 104.595 187.450 111.325 187.590 ;
        RECT 104.595 187.405 104.885 187.450 ;
        RECT 106.880 187.390 107.200 187.450 ;
        RECT 111.035 187.405 111.325 187.450 ;
        RECT 105.975 187.250 106.265 187.295 ;
        RECT 107.340 187.250 107.660 187.310 ;
        RECT 110.115 187.250 110.405 187.295 ;
        RECT 110.560 187.250 110.880 187.310 ;
        RECT 105.975 187.110 110.880 187.250 ;
        RECT 105.975 187.065 106.265 187.110 ;
        RECT 107.340 187.050 107.660 187.110 ;
        RECT 110.115 187.065 110.405 187.110 ;
        RECT 110.560 187.050 110.880 187.110 ;
        RECT 86.730 186.770 87.420 186.910 ;
        RECT 74.335 186.725 74.625 186.770 ;
        RECT 77.455 186.725 77.745 186.770 ;
        RECT 79.345 186.725 79.635 186.770 ;
        RECT 87.100 186.710 87.420 186.770 ;
        RECT 102.755 186.725 103.045 186.955 ;
        RECT 69.160 186.570 69.480 186.630 ;
        RECT 71.475 186.570 71.765 186.615 ;
        RECT 69.160 186.430 71.765 186.570 ;
        RECT 69.160 186.370 69.480 186.430 ;
        RECT 71.475 186.385 71.765 186.430 ;
        RECT 9.290 185.750 129.350 186.230 ;
        RECT 30.075 185.550 30.365 185.595 ;
        RECT 30.980 185.550 31.300 185.610 ;
        RECT 30.075 185.410 31.300 185.550 ;
        RECT 30.075 185.365 30.365 185.410 ;
        RECT 30.980 185.350 31.300 185.410 ;
        RECT 46.635 185.550 46.925 185.595 ;
        RECT 48.000 185.550 48.320 185.610 ;
        RECT 46.635 185.410 48.320 185.550 ;
        RECT 46.635 185.365 46.925 185.410 ;
        RECT 48.000 185.350 48.320 185.410 ;
        RECT 74.695 185.550 74.985 185.595 ;
        RECT 78.820 185.550 79.140 185.610 ;
        RECT 74.695 185.410 79.140 185.550 ;
        RECT 74.695 185.365 74.985 185.410 ;
        RECT 78.820 185.350 79.140 185.410 ;
        RECT 37.075 185.210 37.365 185.255 ;
        RECT 40.195 185.210 40.485 185.255 ;
        RECT 42.085 185.210 42.375 185.255 ;
        RECT 37.075 185.070 42.375 185.210 ;
        RECT 37.075 185.025 37.365 185.070 ;
        RECT 40.195 185.025 40.485 185.070 ;
        RECT 42.085 185.025 42.375 185.070 ;
        RECT 75.600 185.010 75.920 185.270 ;
        RECT 27.315 184.870 27.605 184.915 ;
        RECT 32.360 184.870 32.680 184.930 ;
        RECT 35.580 184.870 35.900 184.930 ;
        RECT 27.315 184.730 35.900 184.870 ;
        RECT 27.315 184.685 27.605 184.730 ;
        RECT 32.360 184.670 32.680 184.730 ;
        RECT 35.580 184.670 35.900 184.730 ;
        RECT 41.100 184.870 41.420 184.930 ;
        RECT 48.935 184.870 49.225 184.915 ;
        RECT 41.100 184.730 49.225 184.870 ;
        RECT 41.100 184.670 41.420 184.730 ;
        RECT 48.935 184.685 49.225 184.730 ;
        RECT 49.395 184.870 49.685 184.915 ;
        RECT 49.840 184.870 50.160 184.930 ;
        RECT 69.160 184.915 69.480 184.930 ;
        RECT 69.050 184.870 69.480 184.915 ;
        RECT 49.395 184.730 50.160 184.870 ;
        RECT 49.395 184.685 49.685 184.730 ;
        RECT 35.995 184.235 36.285 184.550 ;
        RECT 37.075 184.530 37.365 184.575 ;
        RECT 40.655 184.530 40.945 184.575 ;
        RECT 42.490 184.530 42.780 184.575 ;
        RECT 37.075 184.390 42.780 184.530 ;
        RECT 37.075 184.345 37.365 184.390 ;
        RECT 40.655 184.345 40.945 184.390 ;
        RECT 42.490 184.345 42.780 184.390 ;
        RECT 42.955 184.345 43.245 184.575 ;
        RECT 45.700 184.530 46.020 184.590 ;
        RECT 49.470 184.530 49.610 184.685 ;
        RECT 49.840 184.670 50.160 184.730 ;
        RECT 67.410 184.730 69.480 184.870 ;
        RECT 45.700 184.390 49.610 184.530 ;
        RECT 35.695 184.190 36.285 184.235 ;
        RECT 36.500 184.190 36.820 184.250 ;
        RECT 38.935 184.190 39.585 184.235 ;
        RECT 35.695 184.050 39.585 184.190 ;
        RECT 35.695 184.005 35.985 184.050 ;
        RECT 36.500 183.990 36.820 184.050 ;
        RECT 38.935 184.005 39.585 184.050 ;
        RECT 40.180 184.190 40.500 184.250 ;
        RECT 41.575 184.190 41.865 184.235 ;
        RECT 40.180 184.050 41.865 184.190 ;
        RECT 43.030 184.190 43.170 184.345 ;
        RECT 45.700 184.330 46.020 184.390 ;
        RECT 53.520 184.330 53.840 184.590 ;
        RECT 67.410 184.575 67.550 184.730 ;
        RECT 69.050 184.685 69.480 184.730 ;
        RECT 69.160 184.670 69.480 184.685 ;
        RECT 70.080 184.670 70.400 184.930 ;
        RECT 71.000 184.870 71.320 184.930 ;
        RECT 71.475 184.870 71.765 184.915 ;
        RECT 71.000 184.730 71.765 184.870 ;
        RECT 71.000 184.670 71.320 184.730 ;
        RECT 71.475 184.685 71.765 184.730 ;
        RECT 72.840 184.870 73.160 184.930 ;
        RECT 87.100 184.870 87.420 184.930 ;
        RECT 96.300 184.870 96.620 184.930 ;
        RECT 107.340 184.870 107.660 184.930 ;
        RECT 72.840 184.730 76.290 184.870 ;
        RECT 72.840 184.670 73.160 184.730 ;
        RECT 67.335 184.345 67.625 184.575 ;
        RECT 73.760 184.330 74.080 184.590 ;
        RECT 75.600 184.530 75.920 184.590 ;
        RECT 76.150 184.575 76.290 184.730 ;
        RECT 87.100 184.730 107.660 184.870 ;
        RECT 87.100 184.670 87.420 184.730 ;
        RECT 96.300 184.670 96.620 184.730 ;
        RECT 107.340 184.670 107.660 184.730 ;
        RECT 76.075 184.530 76.365 184.575 ;
        RECT 75.600 184.390 76.365 184.530 ;
        RECT 75.600 184.330 75.920 184.390 ;
        RECT 76.075 184.345 76.365 184.390 ;
        RECT 116.080 184.530 116.400 184.590 ;
        RECT 116.555 184.530 116.845 184.575 ;
        RECT 117.935 184.530 118.225 184.575 ;
        RECT 116.080 184.390 118.225 184.530 ;
        RECT 116.080 184.330 116.400 184.390 ;
        RECT 116.555 184.345 116.845 184.390 ;
        RECT 117.935 184.345 118.225 184.390 ;
        RECT 120.235 184.345 120.525 184.575 ;
        RECT 51.220 184.190 51.540 184.250 ;
        RECT 72.380 184.190 72.700 184.250 ;
        RECT 97.235 184.190 97.525 184.235 ;
        RECT 43.030 184.050 51.540 184.190 ;
        RECT 40.180 183.990 40.500 184.050 ;
        RECT 41.575 184.005 41.865 184.050 ;
        RECT 51.220 183.990 51.540 184.050 ;
        RECT 67.870 184.050 72.700 184.190 ;
        RECT 67.870 183.910 68.010 184.050 ;
        RECT 72.380 183.990 72.700 184.050 ;
        RECT 88.570 184.050 97.525 184.190 ;
        RECT 88.570 183.910 88.710 184.050 ;
        RECT 97.235 184.005 97.525 184.050 ;
        RECT 97.695 184.190 97.985 184.235 ;
        RECT 100.900 184.190 101.220 184.250 ;
        RECT 102.280 184.190 102.600 184.250 ;
        RECT 97.695 184.050 102.600 184.190 ;
        RECT 97.695 184.005 97.985 184.050 ;
        RECT 100.900 183.990 101.220 184.050 ;
        RECT 102.280 183.990 102.600 184.050 ;
        RECT 115.620 184.190 115.940 184.250 ;
        RECT 120.310 184.190 120.450 184.345 ;
        RECT 115.620 184.050 120.450 184.190 ;
        RECT 115.620 183.990 115.940 184.050 ;
        RECT 27.760 183.650 28.080 183.910 ;
        RECT 28.220 183.650 28.540 183.910 ;
        RECT 32.820 183.850 33.140 183.910 ;
        RECT 34.215 183.850 34.505 183.895 ;
        RECT 32.820 183.710 34.505 183.850 ;
        RECT 32.820 183.650 33.140 183.710 ;
        RECT 34.215 183.665 34.505 183.710 ;
        RECT 42.940 183.850 43.260 183.910 ;
        RECT 48.475 183.850 48.765 183.895 ;
        RECT 42.940 183.710 48.765 183.850 ;
        RECT 42.940 183.650 43.260 183.710 ;
        RECT 48.475 183.665 48.765 183.710 ;
        RECT 53.060 183.650 53.380 183.910 ;
        RECT 66.400 183.850 66.720 183.910 ;
        RECT 66.875 183.850 67.165 183.895 ;
        RECT 67.780 183.850 68.100 183.910 ;
        RECT 66.400 183.710 68.100 183.850 ;
        RECT 66.400 183.650 66.720 183.710 ;
        RECT 66.875 183.665 67.165 183.710 ;
        RECT 67.780 183.650 68.100 183.710 ;
        RECT 68.240 183.650 68.560 183.910 ;
        RECT 68.700 183.850 69.020 183.910 ;
        RECT 69.635 183.850 69.925 183.895 ;
        RECT 68.700 183.710 69.925 183.850 ;
        RECT 68.700 183.650 69.020 183.710 ;
        RECT 69.635 183.665 69.925 183.710 ;
        RECT 82.500 183.850 82.820 183.910 ;
        RECT 87.560 183.850 87.880 183.910 ;
        RECT 88.035 183.850 88.325 183.895 ;
        RECT 82.500 183.710 88.325 183.850 ;
        RECT 82.500 183.650 82.820 183.710 ;
        RECT 87.560 183.650 87.880 183.710 ;
        RECT 88.035 183.665 88.325 183.710 ;
        RECT 88.480 183.650 88.800 183.910 ;
        RECT 90.320 183.650 90.640 183.910 ;
        RECT 99.520 183.650 99.840 183.910 ;
        RECT 117.000 183.650 117.320 183.910 ;
        RECT 118.380 183.650 118.700 183.910 ;
        RECT 121.155 183.850 121.445 183.895 ;
        RECT 123.900 183.850 124.220 183.910 ;
        RECT 121.155 183.710 124.220 183.850 ;
        RECT 121.155 183.665 121.445 183.710 ;
        RECT 123.900 183.650 124.220 183.710 ;
        RECT 9.290 183.030 129.350 183.510 ;
        RECT 36.500 182.630 36.820 182.890 ;
        RECT 38.355 182.830 38.645 182.875 ;
        RECT 40.180 182.830 40.500 182.890 ;
        RECT 38.355 182.690 40.500 182.830 ;
        RECT 38.355 182.645 38.645 182.690 ;
        RECT 40.180 182.630 40.500 182.690 ;
        RECT 41.100 182.630 41.420 182.890 ;
        RECT 69.160 182.630 69.480 182.890 ;
        RECT 90.795 182.830 91.085 182.875 ;
        RECT 88.570 182.690 91.085 182.830 ;
        RECT 32.820 182.490 33.140 182.550 ;
        RECT 41.575 182.490 41.865 182.535 ;
        RECT 32.820 182.350 41.865 182.490 ;
        RECT 32.820 182.290 33.140 182.350 ;
        RECT 41.575 182.305 41.865 182.350 ;
        RECT 50.875 182.490 51.165 182.535 ;
        RECT 53.060 182.490 53.380 182.550 ;
        RECT 54.115 182.490 54.765 182.535 ;
        RECT 50.875 182.350 54.765 182.490 ;
        RECT 50.875 182.305 51.465 182.350 ;
        RECT 21.335 181.965 21.625 182.195 ;
        RECT 21.410 181.810 21.550 181.965 ;
        RECT 27.300 181.950 27.620 182.210 ;
        RECT 36.055 181.965 36.345 182.195 ;
        RECT 37.435 182.150 37.725 182.195 ;
        RECT 37.435 182.010 39.490 182.150 ;
        RECT 37.435 181.965 37.725 182.010 ;
        RECT 22.700 181.810 23.020 181.870 ;
        RECT 36.130 181.810 36.270 181.965 ;
        RECT 21.410 181.670 36.270 181.810 ;
        RECT 22.700 181.610 23.020 181.670 ;
        RECT 39.350 181.515 39.490 182.010 ;
        RECT 51.175 181.990 51.465 182.305 ;
        RECT 53.060 182.290 53.380 182.350 ;
        RECT 54.115 182.305 54.765 182.350 ;
        RECT 65.940 182.490 66.260 182.550 ;
        RECT 71.000 182.490 71.320 182.550 ;
        RECT 71.475 182.490 71.765 182.535 ;
        RECT 65.940 182.350 68.930 182.490 ;
        RECT 65.940 182.290 66.260 182.350 ;
        RECT 52.255 182.150 52.545 182.195 ;
        RECT 55.835 182.150 56.125 182.195 ;
        RECT 57.670 182.150 57.960 182.195 ;
        RECT 52.255 182.010 57.960 182.150 ;
        RECT 52.255 181.965 52.545 182.010 ;
        RECT 55.835 181.965 56.125 182.010 ;
        RECT 57.670 181.965 57.960 182.010 ;
        RECT 58.120 181.950 58.440 182.210 ;
        RECT 66.875 181.965 67.165 182.195 ;
        RECT 68.790 182.150 68.930 182.350 ;
        RECT 71.000 182.350 71.765 182.490 ;
        RECT 71.000 182.290 71.320 182.350 ;
        RECT 71.475 182.305 71.765 182.350 ;
        RECT 82.615 182.490 82.905 182.535 ;
        RECT 85.855 182.490 86.505 182.535 ;
        RECT 88.020 182.490 88.340 182.550 ;
        RECT 88.570 182.535 88.710 182.690 ;
        RECT 90.795 182.645 91.085 182.690 ;
        RECT 115.620 182.630 115.940 182.890 ;
        RECT 82.615 182.350 88.340 182.490 ;
        RECT 82.615 182.305 83.205 182.350 ;
        RECT 85.855 182.305 86.505 182.350 ;
        RECT 69.160 182.150 69.480 182.210 ;
        RECT 73.315 182.150 73.605 182.195 ;
        RECT 68.790 182.010 73.605 182.150 ;
        RECT 42.035 181.810 42.325 181.855 ;
        RECT 45.700 181.810 46.020 181.870 ;
        RECT 41.190 181.670 46.020 181.810 ;
        RECT 39.275 181.285 39.565 181.515 ;
        RECT 21.780 180.930 22.100 181.190 ;
        RECT 26.380 180.930 26.700 181.190 ;
        RECT 32.360 181.130 32.680 181.190 ;
        RECT 41.190 181.130 41.330 181.670 ;
        RECT 42.035 181.625 42.325 181.670 ;
        RECT 45.700 181.610 46.020 181.670 ;
        RECT 56.740 181.610 57.060 181.870 ;
        RECT 66.950 181.810 67.090 181.965 ;
        RECT 69.160 181.950 69.480 182.010 ;
        RECT 73.315 181.965 73.605 182.010 ;
        RECT 75.600 181.950 75.920 182.210 ;
        RECT 82.915 181.990 83.205 182.305 ;
        RECT 88.020 182.290 88.340 182.350 ;
        RECT 88.495 182.305 88.785 182.535 ;
        RECT 94.115 182.490 94.405 182.535 ;
        RECT 96.300 182.490 96.620 182.550 ;
        RECT 97.355 182.490 98.005 182.535 ;
        RECT 94.115 182.350 98.005 182.490 ;
        RECT 94.115 182.305 94.705 182.350 ;
        RECT 83.995 182.150 84.285 182.195 ;
        RECT 87.575 182.150 87.865 182.195 ;
        RECT 89.410 182.150 89.700 182.195 ;
        RECT 83.995 182.010 89.700 182.150 ;
        RECT 83.995 181.965 84.285 182.010 ;
        RECT 87.575 181.965 87.865 182.010 ;
        RECT 89.410 181.965 89.700 182.010 ;
        RECT 90.320 182.150 90.640 182.210 ;
        RECT 91.715 182.150 92.005 182.195 ;
        RECT 90.320 182.010 92.005 182.150 ;
        RECT 90.320 181.950 90.640 182.010 ;
        RECT 91.715 181.965 92.005 182.010 ;
        RECT 94.415 181.990 94.705 182.305 ;
        RECT 96.300 182.290 96.620 182.350 ;
        RECT 97.355 182.305 98.005 182.350 ;
        RECT 112.860 182.490 113.180 182.550 ;
        RECT 113.795 182.490 114.085 182.535 ;
        RECT 112.860 182.350 114.085 182.490 ;
        RECT 112.860 182.290 113.180 182.350 ;
        RECT 113.795 182.305 114.085 182.350 ;
        RECT 117.000 182.490 117.320 182.550 ;
        RECT 118.035 182.490 118.325 182.535 ;
        RECT 121.275 182.490 121.925 182.535 ;
        RECT 117.000 182.350 121.925 182.490 ;
        RECT 117.000 182.290 117.320 182.350 ;
        RECT 118.035 182.305 118.625 182.350 ;
        RECT 121.275 182.305 121.925 182.350 ;
        RECT 95.495 182.150 95.785 182.195 ;
        RECT 99.075 182.150 99.365 182.195 ;
        RECT 100.910 182.150 101.200 182.195 ;
        RECT 95.495 182.010 101.200 182.150 ;
        RECT 95.495 181.965 95.785 182.010 ;
        RECT 99.075 181.965 99.365 182.010 ;
        RECT 100.910 181.965 101.200 182.010 ;
        RECT 101.375 182.150 101.665 182.195 ;
        RECT 102.740 182.150 103.060 182.210 ;
        RECT 101.375 182.010 103.060 182.150 ;
        RECT 101.375 181.965 101.665 182.010 ;
        RECT 102.740 181.950 103.060 182.010 ;
        RECT 111.020 182.150 111.340 182.210 ;
        RECT 113.335 182.150 113.625 182.195 ;
        RECT 111.020 182.010 116.770 182.150 ;
        RECT 111.020 181.950 111.340 182.010 ;
        RECT 113.335 181.965 113.625 182.010 ;
        RECT 68.700 181.810 69.020 181.870 ;
        RECT 66.950 181.670 69.020 181.810 ;
        RECT 68.700 181.610 69.020 181.670 ;
        RECT 86.640 181.810 86.960 181.870 ;
        RECT 89.875 181.810 90.165 181.855 ;
        RECT 91.240 181.810 91.560 181.870 ;
        RECT 86.640 181.670 91.560 181.810 ;
        RECT 86.640 181.610 86.960 181.670 ;
        RECT 89.875 181.625 90.165 181.670 ;
        RECT 91.240 181.610 91.560 181.670 ;
        RECT 99.980 181.610 100.300 181.870 ;
        RECT 110.560 181.810 110.880 181.870 ;
        RECT 112.400 181.810 112.720 181.870 ;
        RECT 116.630 181.855 116.770 182.010 ;
        RECT 118.335 181.990 118.625 182.305 ;
        RECT 123.900 182.290 124.220 182.550 ;
        RECT 119.415 182.150 119.705 182.195 ;
        RECT 122.995 182.150 123.285 182.195 ;
        RECT 124.830 182.150 125.120 182.195 ;
        RECT 119.415 182.010 125.120 182.150 ;
        RECT 119.415 181.965 119.705 182.010 ;
        RECT 122.995 181.965 123.285 182.010 ;
        RECT 124.830 181.965 125.120 182.010 ;
        RECT 110.560 181.670 112.720 181.810 ;
        RECT 110.560 181.610 110.880 181.670 ;
        RECT 112.400 181.610 112.720 181.670 ;
        RECT 116.555 181.625 116.845 181.855 ;
        RECT 121.140 181.810 121.460 181.870 ;
        RECT 125.295 181.810 125.585 181.855 ;
        RECT 125.740 181.810 126.060 181.870 ;
        RECT 121.140 181.670 126.060 181.810 ;
        RECT 121.140 181.610 121.460 181.670 ;
        RECT 125.295 181.625 125.585 181.670 ;
        RECT 125.740 181.610 126.060 181.670 ;
        RECT 52.255 181.470 52.545 181.515 ;
        RECT 55.375 181.470 55.665 181.515 ;
        RECT 57.265 181.470 57.555 181.515 ;
        RECT 52.255 181.330 57.555 181.470 ;
        RECT 52.255 181.285 52.545 181.330 ;
        RECT 55.375 181.285 55.665 181.330 ;
        RECT 57.265 181.285 57.555 181.330 ;
        RECT 67.320 181.470 67.640 181.530 ;
        RECT 71.460 181.470 71.780 181.530 ;
        RECT 67.320 181.330 71.780 181.470 ;
        RECT 67.320 181.270 67.640 181.330 ;
        RECT 71.460 181.270 71.780 181.330 ;
        RECT 83.995 181.470 84.285 181.515 ;
        RECT 87.115 181.470 87.405 181.515 ;
        RECT 89.005 181.470 89.295 181.515 ;
        RECT 83.995 181.330 89.295 181.470 ;
        RECT 83.995 181.285 84.285 181.330 ;
        RECT 87.115 181.285 87.405 181.330 ;
        RECT 89.005 181.285 89.295 181.330 ;
        RECT 95.495 181.470 95.785 181.515 ;
        RECT 98.615 181.470 98.905 181.515 ;
        RECT 100.505 181.470 100.795 181.515 ;
        RECT 95.495 181.330 100.795 181.470 ;
        RECT 95.495 181.285 95.785 181.330 ;
        RECT 98.615 181.285 98.905 181.330 ;
        RECT 100.505 181.285 100.795 181.330 ;
        RECT 119.415 181.470 119.705 181.515 ;
        RECT 122.535 181.470 122.825 181.515 ;
        RECT 124.425 181.470 124.715 181.515 ;
        RECT 119.415 181.330 124.715 181.470 ;
        RECT 119.415 181.285 119.705 181.330 ;
        RECT 122.535 181.285 122.825 181.330 ;
        RECT 124.425 181.285 124.715 181.330 ;
        RECT 32.360 180.990 41.330 181.130 ;
        RECT 42.940 181.130 43.260 181.190 ;
        RECT 49.395 181.130 49.685 181.175 ;
        RECT 42.940 180.990 49.685 181.130 ;
        RECT 32.360 180.930 32.680 180.990 ;
        RECT 42.940 180.930 43.260 180.990 ;
        RECT 49.395 180.945 49.685 180.990 ;
        RECT 66.400 181.130 66.720 181.190 ;
        RECT 67.795 181.130 68.085 181.175 ;
        RECT 66.400 180.990 68.085 181.130 ;
        RECT 66.400 180.930 66.720 180.990 ;
        RECT 67.795 180.945 68.085 180.990 ;
        RECT 73.760 180.930 74.080 181.190 ;
        RECT 75.140 180.930 75.460 181.190 ;
        RECT 81.135 181.130 81.425 181.175 ;
        RECT 82.500 181.130 82.820 181.190 ;
        RECT 81.135 180.990 82.820 181.130 ;
        RECT 81.135 180.945 81.425 180.990 ;
        RECT 82.500 180.930 82.820 180.990 ;
        RECT 88.480 181.130 88.800 181.190 ;
        RECT 92.635 181.130 92.925 181.175 ;
        RECT 88.480 180.990 92.925 181.130 ;
        RECT 88.480 180.930 88.800 180.990 ;
        RECT 92.635 180.945 92.925 180.990 ;
        RECT 9.290 180.310 129.350 180.790 ;
        RECT 26.395 180.110 26.685 180.155 ;
        RECT 27.300 180.110 27.620 180.170 ;
        RECT 32.360 180.110 32.680 180.170 ;
        RECT 53.995 180.110 54.285 180.155 ;
        RECT 56.740 180.110 57.060 180.170 ;
        RECT 26.395 179.970 27.620 180.110 ;
        RECT 26.395 179.925 26.685 179.970 ;
        RECT 27.300 179.910 27.620 179.970 ;
        RECT 30.150 179.970 32.680 180.110 ;
        RECT 17.605 179.770 17.895 179.815 ;
        RECT 19.495 179.770 19.785 179.815 ;
        RECT 22.615 179.770 22.905 179.815 ;
        RECT 17.605 179.630 22.905 179.770 ;
        RECT 17.605 179.585 17.895 179.630 ;
        RECT 19.495 179.585 19.785 179.630 ;
        RECT 22.615 179.585 22.905 179.630 ;
        RECT 25.475 179.770 25.765 179.815 ;
        RECT 28.220 179.770 28.540 179.830 ;
        RECT 30.150 179.770 30.290 179.970 ;
        RECT 32.360 179.910 32.680 179.970 ;
        RECT 48.090 179.970 53.750 180.110 ;
        RECT 25.475 179.630 28.910 179.770 ;
        RECT 25.475 179.585 25.765 179.630 ;
        RECT 28.220 179.570 28.540 179.630 ;
        RECT 18.115 179.430 18.405 179.475 ;
        RECT 26.380 179.430 26.700 179.490 ;
        RECT 18.115 179.290 26.700 179.430 ;
        RECT 18.115 179.245 18.405 179.290 ;
        RECT 26.380 179.230 26.700 179.290 ;
        RECT 16.720 178.890 17.040 179.150 ;
        RECT 28.770 179.135 28.910 179.630 ;
        RECT 29.690 179.630 30.290 179.770 ;
        RECT 31.900 179.770 32.220 179.830 ;
        RECT 35.580 179.770 35.900 179.830 ;
        RECT 31.900 179.630 35.900 179.770 ;
        RECT 29.690 179.475 29.830 179.630 ;
        RECT 31.900 179.570 32.220 179.630 ;
        RECT 35.580 179.570 35.900 179.630 ;
        RECT 29.615 179.245 29.905 179.475 ;
        RECT 45.700 179.430 46.020 179.490 ;
        RECT 48.090 179.475 48.230 179.970 ;
        RECT 51.235 179.770 51.525 179.815 ;
        RECT 53.610 179.770 53.750 179.970 ;
        RECT 53.995 179.970 57.060 180.110 ;
        RECT 53.995 179.925 54.285 179.970 ;
        RECT 56.740 179.910 57.060 179.970 ;
        RECT 68.255 180.110 68.545 180.155 ;
        RECT 68.700 180.110 69.020 180.170 ;
        RECT 68.255 179.970 69.020 180.110 ;
        RECT 68.255 179.925 68.545 179.970 ;
        RECT 68.700 179.910 69.020 179.970 ;
        RECT 69.620 180.110 69.940 180.170 ;
        RECT 82.975 180.110 83.265 180.155 ;
        RECT 87.100 180.110 87.420 180.170 ;
        RECT 69.620 179.970 81.810 180.110 ;
        RECT 69.620 179.910 69.940 179.970 ;
        RECT 54.915 179.770 55.205 179.815 ;
        RECT 51.235 179.630 52.140 179.770 ;
        RECT 53.610 179.630 55.205 179.770 ;
        RECT 51.235 179.585 51.525 179.630 ;
        RECT 48.015 179.430 48.305 179.475 ;
        RECT 30.150 179.290 33.050 179.430 ;
        RECT 17.200 179.090 17.490 179.135 ;
        RECT 19.035 179.090 19.325 179.135 ;
        RECT 22.615 179.090 22.905 179.135 ;
        RECT 17.200 178.950 22.905 179.090 ;
        RECT 17.200 178.905 17.490 178.950 ;
        RECT 19.035 178.905 19.325 178.950 ;
        RECT 22.615 178.905 22.905 178.950 ;
        RECT 20.395 178.750 21.045 178.795 ;
        RECT 21.780 178.750 22.100 178.810 ;
        RECT 23.695 178.795 23.985 179.110 ;
        RECT 28.695 179.090 28.985 179.135 ;
        RECT 30.150 179.090 30.290 179.290 ;
        RECT 28.695 178.950 30.290 179.090 ;
        RECT 28.695 178.905 28.985 178.950 ;
        RECT 31.900 178.890 32.220 179.150 ;
        RECT 32.910 179.135 33.050 179.290 ;
        RECT 33.830 179.290 37.190 179.430 ;
        RECT 33.830 179.135 33.970 179.290 ;
        RECT 37.050 179.150 37.190 179.290 ;
        RECT 45.700 179.290 48.305 179.430 ;
        RECT 45.700 179.230 46.020 179.290 ;
        RECT 48.015 179.245 48.305 179.290 ;
        RECT 32.375 178.905 32.665 179.135 ;
        RECT 32.835 178.905 33.125 179.135 ;
        RECT 33.755 178.905 34.045 179.135 ;
        RECT 23.695 178.750 24.285 178.795 ;
        RECT 20.395 178.610 24.285 178.750 ;
        RECT 20.395 178.565 21.045 178.610 ;
        RECT 21.780 178.550 22.100 178.610 ;
        RECT 23.995 178.565 24.285 178.610 ;
        RECT 28.220 178.550 28.540 178.810 ;
        RECT 30.520 178.550 30.840 178.810 ;
        RECT 32.450 178.410 32.590 178.905 ;
        RECT 35.580 178.890 35.900 179.150 ;
        RECT 36.040 178.890 36.360 179.150 ;
        RECT 36.500 178.890 36.820 179.150 ;
        RECT 36.960 179.090 37.280 179.150 ;
        RECT 37.435 179.090 37.725 179.135 ;
        RECT 36.960 178.950 37.725 179.090 ;
        RECT 52.000 179.090 52.140 179.630 ;
        RECT 54.915 179.585 55.205 179.630 ;
        RECT 71.115 179.770 71.405 179.815 ;
        RECT 74.235 179.770 74.525 179.815 ;
        RECT 76.125 179.770 76.415 179.815 ;
        RECT 71.115 179.630 76.415 179.770 ;
        RECT 71.115 179.585 71.405 179.630 ;
        RECT 74.235 179.585 74.525 179.630 ;
        RECT 76.125 179.585 76.415 179.630 ;
        RECT 69.620 179.430 69.940 179.490 ;
        RECT 56.370 179.290 69.940 179.430 ;
        RECT 56.370 179.135 56.510 179.290 ;
        RECT 69.620 179.230 69.940 179.290 ;
        RECT 73.760 179.430 74.080 179.490 ;
        RECT 75.615 179.430 75.905 179.475 ;
        RECT 73.760 179.290 75.905 179.430 ;
        RECT 73.760 179.230 74.080 179.290 ;
        RECT 75.615 179.245 75.905 179.290 ;
        RECT 76.995 179.430 77.285 179.475 ;
        RECT 80.660 179.430 80.980 179.490 ;
        RECT 76.995 179.290 80.980 179.430 ;
        RECT 76.995 179.245 77.285 179.290 ;
        RECT 80.660 179.230 80.980 179.290 ;
        RECT 53.075 179.090 53.365 179.135 ;
        RECT 52.000 178.950 53.365 179.090 ;
        RECT 36.960 178.890 37.280 178.950 ;
        RECT 37.435 178.905 37.725 178.950 ;
        RECT 53.075 178.905 53.365 178.950 ;
        RECT 56.295 178.905 56.585 179.135 ;
        RECT 67.780 179.090 68.100 179.150 ;
        RECT 68.700 179.090 69.020 179.150 ;
        RECT 81.670 179.135 81.810 179.970 ;
        RECT 82.975 179.970 87.420 180.110 ;
        RECT 82.975 179.925 83.265 179.970 ;
        RECT 87.100 179.910 87.420 179.970 ;
        RECT 88.020 179.910 88.340 180.170 ;
        RECT 95.855 180.110 96.145 180.155 ;
        RECT 96.300 180.110 96.620 180.170 ;
        RECT 95.855 179.970 96.620 180.110 ;
        RECT 95.855 179.925 96.145 179.970 ;
        RECT 96.300 179.910 96.620 179.970 ;
        RECT 99.980 179.910 100.300 180.170 ;
        RECT 118.955 179.770 119.245 179.815 ;
        RECT 122.075 179.770 122.365 179.815 ;
        RECT 123.965 179.770 124.255 179.815 ;
        RECT 118.955 179.630 124.255 179.770 ;
        RECT 118.955 179.585 119.245 179.630 ;
        RECT 122.075 179.585 122.365 179.630 ;
        RECT 123.965 179.585 124.255 179.630 ;
        RECT 112.400 179.230 112.720 179.490 ;
        RECT 116.095 179.430 116.385 179.475 ;
        RECT 113.410 179.290 116.385 179.430 ;
        RECT 67.780 178.950 69.020 179.090 ;
        RECT 67.780 178.890 68.100 178.950 ;
        RECT 68.700 178.890 69.020 178.950 ;
        RECT 33.280 178.750 33.600 178.810 ;
        RECT 34.215 178.750 34.505 178.795 ;
        RECT 33.280 178.610 34.505 178.750 ;
        RECT 35.670 178.750 35.810 178.890 ;
        RECT 42.940 178.750 43.260 178.810 ;
        RECT 48.935 178.750 49.225 178.795 ;
        RECT 35.670 178.610 37.650 178.750 ;
        RECT 33.280 178.550 33.600 178.610 ;
        RECT 34.215 178.565 34.505 178.610 ;
        RECT 37.510 178.470 37.650 178.610 ;
        RECT 42.940 178.610 49.225 178.750 ;
        RECT 42.940 178.550 43.260 178.610 ;
        RECT 48.935 178.565 49.225 178.610 ;
        RECT 51.220 178.750 51.540 178.810 ;
        RECT 58.120 178.750 58.440 178.810 ;
        RECT 70.035 178.795 70.325 179.110 ;
        RECT 71.115 179.090 71.405 179.135 ;
        RECT 74.695 179.090 74.985 179.135 ;
        RECT 76.530 179.090 76.820 179.135 ;
        RECT 71.115 178.950 76.820 179.090 ;
        RECT 71.115 178.905 71.405 178.950 ;
        RECT 74.695 178.905 74.985 178.950 ;
        RECT 76.530 178.905 76.820 178.950 ;
        RECT 81.595 178.905 81.885 179.135 ;
        RECT 88.495 179.090 88.785 179.135 ;
        RECT 95.840 179.090 96.160 179.150 ;
        RECT 96.315 179.090 96.605 179.135 ;
        RECT 88.495 178.950 96.605 179.090 ;
        RECT 88.495 178.905 88.785 178.950 ;
        RECT 95.840 178.890 96.160 178.950 ;
        RECT 96.315 178.905 96.605 178.950 ;
        RECT 99.075 179.090 99.365 179.135 ;
        RECT 99.520 179.090 99.840 179.150 ;
        RECT 99.075 178.950 99.840 179.090 ;
        RECT 99.075 178.905 99.365 178.950 ;
        RECT 99.520 178.890 99.840 178.950 ;
        RECT 105.960 179.090 106.280 179.150 ;
        RECT 106.895 179.090 107.185 179.135 ;
        RECT 105.960 178.950 107.185 179.090 ;
        RECT 105.960 178.890 106.280 178.950 ;
        RECT 106.895 178.905 107.185 178.950 ;
        RECT 107.340 178.890 107.660 179.150 ;
        RECT 107.800 178.890 108.120 179.150 ;
        RECT 108.735 178.905 109.025 179.135 ;
        RECT 51.220 178.610 58.440 178.750 ;
        RECT 51.220 178.550 51.540 178.610 ;
        RECT 58.120 178.550 58.440 178.610 ;
        RECT 69.735 178.750 70.325 178.795 ;
        RECT 72.975 178.750 73.625 178.795 ;
        RECT 75.140 178.750 75.460 178.810 ;
        RECT 69.735 178.610 75.460 178.750 ;
        RECT 69.735 178.565 70.025 178.610 ;
        RECT 72.975 178.565 73.625 178.610 ;
        RECT 75.140 178.550 75.460 178.610 ;
        RECT 105.040 178.750 105.360 178.810 ;
        RECT 105.515 178.750 105.805 178.795 ;
        RECT 108.810 178.750 108.950 178.905 ;
        RECT 111.480 178.750 111.800 178.810 ;
        RECT 105.040 178.610 105.805 178.750 ;
        RECT 105.040 178.550 105.360 178.610 ;
        RECT 105.515 178.565 105.805 178.610 ;
        RECT 107.890 178.610 111.800 178.750 ;
        RECT 107.890 178.470 108.030 178.610 ;
        RECT 111.480 178.550 111.800 178.610 ;
        RECT 36.040 178.410 36.360 178.470 ;
        RECT 32.450 178.270 36.360 178.410 ;
        RECT 36.040 178.210 36.360 178.270 ;
        RECT 37.420 178.210 37.740 178.470 ;
        RECT 48.000 178.410 48.320 178.470 ;
        RECT 49.395 178.410 49.685 178.455 ;
        RECT 48.000 178.270 49.685 178.410 ;
        RECT 48.000 178.210 48.320 178.270 ;
        RECT 49.395 178.225 49.685 178.270 ;
        RECT 60.880 178.410 61.200 178.470 ;
        RECT 77.440 178.410 77.760 178.470 ;
        RECT 60.880 178.270 77.760 178.410 ;
        RECT 60.880 178.210 61.200 178.270 ;
        RECT 77.440 178.210 77.760 178.270 ;
        RECT 107.800 178.210 108.120 178.470 ;
        RECT 112.860 178.410 113.180 178.470 ;
        RECT 113.410 178.455 113.550 179.290 ;
        RECT 116.095 179.245 116.385 179.290 ;
        RECT 124.835 179.430 125.125 179.475 ;
        RECT 125.740 179.430 126.060 179.490 ;
        RECT 124.835 179.290 126.060 179.430 ;
        RECT 124.835 179.245 125.125 179.290 ;
        RECT 125.740 179.230 126.060 179.290 ;
        RECT 117.875 178.795 118.165 179.110 ;
        RECT 118.955 179.090 119.245 179.135 ;
        RECT 122.535 179.090 122.825 179.135 ;
        RECT 124.370 179.090 124.660 179.135 ;
        RECT 118.955 178.950 124.660 179.090 ;
        RECT 118.955 178.905 119.245 178.950 ;
        RECT 122.535 178.905 122.825 178.950 ;
        RECT 124.370 178.905 124.660 178.950 ;
        RECT 117.575 178.750 118.165 178.795 ;
        RECT 118.380 178.750 118.700 178.810 ;
        RECT 120.815 178.750 121.465 178.795 ;
        RECT 117.575 178.610 121.465 178.750 ;
        RECT 117.575 178.565 117.865 178.610 ;
        RECT 118.380 178.550 118.700 178.610 ;
        RECT 120.815 178.565 121.465 178.610 ;
        RECT 123.440 178.550 123.760 178.810 ;
        RECT 113.335 178.410 113.625 178.455 ;
        RECT 112.860 178.270 113.625 178.410 ;
        RECT 112.860 178.210 113.180 178.270 ;
        RECT 113.335 178.225 113.625 178.270 ;
        RECT 113.780 178.210 114.100 178.470 ;
        RECT 115.620 178.210 115.940 178.470 ;
        RECT 9.290 177.590 129.350 178.070 ;
        RECT 22.715 177.390 23.005 177.435 ;
        RECT 28.220 177.390 28.540 177.450 ;
        RECT 22.715 177.250 28.540 177.390 ;
        RECT 22.715 177.205 23.005 177.250 ;
        RECT 28.220 177.190 28.540 177.250 ;
        RECT 32.820 177.390 33.140 177.450 ;
        RECT 33.755 177.390 34.045 177.435 ;
        RECT 37.880 177.390 38.200 177.450 ;
        RECT 63.195 177.390 63.485 177.435 ;
        RECT 105.960 177.390 106.280 177.450 ;
        RECT 121.615 177.390 121.905 177.435 ;
        RECT 123.440 177.390 123.760 177.450 ;
        RECT 32.820 177.250 38.200 177.390 ;
        RECT 32.820 177.190 33.140 177.250 ;
        RECT 33.755 177.205 34.045 177.250 ;
        RECT 37.880 177.190 38.200 177.250 ;
        RECT 38.890 177.250 113.550 177.390 ;
        RECT 21.795 177.050 22.085 177.095 ;
        RECT 24.195 177.050 24.485 177.095 ;
        RECT 27.435 177.050 28.085 177.095 ;
        RECT 21.795 176.910 28.085 177.050 ;
        RECT 28.310 177.050 28.450 177.190 ;
        RECT 34.215 177.050 34.505 177.095 ;
        RECT 28.310 176.910 34.505 177.050 ;
        RECT 21.795 176.865 22.085 176.910 ;
        RECT 24.195 176.865 24.785 176.910 ;
        RECT 27.435 176.865 28.085 176.910 ;
        RECT 34.215 176.865 34.505 176.910 ;
        RECT 37.420 177.050 37.740 177.110 ;
        RECT 38.890 177.050 39.030 177.250 ;
        RECT 63.195 177.205 63.485 177.250 ;
        RECT 37.420 176.910 39.030 177.050 ;
        RECT 41.100 177.050 41.420 177.110 ;
        RECT 50.875 177.050 51.165 177.095 ;
        RECT 53.060 177.050 53.380 177.110 ;
        RECT 54.115 177.050 54.765 177.095 ;
        RECT 71.000 177.050 71.320 177.110 ;
        RECT 41.100 176.910 44.090 177.050 ;
        RECT 21.335 176.710 21.625 176.755 ;
        RECT 22.700 176.710 23.020 176.770 ;
        RECT 21.335 176.570 23.020 176.710 ;
        RECT 21.335 176.525 21.625 176.570 ;
        RECT 22.700 176.510 23.020 176.570 ;
        RECT 24.495 176.550 24.785 176.865 ;
        RECT 37.420 176.850 37.740 176.910 ;
        RECT 41.100 176.850 41.420 176.910 ;
        RECT 25.575 176.710 25.865 176.755 ;
        RECT 29.155 176.710 29.445 176.755 ;
        RECT 30.990 176.710 31.280 176.755 ;
        RECT 25.575 176.570 31.280 176.710 ;
        RECT 25.575 176.525 25.865 176.570 ;
        RECT 29.155 176.525 29.445 176.570 ;
        RECT 30.990 176.525 31.280 176.570 ;
        RECT 31.440 176.510 31.760 176.770 ;
        RECT 40.640 176.710 40.960 176.770 ;
        RECT 43.950 176.755 44.090 176.910 ;
        RECT 50.875 176.910 54.765 177.050 ;
        RECT 50.875 176.865 51.465 176.910 ;
        RECT 42.955 176.710 43.245 176.755 ;
        RECT 40.640 176.570 43.245 176.710 ;
        RECT 40.640 176.510 40.960 176.570 ;
        RECT 42.955 176.525 43.245 176.570 ;
        RECT 43.415 176.525 43.705 176.755 ;
        RECT 43.875 176.525 44.165 176.755 ;
        RECT 44.795 176.710 45.085 176.755 ;
        RECT 45.240 176.710 45.560 176.770 ;
        RECT 44.795 176.570 45.560 176.710 ;
        RECT 44.795 176.525 45.085 176.570 ;
        RECT 30.060 176.170 30.380 176.430 ;
        RECT 32.360 176.370 32.680 176.430 ;
        RECT 34.675 176.370 34.965 176.415 ;
        RECT 32.360 176.230 34.965 176.370 ;
        RECT 32.360 176.170 32.680 176.230 ;
        RECT 34.675 176.185 34.965 176.230 ;
        RECT 42.480 176.370 42.800 176.430 ;
        RECT 43.490 176.370 43.630 176.525 ;
        RECT 45.240 176.510 45.560 176.570 ;
        RECT 47.095 176.710 47.385 176.755 ;
        RECT 50.300 176.710 50.620 176.770 ;
        RECT 47.095 176.570 50.620 176.710 ;
        RECT 47.095 176.525 47.385 176.570 ;
        RECT 50.300 176.510 50.620 176.570 ;
        RECT 51.175 176.550 51.465 176.865 ;
        RECT 53.060 176.850 53.380 176.910 ;
        RECT 54.115 176.865 54.765 176.910 ;
        RECT 67.410 176.910 71.320 177.050 ;
        RECT 52.255 176.710 52.545 176.755 ;
        RECT 55.835 176.710 56.125 176.755 ;
        RECT 57.670 176.710 57.960 176.755 ;
        RECT 52.255 176.570 57.960 176.710 ;
        RECT 52.255 176.525 52.545 176.570 ;
        RECT 55.835 176.525 56.125 176.570 ;
        RECT 57.670 176.525 57.960 176.570 ;
        RECT 58.120 176.510 58.440 176.770 ;
        RECT 64.115 176.710 64.405 176.755 ;
        RECT 64.005 176.570 64.405 176.710 ;
        RECT 64.115 176.525 64.405 176.570 ;
        RECT 65.940 176.710 66.260 176.770 ;
        RECT 67.410 176.755 67.550 176.910 ;
        RECT 71.000 176.850 71.320 176.910 ;
        RECT 75.600 177.050 75.920 177.110 ;
        RECT 78.835 177.050 79.125 177.095 ;
        RECT 85.275 177.050 85.565 177.095 ;
        RECT 95.840 177.050 96.160 177.110 ;
        RECT 75.600 176.910 79.125 177.050 ;
        RECT 75.600 176.850 75.920 176.910 ;
        RECT 78.835 176.865 79.125 176.910 ;
        RECT 80.290 176.910 84.110 177.050 ;
        RECT 67.335 176.710 67.625 176.755 ;
        RECT 65.940 176.570 67.625 176.710 ;
        RECT 42.480 176.230 43.630 176.370 ;
        RECT 42.480 176.170 42.800 176.230 ;
        RECT 45.700 176.170 46.020 176.430 ;
        RECT 46.635 176.185 46.925 176.415 ;
        RECT 25.575 176.030 25.865 176.075 ;
        RECT 28.695 176.030 28.985 176.075 ;
        RECT 30.585 176.030 30.875 176.075 ;
        RECT 25.575 175.890 30.875 176.030 ;
        RECT 46.710 176.030 46.850 176.185 ;
        RECT 56.740 176.170 57.060 176.430 ;
        RECT 62.720 176.370 63.040 176.430 ;
        RECT 64.190 176.370 64.330 176.525 ;
        RECT 65.940 176.510 66.260 176.570 ;
        RECT 67.335 176.525 67.625 176.570 ;
        RECT 67.780 176.510 68.100 176.770 ;
        RECT 68.715 176.710 69.005 176.755 ;
        RECT 69.160 176.710 69.480 176.770 ;
        RECT 70.080 176.710 70.400 176.770 ;
        RECT 68.715 176.570 70.400 176.710 ;
        RECT 68.715 176.525 69.005 176.570 ;
        RECT 69.160 176.510 69.480 176.570 ;
        RECT 70.080 176.510 70.400 176.570 ;
        RECT 77.440 176.710 77.760 176.770 ;
        RECT 80.290 176.710 80.430 176.910 ;
        RECT 77.440 176.570 80.430 176.710 ;
        RECT 77.440 176.510 77.760 176.570 ;
        RECT 81.580 176.510 81.900 176.770 ;
        RECT 82.040 176.510 82.360 176.770 ;
        RECT 82.515 176.710 82.805 176.755 ;
        RECT 82.960 176.710 83.280 176.770 ;
        RECT 82.515 176.570 83.280 176.710 ;
        RECT 82.515 176.525 82.805 176.570 ;
        RECT 82.960 176.510 83.280 176.570 ;
        RECT 83.420 176.510 83.740 176.770 ;
        RECT 83.970 176.755 84.110 176.910 ;
        RECT 85.275 176.910 96.160 177.050 ;
        RECT 85.275 176.865 85.565 176.910 ;
        RECT 95.840 176.850 96.160 176.910 ;
        RECT 100.070 176.755 100.210 177.250 ;
        RECT 105.960 177.190 106.280 177.250 ;
        RECT 101.910 176.910 107.570 177.050 ;
        RECT 101.910 176.770 102.050 176.910 ;
        RECT 83.895 176.525 84.185 176.755 ;
        RECT 99.995 176.525 100.285 176.755 ;
        RECT 100.455 176.525 100.745 176.755 ;
        RECT 66.415 176.370 66.705 176.415 ;
        RECT 62.720 176.230 66.705 176.370 ;
        RECT 62.720 176.170 63.040 176.230 ;
        RECT 66.415 176.185 66.705 176.230 ;
        RECT 68.255 176.185 68.545 176.415 ;
        RECT 70.540 176.370 70.860 176.430 ;
        RECT 100.530 176.370 100.670 176.525 ;
        RECT 100.900 176.510 101.220 176.770 ;
        RECT 101.820 176.510 102.140 176.770 ;
        RECT 105.960 176.510 106.280 176.770 ;
        RECT 106.435 176.525 106.725 176.755 ;
        RECT 106.510 176.370 106.650 176.525 ;
        RECT 106.880 176.510 107.200 176.770 ;
        RECT 107.430 176.710 107.570 176.910 ;
        RECT 107.800 176.710 108.120 176.770 ;
        RECT 109.730 176.755 109.870 177.250 ;
        RECT 113.410 177.050 113.550 177.250 ;
        RECT 121.615 177.250 123.760 177.390 ;
        RECT 121.615 177.205 121.905 177.250 ;
        RECT 123.440 177.190 123.760 177.250 ;
        RECT 113.410 176.910 114.010 177.050 ;
        RECT 107.430 176.570 108.120 176.710 ;
        RECT 107.800 176.510 108.120 176.570 ;
        RECT 109.655 176.525 109.945 176.755 ;
        RECT 110.100 176.510 110.420 176.770 ;
        RECT 110.575 176.710 110.865 176.755 ;
        RECT 111.020 176.710 111.340 176.770 ;
        RECT 110.575 176.570 111.340 176.710 ;
        RECT 110.575 176.525 110.865 176.570 ;
        RECT 111.020 176.510 111.340 176.570 ;
        RECT 111.480 176.710 111.800 176.770 ;
        RECT 111.955 176.710 112.245 176.755 ;
        RECT 111.480 176.570 112.245 176.710 ;
        RECT 111.480 176.510 111.800 176.570 ;
        RECT 111.955 176.525 112.245 176.570 ;
        RECT 112.860 176.510 113.180 176.770 ;
        RECT 113.870 176.755 114.010 176.910 ;
        RECT 113.335 176.525 113.625 176.755 ;
        RECT 113.795 176.525 114.085 176.755 ;
        RECT 115.620 176.710 115.940 176.770 ;
        RECT 120.695 176.710 120.985 176.755 ;
        RECT 115.620 176.570 120.985 176.710 ;
        RECT 107.340 176.370 107.660 176.430 ;
        RECT 110.190 176.370 110.330 176.510 ;
        RECT 113.410 176.370 113.550 176.525 ;
        RECT 115.620 176.510 115.940 176.570 ;
        RECT 120.695 176.525 120.985 176.570 ;
        RECT 70.540 176.230 113.550 176.370 ;
        RECT 48.000 176.030 48.320 176.090 ;
        RECT 49.395 176.030 49.685 176.075 ;
        RECT 46.710 175.890 49.685 176.030 ;
        RECT 25.575 175.845 25.865 175.890 ;
        RECT 28.695 175.845 28.985 175.890 ;
        RECT 30.585 175.845 30.875 175.890 ;
        RECT 48.000 175.830 48.320 175.890 ;
        RECT 49.395 175.845 49.685 175.890 ;
        RECT 52.255 176.030 52.545 176.075 ;
        RECT 55.375 176.030 55.665 176.075 ;
        RECT 57.265 176.030 57.555 176.075 ;
        RECT 52.255 175.890 57.555 176.030 ;
        RECT 68.330 176.030 68.470 176.185 ;
        RECT 70.540 176.170 70.860 176.230 ;
        RECT 107.340 176.170 107.660 176.230 ;
        RECT 68.700 176.030 69.020 176.090 ;
        RECT 68.330 175.890 69.020 176.030 ;
        RECT 52.255 175.845 52.545 175.890 ;
        RECT 55.375 175.845 55.665 175.890 ;
        RECT 57.265 175.845 57.555 175.890 ;
        RECT 68.700 175.830 69.020 175.890 ;
        RECT 31.900 175.490 32.220 175.750 ;
        RECT 41.100 175.690 41.420 175.750 ;
        RECT 41.575 175.690 41.865 175.735 ;
        RECT 41.100 175.550 41.865 175.690 ;
        RECT 41.100 175.490 41.420 175.550 ;
        RECT 41.575 175.505 41.865 175.550 ;
        RECT 48.935 175.690 49.225 175.735 ;
        RECT 54.900 175.690 55.220 175.750 ;
        RECT 48.935 175.550 55.220 175.690 ;
        RECT 48.935 175.505 49.225 175.550 ;
        RECT 54.900 175.490 55.220 175.550 ;
        RECT 77.440 175.690 77.760 175.750 ;
        RECT 80.215 175.690 80.505 175.735 ;
        RECT 77.440 175.550 80.505 175.690 ;
        RECT 77.440 175.490 77.760 175.550 ;
        RECT 80.215 175.505 80.505 175.550 ;
        RECT 98.600 175.490 98.920 175.750 ;
        RECT 104.120 175.690 104.440 175.750 ;
        RECT 104.595 175.690 104.885 175.735 ;
        RECT 104.120 175.550 104.885 175.690 ;
        RECT 104.120 175.490 104.440 175.550 ;
        RECT 104.595 175.505 104.885 175.550 ;
        RECT 107.800 175.690 108.120 175.750 ;
        RECT 108.275 175.690 108.565 175.735 ;
        RECT 107.800 175.550 108.565 175.690 ;
        RECT 107.800 175.490 108.120 175.550 ;
        RECT 108.275 175.505 108.565 175.550 ;
        RECT 112.860 175.690 113.180 175.750 ;
        RECT 115.175 175.690 115.465 175.735 ;
        RECT 112.860 175.550 115.465 175.690 ;
        RECT 112.860 175.490 113.180 175.550 ;
        RECT 115.175 175.505 115.465 175.550 ;
        RECT 9.290 174.870 129.350 175.350 ;
        RECT 30.060 174.670 30.380 174.730 ;
        RECT 31.455 174.670 31.745 174.715 ;
        RECT 30.060 174.530 31.745 174.670 ;
        RECT 30.060 174.470 30.380 174.530 ;
        RECT 31.455 174.485 31.745 174.530 ;
        RECT 39.810 174.530 52.140 174.670 ;
        RECT 34.200 174.330 34.520 174.390 ;
        RECT 37.420 174.330 37.740 174.390 ;
        RECT 34.200 174.190 37.740 174.330 ;
        RECT 34.200 174.130 34.520 174.190 ;
        RECT 37.420 174.130 37.740 174.190 ;
        RECT 28.220 173.990 28.540 174.050 ;
        RECT 37.880 173.990 38.200 174.050 ;
        RECT 28.220 173.850 35.350 173.990 ;
        RECT 28.220 173.790 28.540 173.850 ;
        RECT 31.900 173.650 32.220 173.710 ;
        RECT 32.375 173.650 32.665 173.695 ;
        RECT 31.900 173.510 32.665 173.650 ;
        RECT 31.900 173.450 32.220 173.510 ;
        RECT 32.375 173.465 32.665 173.510 ;
        RECT 34.200 173.450 34.520 173.710 ;
        RECT 35.210 173.695 35.350 173.850 ;
        RECT 37.880 173.850 39.490 173.990 ;
        RECT 37.880 173.790 38.200 173.850 ;
        RECT 34.675 173.465 34.965 173.695 ;
        RECT 35.135 173.465 35.425 173.695 ;
        RECT 35.580 173.650 35.900 173.710 ;
        RECT 36.055 173.650 36.345 173.695 ;
        RECT 36.960 173.650 37.280 173.710 ;
        RECT 35.580 173.510 37.280 173.650 ;
        RECT 34.750 173.310 34.890 173.465 ;
        RECT 35.580 173.450 35.900 173.510 ;
        RECT 36.055 173.465 36.345 173.510 ;
        RECT 36.960 173.450 37.280 173.510 ;
        RECT 37.420 173.650 37.740 173.710 ;
        RECT 39.350 173.695 39.490 173.850 ;
        RECT 38.355 173.650 38.645 173.695 ;
        RECT 37.420 173.510 38.645 173.650 ;
        RECT 37.420 173.450 37.740 173.510 ;
        RECT 38.355 173.465 38.645 173.510 ;
        RECT 38.815 173.465 39.105 173.695 ;
        RECT 39.275 173.465 39.565 173.695 ;
        RECT 38.890 173.310 39.030 173.465 ;
        RECT 39.810 173.310 39.950 174.530 ;
        RECT 45.240 174.330 45.560 174.390 ;
        RECT 47.540 174.330 47.860 174.390 ;
        RECT 52.000 174.330 52.140 174.530 ;
        RECT 53.060 174.470 53.380 174.730 ;
        RECT 55.835 174.670 56.125 174.715 ;
        RECT 56.740 174.670 57.060 174.730 ;
        RECT 55.835 174.530 57.060 174.670 ;
        RECT 55.835 174.485 56.125 174.530 ;
        RECT 56.740 174.470 57.060 174.530 ;
        RECT 60.435 174.485 60.725 174.715 ;
        RECT 59.960 174.330 60.280 174.390 ;
        RECT 40.730 174.190 50.990 174.330 ;
        RECT 52.000 174.190 60.280 174.330 ;
        RECT 40.730 173.990 40.870 174.190 ;
        RECT 40.270 173.850 40.870 173.990 ;
        RECT 42.110 173.850 43.630 173.990 ;
        RECT 40.270 173.695 40.410 173.850 ;
        RECT 40.195 173.465 40.485 173.695 ;
        RECT 40.640 173.650 40.960 173.710 ;
        RECT 42.110 173.695 42.250 173.850 ;
        RECT 43.490 173.710 43.630 173.850 ;
        RECT 42.035 173.650 42.325 173.695 ;
        RECT 40.640 173.510 42.325 173.650 ;
        RECT 40.640 173.450 40.960 173.510 ;
        RECT 42.035 173.465 42.325 173.510 ;
        RECT 42.480 173.450 42.800 173.710 ;
        RECT 42.940 173.450 43.260 173.710 ;
        RECT 43.400 173.450 43.720 173.710 ;
        RECT 43.875 173.650 44.165 173.695 ;
        RECT 44.410 173.650 44.550 174.190 ;
        RECT 45.240 174.130 45.560 174.190 ;
        RECT 47.540 174.130 47.860 174.190 ;
        RECT 45.790 173.850 49.610 173.990 ;
        RECT 43.875 173.510 44.550 173.650 ;
        RECT 44.780 173.650 45.100 173.710 ;
        RECT 45.790 173.695 45.930 173.850 ;
        RECT 49.470 173.710 49.610 173.850 ;
        RECT 50.850 173.710 50.990 174.190 ;
        RECT 59.960 174.130 60.280 174.190 ;
        RECT 60.510 173.990 60.650 174.485 ;
        RECT 65.480 174.470 65.800 174.730 ;
        RECT 67.780 174.670 68.100 174.730 ;
        RECT 69.160 174.670 69.480 174.730 ;
        RECT 66.950 174.530 69.480 174.670 ;
        RECT 63.640 174.330 63.960 174.390 ;
        RECT 65.570 174.330 65.710 174.470 ;
        RECT 63.640 174.190 64.790 174.330 ;
        RECT 63.640 174.130 63.960 174.190 ;
        RECT 52.000 173.850 63.870 173.990 ;
        RECT 45.715 173.650 46.005 173.695 ;
        RECT 44.780 173.510 46.005 173.650 ;
        RECT 43.875 173.465 44.165 173.510 ;
        RECT 44.780 173.450 45.100 173.510 ;
        RECT 45.715 173.465 46.005 173.510 ;
        RECT 46.175 173.465 46.465 173.695 ;
        RECT 34.750 173.170 39.950 173.310 ;
        RECT 42.570 173.310 42.710 173.450 ;
        RECT 46.250 173.310 46.390 173.465 ;
        RECT 46.620 173.450 46.940 173.710 ;
        RECT 47.540 173.450 47.860 173.710 ;
        RECT 49.380 173.450 49.700 173.710 ;
        RECT 49.855 173.465 50.145 173.695 ;
        RECT 49.930 173.310 50.070 173.465 ;
        RECT 50.300 173.450 50.620 173.710 ;
        RECT 50.760 173.650 51.080 173.710 ;
        RECT 51.235 173.650 51.525 173.695 ;
        RECT 50.760 173.510 51.525 173.650 ;
        RECT 50.760 173.450 51.080 173.510 ;
        RECT 51.235 173.465 51.525 173.510 ;
        RECT 52.000 173.310 52.140 173.850 ;
        RECT 53.520 173.450 53.840 173.710 ;
        RECT 54.900 173.450 55.220 173.710 ;
        RECT 61.340 173.450 61.660 173.710 ;
        RECT 63.180 173.450 63.500 173.710 ;
        RECT 63.730 173.650 63.870 173.850 ;
        RECT 64.100 173.790 64.420 174.050 ;
        RECT 64.650 174.035 64.790 174.190 ;
        RECT 65.110 174.190 65.710 174.330 ;
        RECT 65.110 174.035 65.250 174.190 ;
        RECT 64.575 173.805 64.865 174.035 ;
        RECT 65.035 173.805 65.325 174.035 ;
        RECT 65.495 173.990 65.785 174.035 ;
        RECT 66.950 173.990 67.090 174.530 ;
        RECT 67.780 174.470 68.100 174.530 ;
        RECT 69.160 174.470 69.480 174.530 ;
        RECT 75.600 174.670 75.920 174.730 ;
        RECT 83.895 174.670 84.185 174.715 ;
        RECT 75.600 174.530 84.185 174.670 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 75.600 174.470 75.920 174.530 ;
        RECT 83.895 174.485 84.185 174.530 ;
        RECT 65.495 173.850 67.090 173.990 ;
        RECT 67.410 174.190 85.950 174.330 ;
        RECT 65.495 173.805 65.785 173.850 ;
        RECT 67.410 173.650 67.550 174.190 ;
        RECT 68.700 173.790 69.020 174.050 ;
        RECT 69.160 173.790 69.480 174.050 ;
        RECT 81.670 173.990 81.810 174.190 ;
        RECT 84.800 173.990 85.120 174.050 ;
        RECT 81.670 173.850 82.270 173.990 ;
        RECT 82.130 173.710 82.270 173.850 ;
        RECT 82.590 173.850 85.120 173.990 ;
        RECT 63.730 173.510 67.550 173.650 ;
        RECT 67.780 173.450 68.100 173.710 ;
        RECT 68.255 173.650 68.545 173.695 ;
        RECT 71.000 173.650 71.320 173.710 ;
        RECT 81.580 173.650 81.900 173.710 ;
        RECT 68.255 173.510 71.320 173.650 ;
        RECT 68.255 173.465 68.545 173.510 ;
        RECT 71.000 173.450 71.320 173.510 ;
        RECT 74.310 173.510 81.900 173.650 ;
        RECT 42.570 173.170 52.140 173.310 ;
        RECT 53.610 173.310 53.750 173.450 ;
        RECT 58.120 173.310 58.440 173.370 ;
        RECT 53.610 173.170 58.440 173.310 ;
        RECT 61.430 173.310 61.570 173.450 ;
        RECT 66.415 173.310 66.705 173.355 ;
        RECT 61.430 173.170 66.705 173.310 ;
        RECT 36.130 173.030 36.270 173.170 ;
        RECT 58.120 173.110 58.440 173.170 ;
        RECT 66.415 173.125 66.705 173.170 ;
        RECT 66.875 173.310 67.165 173.355 ;
        RECT 71.460 173.310 71.780 173.370 ;
        RECT 66.875 173.170 71.780 173.310 ;
        RECT 66.875 173.125 67.165 173.170 ;
        RECT 71.460 173.110 71.780 173.170 ;
        RECT 32.360 172.970 32.680 173.030 ;
        RECT 32.835 172.970 33.125 173.015 ;
        RECT 32.360 172.830 33.125 172.970 ;
        RECT 32.360 172.770 32.680 172.830 ;
        RECT 32.835 172.785 33.125 172.830 ;
        RECT 36.040 172.770 36.360 173.030 ;
        RECT 36.975 172.970 37.265 173.015 ;
        RECT 37.420 172.970 37.740 173.030 ;
        RECT 36.975 172.830 37.740 172.970 ;
        RECT 36.975 172.785 37.265 172.830 ;
        RECT 37.420 172.770 37.740 172.830 ;
        RECT 40.655 172.970 40.945 173.015 ;
        RECT 42.480 172.970 42.800 173.030 ;
        RECT 40.655 172.830 42.800 172.970 ;
        RECT 40.655 172.785 40.945 172.830 ;
        RECT 42.480 172.770 42.800 172.830 ;
        RECT 44.320 172.770 44.640 173.030 ;
        RECT 47.540 172.970 47.860 173.030 ;
        RECT 48.015 172.970 48.305 173.015 ;
        RECT 47.540 172.830 48.305 172.970 ;
        RECT 47.540 172.770 47.860 172.830 ;
        RECT 48.015 172.785 48.305 172.830 ;
        RECT 49.380 172.970 49.700 173.030 ;
        RECT 62.275 172.970 62.565 173.015 ;
        RECT 74.310 172.970 74.450 173.510 ;
        RECT 81.580 173.450 81.900 173.510 ;
        RECT 82.040 173.450 82.360 173.710 ;
        RECT 82.590 173.695 82.730 173.850 ;
        RECT 84.800 173.790 85.120 173.850 ;
        RECT 82.515 173.465 82.805 173.695 ;
        RECT 83.420 173.450 83.740 173.710 ;
        RECT 85.810 173.695 85.950 174.190 ;
        RECT 88.480 173.990 88.800 174.050 ;
        RECT 113.780 173.990 114.100 174.050 ;
        RECT 86.270 173.850 88.800 173.990 ;
        RECT 86.270 173.695 86.410 173.850 ;
        RECT 88.480 173.790 88.800 173.850 ;
        RECT 110.650 173.850 114.100 173.990 ;
        RECT 85.275 173.465 85.565 173.695 ;
        RECT 85.735 173.465 86.025 173.695 ;
        RECT 86.195 173.465 86.485 173.695 ;
        RECT 87.115 173.465 87.405 173.695 ;
        RECT 94.475 173.650 94.765 173.695 ;
        RECT 95.840 173.650 96.160 173.710 ;
        RECT 94.475 173.510 96.160 173.650 ;
        RECT 94.475 173.465 94.765 173.510 ;
        RECT 81.670 173.310 81.810 173.450 ;
        RECT 85.350 173.310 85.490 173.465 ;
        RECT 81.670 173.170 85.490 173.310 ;
        RECT 49.380 172.830 74.450 172.970 ;
        RECT 76.520 172.970 76.840 173.030 ;
        RECT 80.215 172.970 80.505 173.015 ;
        RECT 76.520 172.830 80.505 172.970 ;
        RECT 49.380 172.770 49.700 172.830 ;
        RECT 62.275 172.785 62.565 172.830 ;
        RECT 76.520 172.770 76.840 172.830 ;
        RECT 80.215 172.785 80.505 172.830 ;
        RECT 83.420 172.970 83.740 173.030 ;
        RECT 87.190 172.970 87.330 173.465 ;
        RECT 95.840 173.450 96.160 173.510 ;
        RECT 105.960 173.650 106.280 173.710 ;
        RECT 109.655 173.650 109.945 173.695 ;
        RECT 105.960 173.510 109.945 173.650 ;
        RECT 105.960 173.450 106.280 173.510 ;
        RECT 109.655 173.465 109.945 173.510 ;
        RECT 110.100 173.450 110.420 173.710 ;
        RECT 110.650 173.695 110.790 173.850 ;
        RECT 113.780 173.790 114.100 173.850 ;
        RECT 110.575 173.465 110.865 173.695 ;
        RECT 111.480 173.450 111.800 173.710 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 83.420 172.830 87.330 172.970 ;
        RECT 83.420 172.770 83.740 172.830 ;
        RECT 94.920 172.770 95.240 173.030 ;
        RECT 106.420 172.970 106.740 173.030 ;
        RECT 108.275 172.970 108.565 173.015 ;
        RECT 106.420 172.830 108.565 172.970 ;
        RECT 106.420 172.770 106.740 172.830 ;
        RECT 108.275 172.785 108.565 172.830 ;
        RECT 9.290 172.150 129.350 172.630 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 59.960 171.950 60.280 172.010 ;
        RECT 63.655 171.950 63.945 171.995 ;
        RECT 64.100 171.950 64.420 172.010 ;
        RECT 59.960 171.810 64.420 171.950 ;
        RECT 59.960 171.750 60.280 171.810 ;
        RECT 63.655 171.765 63.945 171.810 ;
        RECT 64.100 171.750 64.420 171.810 ;
        RECT 69.160 171.950 69.480 172.010 ;
        RECT 72.395 171.950 72.685 171.995 ;
        RECT 69.160 171.810 72.685 171.950 ;
        RECT 69.160 171.750 69.480 171.810 ;
        RECT 72.395 171.765 72.685 171.810 ;
        RECT 95.840 171.950 96.160 172.010 ;
        RECT 95.840 171.810 100.440 171.950 ;
        RECT 95.840 171.750 96.160 171.810 ;
        RECT 42.020 171.610 42.340 171.670 ;
        RECT 63.180 171.610 63.500 171.670 ;
        RECT 65.035 171.610 65.325 171.655 ;
        RECT 41.190 171.470 48.230 171.610 ;
        RECT 40.640 171.070 40.960 171.330 ;
        RECT 41.190 171.315 41.330 171.470 ;
        RECT 42.020 171.410 42.340 171.470 ;
        RECT 41.115 171.085 41.405 171.315 ;
        RECT 41.575 171.085 41.865 171.315 ;
        RECT 42.495 171.270 42.785 171.315 ;
        RECT 43.860 171.270 44.180 171.330 ;
        RECT 42.495 171.130 44.180 171.270 ;
        RECT 42.495 171.085 42.785 171.130 ;
        RECT 27.760 170.930 28.080 170.990 ;
        RECT 41.650 170.930 41.790 171.085 ;
        RECT 43.860 171.070 44.180 171.130 ;
        RECT 44.780 171.270 45.100 171.330 ;
        RECT 48.090 171.315 48.230 171.470 ;
        RECT 63.180 171.470 65.325 171.610 ;
        RECT 63.180 171.410 63.500 171.470 ;
        RECT 65.035 171.425 65.325 171.470 ;
        RECT 68.715 171.610 69.005 171.655 ;
        RECT 69.620 171.610 69.940 171.670 ;
        RECT 68.715 171.470 69.940 171.610 ;
        RECT 68.715 171.425 69.005 171.470 ;
        RECT 69.620 171.410 69.940 171.470 ;
        RECT 70.095 171.610 70.385 171.655 ;
        RECT 71.000 171.610 71.320 171.670 ;
        RECT 94.920 171.655 95.240 171.670 ;
        RECT 70.095 171.470 71.320 171.610 ;
        RECT 70.095 171.425 70.385 171.470 ;
        RECT 71.000 171.410 71.320 171.470 ;
        RECT 94.915 171.610 95.565 171.655 ;
        RECT 98.515 171.610 98.805 171.655 ;
        RECT 94.915 171.470 98.805 171.610 ;
        RECT 94.915 171.425 95.565 171.470 ;
        RECT 98.215 171.425 98.805 171.470 ;
        RECT 94.920 171.410 95.240 171.425 ;
        RECT 47.555 171.270 47.845 171.315 ;
        RECT 44.780 171.130 47.845 171.270 ;
        RECT 44.780 171.070 45.100 171.130 ;
        RECT 47.555 171.085 47.845 171.130 ;
        RECT 48.015 171.085 48.305 171.315 ;
        RECT 48.460 171.070 48.780 171.330 ;
        RECT 49.380 171.270 49.700 171.330 ;
        RECT 50.760 171.270 51.080 171.330 ;
        RECT 49.380 171.130 51.080 171.270 ;
        RECT 49.380 171.070 49.700 171.130 ;
        RECT 50.760 171.070 51.080 171.130 ;
        RECT 61.340 171.270 61.660 171.330 ;
        RECT 62.735 171.270 63.025 171.315 ;
        RECT 66.415 171.270 66.705 171.315 ;
        RECT 61.340 171.130 66.705 171.270 ;
        RECT 61.340 171.070 61.660 171.130 ;
        RECT 62.735 171.085 63.025 171.130 ;
        RECT 66.415 171.085 66.705 171.130 ;
        RECT 68.255 171.270 68.545 171.315 ;
        RECT 70.540 171.270 70.860 171.330 ;
        RECT 68.255 171.130 70.860 171.270 ;
        RECT 68.255 171.085 68.545 171.130 ;
        RECT 70.540 171.070 70.860 171.130 ;
        RECT 81.580 171.070 81.900 171.330 ;
        RECT 82.040 171.070 82.360 171.330 ;
        RECT 82.500 171.070 82.820 171.330 ;
        RECT 83.420 171.070 83.740 171.330 ;
        RECT 91.240 171.070 91.560 171.330 ;
        RECT 91.720 171.270 92.010 171.315 ;
        RECT 93.555 171.270 93.845 171.315 ;
        RECT 97.135 171.270 97.425 171.315 ;
        RECT 91.720 171.130 97.425 171.270 ;
        RECT 91.720 171.085 92.010 171.130 ;
        RECT 93.555 171.085 93.845 171.130 ;
        RECT 97.135 171.085 97.425 171.130 ;
        RECT 98.215 171.110 98.505 171.425 ;
        RECT 100.300 171.270 100.440 171.810 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 123.915 171.610 124.205 171.655 ;
        RECT 127.580 171.610 127.900 171.670 ;
        RECT 123.915 171.470 127.900 171.610 ;
        RECT 123.915 171.425 124.205 171.470 ;
        RECT 127.580 171.410 127.900 171.470 ;
        RECT 101.835 171.270 102.125 171.315 ;
        RECT 110.115 171.270 110.405 171.315 ;
        RECT 117.015 171.270 117.305 171.315 ;
        RECT 118.395 171.270 118.685 171.315 ;
        RECT 100.300 171.130 118.685 171.270 ;
        RECT 101.835 171.085 102.125 171.130 ;
        RECT 110.115 171.085 110.405 171.130 ;
        RECT 117.015 171.085 117.305 171.130 ;
        RECT 118.395 171.085 118.685 171.130 ;
        RECT 27.760 170.790 41.790 170.930 ;
        RECT 63.640 170.930 63.960 170.990 ;
        RECT 68.700 170.930 69.020 170.990 ;
        RECT 72.840 170.930 73.160 170.990 ;
        RECT 63.640 170.790 73.160 170.930 ;
        RECT 27.760 170.730 28.080 170.790 ;
        RECT 63.640 170.730 63.960 170.790 ;
        RECT 68.700 170.730 69.020 170.790 ;
        RECT 72.840 170.730 73.160 170.790 ;
        RECT 92.620 170.730 92.940 170.990 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 69.175 170.590 69.465 170.635 ;
        RECT 69.620 170.590 69.940 170.650 ;
        RECT 69.175 170.450 69.940 170.590 ;
        RECT 69.175 170.405 69.465 170.450 ;
        RECT 69.620 170.390 69.940 170.450 ;
        RECT 70.080 170.590 70.400 170.650 ;
        RECT 71.920 170.590 72.240 170.650 ;
        RECT 70.080 170.450 72.240 170.590 ;
        RECT 70.080 170.390 70.400 170.450 ;
        RECT 71.920 170.390 72.240 170.450 ;
        RECT 92.125 170.590 92.415 170.635 ;
        RECT 94.015 170.590 94.305 170.635 ;
        RECT 97.135 170.590 97.425 170.635 ;
        RECT 111.020 170.590 111.340 170.650 ;
        RECT 113.780 170.590 114.100 170.650 ;
        RECT 92.125 170.450 97.425 170.590 ;
        RECT 92.125 170.405 92.415 170.450 ;
        RECT 94.015 170.405 94.305 170.450 ;
        RECT 97.135 170.405 97.425 170.450 ;
        RECT 100.070 170.450 114.100 170.590 ;
        RECT 35.580 170.250 35.900 170.310 ;
        RECT 39.275 170.250 39.565 170.295 ;
        RECT 35.580 170.110 39.565 170.250 ;
        RECT 35.580 170.050 35.900 170.110 ;
        RECT 39.275 170.065 39.565 170.110 ;
        RECT 43.400 170.250 43.720 170.310 ;
        RECT 46.175 170.250 46.465 170.295 ;
        RECT 43.400 170.110 46.465 170.250 ;
        RECT 43.400 170.050 43.720 170.110 ;
        RECT 46.175 170.065 46.465 170.110 ;
        RECT 72.380 170.250 72.700 170.310 ;
        RECT 73.775 170.250 74.065 170.295 ;
        RECT 72.380 170.110 74.065 170.250 ;
        RECT 72.380 170.050 72.700 170.110 ;
        RECT 73.775 170.065 74.065 170.110 ;
        RECT 76.060 170.250 76.380 170.310 ;
        RECT 80.215 170.250 80.505 170.295 ;
        RECT 76.060 170.110 80.505 170.250 ;
        RECT 76.060 170.050 76.380 170.110 ;
        RECT 80.215 170.065 80.505 170.110 ;
        RECT 95.380 170.250 95.700 170.310 ;
        RECT 100.070 170.295 100.210 170.450 ;
        RECT 111.020 170.390 111.340 170.450 ;
        RECT 113.780 170.390 114.100 170.450 ;
        RECT 120.680 170.590 121.000 170.650 ;
        RECT 122.995 170.590 123.285 170.635 ;
        RECT 120.680 170.450 123.285 170.590 ;
        RECT 120.680 170.390 121.000 170.450 ;
        RECT 122.995 170.405 123.285 170.450 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 99.995 170.250 100.285 170.295 ;
        RECT 95.380 170.110 100.285 170.250 ;
        RECT 95.380 170.050 95.700 170.110 ;
        RECT 99.995 170.065 100.285 170.110 ;
        RECT 102.280 170.050 102.600 170.310 ;
        RECT 109.655 170.250 109.945 170.295 ;
        RECT 110.560 170.250 110.880 170.310 ;
        RECT 109.655 170.110 110.880 170.250 ;
        RECT 109.655 170.065 109.945 170.110 ;
        RECT 110.560 170.050 110.880 170.110 ;
        RECT 117.460 170.050 117.780 170.310 ;
        RECT 118.380 170.250 118.700 170.310 ;
        RECT 118.855 170.250 119.145 170.295 ;
        RECT 118.380 170.110 119.145 170.250 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 118.380 170.050 118.700 170.110 ;
        RECT 118.855 170.065 119.145 170.110 ;
        RECT 9.290 169.430 129.350 169.910 ;
        RECT 49.380 169.230 49.700 169.290 ;
        RECT 66.875 169.230 67.165 169.275 ;
        RECT 83.420 169.230 83.740 169.290 ;
        RECT 49.380 169.090 83.740 169.230 ;
        RECT 49.380 169.030 49.700 169.090 ;
        RECT 66.875 169.045 67.165 169.090 ;
        RECT 83.420 169.030 83.740 169.090 ;
        RECT 92.620 169.230 92.940 169.290 ;
        RECT 96.775 169.230 97.065 169.275 ;
        RECT 92.620 169.090 97.065 169.230 ;
        RECT 92.620 169.030 92.940 169.090 ;
        RECT 96.775 169.045 97.065 169.090 ;
        RECT 71.000 168.890 71.320 168.950 ;
        RECT 68.790 168.750 71.320 168.890 ;
        RECT 67.780 168.550 68.100 168.610 ;
        RECT 68.790 168.595 68.930 168.750 ;
        RECT 71.000 168.690 71.320 168.750 ;
        RECT 95.855 168.705 96.145 168.935 ;
        RECT 102.755 168.890 103.045 168.935 ;
        RECT 105.960 168.890 106.280 168.950 ;
        RECT 102.755 168.750 106.280 168.890 ;
        RECT 102.755 168.705 103.045 168.750 ;
        RECT 64.650 168.410 68.100 168.550 ;
        RECT 40.640 168.010 40.960 168.270 ;
        RECT 48.000 168.010 48.320 168.270 ;
        RECT 64.650 168.255 64.790 168.410 ;
        RECT 67.780 168.350 68.100 168.410 ;
        RECT 68.715 168.365 69.005 168.595 ;
        RECT 69.160 168.350 69.480 168.610 ;
        RECT 69.635 168.550 69.925 168.595 ;
        RECT 71.920 168.550 72.240 168.610 ;
        RECT 69.635 168.410 72.240 168.550 ;
        RECT 69.635 168.365 69.925 168.410 ;
        RECT 71.920 168.350 72.240 168.410 ;
        RECT 82.040 168.550 82.360 168.610 ;
        RECT 92.635 168.550 92.925 168.595 ;
        RECT 82.040 168.410 92.925 168.550 ;
        RECT 82.040 168.350 82.360 168.410 ;
        RECT 92.635 168.365 92.925 168.410 ;
        RECT 93.555 168.550 93.845 168.595 ;
        RECT 95.380 168.550 95.700 168.610 ;
        RECT 93.555 168.410 95.700 168.550 ;
        RECT 93.555 168.365 93.845 168.410 ;
        RECT 64.575 168.025 64.865 168.255 ;
        RECT 65.955 168.025 66.245 168.255 ;
        RECT 70.095 168.210 70.385 168.255 ;
        RECT 72.840 168.210 73.160 168.270 ;
        RECT 70.095 168.070 73.160 168.210 ;
        RECT 70.095 168.025 70.385 168.070 ;
        RECT 40.180 167.330 40.500 167.590 ;
        RECT 65.035 167.530 65.325 167.575 ;
        RECT 66.030 167.530 66.170 168.025 ;
        RECT 72.840 168.010 73.160 168.070 ;
        RECT 87.100 168.010 87.420 168.270 ;
        RECT 92.710 168.210 92.850 168.365 ;
        RECT 95.380 168.350 95.700 168.410 ;
        RECT 95.930 168.210 96.070 168.705 ;
        RECT 105.960 168.690 106.280 168.750 ;
        RECT 106.535 168.890 106.825 168.935 ;
        RECT 109.655 168.890 109.945 168.935 ;
        RECT 111.545 168.890 111.835 168.935 ;
        RECT 106.535 168.750 111.835 168.890 ;
        RECT 106.535 168.705 106.825 168.750 ;
        RECT 109.655 168.705 109.945 168.750 ;
        RECT 111.545 168.705 111.835 168.750 ;
        RECT 119.875 168.890 120.165 168.935 ;
        RECT 122.995 168.890 123.285 168.935 ;
        RECT 124.885 168.890 125.175 168.935 ;
        RECT 119.875 168.750 125.175 168.890 ;
        RECT 119.875 168.705 120.165 168.750 ;
        RECT 122.995 168.705 123.285 168.750 ;
        RECT 124.885 168.705 125.175 168.750 ;
        RECT 99.535 168.365 99.825 168.595 ;
        RECT 100.455 168.550 100.745 168.595 ;
        RECT 103.660 168.550 103.980 168.610 ;
        RECT 100.455 168.410 103.980 168.550 ;
        RECT 100.455 168.365 100.745 168.410 ;
        RECT 97.695 168.210 97.985 168.255 ;
        RECT 92.710 168.070 95.610 168.210 ;
        RECT 95.930 168.070 97.985 168.210 ;
        RECT 67.795 167.870 68.085 167.915 ;
        RECT 69.160 167.870 69.480 167.930 ;
        RECT 94.015 167.870 94.305 167.915 ;
        RECT 67.795 167.730 69.480 167.870 ;
        RECT 67.795 167.685 68.085 167.730 ;
        RECT 69.160 167.670 69.480 167.730 ;
        RECT 82.590 167.730 94.305 167.870 ;
        RECT 95.470 167.870 95.610 168.070 ;
        RECT 97.695 168.025 97.985 168.070 ;
        RECT 99.610 167.870 99.750 168.365 ;
        RECT 103.660 168.350 103.980 168.410 ;
        RECT 107.340 168.550 107.660 168.610 ;
        RECT 111.035 168.550 111.325 168.595 ;
        RECT 107.340 168.410 111.325 168.550 ;
        RECT 107.340 168.350 107.660 168.410 ;
        RECT 111.035 168.365 111.325 168.410 ;
        RECT 113.795 168.365 114.085 168.595 ;
        RECT 114.255 168.550 114.545 168.595 ;
        RECT 117.000 168.550 117.320 168.610 ;
        RECT 114.255 168.410 117.320 168.550 ;
        RECT 114.255 168.365 114.545 168.410 ;
        RECT 100.915 168.210 101.205 168.255 ;
        RECT 104.580 168.210 104.900 168.270 ;
        RECT 100.915 168.070 104.900 168.210 ;
        RECT 100.915 168.025 101.205 168.070 ;
        RECT 104.580 168.010 104.900 168.070 ;
        RECT 95.470 167.730 99.750 167.870 ;
        RECT 102.280 167.870 102.600 167.930 ;
        RECT 105.455 167.915 105.745 168.230 ;
        RECT 106.535 168.210 106.825 168.255 ;
        RECT 110.115 168.210 110.405 168.255 ;
        RECT 111.950 168.210 112.240 168.255 ;
        RECT 106.535 168.070 112.240 168.210 ;
        RECT 106.535 168.025 106.825 168.070 ;
        RECT 110.115 168.025 110.405 168.070 ;
        RECT 111.950 168.025 112.240 168.070 ;
        RECT 112.415 168.025 112.705 168.255 ;
        RECT 113.870 168.210 114.010 168.365 ;
        RECT 117.000 168.350 117.320 168.410 ;
        RECT 125.740 168.350 126.060 168.610 ;
        RECT 113.870 168.070 114.470 168.210 ;
        RECT 105.155 167.870 105.745 167.915 ;
        RECT 108.395 167.870 109.045 167.915 ;
        RECT 102.280 167.730 109.045 167.870 ;
        RECT 70.080 167.530 70.400 167.590 ;
        RECT 65.035 167.390 70.400 167.530 ;
        RECT 65.035 167.345 65.325 167.390 ;
        RECT 70.080 167.330 70.400 167.390 ;
        RECT 81.580 167.530 81.900 167.590 ;
        RECT 82.590 167.575 82.730 167.730 ;
        RECT 94.015 167.685 94.305 167.730 ;
        RECT 102.280 167.670 102.600 167.730 ;
        RECT 105.155 167.685 105.445 167.730 ;
        RECT 108.395 167.685 109.045 167.730 ;
        RECT 82.515 167.530 82.805 167.575 ;
        RECT 81.580 167.390 82.805 167.530 ;
        RECT 81.580 167.330 81.900 167.390 ;
        RECT 82.515 167.345 82.805 167.390 ;
        RECT 82.960 167.330 83.280 167.590 ;
        RECT 84.800 167.330 85.120 167.590 ;
        RECT 86.180 167.530 86.500 167.590 ;
        RECT 86.655 167.530 86.945 167.575 ;
        RECT 86.180 167.390 86.945 167.530 ;
        RECT 86.180 167.330 86.500 167.390 ;
        RECT 86.655 167.345 86.945 167.390 ;
        RECT 102.740 167.530 103.060 167.590 ;
        RECT 112.490 167.530 112.630 168.025 ;
        RECT 114.330 167.930 114.470 168.070 ;
        RECT 114.240 167.670 114.560 167.930 ;
        RECT 117.460 167.870 117.780 167.930 ;
        RECT 118.795 167.915 119.085 168.230 ;
        RECT 119.875 168.210 120.165 168.255 ;
        RECT 123.455 168.210 123.745 168.255 ;
        RECT 125.290 168.210 125.580 168.255 ;
        RECT 119.875 168.070 125.580 168.210 ;
        RECT 119.875 168.025 120.165 168.070 ;
        RECT 123.455 168.025 123.745 168.070 ;
        RECT 125.290 168.025 125.580 168.070 ;
        RECT 118.495 167.870 119.085 167.915 ;
        RECT 121.735 167.870 122.385 167.915 ;
        RECT 117.460 167.730 122.385 167.870 ;
        RECT 117.460 167.670 117.780 167.730 ;
        RECT 118.495 167.685 118.785 167.730 ;
        RECT 121.735 167.685 122.385 167.730 ;
        RECT 124.360 167.670 124.680 167.930 ;
        RECT 102.740 167.390 112.630 167.530 ;
        RECT 113.780 167.530 114.100 167.590 ;
        RECT 114.715 167.530 115.005 167.575 ;
        RECT 113.780 167.390 115.005 167.530 ;
        RECT 102.740 167.330 103.060 167.390 ;
        RECT 113.780 167.330 114.100 167.390 ;
        RECT 114.715 167.345 115.005 167.390 ;
        RECT 116.555 167.530 116.845 167.575 ;
        RECT 126.660 167.530 126.980 167.590 ;
        RECT 116.555 167.390 126.980 167.530 ;
        RECT 116.555 167.345 116.845 167.390 ;
        RECT 126.660 167.330 126.980 167.390 ;
        RECT 9.290 166.710 129.350 167.190 ;
        RECT 40.640 166.510 40.960 166.570 ;
        RECT 27.850 166.370 40.960 166.510 ;
        RECT 16.260 165.970 16.580 166.230 ;
        RECT 17.640 166.170 17.960 166.230 ;
        RECT 18.555 166.170 19.205 166.215 ;
        RECT 22.155 166.170 22.445 166.215 ;
        RECT 17.640 166.030 22.445 166.170 ;
        RECT 17.640 165.970 17.960 166.030 ;
        RECT 18.555 165.985 19.205 166.030 ;
        RECT 21.855 165.985 22.445 166.030 ;
        RECT 15.360 165.830 15.650 165.875 ;
        RECT 17.195 165.830 17.485 165.875 ;
        RECT 20.775 165.830 21.065 165.875 ;
        RECT 15.360 165.690 21.065 165.830 ;
        RECT 15.360 165.645 15.650 165.690 ;
        RECT 17.195 165.645 17.485 165.690 ;
        RECT 20.775 165.645 21.065 165.690 ;
        RECT 21.855 165.670 22.145 165.985 ;
        RECT 22.700 165.830 23.020 165.890 ;
        RECT 27.850 165.875 27.990 166.370 ;
        RECT 40.640 166.310 40.960 166.370 ;
        RECT 43.860 166.510 44.180 166.570 ;
        RECT 67.320 166.510 67.640 166.570 ;
        RECT 68.715 166.510 69.005 166.555 ;
        RECT 43.860 166.370 69.005 166.510 ;
        RECT 43.860 166.310 44.180 166.370 ;
        RECT 67.320 166.310 67.640 166.370 ;
        RECT 68.715 166.325 69.005 166.370 ;
        RECT 84.800 166.510 85.120 166.570 ;
        RECT 84.800 166.370 91.930 166.510 ;
        RECT 84.800 166.310 85.120 166.370 ;
        RECT 28.235 166.170 28.525 166.215 ;
        RECT 30.635 166.170 30.925 166.215 ;
        RECT 33.875 166.170 34.525 166.215 ;
        RECT 28.235 166.030 34.525 166.170 ;
        RECT 28.235 165.985 28.525 166.030 ;
        RECT 30.635 165.985 31.225 166.030 ;
        RECT 33.875 165.985 34.525 166.030 ;
        RECT 25.015 165.830 25.305 165.875 ;
        RECT 27.775 165.830 28.065 165.875 ;
        RECT 22.700 165.690 28.065 165.830 ;
        RECT 22.700 165.630 23.020 165.690 ;
        RECT 25.015 165.645 25.305 165.690 ;
        RECT 27.775 165.645 28.065 165.690 ;
        RECT 30.935 165.670 31.225 165.985 ;
        RECT 36.500 165.970 36.820 166.230 ;
        RECT 86.180 166.215 86.500 166.230 ;
        RECT 82.910 166.170 83.200 166.215 ;
        RECT 86.170 166.170 86.500 166.215 ;
        RECT 82.910 166.030 86.500 166.170 ;
        RECT 82.910 165.985 83.200 166.030 ;
        RECT 86.170 165.985 86.500 166.030 ;
        RECT 86.180 165.970 86.500 165.985 ;
        RECT 87.090 166.170 87.380 166.215 ;
        RECT 88.950 166.170 89.240 166.215 ;
        RECT 87.090 166.030 89.240 166.170 ;
        RECT 87.090 165.985 87.380 166.030 ;
        RECT 88.950 165.985 89.240 166.030 ;
        RECT 32.015 165.830 32.305 165.875 ;
        RECT 35.595 165.830 35.885 165.875 ;
        RECT 37.430 165.830 37.720 165.875 ;
        RECT 32.015 165.690 37.720 165.830 ;
        RECT 32.015 165.645 32.305 165.690 ;
        RECT 35.595 165.645 35.885 165.690 ;
        RECT 37.430 165.645 37.720 165.690 ;
        RECT 38.340 165.830 38.660 165.890 ;
        RECT 39.735 165.830 40.025 165.875 ;
        RECT 38.340 165.690 40.025 165.830 ;
        RECT 38.340 165.630 38.660 165.690 ;
        RECT 39.735 165.645 40.025 165.690 ;
        RECT 40.640 165.830 40.960 165.890 ;
        RECT 50.315 165.830 50.605 165.875 ;
        RECT 53.535 165.830 53.825 165.875 ;
        RECT 40.640 165.690 53.825 165.830 ;
        RECT 40.640 165.630 40.960 165.690 ;
        RECT 50.315 165.645 50.605 165.690 ;
        RECT 53.535 165.645 53.825 165.690 ;
        RECT 54.915 165.830 55.205 165.875 ;
        RECT 59.040 165.830 59.360 165.890 ;
        RECT 54.915 165.690 59.360 165.830 ;
        RECT 54.915 165.645 55.205 165.690 ;
        RECT 59.040 165.630 59.360 165.690 ;
        RECT 69.635 165.830 69.925 165.875 ;
        RECT 70.080 165.830 70.400 165.890 ;
        RECT 69.635 165.690 70.400 165.830 ;
        RECT 69.635 165.645 69.925 165.690 ;
        RECT 70.080 165.630 70.400 165.690 ;
        RECT 77.900 165.830 78.220 165.890 ;
        RECT 79.295 165.830 79.585 165.875 ;
        RECT 77.900 165.690 79.585 165.830 ;
        RECT 77.900 165.630 78.220 165.690 ;
        RECT 79.295 165.645 79.585 165.690 ;
        RECT 84.770 165.830 85.060 165.875 ;
        RECT 87.090 165.830 87.305 165.985 ;
        RECT 84.770 165.690 87.305 165.830 ;
        RECT 89.875 165.830 90.165 165.875 ;
        RECT 91.240 165.830 91.560 165.890 ;
        RECT 91.790 165.875 91.930 166.370 ;
        RECT 102.740 166.310 103.060 166.570 ;
        RECT 124.360 166.510 124.680 166.570 ;
        RECT 125.755 166.510 126.045 166.555 ;
        RECT 124.360 166.370 126.045 166.510 ;
        RECT 124.360 166.310 124.680 166.370 ;
        RECT 125.755 166.325 126.045 166.370 ;
        RECT 107.915 166.170 108.205 166.215 ;
        RECT 110.560 166.170 110.880 166.230 ;
        RECT 111.155 166.170 111.805 166.215 ;
        RECT 107.915 166.030 111.805 166.170 ;
        RECT 107.915 165.985 108.505 166.030 ;
        RECT 89.875 165.690 91.560 165.830 ;
        RECT 84.770 165.645 85.060 165.690 ;
        RECT 89.875 165.645 90.165 165.690 ;
        RECT 91.240 165.630 91.560 165.690 ;
        RECT 91.715 165.645 92.005 165.875 ;
        RECT 95.395 165.830 95.685 165.875 ;
        RECT 96.300 165.830 96.620 165.890 ;
        RECT 95.395 165.690 96.620 165.830 ;
        RECT 95.395 165.645 95.685 165.690 ;
        RECT 96.300 165.630 96.620 165.690 ;
        RECT 108.215 165.670 108.505 165.985 ;
        RECT 110.560 165.970 110.880 166.030 ;
        RECT 111.155 165.985 111.805 166.030 ;
        RECT 118.035 166.170 118.325 166.215 ;
        RECT 121.275 166.170 121.925 166.215 ;
        RECT 118.035 166.030 121.925 166.170 ;
        RECT 118.035 165.985 118.625 166.030 ;
        RECT 121.275 165.985 121.925 166.030 ;
        RECT 122.520 166.170 122.840 166.230 ;
        RECT 123.915 166.170 124.205 166.215 ;
        RECT 122.520 166.030 124.205 166.170 ;
        RECT 118.335 165.890 118.625 165.985 ;
        RECT 122.520 165.970 122.840 166.030 ;
        RECT 123.915 165.985 124.205 166.030 ;
        RECT 109.295 165.830 109.585 165.875 ;
        RECT 112.875 165.830 113.165 165.875 ;
        RECT 114.710 165.830 115.000 165.875 ;
        RECT 109.295 165.690 115.000 165.830 ;
        RECT 109.295 165.645 109.585 165.690 ;
        RECT 112.875 165.645 113.165 165.690 ;
        RECT 114.710 165.645 115.000 165.690 ;
        RECT 118.335 165.670 118.700 165.890 ;
        RECT 118.380 165.630 118.700 165.670 ;
        RECT 119.415 165.830 119.705 165.875 ;
        RECT 122.995 165.830 123.285 165.875 ;
        RECT 124.830 165.830 125.120 165.875 ;
        RECT 119.415 165.690 125.120 165.830 ;
        RECT 119.415 165.645 119.705 165.690 ;
        RECT 122.995 165.645 123.285 165.690 ;
        RECT 124.830 165.645 125.120 165.690 ;
        RECT 125.295 165.830 125.585 165.875 ;
        RECT 125.740 165.830 126.060 165.890 ;
        RECT 125.295 165.690 126.060 165.830 ;
        RECT 125.295 165.645 125.585 165.690 ;
        RECT 14.895 165.490 15.185 165.535 ;
        RECT 16.720 165.490 17.040 165.550 ;
        RECT 14.895 165.350 17.040 165.490 ;
        RECT 14.895 165.305 15.185 165.350 ;
        RECT 16.720 165.290 17.040 165.350 ;
        RECT 21.320 165.490 21.640 165.550 ;
        RECT 23.635 165.490 23.925 165.535 ;
        RECT 21.320 165.350 23.925 165.490 ;
        RECT 21.320 165.290 21.640 165.350 ;
        RECT 23.635 165.305 23.925 165.350 ;
        RECT 31.440 165.490 31.760 165.550 ;
        RECT 37.895 165.490 38.185 165.535 ;
        RECT 31.440 165.350 38.185 165.490 ;
        RECT 31.440 165.290 31.760 165.350 ;
        RECT 37.895 165.305 38.185 165.350 ;
        RECT 48.000 165.490 48.320 165.550 ;
        RECT 48.475 165.490 48.765 165.535 ;
        RECT 51.220 165.490 51.540 165.550 ;
        RECT 48.000 165.350 51.540 165.490 ;
        RECT 48.000 165.290 48.320 165.350 ;
        RECT 48.475 165.305 48.765 165.350 ;
        RECT 51.220 165.290 51.540 165.350 ;
        RECT 58.120 165.290 58.440 165.550 ;
        RECT 88.035 165.490 88.325 165.535 ;
        RECT 88.035 165.350 91.010 165.490 ;
        RECT 88.035 165.305 88.325 165.350 ;
        RECT 15.765 165.150 16.055 165.195 ;
        RECT 17.655 165.150 17.945 165.195 ;
        RECT 20.775 165.150 21.065 165.195 ;
        RECT 15.765 165.010 21.065 165.150 ;
        RECT 15.765 164.965 16.055 165.010 ;
        RECT 17.655 164.965 17.945 165.010 ;
        RECT 20.775 164.965 21.065 165.010 ;
        RECT 32.015 165.150 32.305 165.195 ;
        RECT 35.135 165.150 35.425 165.195 ;
        RECT 37.025 165.150 37.315 165.195 ;
        RECT 32.015 165.010 37.315 165.150 ;
        RECT 32.015 164.965 32.305 165.010 ;
        RECT 35.135 164.965 35.425 165.010 ;
        RECT 37.025 164.965 37.315 165.010 ;
        RECT 80.905 165.150 81.195 165.195 ;
        RECT 81.580 165.150 81.900 165.210 ;
        RECT 90.870 165.195 91.010 165.350 ;
        RECT 113.780 165.290 114.100 165.550 ;
        RECT 115.175 165.490 115.465 165.535 ;
        RECT 125.370 165.490 125.510 165.645 ;
        RECT 125.740 165.630 126.060 165.690 ;
        RECT 126.660 165.630 126.980 165.890 ;
        RECT 115.175 165.350 125.510 165.490 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 115.175 165.305 115.465 165.350 ;
        RECT 80.905 165.010 81.900 165.150 ;
        RECT 80.905 164.965 81.195 165.010 ;
        RECT 81.580 164.950 81.900 165.010 ;
        RECT 84.770 165.150 85.060 165.195 ;
        RECT 87.550 165.150 87.840 165.195 ;
        RECT 89.410 165.150 89.700 165.195 ;
        RECT 84.770 165.010 89.700 165.150 ;
        RECT 84.770 164.965 85.060 165.010 ;
        RECT 87.550 164.965 87.840 165.010 ;
        RECT 89.410 164.965 89.700 165.010 ;
        RECT 90.795 164.965 91.085 165.195 ;
        RECT 109.295 165.150 109.585 165.195 ;
        RECT 112.415 165.150 112.705 165.195 ;
        RECT 114.305 165.150 114.595 165.195 ;
        RECT 109.295 165.010 114.595 165.150 ;
        RECT 109.295 164.965 109.585 165.010 ;
        RECT 112.415 164.965 112.705 165.010 ;
        RECT 114.305 164.965 114.595 165.010 ;
        RECT 119.415 165.150 119.705 165.195 ;
        RECT 122.535 165.150 122.825 165.195 ;
        RECT 124.425 165.150 124.715 165.195 ;
        RECT 119.415 165.010 124.715 165.150 ;
        RECT 119.415 164.965 119.705 165.010 ;
        RECT 122.535 164.965 122.825 165.010 ;
        RECT 124.425 164.965 124.715 165.010 ;
        RECT 23.620 164.810 23.940 164.870 ;
        RECT 24.555 164.810 24.845 164.855 ;
        RECT 23.620 164.670 24.845 164.810 ;
        RECT 23.620 164.610 23.940 164.670 ;
        RECT 24.555 164.625 24.845 164.670 ;
        RECT 28.680 164.810 29.000 164.870 ;
        RECT 29.155 164.810 29.445 164.855 ;
        RECT 28.680 164.670 29.445 164.810 ;
        RECT 28.680 164.610 29.000 164.670 ;
        RECT 29.155 164.625 29.445 164.670 ;
        RECT 44.780 164.810 45.100 164.870 ;
        RECT 49.855 164.810 50.145 164.855 ;
        RECT 44.780 164.670 50.145 164.810 ;
        RECT 44.780 164.610 45.100 164.670 ;
        RECT 49.855 164.625 50.145 164.670 ;
        RECT 80.215 164.810 80.505 164.855 ;
        RECT 85.260 164.810 85.580 164.870 ;
        RECT 80.215 164.670 85.580 164.810 ;
        RECT 80.215 164.625 80.505 164.670 ;
        RECT 85.260 164.610 85.580 164.670 ;
        RECT 104.580 164.810 104.900 164.870 ;
        RECT 106.435 164.810 106.725 164.855 ;
        RECT 104.580 164.670 106.725 164.810 ;
        RECT 104.580 164.610 104.900 164.670 ;
        RECT 106.435 164.625 106.725 164.670 ;
        RECT 116.540 164.610 116.860 164.870 ;
        RECT 9.290 163.990 129.350 164.470 ;
        RECT 16.260 163.590 16.580 163.850 ;
        RECT 32.835 163.790 33.125 163.835 ;
        RECT 36.500 163.790 36.820 163.850 ;
        RECT 32.835 163.650 36.820 163.790 ;
        RECT 32.835 163.605 33.125 163.650 ;
        RECT 36.500 163.590 36.820 163.650 ;
        RECT 36.960 163.790 37.280 163.850 ;
        RECT 62.260 163.790 62.580 163.850 ;
        RECT 36.960 163.650 62.580 163.790 ;
        RECT 36.960 163.590 37.280 163.650 ;
        RECT 62.260 163.590 62.580 163.650 ;
        RECT 68.240 163.790 68.560 163.850 ;
        RECT 69.635 163.790 69.925 163.835 ;
        RECT 68.240 163.650 69.925 163.790 ;
        RECT 68.240 163.590 68.560 163.650 ;
        RECT 69.635 163.605 69.925 163.650 ;
        RECT 89.875 163.790 90.165 163.835 ;
        RECT 91.240 163.790 91.560 163.850 ;
        RECT 89.875 163.650 91.560 163.790 ;
        RECT 89.875 163.605 90.165 163.650 ;
        RECT 17.605 163.450 17.895 163.495 ;
        RECT 19.495 163.450 19.785 163.495 ;
        RECT 22.615 163.450 22.905 163.495 ;
        RECT 17.605 163.310 22.905 163.450 ;
        RECT 17.605 163.265 17.895 163.310 ;
        RECT 19.495 163.265 19.785 163.310 ;
        RECT 22.615 163.265 22.905 163.310 ;
        RECT 31.440 163.450 31.760 163.510 ;
        RECT 32.360 163.450 32.680 163.510 ;
        RECT 31.440 163.310 32.680 163.450 ;
        RECT 31.440 163.250 31.760 163.310 ;
        RECT 32.360 163.250 32.680 163.310 ;
        RECT 34.165 163.450 34.455 163.495 ;
        RECT 36.055 163.450 36.345 163.495 ;
        RECT 39.175 163.450 39.465 163.495 ;
        RECT 34.165 163.310 39.465 163.450 ;
        RECT 34.165 163.265 34.455 163.310 ;
        RECT 36.055 163.265 36.345 163.310 ;
        RECT 39.175 163.265 39.465 163.310 ;
        RECT 45.355 163.450 45.645 163.495 ;
        RECT 48.475 163.450 48.765 163.495 ;
        RECT 50.365 163.450 50.655 163.495 ;
        RECT 45.355 163.310 50.655 163.450 ;
        RECT 45.355 163.265 45.645 163.310 ;
        RECT 48.475 163.265 48.765 163.310 ;
        RECT 50.365 163.265 50.655 163.310 ;
        RECT 82.010 163.450 82.300 163.495 ;
        RECT 84.790 163.450 85.080 163.495 ;
        RECT 86.650 163.450 86.940 163.495 ;
        RECT 82.010 163.310 86.940 163.450 ;
        RECT 82.010 163.265 82.300 163.310 ;
        RECT 84.790 163.265 85.080 163.310 ;
        RECT 86.650 163.265 86.940 163.310 ;
        RECT 25.475 163.110 25.765 163.155 ;
        RECT 29.140 163.110 29.460 163.170 ;
        RECT 25.475 162.970 29.460 163.110 ;
        RECT 25.475 162.925 25.765 162.970 ;
        RECT 29.140 162.910 29.460 162.970 ;
        RECT 30.075 163.110 30.365 163.155 ;
        RECT 38.340 163.110 38.660 163.170 ;
        RECT 30.075 162.970 38.660 163.110 ;
        RECT 30.075 162.925 30.365 162.970 ;
        RECT 38.340 162.910 38.660 162.970 ;
        RECT 42.035 163.110 42.325 163.155 ;
        RECT 43.860 163.110 44.180 163.170 ;
        RECT 42.035 162.970 44.180 163.110 ;
        RECT 42.035 162.925 42.325 162.970 ;
        RECT 43.860 162.910 44.180 162.970 ;
        RECT 51.220 162.910 51.540 163.170 ;
        RECT 60.880 163.110 61.200 163.170 ;
        RECT 61.355 163.110 61.645 163.155 ;
        RECT 60.880 162.970 61.645 163.110 ;
        RECT 60.880 162.910 61.200 162.970 ;
        RECT 61.355 162.925 61.645 162.970 ;
        RECT 70.540 162.910 70.860 163.170 ;
        RECT 73.775 163.110 74.065 163.155 ;
        RECT 82.500 163.110 82.820 163.170 ;
        RECT 73.775 162.970 82.820 163.110 ;
        RECT 73.775 162.925 74.065 162.970 ;
        RECT 82.500 162.910 82.820 162.970 ;
        RECT 85.260 162.910 85.580 163.170 ;
        RECT 87.115 163.110 87.405 163.155 ;
        RECT 89.400 163.110 89.720 163.170 ;
        RECT 89.950 163.110 90.090 163.605 ;
        RECT 91.240 163.590 91.560 163.650 ;
        RECT 100.530 163.650 106.650 163.790 ;
        RECT 100.530 163.170 100.670 163.650 ;
        RECT 102.755 163.265 103.045 163.495 ;
        RECT 87.115 162.970 90.090 163.110 ;
        RECT 99.995 163.110 100.285 163.155 ;
        RECT 100.440 163.110 100.760 163.170 ;
        RECT 99.995 162.970 100.760 163.110 ;
        RECT 87.115 162.925 87.405 162.970 ;
        RECT 89.400 162.910 89.720 162.970 ;
        RECT 99.995 162.925 100.285 162.970 ;
        RECT 100.440 162.910 100.760 162.970 ;
        RECT 15.340 162.570 15.660 162.830 ;
        RECT 16.720 162.570 17.040 162.830 ;
        RECT 17.200 162.770 17.490 162.815 ;
        RECT 19.035 162.770 19.325 162.815 ;
        RECT 22.615 162.770 22.905 162.815 ;
        RECT 17.200 162.630 22.905 162.770 ;
        RECT 17.200 162.585 17.490 162.630 ;
        RECT 19.035 162.585 19.325 162.630 ;
        RECT 22.615 162.585 22.905 162.630 ;
        RECT 23.620 162.790 23.940 162.830 ;
        RECT 23.620 162.570 23.985 162.790 ;
        RECT 31.915 162.585 32.205 162.815 ;
        RECT 23.695 162.475 23.985 162.570 ;
        RECT 18.115 162.245 18.405 162.475 ;
        RECT 20.395 162.430 21.045 162.475 ;
        RECT 23.695 162.430 24.285 162.475 ;
        RECT 20.395 162.290 24.285 162.430 ;
        RECT 31.990 162.430 32.130 162.585 ;
        RECT 33.280 162.570 33.600 162.830 ;
        RECT 33.760 162.770 34.050 162.815 ;
        RECT 35.595 162.770 35.885 162.815 ;
        RECT 39.175 162.770 39.465 162.815 ;
        RECT 33.760 162.630 39.465 162.770 ;
        RECT 33.760 162.585 34.050 162.630 ;
        RECT 35.595 162.585 35.885 162.630 ;
        RECT 39.175 162.585 39.465 162.630 ;
        RECT 40.180 162.790 40.500 162.830 ;
        RECT 40.180 162.570 40.545 162.790 ;
        RECT 31.990 162.290 33.050 162.430 ;
        RECT 20.395 162.245 21.045 162.290 ;
        RECT 23.995 162.245 24.285 162.290 ;
        RECT 18.190 162.090 18.330 162.245 ;
        RECT 32.910 162.150 33.050 162.290 ;
        RECT 34.660 162.230 34.980 162.490 ;
        RECT 40.255 162.475 40.545 162.570 ;
        RECT 44.275 162.475 44.565 162.790 ;
        RECT 45.355 162.770 45.645 162.815 ;
        RECT 48.935 162.770 49.225 162.815 ;
        RECT 50.770 162.770 51.060 162.815 ;
        RECT 45.355 162.630 51.060 162.770 ;
        RECT 45.355 162.585 45.645 162.630 ;
        RECT 48.935 162.585 49.225 162.630 ;
        RECT 50.770 162.585 51.060 162.630 ;
        RECT 59.040 162.770 59.360 162.830 ;
        RECT 62.735 162.770 63.025 162.815 ;
        RECT 65.480 162.770 65.800 162.830 ;
        RECT 59.040 162.630 65.800 162.770 ;
        RECT 59.040 162.570 59.360 162.630 ;
        RECT 62.735 162.585 63.025 162.630 ;
        RECT 65.480 162.570 65.800 162.630 ;
        RECT 69.160 162.570 69.480 162.830 ;
        RECT 70.080 162.770 70.400 162.830 ;
        RECT 71.015 162.770 71.305 162.815 ;
        RECT 70.080 162.630 71.305 162.770 ;
        RECT 70.080 162.570 70.400 162.630 ;
        RECT 71.015 162.585 71.305 162.630 ;
        RECT 76.980 162.570 77.300 162.830 ;
        RECT 82.010 162.770 82.300 162.815 ;
        RECT 82.010 162.630 84.545 162.770 ;
        RECT 82.010 162.585 82.300 162.630 ;
        RECT 36.955 162.430 37.605 162.475 ;
        RECT 40.255 162.430 40.845 162.475 ;
        RECT 36.955 162.290 40.845 162.430 ;
        RECT 36.955 162.245 37.605 162.290 ;
        RECT 40.555 162.245 40.845 162.290 ;
        RECT 43.975 162.430 44.565 162.475 ;
        RECT 44.780 162.430 45.100 162.490 ;
        RECT 84.330 162.475 84.545 162.630 ;
        RECT 96.300 162.570 96.620 162.830 ;
        RECT 102.830 162.770 102.970 163.265 ;
        RECT 104.580 163.250 104.900 163.510 ;
        RECT 106.510 163.450 106.650 163.650 ;
        RECT 106.880 163.590 107.200 163.850 ;
        RECT 113.780 163.590 114.100 163.850 ;
        RECT 122.075 163.790 122.365 163.835 ;
        RECT 122.520 163.790 122.840 163.850 ;
        RECT 122.075 163.650 122.840 163.790 ;
        RECT 122.075 163.605 122.365 163.650 ;
        RECT 122.520 163.590 122.840 163.650 ;
        RECT 114.240 163.450 114.560 163.510 ;
        RECT 106.510 163.310 108.030 163.450 ;
        RECT 104.670 163.110 104.810 163.250 ;
        RECT 107.890 163.110 108.030 163.310 ;
        RECT 111.110 163.310 115.850 163.450 ;
        RECT 110.115 163.110 110.405 163.155 ;
        RECT 111.110 163.110 111.250 163.310 ;
        RECT 114.240 163.250 114.560 163.310 ;
        RECT 115.710 163.155 115.850 163.310 ;
        RECT 118.855 163.265 119.145 163.495 ;
        RECT 104.670 162.970 107.570 163.110 ;
        RECT 107.890 162.970 111.250 163.110 ;
        RECT 111.570 162.970 115.390 163.110 ;
        RECT 104.595 162.770 104.885 162.815 ;
        RECT 102.830 162.630 104.885 162.770 ;
        RECT 104.595 162.585 104.885 162.630 ;
        RECT 105.960 162.570 106.280 162.830 ;
        RECT 107.430 162.770 107.570 162.970 ;
        RECT 110.115 162.925 110.405 162.970 ;
        RECT 107.430 162.630 111.250 162.770 ;
        RECT 111.110 162.475 111.250 162.630 ;
        RECT 47.215 162.430 47.865 162.475 ;
        RECT 43.975 162.290 47.865 162.430 ;
        RECT 43.975 162.245 44.265 162.290 ;
        RECT 44.780 162.230 45.100 162.290 ;
        RECT 47.215 162.245 47.865 162.290 ;
        RECT 49.855 162.430 50.145 162.475 ;
        RECT 72.395 162.430 72.685 162.475 ;
        RECT 49.855 162.290 50.990 162.430 ;
        RECT 49.855 162.245 50.145 162.290 ;
        RECT 50.850 162.150 50.990 162.290 ;
        RECT 71.090 162.290 72.685 162.430 ;
        RECT 71.090 162.150 71.230 162.290 ;
        RECT 72.395 162.245 72.685 162.290 ;
        RECT 76.535 162.430 76.825 162.475 ;
        RECT 80.150 162.430 80.440 162.475 ;
        RECT 83.410 162.430 83.700 162.475 ;
        RECT 76.535 162.290 83.700 162.430 ;
        RECT 76.535 162.245 76.825 162.290 ;
        RECT 80.150 162.245 80.440 162.290 ;
        RECT 83.410 162.245 83.700 162.290 ;
        RECT 84.330 162.430 84.620 162.475 ;
        RECT 86.190 162.430 86.480 162.475 ;
        RECT 84.330 162.290 86.480 162.430 ;
        RECT 84.330 162.245 84.620 162.290 ;
        RECT 86.190 162.245 86.480 162.290 ;
        RECT 111.035 162.245 111.325 162.475 ;
        RECT 26.380 162.090 26.700 162.150 ;
        RECT 18.190 161.950 26.700 162.090 ;
        RECT 26.380 161.890 26.700 161.950 ;
        RECT 26.840 161.890 27.160 162.150 ;
        RECT 28.680 161.890 29.000 162.150 ;
        RECT 29.140 161.890 29.460 162.150 ;
        RECT 32.820 161.890 33.140 162.150 ;
        RECT 42.495 162.090 42.785 162.135 ;
        RECT 45.240 162.090 45.560 162.150 ;
        RECT 42.495 161.950 45.560 162.090 ;
        RECT 42.495 161.905 42.785 161.950 ;
        RECT 45.240 161.890 45.560 161.950 ;
        RECT 50.760 161.890 51.080 162.150 ;
        RECT 71.000 161.890 71.320 162.150 ;
        RECT 74.680 162.090 75.000 162.150 ;
        RECT 78.145 162.090 78.435 162.135 ;
        RECT 81.120 162.090 81.440 162.150 ;
        RECT 82.960 162.090 83.280 162.150 ;
        RECT 74.680 161.950 83.280 162.090 ;
        RECT 74.680 161.890 75.000 161.950 ;
        RECT 78.145 161.905 78.435 161.950 ;
        RECT 81.120 161.890 81.440 161.950 ;
        RECT 82.960 161.890 83.280 161.950 ;
        RECT 99.980 162.090 100.300 162.150 ;
        RECT 100.455 162.090 100.745 162.135 ;
        RECT 99.980 161.950 100.745 162.090 ;
        RECT 99.980 161.890 100.300 161.950 ;
        RECT 100.455 161.905 100.745 161.950 ;
        RECT 100.915 162.090 101.205 162.135 ;
        RECT 103.660 162.090 103.980 162.150 ;
        RECT 100.915 161.950 103.980 162.090 ;
        RECT 100.915 161.905 101.205 161.950 ;
        RECT 103.660 161.890 103.980 161.950 ;
        RECT 105.500 161.890 105.820 162.150 ;
        RECT 110.560 162.090 110.880 162.150 ;
        RECT 111.570 162.135 111.710 162.970 ;
        RECT 114.715 162.770 115.005 162.815 ;
        RECT 113.410 162.630 115.005 162.770 ;
        RECT 115.250 162.770 115.390 162.970 ;
        RECT 115.635 162.925 115.925 163.155 ;
        RECT 118.930 163.110 119.070 163.265 ;
        RECT 118.930 162.970 121.370 163.110 ;
        RECT 116.540 162.770 116.860 162.830 ;
        RECT 121.230 162.815 121.370 162.970 ;
        RECT 115.250 162.630 116.860 162.770 ;
        RECT 113.410 162.135 113.550 162.630 ;
        RECT 114.715 162.585 115.005 162.630 ;
        RECT 116.540 162.570 116.860 162.630 ;
        RECT 121.195 162.585 121.485 162.815 ;
        RECT 111.495 162.090 111.785 162.135 ;
        RECT 110.560 161.950 111.785 162.090 ;
        RECT 110.560 161.890 110.880 161.950 ;
        RECT 111.495 161.905 111.785 161.950 ;
        RECT 113.335 161.905 113.625 162.135 ;
        RECT 114.240 162.090 114.560 162.150 ;
        RECT 117.000 162.090 117.320 162.150 ;
        RECT 114.240 161.950 117.320 162.090 ;
        RECT 114.240 161.890 114.560 161.950 ;
        RECT 117.000 161.890 117.320 161.950 ;
        RECT 9.290 161.270 129.350 161.750 ;
        RECT 17.640 161.070 17.960 161.130 ;
        RECT 18.115 161.070 18.405 161.115 ;
        RECT 17.640 160.930 18.405 161.070 ;
        RECT 17.640 160.870 17.960 160.930 ;
        RECT 18.115 160.885 18.405 160.930 ;
        RECT 19.035 160.885 19.325 161.115 ;
        RECT 15.340 160.730 15.660 160.790 ;
        RECT 19.110 160.730 19.250 160.885 ;
        RECT 26.380 160.870 26.700 161.130 ;
        RECT 34.660 161.070 34.980 161.130 ;
        RECT 39.735 161.070 40.025 161.115 ;
        RECT 34.660 160.930 40.025 161.070 ;
        RECT 34.660 160.870 34.980 160.930 ;
        RECT 39.735 160.885 40.025 160.930 ;
        RECT 41.115 160.885 41.405 161.115 ;
        RECT 48.935 160.885 49.225 161.115 ;
        RECT 15.340 160.590 19.250 160.730 ;
        RECT 20.875 160.730 21.165 160.775 ;
        RECT 29.140 160.730 29.460 160.790 ;
        RECT 20.875 160.590 29.460 160.730 ;
        RECT 15.340 160.530 15.660 160.590 ;
        RECT 20.875 160.545 21.165 160.590 ;
        RECT 29.140 160.530 29.460 160.590 ;
        RECT 18.575 160.390 18.865 160.435 ;
        RECT 22.700 160.390 23.020 160.450 ;
        RECT 18.575 160.250 23.020 160.390 ;
        RECT 18.575 160.205 18.865 160.250 ;
        RECT 22.700 160.190 23.020 160.250 ;
        RECT 26.840 160.390 27.160 160.450 ;
        RECT 27.315 160.390 27.605 160.435 ;
        RECT 26.840 160.250 27.605 160.390 ;
        RECT 26.840 160.190 27.160 160.250 ;
        RECT 27.315 160.205 27.605 160.250 ;
        RECT 36.500 160.390 36.820 160.450 ;
        RECT 37.880 160.390 38.200 160.450 ;
        RECT 36.500 160.250 38.200 160.390 ;
        RECT 36.500 160.190 36.820 160.250 ;
        RECT 37.880 160.190 38.200 160.250 ;
        RECT 40.655 160.390 40.945 160.435 ;
        RECT 41.190 160.390 41.330 160.885 ;
        RECT 47.095 160.730 47.385 160.775 ;
        RECT 40.655 160.250 41.330 160.390 ;
        RECT 41.650 160.590 47.385 160.730 ;
        RECT 40.655 160.205 40.945 160.250 ;
        RECT 21.320 159.850 21.640 160.110 ;
        RECT 22.240 160.050 22.560 160.110 ;
        RECT 26.380 160.050 26.700 160.110 ;
        RECT 22.240 159.910 26.700 160.050 ;
        RECT 22.240 159.850 22.560 159.910 ;
        RECT 26.380 159.850 26.700 159.910 ;
        RECT 30.980 160.050 31.300 160.110 ;
        RECT 41.650 160.050 41.790 160.590 ;
        RECT 47.095 160.545 47.385 160.590 ;
        RECT 42.955 160.390 43.245 160.435 ;
        RECT 45.240 160.390 45.560 160.450 ;
        RECT 49.010 160.390 49.150 160.885 ;
        RECT 50.760 160.870 51.080 161.130 ;
        RECT 62.260 161.070 62.580 161.130 ;
        RECT 65.495 161.070 65.785 161.115 ;
        RECT 62.260 160.930 65.785 161.070 ;
        RECT 62.260 160.870 62.580 160.930 ;
        RECT 65.495 160.885 65.785 160.930 ;
        RECT 77.900 161.070 78.220 161.130 ;
        RECT 78.835 161.070 79.125 161.115 ;
        RECT 77.900 160.930 79.125 161.070 ;
        RECT 77.900 160.870 78.220 160.930 ;
        RECT 78.835 160.885 79.125 160.930 ;
        RECT 81.120 160.870 81.440 161.130 ;
        RECT 68.715 160.730 69.005 160.775 ;
        RECT 71.000 160.730 71.320 160.790 ;
        RECT 68.715 160.590 71.320 160.730 ;
        RECT 68.715 160.545 69.005 160.590 ;
        RECT 71.000 160.530 71.320 160.590 ;
        RECT 76.980 160.730 77.300 160.790 ;
        RECT 87.100 160.730 87.420 160.790 ;
        RECT 103.200 160.775 103.520 160.790 ;
        RECT 99.930 160.730 100.220 160.775 ;
        RECT 103.190 160.730 103.520 160.775 ;
        RECT 76.980 160.590 95.150 160.730 ;
        RECT 76.980 160.530 77.300 160.590 ;
        RECT 51.695 160.390 51.985 160.435 ;
        RECT 42.955 160.250 46.850 160.390 ;
        RECT 49.010 160.250 51.985 160.390 ;
        RECT 42.955 160.205 43.245 160.250 ;
        RECT 45.240 160.190 45.560 160.250 ;
        RECT 30.980 159.910 41.790 160.050 ;
        RECT 43.415 160.050 43.705 160.095 ;
        RECT 43.860 160.050 44.180 160.110 ;
        RECT 46.710 160.095 46.850 160.250 ;
        RECT 51.695 160.205 51.985 160.250 ;
        RECT 66.415 160.390 66.705 160.435 ;
        RECT 70.080 160.390 70.400 160.450 ;
        RECT 66.415 160.250 70.400 160.390 ;
        RECT 66.415 160.205 66.705 160.250 ;
        RECT 70.080 160.190 70.400 160.250 ;
        RECT 80.660 160.190 80.980 160.450 ;
        RECT 85.350 160.435 85.490 160.590 ;
        RECT 87.100 160.530 87.420 160.590 ;
        RECT 85.275 160.205 85.565 160.435 ;
        RECT 85.720 160.190 86.040 160.450 ;
        RECT 89.400 160.190 89.720 160.450 ;
        RECT 95.010 160.435 95.150 160.590 ;
        RECT 99.930 160.590 103.520 160.730 ;
        RECT 99.930 160.545 100.220 160.590 ;
        RECT 103.190 160.545 103.520 160.590 ;
        RECT 103.200 160.530 103.520 160.545 ;
        RECT 104.110 160.730 104.400 160.775 ;
        RECT 105.970 160.730 106.260 160.775 ;
        RECT 104.110 160.590 106.260 160.730 ;
        RECT 104.110 160.545 104.400 160.590 ;
        RECT 105.970 160.545 106.260 160.590 ;
        RECT 94.935 160.390 95.225 160.435 ;
        RECT 95.380 160.390 95.700 160.450 ;
        RECT 94.935 160.250 95.700 160.390 ;
        RECT 94.935 160.205 95.225 160.250 ;
        RECT 95.380 160.190 95.700 160.250 ;
        RECT 101.790 160.390 102.080 160.435 ;
        RECT 104.110 160.390 104.325 160.545 ;
        RECT 101.790 160.250 104.325 160.390 ;
        RECT 105.055 160.390 105.345 160.435 ;
        RECT 105.500 160.390 105.820 160.450 ;
        RECT 105.055 160.250 105.820 160.390 ;
        RECT 101.790 160.205 102.080 160.250 ;
        RECT 105.055 160.205 105.345 160.250 ;
        RECT 105.500 160.190 105.820 160.250 ;
        RECT 117.920 160.390 118.240 160.450 ;
        RECT 120.680 160.390 121.000 160.450 ;
        RECT 117.920 160.250 121.000 160.390 ;
        RECT 117.920 160.190 118.240 160.250 ;
        RECT 120.680 160.190 121.000 160.250 ;
        RECT 43.415 159.910 44.180 160.050 ;
        RECT 30.980 159.850 31.300 159.910 ;
        RECT 43.415 159.865 43.705 159.910 ;
        RECT 43.860 159.850 44.180 159.910 ;
        RECT 44.335 160.050 44.625 160.095 ;
        RECT 46.175 160.050 46.465 160.095 ;
        RECT 44.335 159.910 46.465 160.050 ;
        RECT 44.335 159.865 44.625 159.910 ;
        RECT 46.175 159.865 46.465 159.910 ;
        RECT 46.635 160.050 46.925 160.095 ;
        RECT 47.540 160.050 47.860 160.110 ;
        RECT 46.635 159.910 47.860 160.050 ;
        RECT 46.635 159.865 46.925 159.910 ;
        RECT 37.880 159.710 38.200 159.770 ;
        RECT 44.410 159.710 44.550 159.865 ;
        RECT 37.880 159.570 44.550 159.710 ;
        RECT 46.250 159.710 46.390 159.865 ;
        RECT 47.540 159.850 47.860 159.910 ;
        RECT 82.055 160.050 82.345 160.095 ;
        RECT 82.500 160.050 82.820 160.110 ;
        RECT 82.055 159.910 82.820 160.050 ;
        RECT 82.055 159.865 82.345 159.910 ;
        RECT 82.500 159.850 82.820 159.910 ;
        RECT 102.740 160.050 103.060 160.110 ;
        RECT 106.895 160.050 107.185 160.095 ;
        RECT 102.740 159.910 107.185 160.050 ;
        RECT 102.740 159.850 103.060 159.910 ;
        RECT 106.895 159.865 107.185 159.910 ;
        RECT 119.300 159.850 119.620 160.110 ;
        RECT 67.335 159.710 67.625 159.755 ;
        RECT 46.250 159.570 67.625 159.710 ;
        RECT 37.880 159.510 38.200 159.570 ;
        RECT 67.335 159.525 67.625 159.570 ;
        RECT 101.790 159.710 102.080 159.755 ;
        RECT 104.570 159.710 104.860 159.755 ;
        RECT 106.430 159.710 106.720 159.755 ;
        RECT 101.790 159.570 106.720 159.710 ;
        RECT 101.790 159.525 102.080 159.570 ;
        RECT 104.570 159.525 104.860 159.570 ;
        RECT 106.430 159.525 106.720 159.570 ;
        RECT 16.720 159.370 17.040 159.430 ;
        RECT 20.400 159.370 20.720 159.430 ;
        RECT 29.155 159.370 29.445 159.415 ;
        RECT 31.900 159.370 32.220 159.430 ;
        RECT 33.280 159.370 33.600 159.430 ;
        RECT 16.720 159.230 33.600 159.370 ;
        RECT 16.720 159.170 17.040 159.230 ;
        RECT 20.400 159.170 20.720 159.230 ;
        RECT 29.155 159.185 29.445 159.230 ;
        RECT 31.900 159.170 32.220 159.230 ;
        RECT 33.280 159.170 33.600 159.230 ;
        RECT 84.800 159.170 85.120 159.430 ;
        RECT 86.655 159.370 86.945 159.415 ;
        RECT 87.560 159.370 87.880 159.430 ;
        RECT 86.655 159.230 87.880 159.370 ;
        RECT 86.655 159.185 86.945 159.230 ;
        RECT 87.560 159.170 87.880 159.230 ;
        RECT 94.475 159.370 94.765 159.415 ;
        RECT 95.840 159.370 96.160 159.430 ;
        RECT 94.475 159.230 96.160 159.370 ;
        RECT 94.475 159.185 94.765 159.230 ;
        RECT 95.840 159.170 96.160 159.230 ;
        RECT 97.925 159.370 98.215 159.415 ;
        RECT 99.980 159.370 100.300 159.430 ;
        RECT 97.925 159.230 100.300 159.370 ;
        RECT 97.925 159.185 98.215 159.230 ;
        RECT 99.980 159.170 100.300 159.230 ;
        RECT 9.290 158.550 129.350 159.030 ;
        RECT 32.820 158.350 33.140 158.410 ;
        RECT 34.675 158.350 34.965 158.395 ;
        RECT 37.880 158.350 38.200 158.410 ;
        RECT 59.960 158.350 60.280 158.410 ;
        RECT 32.820 158.210 34.965 158.350 ;
        RECT 32.820 158.150 33.140 158.210 ;
        RECT 34.675 158.165 34.965 158.210 ;
        RECT 35.210 158.210 38.200 158.350 ;
        RECT 15.310 158.010 15.600 158.055 ;
        RECT 18.090 158.010 18.380 158.055 ;
        RECT 19.950 158.010 20.240 158.055 ;
        RECT 15.310 157.870 20.240 158.010 ;
        RECT 15.310 157.825 15.600 157.870 ;
        RECT 18.090 157.825 18.380 157.870 ;
        RECT 19.950 157.825 20.240 157.870 ;
        RECT 26.380 158.010 26.700 158.070 ;
        RECT 35.210 158.010 35.350 158.210 ;
        RECT 37.880 158.150 38.200 158.210 ;
        RECT 55.450 158.210 60.280 158.350 ;
        RECT 26.380 157.870 35.350 158.010 ;
        RECT 37.510 157.870 38.570 158.010 ;
        RECT 26.380 157.810 26.700 157.870 ;
        RECT 17.640 157.670 17.960 157.730 ;
        RECT 27.390 157.715 27.530 157.870 ;
        RECT 18.575 157.670 18.865 157.715 ;
        RECT 17.640 157.530 18.865 157.670 ;
        RECT 17.640 157.470 17.960 157.530 ;
        RECT 18.575 157.485 18.865 157.530 ;
        RECT 27.315 157.485 27.605 157.715 ;
        RECT 28.680 157.670 29.000 157.730 ;
        RECT 36.975 157.670 37.265 157.715 ;
        RECT 37.510 157.670 37.650 157.870 ;
        RECT 28.680 157.530 37.650 157.670 ;
        RECT 28.680 157.470 29.000 157.530 ;
        RECT 36.975 157.485 37.265 157.530 ;
        RECT 37.880 157.470 38.200 157.730 ;
        RECT 38.430 157.670 38.570 157.870 ;
        RECT 38.800 157.670 39.120 157.730 ;
        RECT 55.450 157.670 55.590 158.210 ;
        RECT 59.960 158.150 60.280 158.210 ;
        RECT 59.155 158.010 59.445 158.055 ;
        RECT 62.275 158.010 62.565 158.055 ;
        RECT 64.165 158.010 64.455 158.055 ;
        RECT 59.155 157.870 64.455 158.010 ;
        RECT 59.155 157.825 59.445 157.870 ;
        RECT 62.275 157.825 62.565 157.870 ;
        RECT 64.165 157.825 64.455 157.870 ;
        RECT 67.335 158.010 67.625 158.055 ;
        RECT 84.310 158.010 84.600 158.055 ;
        RECT 87.090 158.010 87.380 158.055 ;
        RECT 88.950 158.010 89.240 158.055 ;
        RECT 67.335 157.870 71.230 158.010 ;
        RECT 67.335 157.825 67.625 157.870 ;
        RECT 58.580 157.670 58.900 157.730 ;
        RECT 38.430 157.530 39.120 157.670 ;
        RECT 38.800 157.470 39.120 157.530 ;
        RECT 54.530 157.530 55.590 157.670 ;
        RECT 55.910 157.530 58.900 157.670 ;
        RECT 15.310 157.330 15.600 157.375 ;
        RECT 15.310 157.190 17.845 157.330 ;
        RECT 15.310 157.145 15.600 157.190 ;
        RECT 13.450 156.990 13.740 157.035 ;
        RECT 15.800 156.990 16.120 157.050 ;
        RECT 17.630 157.035 17.845 157.190 ;
        RECT 20.400 157.130 20.720 157.390 ;
        RECT 24.080 157.330 24.400 157.390 ;
        RECT 24.555 157.330 24.845 157.375 ;
        RECT 24.080 157.190 24.845 157.330 ;
        RECT 24.080 157.130 24.400 157.190 ;
        RECT 24.555 157.145 24.845 157.190 ;
        RECT 27.760 157.330 28.080 157.390 ;
        RECT 30.980 157.330 31.300 157.390 ;
        RECT 27.760 157.190 31.300 157.330 ;
        RECT 27.760 157.130 28.080 157.190 ;
        RECT 30.980 157.130 31.300 157.190 ;
        RECT 31.900 157.130 32.220 157.390 ;
        RECT 36.515 157.330 36.805 157.375 ;
        RECT 43.860 157.330 44.180 157.390 ;
        RECT 36.515 157.190 44.180 157.330 ;
        RECT 36.515 157.145 36.805 157.190 ;
        RECT 43.860 157.130 44.180 157.190 ;
        RECT 46.160 157.330 46.480 157.390 ;
        RECT 54.530 157.375 54.670 157.530 ;
        RECT 55.910 157.375 56.050 157.530 ;
        RECT 58.580 157.470 58.900 157.530 ;
        RECT 65.940 157.670 66.260 157.730 ;
        RECT 67.410 157.670 67.550 157.825 ;
        RECT 69.160 157.670 69.480 157.730 ;
        RECT 71.090 157.670 71.230 157.870 ;
        RECT 84.310 157.870 89.240 158.010 ;
        RECT 84.310 157.825 84.600 157.870 ;
        RECT 87.090 157.825 87.380 157.870 ;
        RECT 88.950 157.825 89.240 157.870 ;
        RECT 94.430 158.010 94.720 158.055 ;
        RECT 97.210 158.010 97.500 158.055 ;
        RECT 99.070 158.010 99.360 158.055 ;
        RECT 99.995 158.010 100.285 158.055 ;
        RECT 94.430 157.870 99.360 158.010 ;
        RECT 94.430 157.825 94.720 157.870 ;
        RECT 97.210 157.825 97.500 157.870 ;
        RECT 99.070 157.825 99.360 157.870 ;
        RECT 99.610 157.870 100.285 158.010 ;
        RECT 86.640 157.670 86.960 157.730 ;
        RECT 65.940 157.530 67.550 157.670 ;
        RECT 68.330 157.530 70.310 157.670 ;
        RECT 71.090 157.530 86.960 157.670 ;
        RECT 65.940 157.470 66.260 157.530 ;
        RECT 52.155 157.330 52.445 157.375 ;
        RECT 54.455 157.330 54.745 157.375 ;
        RECT 46.160 157.190 54.745 157.330 ;
        RECT 46.160 157.130 46.480 157.190 ;
        RECT 52.155 157.145 52.445 157.190 ;
        RECT 54.455 157.145 54.745 157.190 ;
        RECT 55.835 157.145 56.125 157.375 ;
        RECT 16.710 156.990 17.000 157.035 ;
        RECT 13.450 156.850 17.000 156.990 ;
        RECT 13.450 156.805 13.740 156.850 ;
        RECT 15.800 156.790 16.120 156.850 ;
        RECT 16.710 156.805 17.000 156.850 ;
        RECT 17.630 156.990 17.920 157.035 ;
        RECT 19.490 156.990 19.780 157.035 ;
        RECT 28.235 156.990 28.525 157.035 ;
        RECT 36.960 156.990 37.280 157.050 ;
        RECT 58.075 157.035 58.365 157.350 ;
        RECT 59.155 157.330 59.445 157.375 ;
        RECT 62.735 157.330 63.025 157.375 ;
        RECT 64.570 157.330 64.860 157.375 ;
        RECT 59.155 157.190 64.860 157.330 ;
        RECT 59.155 157.145 59.445 157.190 ;
        RECT 62.735 157.145 63.025 157.190 ;
        RECT 64.570 157.145 64.860 157.190 ;
        RECT 65.020 157.130 65.340 157.390 ;
        RECT 68.330 157.375 68.470 157.530 ;
        RECT 69.160 157.470 69.480 157.530 ;
        RECT 68.255 157.145 68.545 157.375 ;
        RECT 68.700 157.130 69.020 157.390 ;
        RECT 70.170 157.340 70.310 157.530 ;
        RECT 86.640 157.470 86.960 157.530 ;
        RECT 87.560 157.470 87.880 157.730 ;
        RECT 89.400 157.470 89.720 157.730 ;
        RECT 99.610 157.670 99.750 157.870 ;
        RECT 99.995 157.825 100.285 157.870 ;
        RECT 97.770 157.530 99.750 157.670 ;
        RECT 80.660 157.375 80.980 157.390 ;
        RECT 97.770 157.375 97.910 157.530 ;
        RECT 70.555 157.340 70.845 157.375 ;
        RECT 70.170 157.200 70.845 157.340 ;
        RECT 70.555 157.145 70.845 157.200 ;
        RECT 80.445 157.145 80.980 157.375 ;
        RECT 84.310 157.330 84.600 157.375 ;
        RECT 94.430 157.330 94.720 157.375 ;
        RECT 84.310 157.190 86.845 157.330 ;
        RECT 84.310 157.145 84.600 157.190 ;
        RECT 80.660 157.130 80.980 157.145 ;
        RECT 61.340 157.035 61.660 157.050 ;
        RECT 17.630 156.850 19.780 156.990 ;
        RECT 17.630 156.805 17.920 156.850 ;
        RECT 19.490 156.805 19.780 156.850 ;
        RECT 24.400 156.850 37.280 156.990 ;
        RECT 11.445 156.650 11.735 156.695 ;
        RECT 16.260 156.650 16.580 156.710 ;
        RECT 24.400 156.650 24.540 156.850 ;
        RECT 28.235 156.805 28.525 156.850 ;
        RECT 36.960 156.790 37.280 156.850 ;
        RECT 57.775 156.990 58.365 157.035 ;
        RECT 61.015 156.990 61.665 157.035 ;
        RECT 57.775 156.850 61.665 156.990 ;
        RECT 57.775 156.805 58.065 156.850 ;
        RECT 61.015 156.805 61.665 156.850 ;
        RECT 63.655 156.805 63.945 157.035 ;
        RECT 82.450 156.990 82.740 157.035 ;
        RECT 84.800 156.990 85.120 157.050 ;
        RECT 86.630 157.035 86.845 157.190 ;
        RECT 94.430 157.190 96.965 157.330 ;
        RECT 94.430 157.145 94.720 157.190 ;
        RECT 95.840 157.035 96.160 157.050 ;
        RECT 85.710 156.990 86.000 157.035 ;
        RECT 82.450 156.850 86.000 156.990 ;
        RECT 82.450 156.805 82.740 156.850 ;
        RECT 61.340 156.790 61.660 156.805 ;
        RECT 11.445 156.510 24.540 156.650 ;
        RECT 11.445 156.465 11.735 156.510 ;
        RECT 16.260 156.450 16.580 156.510 ;
        RECT 25.000 156.450 25.320 156.710 ;
        RECT 29.600 156.650 29.920 156.710 ;
        RECT 30.075 156.650 30.365 156.695 ;
        RECT 29.600 156.510 30.365 156.650 ;
        RECT 29.600 156.450 29.920 156.510 ;
        RECT 30.075 156.465 30.365 156.510 ;
        RECT 52.615 156.650 52.905 156.695 ;
        RECT 54.440 156.650 54.760 156.710 ;
        RECT 52.615 156.510 54.760 156.650 ;
        RECT 52.615 156.465 52.905 156.510 ;
        RECT 54.440 156.450 54.760 156.510 ;
        RECT 55.820 156.650 56.140 156.710 ;
        RECT 56.295 156.650 56.585 156.695 ;
        RECT 55.820 156.510 56.585 156.650 ;
        RECT 55.820 156.450 56.140 156.510 ;
        RECT 56.295 156.465 56.585 156.510 ;
        RECT 62.720 156.650 63.040 156.710 ;
        RECT 63.730 156.650 63.870 156.805 ;
        RECT 84.800 156.790 85.120 156.850 ;
        RECT 85.710 156.805 86.000 156.850 ;
        RECT 86.630 156.990 86.920 157.035 ;
        RECT 88.490 156.990 88.780 157.035 ;
        RECT 86.630 156.850 88.780 156.990 ;
        RECT 86.630 156.805 86.920 156.850 ;
        RECT 88.490 156.805 88.780 156.850 ;
        RECT 92.570 156.990 92.860 157.035 ;
        RECT 95.830 156.990 96.160 157.035 ;
        RECT 92.570 156.850 96.160 156.990 ;
        RECT 92.570 156.805 92.860 156.850 ;
        RECT 95.830 156.805 96.160 156.850 ;
        RECT 96.750 157.035 96.965 157.190 ;
        RECT 97.695 157.145 97.985 157.375 ;
        RECT 99.520 157.130 99.840 157.390 ;
        RECT 100.900 157.130 101.220 157.390 ;
        RECT 101.835 157.330 102.125 157.375 ;
        RECT 102.740 157.330 103.060 157.390 ;
        RECT 101.835 157.190 103.060 157.330 ;
        RECT 101.835 157.145 102.125 157.190 ;
        RECT 96.750 156.990 97.040 157.035 ;
        RECT 98.610 156.990 98.900 157.035 ;
        RECT 96.750 156.850 98.900 156.990 ;
        RECT 99.610 156.990 99.750 157.130 ;
        RECT 101.910 156.990 102.050 157.145 ;
        RECT 102.740 157.130 103.060 157.190 ;
        RECT 103.200 157.330 103.520 157.390 ;
        RECT 104.135 157.330 104.425 157.375 ;
        RECT 103.200 157.190 104.425 157.330 ;
        RECT 103.200 157.130 103.520 157.190 ;
        RECT 104.135 157.145 104.425 157.190 ;
        RECT 104.595 157.330 104.885 157.375 ;
        RECT 116.540 157.330 116.860 157.390 ;
        RECT 118.395 157.330 118.685 157.375 ;
        RECT 119.300 157.330 119.620 157.390 ;
        RECT 119.775 157.330 120.065 157.375 ;
        RECT 104.595 157.190 120.065 157.330 ;
        RECT 104.595 157.145 104.885 157.190 ;
        RECT 104.670 156.990 104.810 157.145 ;
        RECT 116.540 157.130 116.860 157.190 ;
        RECT 118.395 157.145 118.685 157.190 ;
        RECT 119.300 157.130 119.620 157.190 ;
        RECT 119.775 157.145 120.065 157.190 ;
        RECT 99.610 156.850 102.050 156.990 ;
        RECT 104.210 156.850 104.810 156.990 ;
        RECT 96.750 156.805 97.040 156.850 ;
        RECT 98.610 156.805 98.900 156.850 ;
        RECT 95.840 156.790 96.160 156.805 ;
        RECT 62.720 156.510 63.870 156.650 ;
        RECT 62.720 156.450 63.040 156.510 ;
        RECT 69.620 156.450 69.940 156.710 ;
        RECT 71.000 156.650 71.320 156.710 ;
        RECT 71.475 156.650 71.765 156.695 ;
        RECT 71.000 156.510 71.765 156.650 ;
        RECT 71.000 156.450 71.320 156.510 ;
        RECT 71.475 156.465 71.765 156.510 ;
        RECT 83.420 156.650 83.740 156.710 ;
        RECT 90.565 156.650 90.855 156.695 ;
        RECT 83.420 156.510 90.855 156.650 ;
        RECT 83.420 156.450 83.740 156.510 ;
        RECT 90.565 156.465 90.855 156.510 ;
        RECT 95.380 156.650 95.700 156.710 ;
        RECT 104.210 156.650 104.350 156.850 ;
        RECT 95.380 156.510 104.350 156.650 ;
        RECT 118.855 156.650 119.145 156.695 ;
        RECT 119.760 156.650 120.080 156.710 ;
        RECT 118.855 156.510 120.080 156.650 ;
        RECT 95.380 156.450 95.700 156.510 ;
        RECT 118.855 156.465 119.145 156.510 ;
        RECT 119.760 156.450 120.080 156.510 ;
        RECT 120.235 156.650 120.525 156.695 ;
        RECT 120.680 156.650 121.000 156.710 ;
        RECT 120.235 156.510 121.000 156.650 ;
        RECT 120.235 156.465 120.525 156.510 ;
        RECT 120.680 156.450 121.000 156.510 ;
        RECT 9.290 155.830 129.350 156.310 ;
        RECT 15.800 155.430 16.120 155.690 ;
        RECT 17.640 155.630 17.960 155.690 ;
        RECT 18.575 155.630 18.865 155.675 ;
        RECT 17.640 155.490 18.865 155.630 ;
        RECT 17.640 155.430 17.960 155.490 ;
        RECT 18.575 155.445 18.865 155.490 ;
        RECT 22.945 155.630 23.235 155.675 ;
        RECT 27.760 155.630 28.080 155.690 ;
        RECT 32.820 155.630 33.140 155.690 ;
        RECT 22.945 155.490 33.140 155.630 ;
        RECT 22.945 155.445 23.235 155.490 ;
        RECT 27.760 155.430 28.080 155.490 ;
        RECT 32.820 155.430 33.140 155.490 ;
        RECT 36.040 155.630 36.360 155.690 ;
        RECT 61.340 155.630 61.660 155.690 ;
        RECT 62.275 155.630 62.565 155.675 ;
        RECT 36.040 155.490 38.110 155.630 ;
        RECT 36.040 155.430 36.360 155.490 ;
        RECT 25.000 155.335 25.320 155.350 ;
        RECT 24.950 155.290 25.320 155.335 ;
        RECT 28.210 155.290 28.500 155.335 ;
        RECT 24.950 155.150 28.500 155.290 ;
        RECT 24.950 155.105 25.320 155.150 ;
        RECT 28.210 155.105 28.500 155.150 ;
        RECT 29.130 155.290 29.420 155.335 ;
        RECT 30.990 155.290 31.280 155.335 ;
        RECT 29.130 155.150 31.280 155.290 ;
        RECT 29.130 155.105 29.420 155.150 ;
        RECT 30.990 155.105 31.280 155.150 ;
        RECT 31.530 155.150 37.650 155.290 ;
        RECT 25.000 155.090 25.320 155.105 ;
        RECT 16.275 154.765 16.565 154.995 ;
        RECT 16.350 154.610 16.490 154.765 ;
        RECT 19.480 154.750 19.800 155.010 ;
        RECT 26.810 154.950 27.100 154.995 ;
        RECT 29.130 154.950 29.345 155.105 ;
        RECT 31.530 154.950 31.670 155.150 ;
        RECT 26.810 154.810 29.345 154.950 ;
        RECT 29.690 154.810 31.670 154.950 ;
        RECT 26.810 154.765 27.100 154.810 ;
        RECT 20.860 154.610 21.180 154.670 ;
        RECT 24.080 154.610 24.400 154.670 ;
        RECT 29.690 154.610 29.830 154.810 ;
        RECT 31.900 154.750 32.220 155.010 ;
        RECT 36.040 154.750 36.360 155.010 ;
        RECT 36.515 154.765 36.805 154.995 ;
        RECT 16.350 154.470 29.830 154.610 ;
        RECT 20.860 154.410 21.180 154.470 ;
        RECT 24.080 154.410 24.400 154.470 ;
        RECT 30.060 154.410 30.380 154.670 ;
        RECT 36.590 154.610 36.730 154.765 ;
        RECT 36.960 154.750 37.280 155.010 ;
        RECT 37.510 154.610 37.650 155.150 ;
        RECT 37.970 154.995 38.110 155.490 ;
        RECT 47.170 155.490 61.110 155.630 ;
        RECT 47.170 155.010 47.310 155.490 ;
        RECT 54.440 155.335 54.760 155.350 ;
        RECT 54.390 155.290 54.760 155.335 ;
        RECT 57.650 155.290 57.940 155.335 ;
        RECT 54.390 155.150 57.940 155.290 ;
        RECT 54.390 155.105 54.760 155.150 ;
        RECT 57.650 155.105 57.940 155.150 ;
        RECT 58.570 155.290 58.860 155.335 ;
        RECT 60.430 155.290 60.720 155.335 ;
        RECT 58.570 155.150 60.720 155.290 ;
        RECT 60.970 155.290 61.110 155.490 ;
        RECT 61.340 155.490 62.565 155.630 ;
        RECT 61.340 155.430 61.660 155.490 ;
        RECT 62.275 155.445 62.565 155.490 ;
        RECT 85.260 155.430 85.580 155.690 ;
        RECT 97.695 155.630 97.985 155.675 ;
        RECT 100.900 155.630 101.220 155.690 ;
        RECT 97.695 155.490 101.220 155.630 ;
        RECT 97.695 155.445 97.985 155.490 ;
        RECT 100.900 155.430 101.220 155.490 ;
        RECT 110.190 155.490 114.930 155.630 ;
        RECT 69.620 155.290 69.940 155.350 ;
        RECT 74.220 155.290 74.540 155.350 ;
        RECT 80.660 155.290 80.980 155.350 ;
        RECT 82.975 155.290 83.265 155.335 ;
        RECT 60.970 155.150 79.050 155.290 ;
        RECT 58.570 155.105 58.860 155.150 ;
        RECT 60.430 155.105 60.720 155.150 ;
        RECT 54.440 155.090 54.760 155.105 ;
        RECT 37.895 154.765 38.185 154.995 ;
        RECT 39.720 154.950 40.040 155.010 ;
        RECT 46.620 154.950 46.940 155.010 ;
        RECT 39.720 154.810 46.940 154.950 ;
        RECT 39.720 154.750 40.040 154.810 ;
        RECT 46.620 154.750 46.940 154.810 ;
        RECT 47.080 154.750 47.400 155.010 ;
        RECT 47.540 154.750 47.860 155.010 ;
        RECT 48.445 154.950 48.735 154.995 ;
        RECT 55.360 154.950 55.680 155.010 ;
        RECT 48.090 154.810 55.680 154.950 ;
        RECT 46.160 154.610 46.480 154.670 ;
        RECT 48.090 154.610 48.230 154.810 ;
        RECT 48.445 154.765 48.735 154.810 ;
        RECT 55.360 154.750 55.680 154.810 ;
        RECT 56.250 154.950 56.540 154.995 ;
        RECT 58.570 154.950 58.785 155.105 ;
        RECT 69.620 155.090 69.940 155.150 ;
        RECT 74.220 155.090 74.540 155.150 ;
        RECT 56.250 154.810 58.785 154.950 ;
        RECT 56.250 154.765 56.540 154.810 ;
        RECT 59.500 154.750 59.820 155.010 ;
        RECT 59.960 154.950 60.280 155.010 ;
        RECT 61.815 154.950 62.105 154.995 ;
        RECT 59.960 154.810 62.105 154.950 ;
        RECT 59.960 154.750 60.280 154.810 ;
        RECT 61.815 154.765 62.105 154.810 ;
        RECT 68.240 154.750 68.560 155.010 ;
        RECT 70.080 154.750 70.400 155.010 ;
        RECT 78.360 154.750 78.680 155.010 ;
        RECT 78.910 154.995 79.050 155.150 ;
        RECT 79.370 155.150 83.265 155.290 ;
        RECT 79.370 154.995 79.510 155.150 ;
        RECT 80.660 155.090 80.980 155.150 ;
        RECT 82.975 155.105 83.265 155.150 ;
        RECT 89.860 155.290 90.180 155.350 ;
        RECT 110.190 155.290 110.330 155.490 ;
        RECT 114.240 155.290 114.560 155.350 ;
        RECT 114.790 155.335 114.930 155.490 ;
        RECT 89.860 155.150 110.330 155.290 ;
        RECT 110.650 155.150 114.560 155.290 ;
        RECT 89.860 155.090 90.180 155.150 ;
        RECT 78.835 154.765 79.125 154.995 ;
        RECT 79.295 154.765 79.585 154.995 ;
        RECT 36.590 154.470 37.190 154.610 ;
        RECT 37.510 154.470 46.480 154.610 ;
        RECT 37.050 154.330 37.190 154.470 ;
        RECT 46.160 154.410 46.480 154.470 ;
        RECT 46.710 154.470 48.230 154.610 ;
        RECT 51.220 154.610 51.540 154.670 ;
        RECT 61.355 154.610 61.645 154.655 ;
        RECT 65.020 154.610 65.340 154.670 ;
        RECT 51.220 154.470 65.340 154.610 ;
        RECT 78.910 154.610 79.050 154.765 ;
        RECT 80.200 154.750 80.520 155.010 ;
        RECT 81.120 154.950 81.440 155.010 ;
        RECT 83.420 154.950 83.740 155.010 ;
        RECT 95.395 154.950 95.685 154.995 ;
        RECT 81.120 154.810 95.685 154.950 ;
        RECT 81.120 154.750 81.440 154.810 ;
        RECT 83.420 154.750 83.740 154.810 ;
        RECT 95.395 154.765 95.685 154.810 ;
        RECT 95.840 154.750 96.160 155.010 ;
        RECT 108.260 154.950 108.580 155.010 ;
        RECT 110.650 154.995 110.790 155.150 ;
        RECT 114.240 155.090 114.560 155.150 ;
        RECT 114.715 155.105 115.005 155.335 ;
        RECT 118.495 155.290 118.785 155.335 ;
        RECT 120.680 155.290 121.000 155.350 ;
        RECT 121.735 155.290 122.385 155.335 ;
        RECT 118.495 155.150 122.385 155.290 ;
        RECT 118.495 155.105 119.085 155.150 ;
        RECT 109.655 154.950 109.945 154.995 ;
        RECT 108.260 154.810 109.945 154.950 ;
        RECT 108.260 154.750 108.580 154.810 ;
        RECT 109.655 154.765 109.945 154.810 ;
        RECT 110.115 154.765 110.405 154.995 ;
        RECT 110.575 154.765 110.865 154.995 ;
        RECT 111.495 154.765 111.785 154.995 ;
        RECT 113.335 154.950 113.625 154.995 ;
        RECT 117.920 154.950 118.240 155.010 ;
        RECT 112.030 154.810 118.240 154.950 ;
        RECT 79.740 154.610 80.060 154.670 ;
        RECT 78.910 154.470 80.060 154.610 ;
        RECT 26.810 154.270 27.100 154.315 ;
        RECT 29.590 154.270 29.880 154.315 ;
        RECT 31.450 154.270 31.740 154.315 ;
        RECT 26.810 154.130 31.740 154.270 ;
        RECT 26.810 154.085 27.100 154.130 ;
        RECT 29.590 154.085 29.880 154.130 ;
        RECT 31.450 154.085 31.740 154.130 ;
        RECT 36.960 154.070 37.280 154.330 ;
        RECT 37.880 154.270 38.200 154.330 ;
        RECT 42.020 154.270 42.340 154.330 ;
        RECT 46.710 154.270 46.850 154.470 ;
        RECT 51.220 154.410 51.540 154.470 ;
        RECT 61.355 154.425 61.645 154.470 ;
        RECT 65.020 154.410 65.340 154.470 ;
        RECT 79.740 154.410 80.060 154.470 ;
        RECT 82.500 154.610 82.820 154.670 ;
        RECT 94.475 154.610 94.765 154.655 ;
        RECT 100.440 154.610 100.760 154.670 ;
        RECT 82.500 154.470 100.760 154.610 ;
        RECT 82.500 154.410 82.820 154.470 ;
        RECT 94.475 154.425 94.765 154.470 ;
        RECT 100.440 154.410 100.760 154.470 ;
        RECT 107.340 154.610 107.660 154.670 ;
        RECT 110.190 154.610 110.330 154.765 ;
        RECT 107.340 154.470 110.330 154.610 ;
        RECT 107.340 154.410 107.660 154.470 ;
        RECT 37.880 154.130 46.850 154.270 ;
        RECT 50.760 154.270 51.080 154.330 ;
        RECT 56.250 154.270 56.540 154.315 ;
        RECT 59.030 154.270 59.320 154.315 ;
        RECT 60.890 154.270 61.180 154.315 ;
        RECT 50.760 154.130 56.050 154.270 ;
        RECT 37.880 154.070 38.200 154.130 ;
        RECT 42.020 154.070 42.340 154.130 ;
        RECT 50.760 154.070 51.080 154.130 ;
        RECT 34.675 153.930 34.965 153.975 ;
        RECT 35.580 153.930 35.900 153.990 ;
        RECT 34.675 153.790 35.900 153.930 ;
        RECT 34.675 153.745 34.965 153.790 ;
        RECT 35.580 153.730 35.900 153.790 ;
        RECT 44.780 153.930 45.100 153.990 ;
        RECT 45.255 153.930 45.545 153.975 ;
        RECT 44.780 153.790 45.545 153.930 ;
        RECT 44.780 153.730 45.100 153.790 ;
        RECT 45.255 153.745 45.545 153.790 ;
        RECT 52.385 153.930 52.675 153.975 ;
        RECT 54.440 153.930 54.760 153.990 ;
        RECT 52.385 153.790 54.760 153.930 ;
        RECT 55.910 153.930 56.050 154.130 ;
        RECT 56.250 154.130 61.180 154.270 ;
        RECT 56.250 154.085 56.540 154.130 ;
        RECT 59.030 154.085 59.320 154.130 ;
        RECT 60.890 154.085 61.180 154.130 ;
        RECT 69.160 154.070 69.480 154.330 ;
        RECT 99.060 154.270 99.380 154.330 ;
        RECT 110.100 154.270 110.420 154.330 ;
        RECT 111.570 154.270 111.710 154.765 ;
        RECT 72.010 154.130 99.380 154.270 ;
        RECT 67.335 153.930 67.625 153.975 ;
        RECT 72.010 153.930 72.150 154.130 ;
        RECT 99.060 154.070 99.380 154.130 ;
        RECT 106.510 154.130 109.870 154.270 ;
        RECT 55.910 153.790 72.150 153.930 ;
        RECT 75.600 153.930 75.920 153.990 ;
        RECT 76.995 153.930 77.285 153.975 ;
        RECT 75.600 153.790 77.285 153.930 ;
        RECT 52.385 153.745 52.675 153.790 ;
        RECT 54.440 153.730 54.760 153.790 ;
        RECT 67.335 153.745 67.625 153.790 ;
        RECT 75.600 153.730 75.920 153.790 ;
        RECT 76.995 153.745 77.285 153.790 ;
        RECT 78.820 153.930 79.140 153.990 ;
        RECT 106.510 153.930 106.650 154.130 ;
        RECT 78.820 153.790 106.650 153.930 ;
        RECT 106.880 153.930 107.200 153.990 ;
        RECT 108.275 153.930 108.565 153.975 ;
        RECT 106.880 153.790 108.565 153.930 ;
        RECT 109.730 153.930 109.870 154.130 ;
        RECT 110.100 154.130 111.710 154.270 ;
        RECT 110.100 154.070 110.420 154.130 ;
        RECT 112.030 153.930 112.170 154.810 ;
        RECT 113.335 154.765 113.625 154.810 ;
        RECT 117.920 154.750 118.240 154.810 ;
        RECT 118.795 154.790 119.085 155.105 ;
        RECT 120.680 155.090 121.000 155.150 ;
        RECT 121.735 155.105 122.385 155.150 ;
        RECT 119.875 154.950 120.165 154.995 ;
        RECT 123.455 154.950 123.745 154.995 ;
        RECT 125.290 154.950 125.580 154.995 ;
        RECT 119.875 154.810 125.580 154.950 ;
        RECT 119.875 154.765 120.165 154.810 ;
        RECT 123.455 154.765 123.745 154.810 ;
        RECT 125.290 154.765 125.580 154.810 ;
        RECT 125.740 154.750 126.060 155.010 ;
        RECT 122.520 154.610 122.840 154.670 ;
        RECT 124.375 154.610 124.665 154.655 ;
        RECT 122.520 154.470 124.665 154.610 ;
        RECT 122.520 154.410 122.840 154.470 ;
        RECT 124.375 154.425 124.665 154.470 ;
        RECT 119.875 154.270 120.165 154.315 ;
        RECT 122.995 154.270 123.285 154.315 ;
        RECT 124.885 154.270 125.175 154.315 ;
        RECT 119.875 154.130 125.175 154.270 ;
        RECT 119.875 154.085 120.165 154.130 ;
        RECT 122.995 154.085 123.285 154.130 ;
        RECT 124.885 154.085 125.175 154.130 ;
        RECT 109.730 153.790 112.170 153.930 ;
        RECT 78.820 153.730 79.140 153.790 ;
        RECT 106.880 153.730 107.200 153.790 ;
        RECT 108.275 153.745 108.565 153.790 ;
        RECT 117.000 153.730 117.320 153.990 ;
        RECT 9.290 153.110 129.350 153.590 ;
        RECT 19.480 152.910 19.800 152.970 ;
        RECT 19.955 152.910 20.245 152.955 ;
        RECT 19.480 152.770 20.245 152.910 ;
        RECT 19.480 152.710 19.800 152.770 ;
        RECT 19.955 152.725 20.245 152.770 ;
        RECT 30.060 152.910 30.380 152.970 ;
        RECT 30.535 152.910 30.825 152.955 ;
        RECT 30.060 152.770 30.825 152.910 ;
        RECT 30.060 152.710 30.380 152.770 ;
        RECT 30.535 152.725 30.825 152.770 ;
        RECT 34.200 152.910 34.520 152.970 ;
        RECT 38.340 152.910 38.660 152.970 ;
        RECT 47.080 152.910 47.400 152.970 ;
        RECT 34.200 152.770 38.660 152.910 ;
        RECT 34.200 152.710 34.520 152.770 ;
        RECT 38.340 152.710 38.660 152.770 ;
        RECT 43.030 152.770 47.400 152.910 ;
        RECT 16.260 152.570 16.580 152.630 ;
        RECT 16.260 152.430 17.870 152.570 ;
        RECT 16.260 152.370 16.580 152.430 ;
        RECT 17.730 152.275 17.870 152.430 ;
        RECT 17.195 152.045 17.485 152.275 ;
        RECT 17.655 152.045 17.945 152.275 ;
        RECT 29.140 152.230 29.460 152.290 ;
        RECT 36.960 152.230 37.280 152.290 ;
        RECT 43.030 152.230 43.170 152.770 ;
        RECT 47.080 152.710 47.400 152.770 ;
        RECT 59.055 152.910 59.345 152.955 ;
        RECT 59.500 152.910 59.820 152.970 ;
        RECT 59.055 152.770 59.820 152.910 ;
        RECT 59.055 152.725 59.345 152.770 ;
        RECT 59.500 152.710 59.820 152.770 ;
        RECT 62.720 152.910 63.040 152.970 ;
        RECT 63.655 152.910 63.945 152.955 ;
        RECT 62.720 152.770 63.945 152.910 ;
        RECT 62.720 152.710 63.040 152.770 ;
        RECT 63.655 152.725 63.945 152.770 ;
        RECT 71.475 152.910 71.765 152.955 ;
        RECT 72.380 152.910 72.700 152.970 ;
        RECT 71.475 152.770 72.700 152.910 ;
        RECT 71.475 152.725 71.765 152.770 ;
        RECT 72.380 152.710 72.700 152.770 ;
        RECT 82.960 152.910 83.280 152.970 ;
        RECT 82.960 152.770 100.670 152.910 ;
        RECT 82.960 152.710 83.280 152.770 ;
        RECT 43.860 152.570 44.180 152.630 ;
        RECT 29.140 152.090 35.350 152.230 ;
        RECT 17.270 151.890 17.410 152.045 ;
        RECT 29.140 152.030 29.460 152.090 ;
        RECT 22.240 151.890 22.560 151.950 ;
        RECT 17.270 151.750 22.560 151.890 ;
        RECT 22.240 151.690 22.560 151.750 ;
        RECT 29.600 151.690 29.920 151.950 ;
        RECT 34.200 151.690 34.520 151.950 ;
        RECT 35.210 151.935 35.350 152.090 ;
        RECT 35.670 152.090 43.170 152.230 ;
        RECT 35.670 151.935 35.810 152.090 ;
        RECT 36.960 152.030 37.280 152.090 ;
        RECT 39.350 151.950 39.490 152.090 ;
        RECT 35.135 151.705 35.425 151.935 ;
        RECT 35.595 151.705 35.885 151.935 ;
        RECT 36.055 151.705 36.345 151.935 ;
        RECT 37.895 151.890 38.185 151.935 ;
        RECT 38.340 151.890 38.660 151.950 ;
        RECT 37.895 151.750 38.660 151.890 ;
        RECT 37.895 151.705 38.185 151.750 ;
        RECT 36.130 151.550 36.270 151.705 ;
        RECT 38.340 151.690 38.660 151.750 ;
        RECT 38.800 151.690 39.120 151.950 ;
        RECT 39.260 151.690 39.580 151.950 ;
        RECT 39.720 151.690 40.040 151.950 ;
        RECT 42.020 151.860 42.340 151.950 ;
        RECT 42.495 151.860 42.785 151.935 ;
        RECT 42.020 151.720 42.785 151.860 ;
        RECT 42.020 151.690 42.340 151.720 ;
        RECT 42.495 151.705 42.785 151.720 ;
        RECT 36.960 151.550 37.280 151.610 ;
        RECT 39.810 151.550 39.950 151.690 ;
        RECT 36.130 151.410 39.950 151.550 ;
        RECT 43.030 151.550 43.170 152.090 ;
        RECT 43.490 152.430 44.180 152.570 ;
        RECT 43.490 151.935 43.630 152.430 ;
        RECT 43.860 152.370 44.180 152.430 ;
        RECT 65.480 152.570 65.800 152.630 ;
        RECT 73.760 152.570 74.080 152.630 ;
        RECT 80.200 152.570 80.520 152.630 ;
        RECT 65.480 152.430 73.530 152.570 ;
        RECT 65.480 152.370 65.800 152.430 ;
        RECT 46.620 152.230 46.940 152.290 ;
        RECT 44.410 152.090 46.940 152.230 ;
        RECT 44.410 151.935 44.550 152.090 ;
        RECT 46.620 152.030 46.940 152.090 ;
        RECT 54.915 152.230 55.205 152.275 ;
        RECT 56.280 152.230 56.600 152.290 ;
        RECT 65.940 152.230 66.260 152.290 ;
        RECT 54.915 152.090 56.600 152.230 ;
        RECT 54.915 152.045 55.205 152.090 ;
        RECT 56.280 152.030 56.600 152.090 ;
        RECT 56.830 152.090 66.260 152.230 ;
        RECT 43.390 151.705 43.680 151.935 ;
        RECT 43.875 151.705 44.165 151.935 ;
        RECT 44.335 151.705 44.625 151.935 ;
        RECT 43.950 151.550 44.090 151.705 ;
        RECT 43.030 151.410 44.090 151.550 ;
        RECT 45.240 151.550 45.560 151.610 ;
        RECT 56.830 151.550 56.970 152.090 ;
        RECT 65.940 152.030 66.260 152.090 ;
        RECT 67.780 152.230 68.100 152.290 ;
        RECT 70.540 152.230 70.860 152.290 ;
        RECT 72.395 152.230 72.685 152.275 ;
        RECT 67.780 152.090 72.685 152.230 ;
        RECT 73.390 152.230 73.530 152.430 ;
        RECT 73.760 152.430 82.270 152.570 ;
        RECT 73.760 152.370 74.080 152.430 ;
        RECT 80.200 152.370 80.520 152.430 ;
        RECT 78.820 152.230 79.140 152.290 ;
        RECT 81.580 152.230 81.900 152.290 ;
        RECT 73.390 152.090 79.140 152.230 ;
        RECT 67.780 152.030 68.100 152.090 ;
        RECT 70.540 152.030 70.860 152.090 ;
        RECT 72.395 152.045 72.685 152.090 ;
        RECT 78.820 152.030 79.140 152.090 ;
        RECT 80.290 152.090 81.900 152.230 ;
        RECT 58.135 151.890 58.425 151.935 ;
        RECT 45.240 151.410 56.970 151.550 ;
        RECT 57.750 151.750 58.425 151.890 ;
        RECT 36.960 151.350 37.280 151.410 ;
        RECT 45.240 151.350 45.560 151.410 ;
        RECT 17.640 151.210 17.960 151.270 ;
        RECT 18.115 151.210 18.405 151.255 ;
        RECT 17.640 151.070 18.405 151.210 ;
        RECT 17.640 151.010 17.960 151.070 ;
        RECT 18.115 151.025 18.405 151.070 ;
        RECT 37.435 151.210 37.725 151.255 ;
        RECT 38.800 151.210 39.120 151.270 ;
        RECT 37.435 151.070 39.120 151.210 ;
        RECT 37.435 151.025 37.725 151.070 ;
        RECT 38.800 151.010 39.120 151.070 ;
        RECT 41.115 151.210 41.405 151.255 ;
        RECT 43.860 151.210 44.180 151.270 ;
        RECT 41.115 151.070 44.180 151.210 ;
        RECT 41.115 151.025 41.405 151.070 ;
        RECT 43.860 151.010 44.180 151.070 ;
        RECT 45.715 151.210 46.005 151.255 ;
        RECT 47.540 151.210 47.860 151.270 ;
        RECT 45.715 151.070 47.860 151.210 ;
        RECT 45.715 151.025 46.005 151.070 ;
        RECT 47.540 151.010 47.860 151.070 ;
        RECT 54.440 151.210 54.760 151.270 ;
        RECT 55.375 151.210 55.665 151.255 ;
        RECT 54.440 151.070 55.665 151.210 ;
        RECT 54.440 151.010 54.760 151.070 ;
        RECT 55.375 151.025 55.665 151.070 ;
        RECT 55.820 151.010 56.140 151.270 ;
        RECT 57.750 151.255 57.890 151.750 ;
        RECT 58.135 151.705 58.425 151.750 ;
        RECT 62.720 151.690 63.040 151.950 ;
        RECT 67.335 151.890 67.625 151.935 ;
        RECT 69.175 151.890 69.465 151.935 ;
        RECT 70.080 151.890 70.400 151.950 ;
        RECT 67.335 151.750 70.400 151.890 ;
        RECT 67.335 151.705 67.625 151.750 ;
        RECT 69.175 151.705 69.465 151.750 ;
        RECT 70.080 151.690 70.400 151.750 ;
        RECT 71.000 151.690 71.320 151.950 ;
        RECT 72.855 151.705 73.145 151.935 ;
        RECT 70.170 151.550 70.310 151.690 ;
        RECT 72.930 151.550 73.070 151.705 ;
        RECT 73.760 151.690 74.080 151.950 ;
        RECT 74.680 151.690 75.000 151.950 ;
        RECT 75.155 151.705 75.445 151.935 ;
        RECT 75.615 151.890 75.905 151.935 ;
        RECT 78.360 151.890 78.680 151.950 ;
        RECT 79.295 151.890 79.585 151.935 ;
        RECT 75.615 151.750 79.585 151.890 ;
        RECT 75.615 151.705 75.905 151.750 ;
        RECT 70.170 151.410 73.070 151.550 ;
        RECT 73.300 151.350 73.620 151.610 ;
        RECT 74.220 151.550 74.540 151.610 ;
        RECT 75.230 151.550 75.370 151.705 ;
        RECT 74.220 151.410 75.370 151.550 ;
        RECT 74.220 151.350 74.540 151.410 ;
        RECT 57.675 151.025 57.965 151.255 ;
        RECT 68.240 151.010 68.560 151.270 ;
        RECT 70.080 151.010 70.400 151.270 ;
        RECT 72.840 151.210 73.160 151.270 ;
        RECT 75.690 151.210 75.830 151.705 ;
        RECT 78.360 151.690 78.680 151.750 ;
        RECT 79.295 151.705 79.585 151.750 ;
        RECT 79.740 151.690 80.060 151.950 ;
        RECT 80.290 151.935 80.430 152.090 ;
        RECT 81.580 152.030 81.900 152.090 ;
        RECT 82.130 151.950 82.270 152.430 ;
        RECT 95.840 152.230 96.160 152.290 ;
        RECT 99.980 152.230 100.300 152.290 ;
        RECT 95.840 152.090 100.300 152.230 ;
        RECT 95.840 152.030 96.160 152.090 ;
        RECT 80.215 151.705 80.505 151.935 ;
        RECT 81.135 151.890 81.425 151.935 ;
        RECT 82.040 151.890 82.360 151.950 ;
        RECT 81.135 151.750 82.360 151.890 ;
        RECT 81.135 151.705 81.425 151.750 ;
        RECT 82.040 151.690 82.360 151.750 ;
        RECT 86.640 151.890 86.960 151.950 ;
        RECT 98.615 151.890 98.905 151.935 ;
        RECT 86.640 151.750 98.905 151.890 ;
        RECT 86.640 151.690 86.960 151.750 ;
        RECT 98.615 151.705 98.905 151.750 ;
        RECT 98.690 151.550 98.830 151.705 ;
        RECT 99.060 151.690 99.380 151.950 ;
        RECT 99.610 151.935 99.750 152.090 ;
        RECT 99.980 152.030 100.300 152.090 ;
        RECT 100.530 151.935 100.670 152.770 ;
        RECT 117.015 152.570 117.305 152.615 ;
        RECT 121.570 152.570 121.860 152.615 ;
        RECT 124.350 152.570 124.640 152.615 ;
        RECT 126.210 152.570 126.500 152.615 ;
        RECT 117.015 152.430 121.140 152.570 ;
        RECT 117.015 152.385 117.305 152.430 ;
        RECT 104.580 152.230 104.900 152.290 ;
        RECT 121.000 152.230 121.140 152.430 ;
        RECT 121.570 152.430 126.500 152.570 ;
        RECT 121.570 152.385 121.860 152.430 ;
        RECT 124.350 152.385 124.640 152.430 ;
        RECT 126.210 152.385 126.500 152.430 ;
        RECT 124.835 152.230 125.125 152.275 ;
        RECT 104.580 152.090 107.110 152.230 ;
        RECT 104.580 152.030 104.900 152.090 ;
        RECT 99.535 151.705 99.825 151.935 ;
        RECT 100.455 151.890 100.745 151.935 ;
        RECT 102.740 151.890 103.060 151.950 ;
        RECT 106.970 151.935 107.110 152.090 ;
        RECT 108.350 152.090 111.710 152.230 ;
        RECT 121.000 152.090 125.125 152.230 ;
        RECT 108.350 151.950 108.490 152.090 ;
        RECT 105.975 151.890 106.265 151.935 ;
        RECT 100.455 151.750 106.265 151.890 ;
        RECT 100.455 151.705 100.745 151.750 ;
        RECT 102.740 151.690 103.060 151.750 ;
        RECT 105.975 151.705 106.265 151.750 ;
        RECT 106.895 151.705 107.185 151.935 ;
        RECT 107.340 151.690 107.660 151.950 ;
        RECT 107.815 151.890 108.105 151.935 ;
        RECT 108.260 151.890 108.580 151.950 ;
        RECT 107.815 151.750 108.580 151.890 ;
        RECT 107.815 151.705 108.105 151.750 ;
        RECT 108.260 151.690 108.580 151.750 ;
        RECT 109.655 151.890 109.945 151.935 ;
        RECT 110.100 151.890 110.420 151.950 ;
        RECT 109.655 151.750 110.420 151.890 ;
        RECT 109.655 151.705 109.945 151.750 ;
        RECT 110.100 151.690 110.420 151.750 ;
        RECT 110.560 151.690 110.880 151.950 ;
        RECT 111.570 151.935 111.710 152.090 ;
        RECT 124.835 152.045 125.125 152.090 ;
        RECT 125.740 152.230 126.060 152.290 ;
        RECT 126.675 152.230 126.965 152.275 ;
        RECT 125.740 152.090 126.965 152.230 ;
        RECT 125.740 152.030 126.060 152.090 ;
        RECT 126.675 152.045 126.965 152.090 ;
        RECT 111.035 151.705 111.325 151.935 ;
        RECT 111.495 151.705 111.785 151.935 ;
        RECT 104.580 151.550 104.900 151.610 ;
        RECT 98.690 151.410 104.900 151.550 ;
        RECT 107.430 151.550 107.570 151.690 ;
        RECT 111.110 151.550 111.250 151.705 ;
        RECT 116.080 151.690 116.400 151.950 ;
        RECT 121.570 151.890 121.860 151.935 ;
        RECT 121.570 151.750 124.105 151.890 ;
        RECT 121.570 151.705 121.860 151.750 ;
        RECT 119.760 151.595 120.080 151.610 ;
        RECT 123.890 151.595 124.105 151.750 ;
        RECT 107.430 151.410 111.250 151.550 ;
        RECT 119.710 151.550 120.080 151.595 ;
        RECT 122.970 151.550 123.260 151.595 ;
        RECT 119.710 151.410 123.260 151.550 ;
        RECT 104.580 151.350 104.900 151.410 ;
        RECT 119.710 151.365 120.080 151.410 ;
        RECT 122.970 151.365 123.260 151.410 ;
        RECT 123.890 151.550 124.180 151.595 ;
        RECT 125.750 151.550 126.040 151.595 ;
        RECT 123.890 151.410 126.040 151.550 ;
        RECT 123.890 151.365 124.180 151.410 ;
        RECT 125.750 151.365 126.040 151.410 ;
        RECT 119.760 151.350 120.080 151.365 ;
        RECT 72.840 151.070 75.830 151.210 ;
        RECT 72.840 151.010 73.160 151.070 ;
        RECT 76.980 151.010 77.300 151.270 ;
        RECT 77.900 151.010 78.220 151.270 ;
        RECT 97.235 151.210 97.525 151.255 ;
        RECT 97.680 151.210 98.000 151.270 ;
        RECT 97.235 151.070 98.000 151.210 ;
        RECT 104.670 151.210 104.810 151.350 ;
        RECT 108.260 151.210 108.580 151.270 ;
        RECT 104.670 151.070 108.580 151.210 ;
        RECT 97.235 151.025 97.525 151.070 ;
        RECT 97.680 151.010 98.000 151.070 ;
        RECT 108.260 151.010 108.580 151.070 ;
        RECT 109.195 151.210 109.485 151.255 ;
        RECT 111.480 151.210 111.800 151.270 ;
        RECT 109.195 151.070 111.800 151.210 ;
        RECT 109.195 151.025 109.485 151.070 ;
        RECT 111.480 151.010 111.800 151.070 ;
        RECT 112.875 151.210 113.165 151.255 ;
        RECT 113.320 151.210 113.640 151.270 ;
        RECT 112.875 151.070 113.640 151.210 ;
        RECT 112.875 151.025 113.165 151.070 ;
        RECT 113.320 151.010 113.640 151.070 ;
        RECT 117.705 151.210 117.995 151.255 ;
        RECT 118.840 151.210 119.160 151.270 ;
        RECT 117.705 151.070 119.160 151.210 ;
        RECT 117.705 151.025 117.995 151.070 ;
        RECT 118.840 151.010 119.160 151.070 ;
        RECT 9.290 150.390 129.350 150.870 ;
        RECT 51.235 150.190 51.525 150.235 ;
        RECT 48.550 150.050 51.525 150.190 ;
        RECT 18.115 149.850 18.405 149.895 ;
        RECT 21.320 149.850 21.640 149.910 ;
        RECT 39.260 149.850 39.580 149.910 ;
        RECT 14.510 149.710 16.950 149.850 ;
        RECT 14.510 149.555 14.650 149.710 ;
        RECT 14.435 149.325 14.725 149.555 ;
        RECT 14.895 149.510 15.185 149.555 ;
        RECT 16.810 149.510 16.950 149.710 ;
        RECT 18.115 149.710 36.270 149.850 ;
        RECT 18.115 149.665 18.405 149.710 ;
        RECT 21.320 149.650 21.640 149.710 ;
        RECT 19.940 149.510 20.260 149.570 ;
        RECT 20.860 149.510 21.180 149.570 ;
        RECT 14.895 149.370 16.490 149.510 ;
        RECT 16.810 149.370 21.180 149.510 ;
        RECT 14.895 149.325 15.185 149.370 ;
        RECT 16.350 148.875 16.490 149.370 ;
        RECT 19.940 149.310 20.260 149.370 ;
        RECT 20.860 149.310 21.180 149.370 ;
        RECT 31.440 149.510 31.760 149.570 ;
        RECT 32.835 149.510 33.125 149.555 ;
        RECT 31.440 149.370 33.125 149.510 ;
        RECT 31.440 149.310 31.760 149.370 ;
        RECT 32.835 149.325 33.125 149.370 ;
        RECT 33.295 149.325 33.585 149.555 ;
        RECT 18.560 148.970 18.880 149.230 ;
        RECT 19.495 149.170 19.785 149.215 ;
        RECT 22.240 149.170 22.560 149.230 ;
        RECT 19.495 149.030 22.560 149.170 ;
        RECT 19.495 148.985 19.785 149.030 ;
        RECT 22.240 148.970 22.560 149.030 ;
        RECT 16.275 148.645 16.565 148.875 ;
        RECT 13.960 148.290 14.280 148.550 ;
        RECT 15.800 148.290 16.120 148.550 ;
        RECT 31.440 148.290 31.760 148.550 ;
        RECT 33.370 148.490 33.510 149.325 ;
        RECT 33.740 149.310 34.060 149.570 ;
        RECT 34.675 149.325 34.965 149.555 ;
        RECT 34.750 149.170 34.890 149.325 ;
        RECT 35.120 149.310 35.440 149.570 ;
        RECT 36.130 149.555 36.270 149.710 ;
        RECT 36.590 149.710 39.580 149.850 ;
        RECT 36.590 149.555 36.730 149.710 ;
        RECT 39.260 149.650 39.580 149.710 ;
        RECT 46.175 149.850 46.465 149.895 ;
        RECT 48.550 149.850 48.690 150.050 ;
        RECT 51.235 150.005 51.525 150.050 ;
        RECT 55.820 150.190 56.140 150.250 ;
        RECT 60.895 150.190 61.185 150.235 ;
        RECT 55.820 150.050 61.185 150.190 ;
        RECT 55.820 149.990 56.140 150.050 ;
        RECT 60.895 150.005 61.185 150.050 ;
        RECT 62.720 150.190 63.040 150.250 ;
        RECT 63.195 150.190 63.485 150.235 ;
        RECT 62.720 150.050 63.485 150.190 ;
        RECT 62.720 149.990 63.040 150.050 ;
        RECT 63.195 150.005 63.485 150.050 ;
        RECT 68.240 150.190 68.560 150.250 ;
        RECT 82.960 150.190 83.280 150.250 ;
        RECT 68.240 150.050 83.280 150.190 ;
        RECT 68.240 149.990 68.560 150.050 ;
        RECT 82.960 149.990 83.280 150.050 ;
        RECT 116.080 150.190 116.400 150.250 ;
        RECT 117.475 150.190 117.765 150.235 ;
        RECT 116.080 150.050 117.765 150.190 ;
        RECT 116.080 149.990 116.400 150.050 ;
        RECT 117.475 150.005 117.765 150.050 ;
        RECT 122.520 149.990 122.840 150.250 ;
        RECT 55.910 149.850 56.050 149.990 ;
        RECT 46.175 149.710 48.690 149.850 ;
        RECT 53.610 149.710 56.050 149.850 ;
        RECT 56.280 149.850 56.600 149.910 ;
        RECT 68.715 149.850 69.005 149.895 ;
        RECT 56.280 149.710 69.005 149.850 ;
        RECT 46.175 149.665 46.465 149.710 ;
        RECT 36.055 149.325 36.345 149.555 ;
        RECT 36.515 149.325 36.805 149.555 ;
        RECT 36.960 149.310 37.280 149.570 ;
        RECT 44.780 149.310 45.100 149.570 ;
        RECT 47.540 149.310 47.860 149.570 ;
        RECT 48.000 149.310 48.320 149.570 ;
        RECT 48.935 149.510 49.225 149.555 ;
        RECT 52.140 149.510 52.460 149.570 ;
        RECT 53.610 149.555 53.750 149.710 ;
        RECT 56.280 149.650 56.600 149.710 ;
        RECT 48.935 149.370 52.460 149.510 ;
        RECT 48.935 149.325 49.225 149.370 ;
        RECT 52.140 149.310 52.460 149.370 ;
        RECT 52.615 149.325 52.905 149.555 ;
        RECT 53.075 149.325 53.365 149.555 ;
        RECT 53.535 149.325 53.825 149.555 ;
        RECT 54.455 149.510 54.745 149.555 ;
        RECT 55.360 149.510 55.680 149.570 ;
        RECT 54.455 149.370 55.680 149.510 ;
        RECT 54.455 149.325 54.745 149.370 ;
        RECT 44.320 149.170 44.640 149.230 ;
        RECT 45.255 149.170 45.545 149.215 ;
        RECT 34.750 149.030 36.730 149.170 ;
        RECT 36.590 148.890 36.730 149.030 ;
        RECT 44.320 149.030 45.545 149.170 ;
        RECT 44.320 148.970 44.640 149.030 ;
        RECT 45.255 148.985 45.545 149.030 ;
        RECT 51.680 149.170 52.000 149.230 ;
        RECT 52.690 149.170 52.830 149.325 ;
        RECT 51.680 149.030 52.830 149.170 ;
        RECT 53.150 149.170 53.290 149.325 ;
        RECT 55.360 149.310 55.680 149.370 ;
        RECT 53.980 149.170 54.300 149.230 ;
        RECT 53.150 149.030 54.300 149.170 ;
        RECT 51.680 148.970 52.000 149.030 ;
        RECT 53.980 148.970 54.300 149.030 ;
        RECT 60.435 149.170 60.725 149.215 ;
        RECT 60.970 149.170 61.110 149.710 ;
        RECT 68.715 149.665 69.005 149.710 ;
        RECT 70.555 149.850 70.845 149.895 ;
        RECT 73.300 149.850 73.620 149.910 ;
        RECT 76.075 149.850 76.365 149.895 ;
        RECT 95.380 149.850 95.700 149.910 ;
        RECT 70.555 149.710 76.365 149.850 ;
        RECT 70.555 149.665 70.845 149.710 ;
        RECT 73.300 149.650 73.620 149.710 ;
        RECT 76.075 149.665 76.365 149.710 ;
        RECT 93.630 149.710 95.700 149.850 ;
        RECT 61.340 149.310 61.660 149.570 ;
        RECT 66.415 149.325 66.705 149.555 ;
        RECT 66.860 149.510 67.180 149.570 ;
        RECT 68.255 149.510 68.545 149.555 ;
        RECT 71.000 149.510 71.320 149.570 ;
        RECT 71.475 149.510 71.765 149.555 ;
        RECT 66.860 149.370 71.765 149.510 ;
        RECT 60.435 149.030 61.110 149.170 ;
        RECT 66.490 149.170 66.630 149.325 ;
        RECT 66.860 149.310 67.180 149.370 ;
        RECT 68.255 149.325 68.545 149.370 ;
        RECT 71.000 149.310 71.320 149.370 ;
        RECT 71.475 149.325 71.765 149.370 ;
        RECT 72.840 149.510 73.160 149.570 ;
        RECT 79.755 149.510 80.045 149.555 ;
        RECT 72.840 149.370 80.045 149.510 ;
        RECT 72.840 149.310 73.160 149.370 ;
        RECT 79.755 149.325 80.045 149.370 ;
        RECT 80.200 149.310 80.520 149.570 ;
        RECT 80.675 149.510 80.965 149.555 ;
        RECT 81.120 149.510 81.440 149.570 ;
        RECT 80.675 149.370 81.440 149.510 ;
        RECT 80.675 149.325 80.965 149.370 ;
        RECT 81.120 149.310 81.440 149.370 ;
        RECT 81.595 149.510 81.885 149.555 ;
        RECT 82.040 149.510 82.360 149.570 ;
        RECT 81.595 149.370 82.360 149.510 ;
        RECT 81.595 149.325 81.885 149.370 ;
        RECT 82.040 149.310 82.360 149.370 ;
        RECT 86.180 149.510 86.500 149.570 ;
        RECT 93.630 149.555 93.770 149.710 ;
        RECT 95.380 149.650 95.700 149.710 ;
        RECT 99.060 149.850 99.380 149.910 ;
        RECT 107.340 149.850 107.660 149.910 ;
        RECT 111.020 149.850 111.340 149.910 ;
        RECT 99.060 149.710 108.490 149.850 ;
        RECT 99.060 149.650 99.380 149.710 ;
        RECT 88.035 149.510 88.325 149.555 ;
        RECT 86.180 149.370 88.325 149.510 ;
        RECT 86.180 149.310 86.500 149.370 ;
        RECT 88.035 149.325 88.325 149.370 ;
        RECT 93.555 149.325 93.845 149.555 ;
        RECT 94.475 149.325 94.765 149.555 ;
        RECT 71.920 149.170 72.240 149.230 ;
        RECT 66.490 149.030 72.240 149.170 ;
        RECT 60.435 148.985 60.725 149.030 ;
        RECT 71.920 148.970 72.240 149.030 ;
        RECT 77.455 149.170 77.745 149.215 ;
        RECT 86.640 149.170 86.960 149.230 ;
        RECT 77.455 149.030 86.960 149.170 ;
        RECT 77.455 148.985 77.745 149.030 ;
        RECT 86.640 148.970 86.960 149.030 ;
        RECT 87.560 148.970 87.880 149.230 ;
        RECT 94.550 149.170 94.690 149.325 ;
        RECT 102.740 149.310 103.060 149.570 ;
        RECT 103.660 149.310 103.980 149.570 ;
        RECT 104.210 149.555 104.350 149.710 ;
        RECT 107.340 149.650 107.660 149.710 ;
        RECT 104.135 149.325 104.425 149.555 ;
        RECT 104.580 149.510 104.900 149.570 ;
        RECT 108.350 149.555 108.490 149.710 ;
        RECT 108.810 149.710 111.340 149.850 ;
        RECT 108.810 149.555 108.950 149.710 ;
        RECT 111.020 149.650 111.340 149.710 ;
        RECT 114.240 149.850 114.560 149.910 ;
        RECT 114.240 149.710 120.450 149.850 ;
        RECT 114.240 149.650 114.560 149.710 ;
        RECT 107.815 149.510 108.105 149.555 ;
        RECT 104.580 149.370 108.105 149.510 ;
        RECT 104.580 149.310 104.900 149.370 ;
        RECT 107.815 149.325 108.105 149.370 ;
        RECT 108.275 149.325 108.565 149.555 ;
        RECT 108.735 149.325 109.025 149.555 ;
        RECT 109.655 149.325 109.945 149.555 ;
        RECT 110.100 149.510 110.420 149.570 ;
        RECT 113.795 149.510 114.085 149.555 ;
        RECT 110.100 149.370 114.085 149.510 ;
        RECT 89.950 149.030 94.690 149.170 ;
        RECT 102.830 149.170 102.970 149.310 ;
        RECT 109.730 149.170 109.870 149.325 ;
        RECT 110.100 149.310 110.420 149.370 ;
        RECT 113.795 149.325 114.085 149.370 ;
        RECT 119.315 149.325 119.605 149.555 ;
        RECT 110.560 149.170 110.880 149.230 ;
        RECT 102.830 149.030 110.880 149.170 ;
        RECT 36.500 148.630 36.820 148.890 ;
        RECT 46.635 148.830 46.925 148.875 ;
        RECT 57.200 148.830 57.520 148.890 ;
        RECT 46.635 148.690 57.520 148.830 ;
        RECT 46.635 148.645 46.925 148.690 ;
        RECT 57.200 148.630 57.520 148.690 ;
        RECT 61.800 148.830 62.120 148.890 ;
        RECT 67.335 148.830 67.625 148.875 ;
        RECT 61.800 148.690 67.625 148.830 ;
        RECT 61.800 148.630 62.120 148.690 ;
        RECT 67.335 148.645 67.625 148.690 ;
        RECT 72.395 148.830 72.685 148.875 ;
        RECT 82.040 148.830 82.360 148.890 ;
        RECT 89.950 148.875 90.090 149.030 ;
        RECT 110.560 148.970 110.880 149.030 ;
        RECT 112.875 148.985 113.165 149.215 ;
        RECT 113.335 149.170 113.625 149.215 ;
        RECT 114.240 149.170 114.560 149.230 ;
        RECT 117.000 149.170 117.320 149.230 ;
        RECT 119.390 149.170 119.530 149.325 ;
        RECT 113.335 149.030 119.530 149.170 ;
        RECT 113.335 148.985 113.625 149.030 ;
        RECT 72.395 148.690 82.360 148.830 ;
        RECT 72.395 148.645 72.685 148.690 ;
        RECT 82.040 148.630 82.360 148.690 ;
        RECT 89.875 148.645 90.165 148.875 ;
        RECT 112.950 148.830 113.090 148.985 ;
        RECT 114.240 148.970 114.560 149.030 ;
        RECT 117.000 148.970 117.320 149.030 ;
        RECT 119.760 148.970 120.080 149.230 ;
        RECT 120.310 149.215 120.450 149.710 ;
        RECT 121.615 149.325 121.905 149.555 ;
        RECT 120.235 148.985 120.525 149.215 ;
        RECT 113.780 148.830 114.100 148.890 ;
        RECT 112.950 148.690 114.100 148.830 ;
        RECT 113.780 148.630 114.100 148.690 ;
        RECT 115.635 148.830 115.925 148.875 ;
        RECT 121.690 148.830 121.830 149.325 ;
        RECT 115.635 148.690 121.830 148.830 ;
        RECT 115.635 148.645 115.925 148.690 ;
        RECT 36.960 148.490 37.280 148.550 ;
        RECT 33.370 148.350 37.280 148.490 ;
        RECT 36.960 148.290 37.280 148.350 ;
        RECT 38.355 148.490 38.645 148.535 ;
        RECT 40.180 148.490 40.500 148.550 ;
        RECT 38.355 148.350 40.500 148.490 ;
        RECT 38.355 148.305 38.645 148.350 ;
        RECT 40.180 148.290 40.500 148.350 ;
        RECT 43.875 148.490 44.165 148.535 ;
        RECT 44.320 148.490 44.640 148.550 ;
        RECT 43.875 148.350 44.640 148.490 ;
        RECT 43.875 148.305 44.165 148.350 ;
        RECT 44.320 148.290 44.640 148.350 ;
        RECT 45.700 148.290 46.020 148.550 ;
        RECT 47.080 148.490 47.400 148.550 ;
        RECT 47.555 148.490 47.845 148.535 ;
        RECT 47.080 148.350 47.845 148.490 ;
        RECT 47.080 148.290 47.400 148.350 ;
        RECT 47.555 148.305 47.845 148.350 ;
        RECT 62.720 148.490 63.040 148.550 ;
        RECT 65.495 148.490 65.785 148.535 ;
        RECT 62.720 148.350 65.785 148.490 ;
        RECT 62.720 148.290 63.040 148.350 ;
        RECT 65.495 148.305 65.785 148.350 ;
        RECT 78.360 148.290 78.680 148.550 ;
        RECT 92.160 148.490 92.480 148.550 ;
        RECT 93.095 148.490 93.385 148.535 ;
        RECT 92.160 148.350 93.385 148.490 ;
        RECT 92.160 148.290 92.480 148.350 ;
        RECT 93.095 148.305 93.385 148.350 ;
        RECT 95.380 148.290 95.700 148.550 ;
        RECT 104.580 148.490 104.900 148.550 ;
        RECT 105.975 148.490 106.265 148.535 ;
        RECT 104.580 148.350 106.265 148.490 ;
        RECT 104.580 148.290 104.900 148.350 ;
        RECT 105.975 148.305 106.265 148.350 ;
        RECT 106.420 148.290 106.740 148.550 ;
        RECT 9.290 147.670 129.350 148.150 ;
        RECT 10.985 147.470 11.275 147.515 ;
        RECT 18.560 147.470 18.880 147.530 ;
        RECT 32.820 147.470 33.140 147.530 ;
        RECT 33.295 147.470 33.585 147.515 ;
        RECT 10.985 147.330 30.290 147.470 ;
        RECT 10.985 147.285 11.275 147.330 ;
        RECT 18.560 147.270 18.880 147.330 ;
        RECT 14.850 147.130 15.140 147.175 ;
        RECT 17.630 147.130 17.920 147.175 ;
        RECT 19.490 147.130 19.780 147.175 ;
        RECT 20.400 147.130 20.720 147.190 ;
        RECT 14.850 146.990 19.780 147.130 ;
        RECT 14.850 146.945 15.140 146.990 ;
        RECT 17.630 146.945 17.920 146.990 ;
        RECT 19.490 146.945 19.780 146.990 ;
        RECT 20.030 146.990 20.720 147.130 ;
        RECT 15.800 146.790 16.120 146.850 ;
        RECT 20.030 146.835 20.170 146.990 ;
        RECT 20.400 146.930 20.720 146.990 ;
        RECT 18.115 146.790 18.405 146.835 ;
        RECT 15.800 146.650 18.405 146.790 ;
        RECT 15.800 146.590 16.120 146.650 ;
        RECT 18.115 146.605 18.405 146.650 ;
        RECT 19.955 146.605 20.245 146.835 ;
        RECT 22.240 146.590 22.560 146.850 ;
        RECT 14.850 146.450 15.140 146.495 ;
        RECT 14.850 146.310 17.385 146.450 ;
        RECT 14.850 146.265 15.140 146.310 ;
        RECT 12.990 146.110 13.280 146.155 ;
        RECT 13.960 146.110 14.280 146.170 ;
        RECT 17.170 146.155 17.385 146.310 ;
        RECT 20.400 146.250 20.720 146.510 ;
        RECT 23.710 146.495 23.850 147.330 ;
        RECT 25.475 146.945 25.765 147.175 ;
        RECT 30.150 147.130 30.290 147.330 ;
        RECT 32.820 147.330 33.585 147.470 ;
        RECT 32.820 147.270 33.140 147.330 ;
        RECT 33.295 147.285 33.585 147.330 ;
        RECT 52.140 147.270 52.460 147.530 ;
        RECT 53.980 147.470 54.300 147.530 ;
        RECT 80.215 147.470 80.505 147.515 ;
        RECT 81.580 147.470 81.900 147.530 ;
        RECT 53.980 147.330 70.770 147.470 ;
        RECT 53.980 147.270 54.300 147.330 ;
        RECT 30.150 146.990 36.270 147.130 ;
        RECT 23.635 146.265 23.925 146.495 ;
        RECT 25.550 146.450 25.690 146.945 ;
        RECT 32.360 146.790 32.680 146.850 ;
        RECT 33.755 146.790 34.045 146.835 ;
        RECT 32.360 146.650 34.045 146.790 ;
        RECT 32.360 146.590 32.680 146.650 ;
        RECT 33.755 146.605 34.045 146.650 ;
        RECT 26.855 146.450 27.145 146.495 ;
        RECT 25.550 146.310 27.145 146.450 ;
        RECT 26.855 146.265 27.145 146.310 ;
        RECT 31.440 146.450 31.760 146.510 ;
        RECT 33.295 146.450 33.585 146.495 ;
        RECT 31.440 146.310 33.585 146.450 ;
        RECT 31.440 146.250 31.760 146.310 ;
        RECT 33.295 146.265 33.585 146.310 ;
        RECT 35.120 146.250 35.440 146.510 ;
        RECT 36.130 146.495 36.270 146.990 ;
        RECT 36.960 146.930 37.280 147.190 ;
        RECT 50.760 147.130 51.080 147.190 ;
        RECT 38.200 146.990 51.080 147.130 ;
        RECT 37.050 146.790 37.190 146.930 ;
        RECT 38.200 146.790 38.340 146.990 ;
        RECT 50.760 146.930 51.080 146.990 ;
        RECT 51.220 147.130 51.540 147.190 ;
        RECT 54.070 147.130 54.210 147.270 ;
        RECT 51.220 146.990 54.210 147.130 ;
        RECT 51.220 146.930 51.540 146.990 ;
        RECT 62.260 146.930 62.580 147.190 ;
        RECT 70.630 147.175 70.770 147.330 ;
        RECT 80.215 147.330 81.900 147.470 ;
        RECT 80.215 147.285 80.505 147.330 ;
        RECT 81.580 147.270 81.900 147.330 ;
        RECT 87.560 147.470 87.880 147.530 ;
        RECT 89.875 147.470 90.165 147.515 ;
        RECT 103.660 147.470 103.980 147.530 ;
        RECT 104.595 147.470 104.885 147.515 ;
        RECT 87.560 147.330 100.210 147.470 ;
        RECT 87.560 147.270 87.880 147.330 ;
        RECT 89.875 147.285 90.165 147.330 ;
        RECT 70.555 147.130 70.845 147.175 ;
        RECT 74.680 147.130 75.000 147.190 ;
        RECT 70.555 146.990 75.000 147.130 ;
        RECT 70.555 146.945 70.845 146.990 ;
        RECT 74.680 146.930 75.000 146.990 ;
        RECT 92.735 147.130 93.025 147.175 ;
        RECT 95.855 147.130 96.145 147.175 ;
        RECT 97.745 147.130 98.035 147.175 ;
        RECT 92.735 146.990 98.035 147.130 ;
        RECT 100.070 147.130 100.210 147.330 ;
        RECT 103.660 147.330 104.885 147.470 ;
        RECT 103.660 147.270 103.980 147.330 ;
        RECT 104.595 147.285 104.885 147.330 ;
        RECT 107.340 147.470 107.660 147.530 ;
        RECT 111.020 147.470 111.340 147.530 ;
        RECT 107.340 147.330 111.340 147.470 ;
        RECT 107.340 147.270 107.660 147.330 ;
        RECT 111.020 147.270 111.340 147.330 ;
        RECT 109.180 147.130 109.500 147.190 ;
        RECT 100.070 146.990 108.950 147.130 ;
        RECT 92.735 146.945 93.025 146.990 ;
        RECT 95.855 146.945 96.145 146.990 ;
        RECT 97.745 146.945 98.035 146.990 ;
        RECT 45.240 146.790 45.560 146.850 ;
        RECT 36.590 146.650 38.340 146.790 ;
        RECT 43.030 146.650 45.560 146.790 ;
        RECT 36.590 146.495 36.730 146.650 ;
        RECT 36.055 146.265 36.345 146.495 ;
        RECT 36.515 146.265 36.805 146.495 ;
        RECT 36.975 146.450 37.265 146.495 ;
        RECT 37.880 146.450 38.200 146.510 ;
        RECT 43.030 146.450 43.170 146.650 ;
        RECT 45.240 146.590 45.560 146.650 ;
        RECT 48.475 146.790 48.765 146.835 ;
        RECT 56.280 146.790 56.600 146.850 ;
        RECT 70.080 146.790 70.400 146.850 ;
        RECT 48.475 146.650 56.600 146.790 ;
        RECT 48.475 146.605 48.765 146.650 ;
        RECT 56.280 146.590 56.600 146.650 ;
        RECT 56.830 146.650 70.400 146.790 ;
        RECT 36.975 146.310 43.170 146.450 ;
        RECT 36.975 146.265 37.265 146.310 ;
        RECT 37.880 146.250 38.200 146.310 ;
        RECT 46.160 146.250 46.480 146.510 ;
        RECT 51.680 146.450 52.000 146.510 ;
        RECT 53.535 146.450 53.825 146.495 ;
        RECT 47.170 146.310 53.825 146.450 ;
        RECT 16.250 146.110 16.540 146.155 ;
        RECT 12.990 145.970 16.540 146.110 ;
        RECT 12.990 145.925 13.280 145.970 ;
        RECT 13.960 145.910 14.280 145.970 ;
        RECT 16.250 145.925 16.540 145.970 ;
        RECT 17.170 146.110 17.460 146.155 ;
        RECT 19.030 146.110 19.320 146.155 ;
        RECT 17.170 145.970 19.320 146.110 ;
        RECT 17.170 145.925 17.460 145.970 ;
        RECT 19.030 145.925 19.320 145.970 ;
        RECT 21.780 146.110 22.100 146.170 ;
        RECT 34.675 146.110 34.965 146.155 ;
        RECT 44.780 146.110 45.100 146.170 ;
        RECT 21.780 145.970 32.590 146.110 ;
        RECT 21.780 145.910 22.100 145.970 ;
        RECT 20.875 145.770 21.165 145.815 ;
        RECT 22.700 145.770 23.020 145.830 ;
        RECT 20.875 145.630 23.020 145.770 ;
        RECT 20.875 145.585 21.165 145.630 ;
        RECT 22.700 145.570 23.020 145.630 ;
        RECT 23.160 145.570 23.480 145.830 ;
        RECT 27.760 145.570 28.080 145.830 ;
        RECT 32.450 145.815 32.590 145.970 ;
        RECT 34.675 145.970 45.100 146.110 ;
        RECT 34.675 145.925 34.965 145.970 ;
        RECT 44.780 145.910 45.100 145.970 ;
        RECT 45.240 146.110 45.560 146.170 ;
        RECT 47.170 146.110 47.310 146.310 ;
        RECT 51.680 146.250 52.000 146.310 ;
        RECT 53.535 146.265 53.825 146.310 ;
        RECT 53.980 146.250 54.300 146.510 ;
        RECT 54.440 146.250 54.760 146.510 ;
        RECT 55.360 146.450 55.680 146.510 ;
        RECT 56.830 146.450 56.970 146.650 ;
        RECT 70.080 146.590 70.400 146.650 ;
        RECT 77.440 146.790 77.760 146.850 ;
        RECT 79.295 146.790 79.585 146.835 ;
        RECT 77.440 146.650 79.585 146.790 ;
        RECT 77.440 146.590 77.760 146.650 ;
        RECT 79.295 146.605 79.585 146.650 ;
        RECT 86.195 146.790 86.485 146.835 ;
        RECT 86.640 146.790 86.960 146.850 ;
        RECT 86.195 146.650 86.960 146.790 ;
        RECT 86.195 146.605 86.485 146.650 ;
        RECT 86.640 146.590 86.960 146.650 ;
        RECT 95.380 146.790 95.700 146.850 ;
        RECT 97.235 146.790 97.525 146.835 ;
        RECT 95.380 146.650 97.525 146.790 ;
        RECT 95.380 146.590 95.700 146.650 ;
        RECT 97.235 146.605 97.525 146.650 ;
        RECT 98.615 146.790 98.905 146.835 ;
        RECT 99.520 146.790 99.840 146.850 ;
        RECT 98.615 146.650 99.840 146.790 ;
        RECT 98.615 146.605 98.905 146.650 ;
        RECT 99.520 146.590 99.840 146.650 ;
        RECT 105.515 146.790 105.805 146.835 ;
        RECT 105.960 146.790 106.280 146.850 ;
        RECT 105.515 146.650 106.280 146.790 ;
        RECT 105.515 146.605 105.805 146.650 ;
        RECT 105.960 146.590 106.280 146.650 ;
        RECT 108.810 146.790 108.950 146.990 ;
        RECT 109.180 146.990 112.170 147.130 ;
        RECT 109.180 146.930 109.500 146.990 ;
        RECT 110.100 146.790 110.420 146.850 ;
        RECT 108.810 146.650 110.420 146.790 ;
        RECT 55.360 146.310 56.970 146.450 ;
        RECT 69.635 146.450 69.925 146.495 ;
        RECT 72.380 146.450 72.700 146.510 ;
        RECT 69.635 146.310 72.700 146.450 ;
        RECT 55.360 146.250 55.680 146.310 ;
        RECT 69.635 146.265 69.925 146.310 ;
        RECT 72.380 146.250 72.700 146.310 ;
        RECT 77.900 146.450 78.220 146.510 ;
        RECT 78.835 146.450 79.125 146.495 ;
        RECT 77.900 146.310 79.125 146.450 ;
        RECT 77.900 146.250 78.220 146.310 ;
        RECT 78.835 146.265 79.125 146.310 ;
        RECT 84.815 146.450 85.105 146.495 ;
        RECT 89.860 146.450 90.180 146.510 ;
        RECT 84.815 146.310 90.180 146.450 ;
        RECT 84.815 146.265 85.105 146.310 ;
        RECT 89.860 146.250 90.180 146.310 ;
        RECT 45.240 145.970 47.310 146.110 ;
        RECT 47.540 146.110 47.860 146.170 ;
        RECT 48.935 146.110 49.225 146.155 ;
        RECT 47.540 145.970 49.225 146.110 ;
        RECT 45.240 145.910 45.560 145.970 ;
        RECT 47.540 145.910 47.860 145.970 ;
        RECT 48.935 145.925 49.225 145.970 ;
        RECT 49.395 146.110 49.685 146.155 ;
        RECT 54.530 146.110 54.670 146.250 ;
        RECT 49.395 145.970 54.670 146.110 ;
        RECT 49.395 145.925 49.685 145.970 ;
        RECT 68.700 145.910 69.020 146.170 ;
        RECT 80.215 146.110 80.505 146.155 ;
        RECT 80.660 146.110 80.980 146.170 ;
        RECT 80.215 145.970 80.980 146.110 ;
        RECT 80.215 145.925 80.505 145.970 ;
        RECT 80.660 145.910 80.980 145.970 ;
        RECT 86.180 146.110 86.500 146.170 ;
        RECT 91.655 146.155 91.945 146.470 ;
        RECT 92.735 146.450 93.025 146.495 ;
        RECT 96.315 146.450 96.605 146.495 ;
        RECT 98.150 146.450 98.440 146.495 ;
        RECT 92.735 146.310 98.440 146.450 ;
        RECT 92.735 146.265 93.025 146.310 ;
        RECT 96.315 146.265 96.605 146.310 ;
        RECT 98.150 146.265 98.440 146.310 ;
        RECT 104.595 146.450 104.885 146.495 ;
        RECT 106.880 146.450 107.200 146.510 ;
        RECT 104.595 146.310 107.200 146.450 ;
        RECT 104.595 146.265 104.885 146.310 ;
        RECT 106.880 146.250 107.200 146.310 ;
        RECT 107.340 146.450 107.660 146.510 ;
        RECT 107.815 146.450 108.105 146.495 ;
        RECT 107.340 146.310 108.105 146.450 ;
        RECT 107.340 146.250 107.660 146.310 ;
        RECT 107.815 146.265 108.105 146.310 ;
        RECT 108.260 146.250 108.580 146.510 ;
        RECT 108.810 146.495 108.950 146.650 ;
        RECT 110.100 146.590 110.420 146.650 ;
        RECT 112.030 146.510 112.170 146.990 ;
        RECT 114.240 146.790 114.560 146.850 ;
        RECT 112.490 146.650 114.560 146.790 ;
        RECT 108.735 146.265 109.025 146.495 ;
        RECT 109.655 146.450 109.945 146.495 ;
        RECT 110.560 146.450 110.880 146.510 ;
        RECT 109.655 146.310 110.880 146.450 ;
        RECT 109.655 146.265 109.945 146.310 ;
        RECT 110.560 146.250 110.880 146.310 ;
        RECT 111.020 146.450 111.340 146.510 ;
        RECT 111.495 146.450 111.785 146.495 ;
        RECT 111.020 146.310 111.785 146.450 ;
        RECT 111.020 146.250 111.340 146.310 ;
        RECT 111.495 146.265 111.785 146.310 ;
        RECT 111.940 146.250 112.260 146.510 ;
        RECT 112.490 146.495 112.630 146.650 ;
        RECT 114.240 146.590 114.560 146.650 ;
        RECT 112.415 146.265 112.705 146.495 ;
        RECT 113.335 146.265 113.625 146.495 ;
        RECT 86.655 146.110 86.945 146.155 ;
        RECT 86.180 145.970 86.945 146.110 ;
        RECT 86.180 145.910 86.500 145.970 ;
        RECT 86.655 145.925 86.945 145.970 ;
        RECT 91.355 146.110 91.945 146.155 ;
        RECT 92.160 146.110 92.480 146.170 ;
        RECT 94.595 146.110 95.245 146.155 ;
        RECT 91.355 145.970 95.245 146.110 ;
        RECT 91.355 145.925 91.645 145.970 ;
        RECT 92.160 145.910 92.480 145.970 ;
        RECT 94.595 145.925 95.245 145.970 ;
        RECT 105.975 146.110 106.265 146.155 ;
        RECT 110.115 146.110 110.405 146.155 ;
        RECT 105.975 145.970 110.405 146.110 ;
        RECT 110.650 146.110 110.790 146.250 ;
        RECT 113.410 146.110 113.550 146.265 ;
        RECT 110.650 145.970 113.550 146.110 ;
        RECT 105.975 145.925 106.265 145.970 ;
        RECT 110.115 145.925 110.405 145.970 ;
        RECT 32.375 145.585 32.665 145.815 ;
        RECT 38.340 145.570 38.660 145.830 ;
        RECT 46.635 145.770 46.925 145.815 ;
        RECT 48.000 145.770 48.320 145.830 ;
        RECT 46.635 145.630 48.320 145.770 ;
        RECT 46.635 145.585 46.925 145.630 ;
        RECT 48.000 145.570 48.320 145.630 ;
        RECT 51.235 145.770 51.525 145.815 ;
        RECT 51.680 145.770 52.000 145.830 ;
        RECT 51.235 145.630 52.000 145.770 ;
        RECT 51.235 145.585 51.525 145.630 ;
        RECT 51.680 145.570 52.000 145.630 ;
        RECT 77.440 145.770 77.760 145.830 ;
        RECT 77.915 145.770 78.205 145.815 ;
        RECT 77.440 145.630 78.205 145.770 ;
        RECT 77.440 145.570 77.760 145.630 ;
        RECT 77.915 145.585 78.205 145.630 ;
        RECT 84.340 145.570 84.660 145.830 ;
        RECT 85.720 145.770 86.040 145.830 ;
        RECT 87.115 145.770 87.405 145.815 ;
        RECT 85.720 145.630 87.405 145.770 ;
        RECT 85.720 145.570 86.040 145.630 ;
        RECT 87.115 145.585 87.405 145.630 ;
        RECT 88.955 145.770 89.245 145.815 ;
        RECT 90.780 145.770 91.100 145.830 ;
        RECT 88.955 145.630 91.100 145.770 ;
        RECT 88.955 145.585 89.245 145.630 ;
        RECT 90.780 145.570 91.100 145.630 ;
        RECT 102.280 145.770 102.600 145.830 ;
        RECT 103.675 145.770 103.965 145.815 ;
        RECT 102.280 145.630 103.965 145.770 ;
        RECT 102.280 145.570 102.600 145.630 ;
        RECT 103.675 145.585 103.965 145.630 ;
        RECT 105.040 145.770 105.360 145.830 ;
        RECT 106.435 145.770 106.725 145.815 ;
        RECT 105.040 145.630 106.725 145.770 ;
        RECT 105.040 145.570 105.360 145.630 ;
        RECT 106.435 145.585 106.725 145.630 ;
        RECT 107.340 145.770 107.660 145.830 ;
        RECT 122.980 145.770 123.300 145.830 ;
        RECT 107.340 145.630 123.300 145.770 ;
        RECT 107.340 145.570 107.660 145.630 ;
        RECT 122.980 145.570 123.300 145.630 ;
        RECT 9.290 144.950 129.350 145.430 ;
        RECT 16.275 144.565 16.565 144.795 ;
        RECT 23.160 144.750 23.480 144.810 ;
        RECT 42.480 144.750 42.800 144.810 ;
        RECT 42.955 144.750 43.245 144.795 ;
        RECT 22.330 144.610 34.890 144.750 ;
        RECT 14.895 144.070 15.185 144.115 ;
        RECT 16.350 144.070 16.490 144.565 ;
        RECT 18.115 144.410 18.405 144.455 ;
        RECT 20.645 144.410 20.935 144.455 ;
        RECT 22.330 144.410 22.470 144.610 ;
        RECT 23.160 144.550 23.480 144.610 ;
        RECT 22.700 144.455 23.020 144.470 ;
        RECT 18.115 144.270 22.470 144.410 ;
        RECT 22.650 144.410 23.020 144.455 ;
        RECT 25.910 144.410 26.200 144.455 ;
        RECT 22.650 144.270 26.200 144.410 ;
        RECT 18.115 144.225 18.405 144.270 ;
        RECT 20.645 144.225 20.935 144.270 ;
        RECT 22.650 144.225 23.020 144.270 ;
        RECT 25.910 144.225 26.200 144.270 ;
        RECT 26.830 144.410 27.120 144.455 ;
        RECT 28.690 144.410 28.980 144.455 ;
        RECT 26.830 144.270 28.980 144.410 ;
        RECT 26.830 144.225 27.120 144.270 ;
        RECT 28.690 144.225 28.980 144.270 ;
        RECT 30.980 144.410 31.300 144.470 ;
        RECT 32.375 144.410 32.665 144.455 ;
        RECT 30.980 144.270 32.665 144.410 ;
        RECT 22.700 144.210 23.020 144.225 ;
        RECT 14.895 143.930 16.490 144.070 ;
        RECT 24.510 144.070 24.800 144.115 ;
        RECT 26.830 144.070 27.045 144.225 ;
        RECT 30.980 144.210 31.300 144.270 ;
        RECT 32.375 144.225 32.665 144.270 ;
        RECT 24.510 143.930 27.045 144.070 ;
        RECT 14.895 143.885 15.185 143.930 ;
        RECT 24.510 143.885 24.800 143.930 ;
        RECT 27.760 143.870 28.080 144.130 ;
        RECT 34.750 144.115 34.890 144.610 ;
        RECT 42.480 144.610 43.245 144.750 ;
        RECT 42.480 144.550 42.800 144.610 ;
        RECT 42.955 144.565 43.245 144.610 ;
        RECT 44.780 144.750 45.100 144.810 ;
        RECT 60.895 144.750 61.185 144.795 ;
        RECT 81.120 144.750 81.440 144.810 ;
        RECT 44.780 144.610 61.185 144.750 ;
        RECT 44.780 144.550 45.100 144.610 ;
        RECT 60.895 144.565 61.185 144.610 ;
        RECT 78.450 144.610 81.440 144.750 ;
        RECT 48.000 144.455 48.320 144.470 ;
        RECT 47.950 144.410 48.320 144.455 ;
        RECT 51.210 144.410 51.500 144.455 ;
        RECT 47.950 144.270 51.500 144.410 ;
        RECT 47.950 144.225 48.320 144.270 ;
        RECT 51.210 144.225 51.500 144.270 ;
        RECT 52.130 144.410 52.420 144.455 ;
        RECT 53.990 144.410 54.280 144.455 ;
        RECT 63.640 144.410 63.960 144.470 ;
        RECT 52.130 144.270 54.280 144.410 ;
        RECT 52.130 144.225 52.420 144.270 ;
        RECT 53.990 144.225 54.280 144.270 ;
        RECT 60.970 144.270 63.960 144.410 ;
        RECT 48.000 144.210 48.320 144.225 ;
        RECT 33.755 143.885 34.045 144.115 ;
        RECT 34.215 143.885 34.505 144.115 ;
        RECT 34.675 143.885 34.965 144.115 ;
        RECT 35.595 144.070 35.885 144.115 ;
        RECT 36.500 144.070 36.820 144.130 ;
        RECT 35.595 143.930 36.820 144.070 ;
        RECT 35.595 143.885 35.885 143.930 ;
        RECT 17.640 143.730 17.960 143.790 ;
        RECT 18.575 143.730 18.865 143.775 ;
        RECT 17.640 143.590 18.865 143.730 ;
        RECT 17.640 143.530 17.960 143.590 ;
        RECT 18.575 143.545 18.865 143.590 ;
        RECT 19.495 143.545 19.785 143.775 ;
        RECT 21.320 143.730 21.640 143.790 ;
        RECT 29.615 143.730 29.905 143.775 ;
        RECT 21.320 143.590 29.905 143.730 ;
        RECT 19.570 143.390 19.710 143.545 ;
        RECT 21.320 143.530 21.640 143.590 ;
        RECT 29.615 143.545 29.905 143.590 ;
        RECT 22.240 143.390 22.560 143.450 ;
        RECT 19.570 143.250 22.560 143.390 ;
        RECT 22.240 143.190 22.560 143.250 ;
        RECT 24.510 143.390 24.800 143.435 ;
        RECT 27.290 143.390 27.580 143.435 ;
        RECT 29.150 143.390 29.440 143.435 ;
        RECT 24.510 143.250 29.440 143.390 ;
        RECT 24.510 143.205 24.800 143.250 ;
        RECT 27.290 143.205 27.580 143.250 ;
        RECT 29.150 143.205 29.440 143.250 ;
        RECT 31.440 143.390 31.760 143.450 ;
        RECT 32.360 143.390 32.680 143.450 ;
        RECT 33.830 143.390 33.970 143.885 ;
        RECT 34.290 143.730 34.430 143.885 ;
        RECT 36.500 143.870 36.820 143.930 ;
        RECT 43.860 143.870 44.180 144.130 ;
        RECT 45.255 144.070 45.545 144.115 ;
        RECT 46.620 144.070 46.940 144.130 ;
        RECT 45.255 143.930 46.940 144.070 ;
        RECT 45.255 143.885 45.545 143.930 ;
        RECT 46.620 143.870 46.940 143.930 ;
        RECT 49.810 144.070 50.100 144.115 ;
        RECT 52.130 144.070 52.345 144.225 ;
        RECT 55.360 144.070 55.680 144.130 ;
        RECT 49.810 143.930 52.345 144.070 ;
        RECT 52.690 143.930 55.680 144.070 ;
        RECT 49.810 143.885 50.100 143.930 ;
        RECT 36.960 143.730 37.280 143.790 ;
        RECT 34.290 143.590 37.280 143.730 ;
        RECT 36.960 143.530 37.280 143.590 ;
        RECT 43.400 143.730 43.720 143.790 ;
        RECT 44.335 143.730 44.625 143.775 ;
        RECT 43.400 143.590 44.625 143.730 ;
        RECT 43.400 143.530 43.720 143.590 ;
        RECT 44.335 143.545 44.625 143.590 ;
        RECT 50.300 143.730 50.620 143.790 ;
        RECT 52.690 143.730 52.830 143.930 ;
        RECT 55.360 143.870 55.680 143.930 ;
        RECT 59.515 143.885 59.805 144.115 ;
        RECT 50.300 143.590 52.830 143.730 ;
        RECT 50.300 143.530 50.620 143.590 ;
        RECT 53.060 143.530 53.380 143.790 ;
        RECT 54.915 143.730 55.205 143.775 ;
        RECT 59.040 143.730 59.360 143.790 ;
        RECT 54.915 143.590 59.360 143.730 ;
        RECT 59.590 143.730 59.730 143.885 ;
        RECT 60.970 143.790 61.110 144.270 ;
        RECT 63.640 144.210 63.960 144.270 ;
        RECT 74.680 144.410 75.000 144.470 ;
        RECT 78.450 144.410 78.590 144.610 ;
        RECT 81.120 144.550 81.440 144.610 ;
        RECT 90.795 144.565 91.085 144.795 ;
        RECT 74.680 144.270 78.590 144.410 ;
        RECT 74.680 144.210 75.000 144.270 ;
        RECT 61.800 144.070 62.120 144.130 ;
        RECT 62.275 144.070 62.565 144.115 ;
        RECT 61.800 143.930 62.565 144.070 ;
        RECT 61.800 143.870 62.120 143.930 ;
        RECT 62.275 143.885 62.565 143.930 ;
        RECT 62.720 143.870 63.040 144.130 ;
        RECT 63.195 143.885 63.485 144.115 ;
        RECT 64.115 144.070 64.405 144.115 ;
        RECT 67.320 144.070 67.640 144.130 ;
        RECT 78.450 144.115 78.590 144.270 ;
        RECT 80.215 144.225 80.505 144.455 ;
        RECT 82.910 144.410 83.200 144.455 ;
        RECT 84.340 144.410 84.660 144.470 ;
        RECT 86.170 144.410 86.460 144.455 ;
        RECT 82.910 144.270 86.460 144.410 ;
        RECT 82.910 144.225 83.200 144.270 ;
        RECT 64.115 143.930 67.640 144.070 ;
        RECT 64.115 143.885 64.405 143.930 ;
        RECT 60.880 143.730 61.200 143.790 ;
        RECT 59.590 143.590 61.200 143.730 ;
        RECT 54.915 143.545 55.205 143.590 ;
        RECT 37.880 143.390 38.200 143.450 ;
        RECT 31.440 143.250 38.200 143.390 ;
        RECT 31.440 143.190 31.760 143.250 ;
        RECT 32.360 143.190 32.680 143.250 ;
        RECT 37.880 143.190 38.200 143.250 ;
        RECT 49.810 143.390 50.100 143.435 ;
        RECT 52.590 143.390 52.880 143.435 ;
        RECT 54.450 143.390 54.740 143.435 ;
        RECT 49.810 143.250 54.740 143.390 ;
        RECT 49.810 143.205 50.100 143.250 ;
        RECT 52.590 143.205 52.880 143.250 ;
        RECT 54.450 143.205 54.740 143.250 ;
        RECT 15.815 143.050 16.105 143.095 ;
        RECT 16.260 143.050 16.580 143.110 ;
        RECT 15.815 142.910 16.580 143.050 ;
        RECT 15.815 142.865 16.105 142.910 ;
        RECT 16.260 142.850 16.580 142.910 ;
        RECT 44.780 142.850 45.100 143.110 ;
        RECT 45.945 143.050 46.235 143.095 ;
        RECT 48.000 143.050 48.320 143.110 ;
        RECT 45.945 142.910 48.320 143.050 ;
        RECT 45.945 142.865 46.235 142.910 ;
        RECT 48.000 142.850 48.320 142.910 ;
        RECT 50.760 143.050 51.080 143.110 ;
        RECT 54.990 143.050 55.130 143.545 ;
        RECT 59.040 143.530 59.360 143.590 ;
        RECT 60.880 143.530 61.200 143.590 ;
        RECT 61.340 143.730 61.660 143.790 ;
        RECT 63.270 143.730 63.410 143.885 ;
        RECT 67.320 143.870 67.640 143.930 ;
        RECT 76.995 143.885 77.285 144.115 ;
        RECT 77.915 143.885 78.205 144.115 ;
        RECT 78.375 143.885 78.665 144.115 ;
        RECT 78.835 144.070 79.125 144.115 ;
        RECT 79.740 144.070 80.060 144.130 ;
        RECT 78.835 143.930 80.060 144.070 ;
        RECT 80.290 144.070 80.430 144.225 ;
        RECT 84.340 144.210 84.660 144.270 ;
        RECT 86.170 144.225 86.460 144.270 ;
        RECT 87.090 144.410 87.380 144.455 ;
        RECT 88.950 144.410 89.240 144.455 ;
        RECT 87.090 144.270 89.240 144.410 ;
        RECT 87.090 144.225 87.380 144.270 ;
        RECT 88.950 144.225 89.240 144.270 ;
        RECT 80.660 144.070 80.980 144.130 ;
        RECT 80.290 143.930 80.980 144.070 ;
        RECT 78.835 143.885 79.125 143.930 ;
        RECT 61.340 143.590 63.410 143.730 ;
        RECT 61.340 143.530 61.660 143.590 ;
        RECT 63.270 143.390 63.410 143.590 ;
        RECT 70.080 143.730 70.400 143.790 ;
        RECT 77.070 143.730 77.210 143.885 ;
        RECT 70.080 143.590 77.210 143.730 ;
        RECT 77.990 143.730 78.130 143.885 ;
        RECT 79.740 143.870 80.060 143.930 ;
        RECT 80.660 143.870 80.980 143.930 ;
        RECT 84.770 144.070 85.060 144.115 ;
        RECT 87.090 144.070 87.305 144.225 ;
        RECT 84.770 143.930 87.305 144.070 ;
        RECT 88.035 144.070 88.325 144.115 ;
        RECT 90.870 144.070 91.010 144.565 ;
        RECT 107.340 144.550 107.660 144.810 ;
        RECT 113.780 144.750 114.100 144.810 ;
        RECT 115.175 144.750 115.465 144.795 ;
        RECT 113.780 144.610 115.465 144.750 ;
        RECT 113.780 144.550 114.100 144.610 ;
        RECT 115.175 144.565 115.465 144.610 ;
        RECT 105.040 144.210 105.360 144.470 ;
        RECT 112.415 144.410 112.705 144.455 ;
        RECT 112.875 144.410 113.165 144.455 ;
        RECT 110.190 144.270 112.170 144.410 ;
        RECT 88.035 143.930 91.010 144.070 ;
        RECT 91.240 144.070 91.560 144.130 ;
        RECT 91.715 144.070 92.005 144.115 ;
        RECT 91.240 143.930 92.005 144.070 ;
        RECT 84.770 143.885 85.060 143.930 ;
        RECT 88.035 143.885 88.325 143.930 ;
        RECT 91.240 143.870 91.560 143.930 ;
        RECT 91.715 143.885 92.005 143.930 ;
        RECT 106.420 143.870 106.740 144.130 ;
        RECT 110.190 144.115 110.330 144.270 ;
        RECT 109.195 143.885 109.485 144.115 ;
        RECT 110.115 143.885 110.405 144.115 ;
        RECT 110.575 143.885 110.865 144.115 ;
        RECT 89.875 143.730 90.165 143.775 ;
        RECT 92.620 143.730 92.940 143.790 ;
        RECT 77.990 143.590 81.120 143.730 ;
        RECT 70.080 143.530 70.400 143.590 ;
        RECT 65.480 143.390 65.800 143.450 ;
        RECT 63.270 143.250 65.800 143.390 ;
        RECT 77.070 143.390 77.210 143.590 ;
        RECT 79.740 143.390 80.060 143.450 ;
        RECT 77.070 143.250 80.060 143.390 ;
        RECT 65.480 143.190 65.800 143.250 ;
        RECT 79.740 143.190 80.060 143.250 ;
        RECT 50.760 142.910 55.130 143.050 ;
        RECT 59.975 143.050 60.265 143.095 ;
        RECT 62.720 143.050 63.040 143.110 ;
        RECT 59.975 142.910 63.040 143.050 ;
        RECT 50.760 142.850 51.080 142.910 ;
        RECT 59.975 142.865 60.265 142.910 ;
        RECT 62.720 142.850 63.040 142.910 ;
        RECT 63.640 143.050 63.960 143.110 ;
        RECT 72.380 143.050 72.700 143.110 ;
        RECT 80.980 143.095 81.120 143.590 ;
        RECT 89.875 143.590 92.940 143.730 ;
        RECT 89.875 143.545 90.165 143.590 ;
        RECT 92.620 143.530 92.940 143.590 ;
        RECT 105.500 143.530 105.820 143.790 ;
        RECT 84.770 143.390 85.060 143.435 ;
        RECT 87.550 143.390 87.840 143.435 ;
        RECT 89.410 143.390 89.700 143.435 ;
        RECT 84.770 143.250 89.700 143.390 ;
        RECT 109.270 143.390 109.410 143.885 ;
        RECT 109.640 143.730 109.960 143.790 ;
        RECT 110.650 143.730 110.790 143.885 ;
        RECT 111.020 143.870 111.340 144.130 ;
        RECT 112.030 144.070 112.170 144.270 ;
        RECT 112.415 144.270 113.165 144.410 ;
        RECT 112.415 144.225 112.705 144.270 ;
        RECT 112.875 144.225 113.165 144.270 ;
        RECT 113.320 144.410 113.640 144.470 ;
        RECT 113.320 144.270 114.470 144.410 ;
        RECT 113.320 144.210 113.640 144.270 ;
        RECT 114.330 144.115 114.470 144.270 ;
        RECT 112.030 143.930 114.010 144.070 ;
        RECT 109.640 143.590 110.790 143.730 ;
        RECT 112.860 143.730 113.180 143.790 ;
        RECT 113.335 143.730 113.625 143.775 ;
        RECT 112.860 143.590 113.625 143.730 ;
        RECT 113.870 143.730 114.010 143.930 ;
        RECT 114.255 143.885 114.545 144.115 ;
        RECT 119.760 143.730 120.080 143.790 ;
        RECT 113.870 143.590 120.080 143.730 ;
        RECT 109.640 143.530 109.960 143.590 ;
        RECT 112.860 143.530 113.180 143.590 ;
        RECT 113.335 143.545 113.625 143.590 ;
        RECT 119.760 143.530 120.080 143.590 ;
        RECT 110.560 143.390 110.880 143.450 ;
        RECT 111.940 143.390 112.260 143.450 ;
        RECT 109.270 143.250 112.260 143.390 ;
        RECT 84.770 143.205 85.060 143.250 ;
        RECT 87.550 143.205 87.840 143.250 ;
        RECT 89.410 143.205 89.700 143.250 ;
        RECT 110.560 143.190 110.880 143.250 ;
        RECT 111.940 143.190 112.260 143.250 ;
        RECT 63.640 142.910 72.700 143.050 ;
        RECT 63.640 142.850 63.960 142.910 ;
        RECT 72.380 142.850 72.700 142.910 ;
        RECT 80.905 143.050 81.195 143.095 ;
        RECT 86.180 143.050 86.500 143.110 ;
        RECT 80.905 142.910 86.500 143.050 ;
        RECT 80.905 142.865 81.195 142.910 ;
        RECT 86.180 142.850 86.500 142.910 ;
        RECT 106.420 142.850 106.740 143.110 ;
        RECT 113.780 142.850 114.100 143.110 ;
        RECT 9.290 142.230 129.350 142.710 ;
        RECT 17.640 142.030 17.960 142.090 ;
        RECT 23.405 142.030 23.695 142.075 ;
        RECT 17.640 141.890 24.540 142.030 ;
        RECT 17.640 141.830 17.960 141.890 ;
        RECT 23.405 141.845 23.695 141.890 ;
        RECT 14.900 141.690 15.190 141.735 ;
        RECT 16.760 141.690 17.050 141.735 ;
        RECT 19.540 141.690 19.830 141.735 ;
        RECT 14.900 141.550 19.830 141.690 ;
        RECT 24.400 141.690 24.540 141.890 ;
        RECT 46.620 141.830 46.940 142.090 ;
        RECT 53.060 142.030 53.380 142.090 ;
        RECT 53.535 142.030 53.825 142.075 ;
        RECT 65.480 142.030 65.800 142.090 ;
        RECT 68.025 142.030 68.315 142.075 ;
        RECT 80.215 142.030 80.505 142.075 ;
        RECT 82.960 142.030 83.280 142.090 ;
        RECT 53.060 141.890 53.825 142.030 ;
        RECT 53.060 141.830 53.380 141.890 ;
        RECT 53.535 141.845 53.825 141.890 ;
        RECT 55.910 141.890 68.315 142.030 ;
        RECT 51.220 141.690 51.540 141.750 ;
        RECT 24.400 141.550 34.890 141.690 ;
        RECT 14.900 141.505 15.190 141.550 ;
        RECT 16.760 141.505 17.050 141.550 ;
        RECT 19.540 141.505 19.830 141.550 ;
        RECT 16.260 141.150 16.580 141.410 ;
        RECT 21.320 141.350 21.640 141.410 ;
        RECT 16.810 141.210 21.640 141.350 ;
        RECT 14.435 141.010 14.725 141.055 ;
        RECT 16.810 141.010 16.950 141.210 ;
        RECT 21.320 141.150 21.640 141.210 ;
        RECT 19.540 141.010 19.830 141.055 ;
        RECT 14.435 140.870 16.950 141.010 ;
        RECT 17.295 140.870 19.830 141.010 ;
        RECT 14.435 140.825 14.725 140.870 ;
        RECT 17.295 140.715 17.510 140.870 ;
        RECT 19.540 140.825 19.830 140.870 ;
        RECT 32.360 141.010 32.680 141.070 ;
        RECT 34.750 141.055 34.890 141.550 ;
        RECT 48.550 141.550 51.540 141.690 ;
        RECT 46.620 141.350 46.940 141.410 ;
        RECT 48.550 141.350 48.690 141.550 ;
        RECT 51.220 141.490 51.540 141.550 ;
        RECT 46.620 141.210 48.690 141.350 ;
        RECT 46.620 141.150 46.940 141.210 ;
        RECT 33.755 141.010 34.045 141.055 ;
        RECT 32.360 140.870 34.045 141.010 ;
        RECT 32.360 140.810 32.680 140.870 ;
        RECT 33.755 140.825 34.045 140.870 ;
        RECT 34.215 140.825 34.505 141.055 ;
        RECT 34.675 140.825 34.965 141.055 ;
        RECT 35.595 141.010 35.885 141.055 ;
        RECT 36.500 141.010 36.820 141.070 ;
        RECT 35.595 140.870 36.820 141.010 ;
        RECT 35.595 140.825 35.885 140.870 ;
        RECT 15.360 140.670 15.650 140.715 ;
        RECT 17.220 140.670 17.510 140.715 ;
        RECT 18.140 140.670 18.430 140.715 ;
        RECT 21.400 140.670 21.690 140.715 ;
        RECT 15.360 140.530 17.510 140.670 ;
        RECT 15.360 140.485 15.650 140.530 ;
        RECT 17.220 140.485 17.510 140.530 ;
        RECT 17.730 140.530 21.690 140.670 ;
        RECT 34.290 140.670 34.430 140.825 ;
        RECT 36.500 140.810 36.820 140.870 ;
        RECT 45.240 141.010 45.560 141.070 ;
        RECT 48.550 141.055 48.690 141.210 ;
        RECT 48.015 141.010 48.305 141.055 ;
        RECT 45.240 140.870 48.305 141.010 ;
        RECT 45.240 140.810 45.560 140.870 ;
        RECT 48.015 140.825 48.305 140.870 ;
        RECT 48.475 140.825 48.765 141.055 ;
        RECT 48.935 140.825 49.225 141.055 ;
        RECT 49.855 141.010 50.145 141.055 ;
        RECT 50.300 141.010 50.620 141.070 ;
        RECT 51.220 141.010 51.540 141.070 ;
        RECT 49.855 140.870 51.540 141.010 ;
        RECT 49.855 140.825 50.145 140.870 ;
        RECT 36.960 140.670 37.280 140.730 ;
        RECT 49.010 140.670 49.150 140.825 ;
        RECT 50.300 140.810 50.620 140.870 ;
        RECT 51.220 140.810 51.540 140.870 ;
        RECT 51.680 141.010 52.000 141.070 ;
        RECT 55.910 141.055 56.050 141.890 ;
        RECT 65.480 141.830 65.800 141.890 ;
        RECT 68.025 141.845 68.315 141.890 ;
        RECT 72.010 141.890 79.970 142.030 ;
        RECT 58.595 141.505 58.885 141.735 ;
        RECT 59.520 141.690 59.810 141.735 ;
        RECT 61.380 141.690 61.670 141.735 ;
        RECT 64.160 141.690 64.450 141.735 ;
        RECT 59.520 141.550 64.450 141.690 ;
        RECT 59.520 141.505 59.810 141.550 ;
        RECT 61.380 141.505 61.670 141.550 ;
        RECT 64.160 141.505 64.450 141.550 ;
        RECT 67.320 141.690 67.640 141.750 ;
        RECT 72.010 141.690 72.150 141.890 ;
        RECT 67.320 141.550 72.150 141.690 ;
        RECT 72.380 141.690 72.700 141.750 ;
        RECT 72.380 141.550 73.530 141.690 ;
        RECT 52.615 141.010 52.905 141.055 ;
        RECT 51.680 140.870 52.905 141.010 ;
        RECT 51.680 140.810 52.000 140.870 ;
        RECT 52.615 140.825 52.905 140.870 ;
        RECT 55.835 140.825 56.125 141.055 ;
        RECT 56.280 141.010 56.600 141.070 ;
        RECT 56.755 141.010 57.045 141.055 ;
        RECT 56.280 140.870 57.045 141.010 ;
        RECT 56.280 140.810 56.600 140.870 ;
        RECT 56.755 140.825 57.045 140.870 ;
        RECT 57.660 140.810 57.980 141.070 ;
        RECT 58.670 141.010 58.810 141.505 ;
        RECT 67.320 141.490 67.640 141.550 ;
        RECT 72.380 141.490 72.700 141.550 ;
        RECT 59.040 141.150 59.360 141.410 ;
        RECT 61.800 141.350 62.120 141.410 ;
        RECT 65.480 141.350 65.800 141.410 ;
        RECT 71.460 141.350 71.780 141.410 ;
        RECT 61.800 141.210 71.780 141.350 ;
        RECT 61.800 141.150 62.120 141.210 ;
        RECT 65.480 141.150 65.800 141.210 ;
        RECT 70.170 141.055 70.310 141.210 ;
        RECT 71.460 141.150 71.780 141.210 ;
        RECT 60.895 141.010 61.185 141.055 ;
        RECT 64.160 141.010 64.450 141.055 ;
        RECT 58.670 140.870 61.185 141.010 ;
        RECT 60.895 140.825 61.185 140.870 ;
        RECT 61.915 140.870 64.450 141.010 ;
        RECT 57.215 140.670 57.505 140.715 ;
        RECT 34.290 140.530 37.280 140.670 ;
        RECT 17.730 140.390 17.870 140.530 ;
        RECT 18.140 140.485 18.430 140.530 ;
        RECT 21.400 140.485 21.690 140.530 ;
        RECT 36.960 140.470 37.280 140.530 ;
        RECT 48.090 140.530 49.150 140.670 ;
        RECT 56.830 140.530 57.505 140.670 ;
        RECT 57.750 140.670 57.890 140.810 ;
        RECT 61.915 140.715 62.130 140.870 ;
        RECT 64.160 140.825 64.450 140.870 ;
        RECT 70.095 140.825 70.385 141.055 ;
        RECT 70.540 140.810 70.860 141.070 ;
        RECT 71.015 140.825 71.305 141.055 ;
        RECT 59.980 140.670 60.270 140.715 ;
        RECT 61.840 140.670 62.130 140.715 ;
        RECT 57.750 140.530 59.270 140.670 ;
        RECT 48.090 140.390 48.230 140.530 ;
        RECT 56.830 140.390 56.970 140.530 ;
        RECT 57.215 140.485 57.505 140.530 ;
        RECT 17.640 140.130 17.960 140.390 ;
        RECT 28.220 140.330 28.540 140.390 ;
        RECT 32.375 140.330 32.665 140.375 ;
        RECT 28.220 140.190 32.665 140.330 ;
        RECT 28.220 140.130 28.540 140.190 ;
        RECT 32.375 140.145 32.665 140.190 ;
        RECT 48.000 140.130 48.320 140.390 ;
        RECT 56.740 140.130 57.060 140.390 ;
        RECT 59.130 140.330 59.270 140.530 ;
        RECT 59.980 140.530 62.130 140.670 ;
        RECT 59.980 140.485 60.270 140.530 ;
        RECT 61.840 140.485 62.130 140.530 ;
        RECT 62.720 140.715 63.040 140.730 ;
        RECT 62.720 140.670 63.050 140.715 ;
        RECT 66.020 140.670 66.310 140.715 ;
        RECT 62.720 140.530 66.310 140.670 ;
        RECT 62.720 140.485 63.050 140.530 ;
        RECT 66.020 140.485 66.310 140.530 ;
        RECT 69.160 140.670 69.480 140.730 ;
        RECT 71.090 140.670 71.230 140.825 ;
        RECT 71.920 140.810 72.240 141.070 ;
        RECT 73.390 141.055 73.530 141.550 ;
        RECT 76.520 141.350 76.840 141.410 ;
        RECT 79.295 141.350 79.585 141.395 ;
        RECT 76.520 141.210 79.585 141.350 ;
        RECT 76.520 141.150 76.840 141.210 ;
        RECT 79.295 141.165 79.585 141.210 ;
        RECT 73.315 140.825 73.605 141.055 ;
        RECT 76.980 141.010 77.300 141.070 ;
        RECT 78.835 141.010 79.125 141.055 ;
        RECT 76.980 140.870 79.125 141.010 ;
        RECT 79.830 141.010 79.970 141.890 ;
        RECT 80.215 141.890 83.280 142.030 ;
        RECT 80.215 141.845 80.505 141.890 ;
        RECT 82.960 141.830 83.280 141.890 ;
        RECT 111.020 141.690 111.340 141.750 ;
        RECT 110.190 141.550 111.340 141.690 ;
        RECT 80.200 141.350 80.520 141.410 ;
        RECT 82.040 141.350 82.360 141.410 ;
        RECT 80.200 141.210 82.360 141.350 ;
        RECT 80.200 141.150 80.520 141.210 ;
        RECT 82.040 141.150 82.360 141.210 ;
        RECT 102.740 141.010 103.060 141.070 ;
        RECT 79.830 140.870 103.060 141.010 ;
        RECT 76.980 140.810 77.300 140.870 ;
        RECT 78.835 140.825 79.125 140.870 ;
        RECT 102.740 140.810 103.060 140.870 ;
        RECT 107.340 141.010 107.660 141.070 ;
        RECT 110.190 141.055 110.330 141.550 ;
        RECT 111.020 141.490 111.340 141.550 ;
        RECT 121.615 141.505 121.905 141.735 ;
        RECT 114.240 141.350 114.560 141.410 ;
        RECT 118.395 141.350 118.685 141.395 ;
        RECT 114.240 141.210 118.685 141.350 ;
        RECT 114.240 141.150 114.560 141.210 ;
        RECT 118.395 141.165 118.685 141.210 ;
        RECT 110.115 141.010 110.405 141.055 ;
        RECT 107.340 140.870 110.405 141.010 ;
        RECT 107.340 140.810 107.660 140.870 ;
        RECT 110.115 140.825 110.405 140.870 ;
        RECT 110.575 140.825 110.865 141.055 ;
        RECT 69.160 140.530 71.230 140.670 ;
        RECT 80.215 140.670 80.505 140.715 ;
        RECT 80.660 140.670 80.980 140.730 ;
        RECT 80.215 140.530 80.980 140.670 ;
        RECT 62.720 140.470 63.040 140.485 ;
        RECT 69.160 140.470 69.480 140.530 ;
        RECT 80.215 140.485 80.505 140.530 ;
        RECT 80.660 140.470 80.980 140.530 ;
        RECT 109.640 140.670 109.960 140.730 ;
        RECT 110.650 140.670 110.790 140.825 ;
        RECT 111.020 140.810 111.340 141.070 ;
        RECT 111.940 140.810 112.260 141.070 ;
        RECT 116.540 140.810 116.860 141.070 ;
        RECT 119.760 140.810 120.080 141.070 ;
        RECT 121.690 141.010 121.830 141.505 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 122.995 141.010 123.285 141.055 ;
        RECT 121.690 140.870 123.285 141.010 ;
        RECT 122.995 140.825 123.285 140.870 ;
        RECT 112.400 140.670 112.720 140.730 ;
        RECT 109.640 140.530 112.720 140.670 ;
        RECT 109.640 140.470 109.960 140.530 ;
        RECT 112.400 140.470 112.720 140.530 ;
        RECT 68.715 140.330 69.005 140.375 ;
        RECT 59.130 140.190 69.005 140.330 ;
        RECT 68.715 140.145 69.005 140.190 ;
        RECT 72.840 140.130 73.160 140.390 ;
        RECT 76.520 140.330 76.840 140.390 ;
        RECT 77.915 140.330 78.205 140.375 ;
        RECT 76.520 140.190 78.205 140.330 ;
        RECT 76.520 140.130 76.840 140.190 ;
        RECT 77.915 140.145 78.205 140.190 ;
        RECT 79.740 140.330 80.060 140.390 ;
        RECT 82.500 140.330 82.820 140.390 ;
        RECT 79.740 140.190 82.820 140.330 ;
        RECT 79.740 140.130 80.060 140.190 ;
        RECT 82.500 140.130 82.820 140.190 ;
        RECT 108.735 140.330 109.025 140.375 ;
        RECT 110.560 140.330 110.880 140.390 ;
        RECT 108.735 140.190 110.880 140.330 ;
        RECT 108.735 140.145 109.025 140.190 ;
        RECT 110.560 140.130 110.880 140.190 ;
        RECT 117.000 140.130 117.320 140.390 ;
        RECT 119.300 140.130 119.620 140.390 ;
        RECT 123.915 140.330 124.205 140.375 ;
        RECT 125.280 140.330 125.600 140.390 ;
        RECT 123.915 140.190 125.600 140.330 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 123.915 140.145 124.205 140.190 ;
        RECT 125.280 140.130 125.600 140.190 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 9.290 139.510 129.350 139.990 ;
        RECT 17.640 139.310 17.960 139.370 ;
        RECT 18.115 139.310 18.405 139.355 ;
        RECT 17.640 139.170 18.405 139.310 ;
        RECT 17.640 139.110 17.960 139.170 ;
        RECT 18.115 139.125 18.405 139.170 ;
        RECT 28.680 139.310 29.000 139.370 ;
        RECT 30.075 139.310 30.365 139.355 ;
        RECT 28.680 139.170 30.365 139.310 ;
        RECT 28.680 139.110 29.000 139.170 ;
        RECT 30.075 139.125 30.365 139.170 ;
        RECT 32.835 139.125 33.125 139.355 ;
        RECT 43.860 139.310 44.180 139.370 ;
        RECT 46.160 139.310 46.480 139.370 ;
        RECT 43.860 139.170 46.480 139.310 ;
        RECT 27.760 138.970 28.080 139.030 ;
        RECT 32.910 138.970 33.050 139.125 ;
        RECT 43.860 139.110 44.180 139.170 ;
        RECT 46.160 139.110 46.480 139.170 ;
        RECT 48.000 139.310 48.320 139.370 ;
        RECT 49.855 139.310 50.145 139.355 ;
        RECT 48.000 139.170 50.145 139.310 ;
        RECT 48.000 139.110 48.320 139.170 ;
        RECT 49.855 139.125 50.145 139.170 ;
        RECT 62.260 139.310 62.580 139.370 ;
        RECT 71.460 139.310 71.780 139.370 ;
        RECT 79.295 139.310 79.585 139.355 ;
        RECT 80.660 139.310 80.980 139.370 ;
        RECT 102.740 139.310 103.060 139.370 ;
        RECT 111.940 139.310 112.260 139.370 ;
        RECT 118.165 139.310 118.455 139.355 ;
        RECT 119.300 139.310 119.620 139.370 ;
        RECT 62.260 139.170 62.950 139.310 ;
        RECT 62.260 139.110 62.580 139.170 ;
        RECT 27.760 138.830 33.050 138.970 ;
        RECT 35.135 138.970 35.425 139.015 ;
        RECT 36.040 138.970 36.360 139.030 ;
        RECT 35.135 138.830 36.360 138.970 ;
        RECT 27.760 138.770 28.080 138.830 ;
        RECT 35.135 138.785 35.425 138.830 ;
        RECT 36.040 138.770 36.360 138.830 ;
        RECT 36.500 138.970 36.820 139.030 ;
        RECT 36.500 138.830 61.570 138.970 ;
        RECT 36.500 138.770 36.820 138.830 ;
        RECT 17.655 138.630 17.945 138.675 ;
        RECT 20.400 138.630 20.720 138.690 ;
        RECT 17.655 138.490 20.720 138.630 ;
        RECT 17.655 138.445 17.945 138.490 ;
        RECT 20.400 138.430 20.720 138.490 ;
        RECT 28.220 138.430 28.540 138.690 ;
        RECT 29.600 138.430 29.920 138.690 ;
        RECT 30.980 138.430 31.300 138.690 ;
        RECT 32.375 138.445 32.665 138.675 ;
        RECT 33.755 138.630 34.045 138.675 ;
        RECT 57.660 138.630 57.980 138.690 ;
        RECT 33.755 138.490 57.980 138.630 ;
        RECT 33.755 138.445 34.045 138.490 ;
        RECT 29.155 138.290 29.445 138.335 ;
        RECT 30.520 138.290 30.840 138.350 ;
        RECT 29.155 138.150 30.840 138.290 ;
        RECT 29.155 138.105 29.445 138.150 ;
        RECT 30.520 138.090 30.840 138.150 ;
        RECT 31.900 138.090 32.220 138.350 ;
        RECT 32.450 137.950 32.590 138.445 ;
        RECT 57.660 138.430 57.980 138.490 ;
        RECT 34.675 138.290 34.965 138.335 ;
        RECT 35.580 138.290 35.900 138.350 ;
        RECT 34.675 138.150 35.900 138.290 ;
        RECT 34.675 138.105 34.965 138.150 ;
        RECT 35.580 138.090 35.900 138.150 ;
        RECT 46.160 138.290 46.480 138.350 ;
        RECT 50.315 138.290 50.605 138.335 ;
        RECT 46.160 138.150 50.605 138.290 ;
        RECT 46.160 138.090 46.480 138.150 ;
        RECT 50.315 138.105 50.605 138.150 ;
        RECT 51.235 138.290 51.525 138.335 ;
        RECT 51.680 138.290 52.000 138.350 ;
        RECT 56.280 138.290 56.600 138.350 ;
        RECT 51.235 138.150 56.600 138.290 ;
        RECT 51.235 138.105 51.525 138.150 ;
        RECT 51.680 138.090 52.000 138.150 ;
        RECT 56.280 138.090 56.600 138.150 ;
        RECT 60.895 137.950 61.185 137.995 ;
        RECT 32.450 137.810 61.185 137.950 ;
        RECT 61.430 137.950 61.570 138.830 ;
        RECT 61.800 138.770 62.120 139.030 ;
        RECT 62.810 138.970 62.950 139.170 ;
        RECT 71.460 139.170 79.050 139.310 ;
        RECT 71.460 139.110 71.780 139.170 ;
        RECT 65.940 138.970 66.260 139.030 ;
        RECT 62.810 138.830 66.260 138.970 ;
        RECT 61.890 138.630 62.030 138.770 ;
        RECT 62.810 138.675 62.950 138.830 ;
        RECT 65.940 138.770 66.260 138.830 ;
        RECT 70.490 138.970 70.780 139.015 ;
        RECT 72.840 138.970 73.160 139.030 ;
        RECT 73.750 138.970 74.040 139.015 ;
        RECT 70.490 138.830 74.040 138.970 ;
        RECT 70.490 138.785 70.780 138.830 ;
        RECT 72.840 138.770 73.160 138.830 ;
        RECT 73.750 138.785 74.040 138.830 ;
        RECT 74.670 138.970 74.960 139.015 ;
        RECT 76.530 138.970 76.820 139.015 ;
        RECT 74.670 138.830 76.820 138.970 ;
        RECT 78.910 138.970 79.050 139.170 ;
        RECT 79.295 139.170 80.980 139.310 ;
        RECT 79.295 139.125 79.585 139.170 ;
        RECT 80.660 139.110 80.980 139.170 ;
        RECT 81.210 139.170 101.130 139.310 ;
        RECT 81.210 138.970 81.350 139.170 ;
        RECT 85.720 138.970 86.040 139.030 ;
        RECT 78.910 138.830 81.350 138.970 ;
        RECT 81.670 138.830 86.040 138.970 ;
        RECT 74.670 138.785 74.960 138.830 ;
        RECT 76.530 138.785 76.820 138.830 ;
        RECT 62.275 138.630 62.565 138.675 ;
        RECT 61.890 138.490 62.565 138.630 ;
        RECT 62.275 138.445 62.565 138.490 ;
        RECT 62.735 138.445 63.025 138.675 ;
        RECT 63.195 138.445 63.485 138.675 ;
        RECT 64.115 138.630 64.405 138.675 ;
        RECT 67.320 138.630 67.640 138.690 ;
        RECT 64.115 138.490 67.640 138.630 ;
        RECT 64.115 138.445 64.405 138.490 ;
        RECT 61.800 138.290 62.120 138.350 ;
        RECT 63.270 138.290 63.410 138.445 ;
        RECT 67.320 138.430 67.640 138.490 ;
        RECT 72.350 138.630 72.640 138.675 ;
        RECT 74.670 138.630 74.885 138.785 ;
        RECT 72.350 138.490 74.885 138.630 ;
        RECT 72.350 138.445 72.640 138.490 ;
        RECT 80.660 138.430 80.980 138.690 ;
        RECT 81.120 138.430 81.440 138.690 ;
        RECT 81.670 138.675 81.810 138.830 ;
        RECT 85.720 138.770 86.040 138.830 ;
        RECT 99.075 138.970 99.365 139.015 ;
        RECT 99.535 138.970 99.825 139.015 ;
        RECT 99.075 138.830 99.825 138.970 ;
        RECT 99.075 138.785 99.365 138.830 ;
        RECT 99.535 138.785 99.825 138.830 ;
        RECT 100.990 138.970 101.130 139.170 ;
        RECT 102.740 139.170 112.260 139.310 ;
        RECT 102.740 139.110 103.060 139.170 ;
        RECT 105.975 138.970 106.265 139.015 ;
        RECT 106.435 138.970 106.725 139.015 ;
        RECT 100.990 138.830 105.270 138.970 ;
        RECT 81.595 138.445 81.885 138.675 ;
        RECT 82.500 138.430 82.820 138.690 ;
        RECT 89.860 138.430 90.180 138.690 ;
        RECT 97.680 138.430 98.000 138.690 ;
        RECT 100.990 138.675 101.130 138.830 ;
        RECT 100.915 138.445 101.205 138.675 ;
        RECT 101.375 138.445 101.665 138.675 ;
        RECT 61.800 138.150 63.410 138.290 ;
        RECT 61.800 138.090 62.120 138.150 ;
        RECT 68.240 138.090 68.560 138.350 ;
        RECT 71.920 138.290 72.240 138.350 ;
        RECT 71.550 138.150 72.240 138.290 ;
        RECT 68.330 137.950 68.470 138.090 ;
        RECT 71.550 137.950 71.690 138.150 ;
        RECT 71.920 138.090 72.240 138.150 ;
        RECT 74.220 138.290 74.540 138.350 ;
        RECT 75.615 138.290 75.905 138.335 ;
        RECT 74.220 138.150 75.905 138.290 ;
        RECT 74.220 138.090 74.540 138.150 ;
        RECT 75.615 138.105 75.905 138.150 ;
        RECT 77.455 138.290 77.745 138.335 ;
        RECT 92.620 138.290 92.940 138.350 ;
        RECT 77.455 138.150 92.940 138.290 ;
        RECT 77.455 138.105 77.745 138.150 ;
        RECT 92.620 138.090 92.940 138.150 ;
        RECT 98.600 138.090 98.920 138.350 ;
        RECT 61.430 137.810 71.690 137.950 ;
        RECT 72.350 137.950 72.640 137.995 ;
        RECT 75.130 137.950 75.420 137.995 ;
        RECT 76.990 137.950 77.280 137.995 ;
        RECT 72.350 137.810 77.280 137.950 ;
        RECT 60.895 137.765 61.185 137.810 ;
        RECT 72.350 137.765 72.640 137.810 ;
        RECT 75.130 137.765 75.420 137.810 ;
        RECT 76.990 137.765 77.280 137.810 ;
        RECT 80.660 137.950 80.980 138.010 ;
        RECT 82.040 137.950 82.360 138.010 ;
        RECT 101.450 137.950 101.590 138.445 ;
        RECT 101.820 138.430 102.140 138.690 ;
        RECT 102.740 138.430 103.060 138.690 ;
        RECT 104.580 138.430 104.900 138.690 ;
        RECT 105.130 138.630 105.270 138.830 ;
        RECT 105.975 138.830 106.725 138.970 ;
        RECT 105.975 138.785 106.265 138.830 ;
        RECT 106.435 138.785 106.725 138.830 ;
        RECT 107.340 138.630 107.660 138.690 ;
        RECT 109.730 138.675 109.870 139.170 ;
        RECT 111.940 139.110 112.260 139.170 ;
        RECT 113.870 139.170 119.620 139.310 ;
        RECT 111.020 138.970 111.340 139.030 ;
        RECT 113.870 139.015 114.010 139.170 ;
        RECT 118.165 139.125 118.455 139.170 ;
        RECT 119.300 139.110 119.620 139.170 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 113.795 138.970 114.085 139.015 ;
        RECT 111.020 138.830 114.085 138.970 ;
        RECT 111.020 138.770 111.340 138.830 ;
        RECT 113.795 138.785 114.085 138.830 ;
        RECT 117.000 138.970 117.320 139.030 ;
        RECT 120.170 138.970 120.460 139.015 ;
        RECT 123.430 138.970 123.720 139.015 ;
        RECT 117.000 138.830 123.720 138.970 ;
        RECT 117.000 138.770 117.320 138.830 ;
        RECT 120.170 138.785 120.460 138.830 ;
        RECT 123.430 138.785 123.720 138.830 ;
        RECT 124.350 138.970 124.640 139.015 ;
        RECT 126.210 138.970 126.500 139.015 ;
        RECT 124.350 138.830 126.500 138.970 ;
        RECT 124.350 138.785 124.640 138.830 ;
        RECT 126.210 138.785 126.500 138.830 ;
        RECT 107.815 138.630 108.105 138.675 ;
        RECT 105.130 138.490 108.105 138.630 ;
        RECT 107.340 138.430 107.660 138.490 ;
        RECT 107.815 138.445 108.105 138.490 ;
        RECT 108.275 138.445 108.565 138.675 ;
        RECT 108.735 138.445 109.025 138.675 ;
        RECT 109.655 138.445 109.945 138.675 ;
        RECT 114.240 138.630 114.560 138.690 ;
        RECT 112.950 138.490 114.560 138.630 ;
        RECT 104.120 138.290 104.440 138.350 ;
        RECT 105.055 138.290 105.345 138.335 ;
        RECT 104.120 138.150 105.345 138.290 ;
        RECT 104.120 138.090 104.440 138.150 ;
        RECT 105.055 138.105 105.345 138.150 ;
        RECT 108.350 137.950 108.490 138.445 ;
        RECT 80.660 137.810 82.360 137.950 ;
        RECT 80.660 137.750 80.980 137.810 ;
        RECT 82.040 137.750 82.360 137.810 ;
        RECT 89.030 137.810 108.490 137.950 ;
        RECT 108.810 137.950 108.950 138.445 ;
        RECT 111.020 138.290 111.340 138.350 ;
        RECT 112.415 138.290 112.705 138.335 ;
        RECT 112.950 138.290 113.090 138.490 ;
        RECT 114.240 138.430 114.560 138.490 ;
        RECT 116.540 138.430 116.860 138.690 ;
        RECT 122.030 138.630 122.320 138.675 ;
        RECT 124.350 138.630 124.565 138.785 ;
        RECT 122.030 138.490 124.565 138.630 ;
        RECT 122.030 138.445 122.320 138.490 ;
        RECT 125.280 138.430 125.600 138.690 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 111.020 138.150 113.090 138.290 ;
        RECT 111.020 138.090 111.340 138.150 ;
        RECT 112.415 138.105 112.705 138.150 ;
        RECT 113.320 138.090 113.640 138.350 ;
        RECT 127.120 138.090 127.440 138.350 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 113.410 137.950 113.550 138.090 ;
        RECT 108.810 137.810 113.550 137.950 ;
        RECT 122.030 137.950 122.320 137.995 ;
        RECT 124.810 137.950 125.100 137.995 ;
        RECT 126.670 137.950 126.960 137.995 ;
        RECT 122.030 137.810 126.960 137.950 ;
        RECT 27.300 137.410 27.620 137.670 ;
        RECT 28.220 137.410 28.540 137.670 ;
        RECT 30.060 137.610 30.380 137.670 ;
        RECT 31.455 137.610 31.745 137.655 ;
        RECT 30.060 137.470 31.745 137.610 ;
        RECT 30.060 137.410 30.380 137.470 ;
        RECT 31.455 137.425 31.745 137.470 ;
        RECT 32.360 137.610 32.680 137.670 ;
        RECT 33.755 137.610 34.045 137.655 ;
        RECT 32.360 137.470 34.045 137.610 ;
        RECT 32.360 137.410 32.680 137.470 ;
        RECT 33.755 137.425 34.045 137.470 ;
        RECT 47.540 137.610 47.860 137.670 ;
        RECT 48.015 137.610 48.305 137.655 ;
        RECT 47.540 137.470 48.305 137.610 ;
        RECT 47.540 137.410 47.860 137.470 ;
        RECT 48.015 137.425 48.305 137.470 ;
        RECT 56.740 137.610 57.060 137.670 ;
        RECT 66.400 137.610 66.720 137.670 ;
        RECT 67.780 137.610 68.100 137.670 ;
        RECT 56.740 137.470 68.100 137.610 ;
        RECT 56.740 137.410 57.060 137.470 ;
        RECT 66.400 137.410 66.720 137.470 ;
        RECT 67.780 137.410 68.100 137.470 ;
        RECT 68.485 137.610 68.775 137.655 ;
        RECT 69.160 137.610 69.480 137.670 ;
        RECT 68.485 137.470 69.480 137.610 ;
        RECT 68.485 137.425 68.775 137.470 ;
        RECT 69.160 137.410 69.480 137.470 ;
        RECT 70.540 137.610 70.860 137.670 ;
        RECT 89.030 137.610 89.170 137.810 ;
        RECT 70.540 137.470 89.170 137.610 ;
        RECT 89.415 137.610 89.705 137.655 ;
        RECT 89.860 137.610 90.180 137.670 ;
        RECT 89.415 137.470 90.180 137.610 ;
        RECT 70.540 137.410 70.860 137.470 ;
        RECT 89.415 137.425 89.705 137.470 ;
        RECT 89.860 137.410 90.180 137.470 ;
        RECT 96.775 137.610 97.065 137.655 ;
        RECT 97.220 137.610 97.540 137.670 ;
        RECT 96.775 137.470 97.540 137.610 ;
        RECT 96.775 137.425 97.065 137.470 ;
        RECT 97.220 137.410 97.540 137.470 ;
        RECT 98.600 137.410 98.920 137.670 ;
        RECT 103.675 137.610 103.965 137.655 ;
        RECT 104.120 137.610 104.440 137.670 ;
        RECT 103.675 137.470 104.440 137.610 ;
        RECT 103.675 137.425 103.965 137.470 ;
        RECT 104.120 137.410 104.440 137.470 ;
        RECT 105.960 137.410 106.280 137.670 ;
        RECT 108.350 137.610 108.490 137.810 ;
        RECT 122.030 137.765 122.320 137.810 ;
        RECT 124.810 137.765 125.100 137.810 ;
        RECT 126.670 137.765 126.960 137.810 ;
        RECT 112.400 137.610 112.720 137.670 ;
        RECT 108.350 137.470 112.720 137.610 ;
        RECT 112.400 137.410 112.720 137.470 ;
        RECT 115.620 137.410 115.940 137.670 ;
        RECT 117.000 137.410 117.320 137.670 ;
        RECT 9.290 136.790 129.350 137.270 ;
        RECT 64.115 136.590 64.405 136.635 ;
        RECT 42.110 136.450 64.405 136.590 ;
        RECT 29.600 136.250 29.920 136.310 ;
        RECT 42.110 136.250 42.250 136.450 ;
        RECT 64.115 136.405 64.405 136.450 ;
        RECT 74.220 136.390 74.540 136.650 ;
        RECT 84.585 136.590 84.875 136.635 ;
        RECT 85.720 136.590 86.040 136.650 ;
        RECT 84.585 136.450 86.040 136.590 ;
        RECT 84.585 136.405 84.875 136.450 ;
        RECT 85.720 136.390 86.040 136.450 ;
        RECT 107.800 136.390 108.120 136.650 ;
        RECT 113.320 136.590 113.640 136.650 ;
        RECT 117.245 136.590 117.535 136.635 ;
        RECT 113.320 136.450 117.535 136.590 ;
        RECT 113.320 136.390 113.640 136.450 ;
        RECT 117.245 136.405 117.535 136.450 ;
        RECT 29.600 136.110 42.250 136.250 ;
        RECT 45.210 136.250 45.500 136.295 ;
        RECT 47.990 136.250 48.280 136.295 ;
        RECT 49.850 136.250 50.140 136.295 ;
        RECT 45.210 136.110 50.140 136.250 ;
        RECT 29.600 136.050 29.920 136.110 ;
        RECT 45.210 136.065 45.500 136.110 ;
        RECT 47.990 136.065 48.280 136.110 ;
        RECT 49.850 136.065 50.140 136.110 ;
        RECT 71.475 136.250 71.765 136.295 ;
        RECT 88.450 136.250 88.740 136.295 ;
        RECT 91.230 136.250 91.520 136.295 ;
        RECT 93.090 136.250 93.380 136.295 ;
        RECT 71.475 136.110 72.840 136.250 ;
        RECT 71.475 136.065 71.765 136.110 ;
        RECT 50.315 135.910 50.605 135.955 ;
        RECT 50.760 135.910 51.080 135.970 ;
        RECT 43.950 135.770 50.070 135.910 ;
        RECT 43.950 135.630 44.090 135.770 ;
        RECT 39.735 135.570 40.025 135.615 ;
        RECT 43.860 135.570 44.180 135.630 ;
        RECT 39.735 135.430 44.180 135.570 ;
        RECT 39.735 135.385 40.025 135.430 ;
        RECT 43.860 135.370 44.180 135.430 ;
        RECT 45.210 135.570 45.500 135.615 ;
        RECT 48.000 135.570 48.320 135.630 ;
        RECT 48.475 135.570 48.765 135.615 ;
        RECT 45.210 135.430 47.745 135.570 ;
        RECT 45.210 135.385 45.500 135.430 ;
        RECT 47.530 135.275 47.745 135.430 ;
        RECT 48.000 135.430 48.765 135.570 ;
        RECT 49.930 135.570 50.070 135.770 ;
        RECT 50.315 135.770 51.080 135.910 ;
        RECT 50.315 135.725 50.605 135.770 ;
        RECT 50.760 135.710 51.080 135.770 ;
        RECT 56.280 135.910 56.600 135.970 ;
        RECT 65.020 135.910 65.340 135.970 ;
        RECT 68.255 135.910 68.545 135.955 ;
        RECT 56.280 135.770 68.545 135.910 ;
        RECT 56.280 135.710 56.600 135.770 ;
        RECT 65.020 135.710 65.340 135.770 ;
        RECT 68.255 135.725 68.545 135.770 ;
        RECT 69.160 135.710 69.480 135.970 ;
        RECT 55.360 135.570 55.680 135.630 ;
        RECT 49.930 135.430 55.680 135.570 ;
        RECT 48.000 135.370 48.320 135.430 ;
        RECT 48.475 135.385 48.765 135.430 ;
        RECT 55.360 135.370 55.680 135.430 ;
        RECT 65.480 135.370 65.800 135.630 ;
        RECT 65.940 135.370 66.260 135.630 ;
        RECT 66.415 135.570 66.705 135.615 ;
        RECT 66.860 135.570 67.180 135.630 ;
        RECT 66.415 135.430 67.180 135.570 ;
        RECT 66.415 135.385 66.705 135.430 ;
        RECT 66.860 135.370 67.180 135.430 ;
        RECT 67.320 135.370 67.640 135.630 ;
        RECT 72.700 135.570 72.840 136.110 ;
        RECT 88.450 136.110 93.380 136.250 ;
        RECT 88.450 136.065 88.740 136.110 ;
        RECT 91.230 136.065 91.520 136.110 ;
        RECT 93.090 136.065 93.380 136.110 ;
        RECT 121.110 136.250 121.400 136.295 ;
        RECT 123.890 136.250 124.180 136.295 ;
        RECT 125.750 136.250 126.040 136.295 ;
        RECT 121.110 136.110 126.040 136.250 ;
        RECT 121.110 136.065 121.400 136.110 ;
        RECT 123.890 136.065 124.180 136.110 ;
        RECT 125.750 136.065 126.040 136.110 ;
        RECT 92.620 135.910 92.940 135.970 ;
        RECT 93.555 135.910 93.845 135.955 ;
        RECT 92.620 135.770 93.845 135.910 ;
        RECT 92.620 135.710 92.940 135.770 ;
        RECT 93.555 135.725 93.845 135.770 ;
        RECT 108.260 135.710 108.580 135.970 ;
        RECT 111.480 135.910 111.800 135.970 ;
        RECT 108.810 135.770 111.800 135.910 ;
        RECT 73.315 135.570 73.605 135.615 ;
        RECT 72.700 135.430 73.605 135.570 ;
        RECT 73.315 135.385 73.605 135.430 ;
        RECT 88.450 135.570 88.740 135.615 ;
        RECT 88.450 135.430 90.985 135.570 ;
        RECT 88.450 135.385 88.740 135.430 ;
        RECT 40.195 135.230 40.485 135.275 ;
        RECT 43.350 135.230 43.640 135.275 ;
        RECT 46.610 135.230 46.900 135.275 ;
        RECT 40.195 135.090 46.900 135.230 ;
        RECT 40.195 135.045 40.485 135.090 ;
        RECT 43.350 135.045 43.640 135.090 ;
        RECT 46.610 135.045 46.900 135.090 ;
        RECT 47.530 135.230 47.820 135.275 ;
        RECT 49.390 135.230 49.680 135.275 ;
        RECT 47.530 135.090 49.680 135.230 ;
        RECT 47.530 135.045 47.820 135.090 ;
        RECT 49.390 135.045 49.680 135.090 ;
        RECT 41.345 134.890 41.635 134.935 ;
        RECT 46.160 134.890 46.480 134.950 ;
        RECT 41.345 134.750 46.480 134.890 ;
        RECT 66.030 134.890 66.170 135.370 ;
        RECT 66.950 135.230 67.090 135.370 ;
        RECT 89.860 135.275 90.180 135.290 ;
        RECT 69.635 135.230 69.925 135.275 ;
        RECT 66.950 135.090 69.925 135.230 ;
        RECT 69.635 135.045 69.925 135.090 ;
        RECT 86.590 135.230 86.880 135.275 ;
        RECT 89.850 135.230 90.180 135.275 ;
        RECT 86.590 135.090 90.180 135.230 ;
        RECT 86.590 135.045 86.880 135.090 ;
        RECT 89.850 135.045 90.180 135.090 ;
        RECT 90.770 135.275 90.985 135.430 ;
        RECT 91.700 135.370 92.020 135.630 ;
        RECT 107.815 135.570 108.105 135.615 ;
        RECT 108.810 135.570 108.950 135.770 ;
        RECT 111.480 135.710 111.800 135.770 ;
        RECT 126.215 135.910 126.505 135.955 ;
        RECT 127.120 135.910 127.440 135.970 ;
        RECT 126.215 135.770 127.440 135.910 ;
        RECT 126.215 135.725 126.505 135.770 ;
        RECT 127.120 135.710 127.440 135.770 ;
        RECT 107.815 135.430 108.950 135.570 ;
        RECT 109.195 135.570 109.485 135.615 ;
        RECT 110.560 135.570 110.880 135.630 ;
        RECT 109.195 135.430 110.880 135.570 ;
        RECT 107.815 135.385 108.105 135.430 ;
        RECT 109.195 135.385 109.485 135.430 ;
        RECT 110.560 135.370 110.880 135.430 ;
        RECT 121.110 135.570 121.400 135.615 ;
        RECT 121.110 135.430 123.645 135.570 ;
        RECT 121.110 135.385 121.400 135.430 ;
        RECT 90.770 135.230 91.060 135.275 ;
        RECT 92.630 135.230 92.920 135.275 ;
        RECT 90.770 135.090 92.920 135.230 ;
        RECT 90.770 135.045 91.060 135.090 ;
        RECT 92.630 135.045 92.920 135.090 ;
        RECT 117.000 135.230 117.320 135.290 ;
        RECT 123.430 135.275 123.645 135.430 ;
        RECT 124.360 135.370 124.680 135.630 ;
        RECT 119.250 135.230 119.540 135.275 ;
        RECT 122.510 135.230 122.800 135.275 ;
        RECT 117.000 135.090 122.800 135.230 ;
        RECT 89.860 135.030 90.180 135.045 ;
        RECT 117.000 135.030 117.320 135.090 ;
        RECT 119.250 135.045 119.540 135.090 ;
        RECT 122.510 135.045 122.800 135.090 ;
        RECT 123.430 135.230 123.720 135.275 ;
        RECT 125.290 135.230 125.580 135.275 ;
        RECT 123.430 135.090 125.580 135.230 ;
        RECT 123.430 135.045 123.720 135.090 ;
        RECT 125.290 135.045 125.580 135.090 ;
        RECT 70.540 134.890 70.860 134.950 ;
        RECT 66.030 134.750 70.860 134.890 ;
        RECT 41.345 134.705 41.635 134.750 ;
        RECT 46.160 134.690 46.480 134.750 ;
        RECT 70.540 134.690 70.860 134.750 ;
        RECT 106.880 134.690 107.200 134.950 ;
        RECT 9.290 134.070 129.350 134.550 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 27.775 133.870 28.065 133.915 ;
        RECT 28.220 133.870 28.540 133.930 ;
        RECT 27.775 133.730 28.540 133.870 ;
        RECT 27.775 133.685 28.065 133.730 ;
        RECT 28.220 133.670 28.540 133.730 ;
        RECT 30.060 133.670 30.380 133.930 ;
        RECT 32.360 133.670 32.680 133.930 ;
        RECT 47.540 133.670 47.860 133.930 ;
        RECT 48.000 133.870 48.320 133.930 ;
        RECT 49.395 133.870 49.685 133.915 ;
        RECT 48.000 133.730 49.685 133.870 ;
        RECT 48.000 133.670 48.320 133.730 ;
        RECT 49.395 133.685 49.685 133.730 ;
        RECT 82.500 133.670 82.820 133.930 ;
        RECT 85.720 133.670 86.040 133.930 ;
        RECT 89.875 133.870 90.165 133.915 ;
        RECT 91.700 133.870 92.020 133.930 ;
        RECT 89.875 133.730 92.020 133.870 ;
        RECT 89.875 133.685 90.165 133.730 ;
        RECT 91.700 133.670 92.020 133.730 ;
        RECT 110.115 133.870 110.405 133.915 ;
        RECT 113.320 133.870 113.640 133.930 ;
        RECT 110.115 133.730 113.640 133.870 ;
        RECT 110.115 133.685 110.405 133.730 ;
        RECT 113.320 133.670 113.640 133.730 ;
        RECT 123.455 133.870 123.745 133.915 ;
        RECT 124.360 133.870 124.680 133.930 ;
        RECT 123.455 133.730 124.680 133.870 ;
        RECT 123.455 133.685 123.745 133.730 ;
        RECT 124.360 133.670 124.680 133.730 ;
        RECT 17.655 133.530 17.945 133.575 ;
        RECT 22.700 133.530 23.020 133.590 ;
        RECT 43.415 133.530 43.705 133.575 ;
        RECT 45.715 133.530 46.005 133.575 ;
        RECT 17.655 133.390 27.530 133.530 ;
        RECT 17.655 133.345 17.945 133.390 ;
        RECT 22.700 133.330 23.020 133.390 ;
        RECT 18.115 133.190 18.405 133.235 ;
        RECT 20.400 133.190 20.720 133.250 ;
        RECT 25.935 133.190 26.225 133.235 ;
        RECT 18.115 133.050 26.225 133.190 ;
        RECT 18.115 133.005 18.405 133.050 ;
        RECT 20.400 132.990 20.720 133.050 ;
        RECT 25.935 133.005 26.225 133.050 ;
        RECT 26.840 132.990 27.160 133.250 ;
        RECT 27.390 133.190 27.530 133.390 ;
        RECT 43.415 133.390 46.005 133.530 ;
        RECT 47.630 133.530 47.770 133.670 ;
        RECT 51.220 133.530 51.540 133.590 ;
        RECT 47.630 133.390 50.530 133.530 ;
        RECT 43.415 133.345 43.705 133.390 ;
        RECT 45.715 133.345 46.005 133.390 ;
        RECT 27.390 133.180 27.990 133.190 ;
        RECT 28.695 133.180 28.985 133.235 ;
        RECT 27.390 133.050 28.985 133.180 ;
        RECT 27.850 133.040 28.985 133.050 ;
        RECT 28.695 133.005 28.985 133.040 ;
        RECT 29.155 133.190 29.445 133.235 ;
        RECT 31.440 133.190 31.760 133.250 ;
        RECT 29.155 133.050 31.760 133.190 ;
        RECT 29.155 133.005 29.445 133.050 ;
        RECT 17.195 132.850 17.485 132.895 ;
        RECT 17.640 132.850 17.960 132.910 ;
        RECT 17.195 132.710 17.960 132.850 ;
        RECT 17.195 132.665 17.485 132.710 ;
        RECT 17.640 132.650 17.960 132.710 ;
        RECT 30.520 132.650 30.840 132.910 ;
        RECT 26.840 132.510 27.160 132.570 ;
        RECT 31.070 132.510 31.210 133.050 ;
        RECT 31.440 132.990 31.760 133.050 ;
        RECT 38.800 133.190 39.120 133.250 ;
        RECT 42.035 133.190 42.325 133.235 ;
        RECT 38.800 133.050 42.325 133.190 ;
        RECT 38.800 132.990 39.120 133.050 ;
        RECT 42.035 133.005 42.325 133.050 ;
        RECT 45.240 133.190 45.560 133.250 ;
        RECT 47.095 133.190 47.385 133.235 ;
        RECT 45.240 133.050 47.385 133.190 ;
        RECT 45.240 132.990 45.560 133.050 ;
        RECT 47.095 133.005 47.385 133.050 ;
        RECT 47.540 132.990 47.860 133.250 ;
        RECT 48.015 133.005 48.305 133.235 ;
        RECT 48.920 133.190 49.240 133.250 ;
        RECT 50.390 133.235 50.530 133.390 ;
        RECT 50.850 133.390 51.540 133.530 ;
        RECT 48.920 133.050 50.070 133.190 ;
        RECT 42.940 132.650 43.260 132.910 ;
        RECT 46.160 132.850 46.480 132.910 ;
        RECT 48.090 132.850 48.230 133.005 ;
        RECT 48.920 132.990 49.240 133.050 ;
        RECT 49.380 132.850 49.700 132.910 ;
        RECT 46.160 132.710 49.700 132.850 ;
        RECT 49.930 132.850 50.070 133.050 ;
        RECT 50.315 133.005 50.605 133.235 ;
        RECT 50.850 132.850 50.990 133.390 ;
        RECT 51.220 133.330 51.540 133.390 ;
        RECT 81.120 133.530 81.440 133.590 ;
        RECT 82.590 133.530 82.730 133.670 ;
        RECT 86.640 133.530 86.960 133.590 ;
        RECT 81.120 133.390 82.270 133.530 ;
        RECT 82.590 133.390 83.650 133.530 ;
        RECT 81.120 133.330 81.440 133.390 ;
        RECT 55.360 132.990 55.680 133.250 ;
        RECT 56.755 133.005 57.045 133.235 ;
        RECT 80.200 133.190 80.520 133.250 ;
        RECT 82.130 133.235 82.270 133.390 ;
        RECT 83.510 133.250 83.650 133.390 ;
        RECT 86.640 133.390 97.910 133.530 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 86.640 133.330 86.960 133.390 ;
        RECT 81.595 133.190 81.885 133.235 ;
        RECT 80.200 133.050 81.885 133.190 ;
        RECT 49.930 132.710 50.990 132.850 ;
        RECT 51.220 132.850 51.540 132.910 ;
        RECT 56.830 132.850 56.970 133.005 ;
        RECT 80.200 132.990 80.520 133.050 ;
        RECT 81.595 133.005 81.885 133.050 ;
        RECT 82.055 133.005 82.345 133.235 ;
        RECT 82.500 132.990 82.820 133.250 ;
        RECT 83.420 132.990 83.740 133.250 ;
        RECT 86.180 132.990 86.500 133.250 ;
        RECT 88.955 133.190 89.245 133.235 ;
        RECT 88.110 133.050 89.245 133.190 ;
        RECT 51.220 132.710 56.970 132.850 ;
        RECT 85.275 132.850 85.565 132.895 ;
        RECT 86.640 132.850 86.960 132.910 ;
        RECT 85.275 132.710 86.960 132.850 ;
        RECT 46.160 132.650 46.480 132.710 ;
        RECT 49.380 132.650 49.700 132.710 ;
        RECT 51.220 132.650 51.540 132.710 ;
        RECT 85.275 132.665 85.565 132.710 ;
        RECT 86.640 132.650 86.960 132.710 ;
        RECT 26.840 132.370 31.210 132.510 ;
        RECT 41.115 132.510 41.405 132.555 ;
        RECT 43.400 132.510 43.720 132.570 ;
        RECT 41.115 132.370 43.720 132.510 ;
        RECT 26.840 132.310 27.160 132.370 ;
        RECT 41.115 132.325 41.405 132.370 ;
        RECT 43.400 132.310 43.720 132.370 ;
        RECT 46.620 132.510 46.940 132.570 ;
        RECT 47.540 132.510 47.860 132.570 ;
        RECT 88.110 132.555 88.250 133.050 ;
        RECT 88.955 133.005 89.245 133.050 ;
        RECT 90.320 133.190 90.640 133.250 ;
        RECT 96.315 133.190 96.605 133.235 ;
        RECT 90.320 133.050 96.605 133.190 ;
        RECT 90.320 132.990 90.640 133.050 ;
        RECT 96.315 133.005 96.605 133.050 ;
        RECT 97.770 132.850 97.910 133.390 ;
        RECT 99.535 133.190 99.825 133.235 ;
        RECT 101.820 133.190 102.140 133.250 ;
        RECT 105.500 133.190 105.820 133.250 ;
        RECT 109.655 133.190 109.945 133.235 ;
        RECT 112.415 133.190 112.705 133.235 ;
        RECT 99.535 133.050 109.945 133.190 ;
        RECT 99.535 133.005 99.825 133.050 ;
        RECT 101.820 132.990 102.140 133.050 ;
        RECT 105.500 132.990 105.820 133.050 ;
        RECT 109.655 133.005 109.945 133.050 ;
        RECT 112.030 133.050 112.705 133.190 ;
        RECT 98.155 132.850 98.445 132.895 ;
        RECT 97.770 132.710 98.445 132.850 ;
        RECT 98.155 132.665 98.445 132.710 ;
        RECT 46.620 132.370 47.860 132.510 ;
        RECT 46.620 132.310 46.940 132.370 ;
        RECT 47.540 132.310 47.860 132.370 ;
        RECT 88.035 132.325 88.325 132.555 ;
        RECT 98.230 132.510 98.370 132.665 ;
        RECT 99.060 132.650 99.380 132.910 ;
        RECT 108.735 132.850 109.025 132.895 ;
        RECT 111.020 132.850 111.340 132.910 ;
        RECT 108.735 132.710 111.340 132.850 ;
        RECT 108.735 132.665 109.025 132.710 ;
        RECT 108.810 132.510 108.950 132.665 ;
        RECT 111.020 132.650 111.340 132.710 ;
        RECT 112.030 132.555 112.170 133.050 ;
        RECT 112.415 133.005 112.705 133.050 ;
        RECT 115.620 133.190 115.940 133.250 ;
        RECT 122.535 133.190 122.825 133.235 ;
        RECT 115.620 133.050 122.825 133.190 ;
        RECT 115.620 132.990 115.940 133.050 ;
        RECT 122.535 133.005 122.825 133.050 ;
        RECT 98.230 132.370 108.950 132.510 ;
        RECT 111.955 132.325 112.245 132.555 ;
        RECT 19.955 132.170 20.245 132.215 ;
        RECT 22.240 132.170 22.560 132.230 ;
        RECT 19.955 132.030 22.560 132.170 ;
        RECT 19.955 131.985 20.245 132.030 ;
        RECT 22.240 131.970 22.560 132.030 ;
        RECT 42.020 131.970 42.340 132.230 ;
        RECT 55.820 131.970 56.140 132.230 ;
        RECT 57.660 131.970 57.980 132.230 ;
        RECT 80.215 132.170 80.505 132.215 ;
        RECT 80.660 132.170 80.980 132.230 ;
        RECT 80.215 132.030 80.980 132.170 ;
        RECT 80.215 131.985 80.505 132.030 ;
        RECT 80.660 131.970 80.980 132.030 ;
        RECT 96.760 131.970 97.080 132.230 ;
        RECT 101.360 131.970 101.680 132.230 ;
        RECT 113.320 131.970 113.640 132.230 ;
        RECT 9.290 131.350 129.350 131.830 ;
        RECT 24.540 131.150 24.860 131.210 ;
        RECT 30.520 131.150 30.840 131.210 ;
        RECT 24.540 131.010 30.840 131.150 ;
        RECT 24.540 130.950 24.860 131.010 ;
        RECT 30.520 130.950 30.840 131.010 ;
        RECT 38.800 130.950 39.120 131.210 ;
        RECT 40.640 130.950 40.960 131.210 ;
        RECT 51.220 130.950 51.540 131.210 ;
        RECT 76.980 130.950 77.300 131.210 ;
        RECT 82.500 131.150 82.820 131.210 ;
        RECT 93.785 131.150 94.075 131.195 ;
        RECT 99.060 131.150 99.380 131.210 ;
        RECT 82.500 131.010 99.380 131.150 ;
        RECT 82.500 130.950 82.820 131.010 ;
        RECT 15.770 130.810 16.060 130.855 ;
        RECT 18.550 130.810 18.840 130.855 ;
        RECT 20.410 130.810 20.700 130.855 ;
        RECT 15.770 130.670 20.700 130.810 ;
        RECT 15.770 130.625 16.060 130.670 ;
        RECT 18.550 130.625 18.840 130.670 ;
        RECT 20.410 130.625 20.700 130.670 ;
        RECT 56.250 130.810 56.540 130.855 ;
        RECT 59.030 130.810 59.320 130.855 ;
        RECT 60.890 130.810 61.180 130.855 ;
        RECT 56.250 130.670 61.180 130.810 ;
        RECT 56.250 130.625 56.540 130.670 ;
        RECT 59.030 130.625 59.320 130.670 ;
        RECT 60.890 130.625 61.180 130.670 ;
        RECT 81.120 130.610 81.440 130.870 ;
        RECT 11.905 130.285 12.195 130.515 ;
        RECT 32.375 130.470 32.665 130.515 ;
        RECT 35.580 130.470 35.900 130.530 ;
        RECT 46.620 130.470 46.940 130.530 ;
        RECT 32.375 130.330 35.900 130.470 ;
        RECT 32.375 130.285 32.665 130.330 ;
        RECT 11.980 130.130 12.120 130.285 ;
        RECT 35.580 130.270 35.900 130.330 ;
        RECT 45.790 130.330 46.940 130.470 ;
        RECT 11.750 129.990 12.120 130.130 ;
        RECT 15.770 130.130 16.060 130.175 ;
        RECT 19.035 130.130 19.325 130.175 ;
        RECT 15.770 129.990 18.305 130.130 ;
        RECT 11.750 129.450 11.890 129.990 ;
        RECT 15.770 129.945 16.060 129.990 ;
        RECT 12.120 129.790 12.440 129.850 ;
        RECT 18.090 129.835 18.305 129.990 ;
        RECT 19.035 129.990 20.630 130.130 ;
        RECT 19.035 129.945 19.325 129.990 ;
        RECT 13.910 129.790 14.200 129.835 ;
        RECT 17.170 129.790 17.460 129.835 ;
        RECT 12.120 129.650 17.460 129.790 ;
        RECT 12.120 129.590 12.440 129.650 ;
        RECT 13.910 129.605 14.200 129.650 ;
        RECT 17.170 129.605 17.460 129.650 ;
        RECT 18.090 129.790 18.380 129.835 ;
        RECT 19.950 129.790 20.240 129.835 ;
        RECT 18.090 129.650 20.240 129.790 ;
        RECT 20.490 129.790 20.630 129.990 ;
        RECT 20.860 129.930 21.180 130.190 ;
        RECT 22.240 129.930 22.560 130.190 ;
        RECT 24.080 129.930 24.400 130.190 ;
        RECT 30.980 129.930 31.300 130.190 ;
        RECT 31.440 130.130 31.760 130.190 ;
        RECT 33.295 130.130 33.585 130.175 ;
        RECT 36.960 130.130 37.280 130.190 ;
        RECT 31.440 129.990 37.280 130.130 ;
        RECT 31.440 129.930 31.760 129.990 ;
        RECT 33.295 129.945 33.585 129.990 ;
        RECT 36.960 129.930 37.280 129.990 ;
        RECT 37.435 129.945 37.725 130.175 ;
        RECT 32.820 129.790 33.140 129.850 ;
        RECT 34.215 129.790 34.505 129.835 ;
        RECT 20.490 129.650 21.550 129.790 ;
        RECT 18.090 129.605 18.380 129.650 ;
        RECT 19.950 129.605 20.240 129.650 ;
        RECT 20.400 129.450 20.720 129.510 ;
        RECT 21.410 129.495 21.550 129.650 ;
        RECT 32.820 129.650 34.505 129.790 ;
        RECT 37.510 129.790 37.650 129.945 ;
        RECT 37.880 129.930 38.200 130.190 ;
        RECT 40.180 129.930 40.500 130.190 ;
        RECT 40.655 130.130 40.945 130.175 ;
        RECT 41.100 130.130 41.420 130.190 ;
        RECT 40.655 129.990 41.420 130.130 ;
        RECT 40.655 129.945 40.945 129.990 ;
        RECT 41.100 129.930 41.420 129.990 ;
        RECT 45.240 129.930 45.560 130.190 ;
        RECT 45.790 130.175 45.930 130.330 ;
        RECT 46.620 130.270 46.940 130.330 ;
        RECT 48.475 130.470 48.765 130.515 ;
        RECT 51.680 130.470 52.000 130.530 ;
        RECT 48.475 130.330 52.000 130.470 ;
        RECT 48.475 130.285 48.765 130.330 ;
        RECT 51.680 130.270 52.000 130.330 ;
        RECT 57.660 130.470 57.980 130.530 ;
        RECT 65.480 130.470 65.800 130.530 ;
        RECT 66.415 130.470 66.705 130.515 ;
        RECT 57.660 130.330 59.270 130.470 ;
        RECT 57.660 130.270 57.980 130.330 ;
        RECT 45.715 129.945 46.005 130.175 ;
        RECT 46.175 129.945 46.465 130.175 ;
        RECT 47.095 130.130 47.385 130.175 ;
        RECT 47.540 130.130 47.860 130.190 ;
        RECT 48.920 130.130 49.240 130.190 ;
        RECT 47.095 129.990 49.240 130.130 ;
        RECT 47.095 129.945 47.385 129.990 ;
        RECT 38.340 129.790 38.660 129.850 ;
        RECT 37.510 129.650 38.660 129.790 ;
        RECT 32.820 129.590 33.140 129.650 ;
        RECT 34.215 129.605 34.505 129.650 ;
        RECT 38.340 129.590 38.660 129.650 ;
        RECT 38.815 129.790 39.105 129.835 ;
        RECT 41.575 129.790 41.865 129.835 ;
        RECT 43.875 129.790 44.165 129.835 ;
        RECT 38.815 129.650 41.330 129.790 ;
        RECT 38.815 129.605 39.105 129.650 ;
        RECT 11.750 129.310 20.720 129.450 ;
        RECT 20.400 129.250 20.720 129.310 ;
        RECT 21.335 129.265 21.625 129.495 ;
        RECT 23.160 129.250 23.480 129.510 ;
        RECT 31.900 129.250 32.220 129.510 ;
        RECT 36.515 129.450 36.805 129.495 ;
        RECT 37.880 129.450 38.200 129.510 ;
        RECT 36.515 129.310 38.200 129.450 ;
        RECT 36.515 129.265 36.805 129.310 ;
        RECT 37.880 129.250 38.200 129.310 ;
        RECT 39.275 129.450 39.565 129.495 ;
        RECT 39.720 129.450 40.040 129.510 ;
        RECT 39.275 129.310 40.040 129.450 ;
        RECT 41.190 129.450 41.330 129.650 ;
        RECT 41.575 129.650 44.165 129.790 ;
        RECT 46.250 129.790 46.390 129.945 ;
        RECT 47.540 129.930 47.860 129.990 ;
        RECT 48.920 129.930 49.240 129.990 ;
        RECT 49.380 129.930 49.700 130.190 ;
        RECT 56.250 130.130 56.540 130.175 ;
        RECT 59.130 130.130 59.270 130.330 ;
        RECT 65.480 130.330 66.705 130.470 ;
        RECT 81.210 130.470 81.350 130.610 ;
        RECT 86.195 130.470 86.485 130.515 ;
        RECT 86.640 130.470 86.960 130.530 ;
        RECT 81.210 130.330 81.810 130.470 ;
        RECT 65.480 130.270 65.800 130.330 ;
        RECT 66.415 130.285 66.705 130.330 ;
        RECT 59.515 130.130 59.805 130.175 ;
        RECT 56.250 129.990 58.785 130.130 ;
        RECT 59.130 129.990 59.805 130.130 ;
        RECT 56.250 129.945 56.540 129.990 ;
        RECT 54.390 129.790 54.680 129.835 ;
        RECT 55.820 129.790 56.140 129.850 ;
        RECT 58.570 129.835 58.785 129.990 ;
        RECT 59.515 129.945 59.805 129.990 ;
        RECT 61.355 130.130 61.645 130.175 ;
        RECT 62.720 130.130 63.040 130.190 ;
        RECT 70.555 130.130 70.845 130.175 ;
        RECT 61.355 129.990 63.040 130.130 ;
        RECT 61.355 129.945 61.645 129.990 ;
        RECT 62.720 129.930 63.040 129.990 ;
        RECT 69.710 129.990 70.845 130.130 ;
        RECT 57.650 129.790 57.940 129.835 ;
        RECT 46.250 129.650 49.150 129.790 ;
        RECT 41.575 129.605 41.865 129.650 ;
        RECT 43.875 129.605 44.165 129.650 ;
        RECT 48.000 129.450 48.320 129.510 ;
        RECT 49.010 129.495 49.150 129.650 ;
        RECT 54.390 129.650 57.940 129.790 ;
        RECT 54.390 129.605 54.680 129.650 ;
        RECT 55.820 129.590 56.140 129.650 ;
        RECT 57.650 129.605 57.940 129.650 ;
        RECT 58.570 129.790 58.860 129.835 ;
        RECT 60.430 129.790 60.720 129.835 ;
        RECT 58.570 129.650 60.720 129.790 ;
        RECT 58.570 129.605 58.860 129.650 ;
        RECT 60.430 129.605 60.720 129.650 ;
        RECT 61.800 129.790 62.120 129.850 ;
        RECT 67.795 129.790 68.085 129.835 ;
        RECT 61.800 129.650 68.085 129.790 ;
        RECT 61.800 129.590 62.120 129.650 ;
        RECT 67.795 129.605 68.085 129.650 ;
        RECT 52.140 129.495 52.460 129.510 ;
        RECT 41.190 129.310 48.320 129.450 ;
        RECT 39.275 129.265 39.565 129.310 ;
        RECT 39.720 129.250 40.040 129.310 ;
        RECT 48.000 129.250 48.320 129.310 ;
        RECT 48.935 129.450 49.225 129.495 ;
        RECT 52.140 129.450 52.675 129.495 ;
        RECT 66.860 129.450 67.180 129.510 ;
        RECT 69.710 129.495 69.850 129.990 ;
        RECT 70.555 129.945 70.845 129.990 ;
        RECT 75.600 129.930 75.920 130.190 ;
        RECT 76.060 129.930 76.380 130.190 ;
        RECT 80.200 130.130 80.520 130.190 ;
        RECT 81.670 130.175 81.810 130.330 ;
        RECT 86.195 130.330 86.960 130.470 ;
        RECT 86.195 130.285 86.485 130.330 ;
        RECT 86.640 130.270 86.960 130.330 ;
        RECT 81.135 130.130 81.425 130.175 ;
        RECT 80.200 129.990 81.425 130.130 ;
        RECT 80.200 129.930 80.520 129.990 ;
        RECT 81.135 129.945 81.425 129.990 ;
        RECT 81.595 129.945 81.885 130.175 ;
        RECT 82.040 129.930 82.360 130.190 ;
        RECT 82.975 130.130 83.265 130.175 ;
        RECT 83.420 130.130 83.740 130.190 ;
        RECT 82.975 129.990 83.740 130.130 ;
        RECT 82.975 129.945 83.265 129.990 ;
        RECT 83.420 129.930 83.740 129.990 ;
        RECT 87.115 130.130 87.405 130.175 ;
        RECT 88.570 130.130 88.710 131.010 ;
        RECT 93.785 130.965 94.075 131.010 ;
        RECT 99.060 130.950 99.380 131.010 ;
        RECT 97.650 130.810 97.940 130.855 ;
        RECT 100.430 130.810 100.720 130.855 ;
        RECT 102.290 130.810 102.580 130.855 ;
        RECT 97.650 130.670 102.580 130.810 ;
        RECT 97.650 130.625 97.940 130.670 ;
        RECT 100.430 130.625 100.720 130.670 ;
        RECT 102.290 130.625 102.580 130.670 ;
        RECT 110.070 130.810 110.360 130.855 ;
        RECT 112.850 130.810 113.140 130.855 ;
        RECT 114.710 130.810 115.000 130.855 ;
        RECT 110.070 130.670 115.000 130.810 ;
        RECT 110.070 130.625 110.360 130.670 ;
        RECT 112.850 130.625 113.140 130.670 ;
        RECT 114.710 130.625 115.000 130.670 ;
        RECT 113.320 130.270 113.640 130.530 ;
        RECT 90.335 130.130 90.625 130.175 ;
        RECT 87.115 129.990 88.710 130.130 ;
        RECT 89.030 129.990 90.625 130.130 ;
        RECT 87.115 129.945 87.405 129.990 ;
        RECT 76.995 129.790 77.285 129.835 ;
        RECT 79.755 129.790 80.045 129.835 ;
        RECT 76.995 129.650 80.045 129.790 ;
        RECT 82.130 129.790 82.270 129.930 ;
        RECT 86.180 129.790 86.500 129.850 ;
        RECT 86.655 129.790 86.945 129.835 ;
        RECT 82.130 129.650 86.945 129.790 ;
        RECT 76.995 129.605 77.285 129.650 ;
        RECT 79.755 129.605 80.045 129.650 ;
        RECT 86.180 129.590 86.500 129.650 ;
        RECT 86.655 129.605 86.945 129.650 ;
        RECT 67.335 129.450 67.625 129.495 ;
        RECT 48.935 129.310 52.895 129.450 ;
        RECT 66.860 129.310 67.625 129.450 ;
        RECT 48.935 129.265 49.225 129.310 ;
        RECT 52.140 129.265 52.675 129.310 ;
        RECT 52.140 129.250 52.460 129.265 ;
        RECT 66.860 129.250 67.180 129.310 ;
        RECT 67.335 129.265 67.625 129.310 ;
        RECT 69.635 129.265 69.925 129.495 ;
        RECT 71.475 129.450 71.765 129.495 ;
        RECT 72.840 129.450 73.160 129.510 ;
        RECT 71.475 129.310 73.160 129.450 ;
        RECT 71.475 129.265 71.765 129.310 ;
        RECT 72.840 129.250 73.160 129.310 ;
        RECT 74.695 129.450 74.985 129.495 ;
        RECT 76.060 129.450 76.380 129.510 ;
        RECT 89.030 129.495 89.170 129.990 ;
        RECT 90.335 129.945 90.625 129.990 ;
        RECT 97.650 130.130 97.940 130.175 ;
        RECT 97.650 129.990 100.185 130.130 ;
        RECT 97.650 129.945 97.940 129.990 ;
        RECT 95.790 129.790 96.080 129.835 ;
        RECT 96.760 129.790 97.080 129.850 ;
        RECT 99.970 129.835 100.185 129.990 ;
        RECT 100.900 129.930 101.220 130.190 ;
        RECT 102.740 129.930 103.060 130.190 ;
        RECT 105.500 130.130 105.820 130.190 ;
        RECT 106.205 130.130 106.495 130.175 ;
        RECT 105.500 129.990 106.495 130.130 ;
        RECT 105.500 129.930 105.820 129.990 ;
        RECT 106.205 129.945 106.495 129.990 ;
        RECT 110.070 130.130 110.360 130.175 ;
        RECT 115.175 130.130 115.465 130.175 ;
        RECT 127.120 130.130 127.440 130.190 ;
        RECT 110.070 129.990 112.605 130.130 ;
        RECT 110.070 129.945 110.360 129.990 ;
        RECT 99.050 129.790 99.340 129.835 ;
        RECT 95.790 129.650 99.340 129.790 ;
        RECT 95.790 129.605 96.080 129.650 ;
        RECT 96.760 129.590 97.080 129.650 ;
        RECT 99.050 129.605 99.340 129.650 ;
        RECT 99.970 129.790 100.260 129.835 ;
        RECT 101.830 129.790 102.120 129.835 ;
        RECT 99.970 129.650 102.120 129.790 ;
        RECT 99.970 129.605 100.260 129.650 ;
        RECT 101.830 129.605 102.120 129.650 ;
        RECT 107.340 129.790 107.660 129.850 ;
        RECT 112.390 129.835 112.605 129.990 ;
        RECT 115.175 129.990 127.440 130.130 ;
        RECT 115.175 129.945 115.465 129.990 ;
        RECT 127.120 129.930 127.440 129.990 ;
        RECT 108.210 129.790 108.500 129.835 ;
        RECT 111.470 129.790 111.760 129.835 ;
        RECT 107.340 129.650 111.760 129.790 ;
        RECT 107.340 129.590 107.660 129.650 ;
        RECT 108.210 129.605 108.500 129.650 ;
        RECT 111.470 129.605 111.760 129.650 ;
        RECT 112.390 129.790 112.680 129.835 ;
        RECT 114.250 129.790 114.540 129.835 ;
        RECT 112.390 129.650 114.540 129.790 ;
        RECT 112.390 129.605 112.680 129.650 ;
        RECT 114.250 129.605 114.540 129.650 ;
        RECT 74.695 129.310 76.380 129.450 ;
        RECT 74.695 129.265 74.985 129.310 ;
        RECT 76.060 129.250 76.380 129.310 ;
        RECT 88.955 129.265 89.245 129.495 ;
        RECT 89.400 129.250 89.720 129.510 ;
        RECT 9.290 128.630 129.350 129.110 ;
        RECT 12.120 128.230 12.440 128.490 ;
        RECT 13.745 128.430 14.035 128.475 ;
        RECT 24.540 128.430 24.860 128.490 ;
        RECT 13.745 128.290 24.860 128.430 ;
        RECT 13.745 128.245 14.035 128.290 ;
        RECT 24.540 128.230 24.860 128.290 ;
        RECT 26.855 128.430 27.145 128.475 ;
        RECT 30.980 128.430 31.300 128.490 ;
        RECT 26.855 128.290 31.300 128.430 ;
        RECT 26.855 128.245 27.145 128.290 ;
        RECT 30.980 128.230 31.300 128.290 ;
        RECT 45.700 128.230 46.020 128.490 ;
        RECT 46.620 128.230 46.940 128.490 ;
        RECT 48.000 128.230 48.320 128.490 ;
        RECT 49.380 128.430 49.700 128.490 ;
        RECT 51.220 128.430 51.540 128.490 ;
        RECT 49.380 128.290 51.540 128.430 ;
        RECT 49.380 128.230 49.700 128.290 ;
        RECT 51.220 128.230 51.540 128.290 ;
        RECT 65.725 128.430 66.015 128.475 ;
        RECT 66.860 128.430 67.180 128.490 ;
        RECT 65.725 128.290 67.180 128.430 ;
        RECT 65.725 128.245 66.015 128.290 ;
        RECT 66.860 128.230 67.180 128.290 ;
        RECT 80.905 128.430 81.195 128.475 ;
        RECT 82.040 128.430 82.360 128.490 ;
        RECT 91.255 128.430 91.545 128.475 ;
        RECT 80.905 128.290 82.360 128.430 ;
        RECT 80.905 128.245 81.195 128.290 ;
        RECT 82.040 128.230 82.360 128.290 ;
        RECT 86.730 128.290 91.545 128.430 ;
        RECT 15.800 128.135 16.120 128.150 ;
        RECT 15.750 128.090 16.120 128.135 ;
        RECT 19.010 128.090 19.300 128.135 ;
        RECT 15.750 127.950 19.300 128.090 ;
        RECT 15.750 127.905 16.120 127.950 ;
        RECT 19.010 127.905 19.300 127.950 ;
        RECT 19.930 128.090 20.220 128.135 ;
        RECT 21.790 128.090 22.080 128.135 ;
        RECT 19.930 127.950 22.080 128.090 ;
        RECT 19.930 127.905 20.220 127.950 ;
        RECT 21.790 127.905 22.080 127.950 ;
        RECT 15.800 127.890 16.120 127.905 ;
        RECT 12.580 127.550 12.900 127.810 ;
        RECT 17.610 127.750 17.900 127.795 ;
        RECT 19.930 127.750 20.145 127.905 ;
        RECT 25.000 127.890 25.320 128.150 ;
        RECT 46.710 128.090 46.850 128.230 ;
        RECT 52.140 128.090 52.460 128.150 ;
        RECT 55.835 128.090 56.125 128.135 ;
        RECT 46.710 127.950 50.070 128.090 ;
        RECT 17.610 127.610 20.145 127.750 ;
        RECT 21.320 127.750 21.640 127.810 ;
        RECT 22.715 127.750 23.005 127.795 ;
        RECT 21.320 127.610 29.830 127.750 ;
        RECT 17.610 127.565 17.900 127.610 ;
        RECT 21.320 127.550 21.640 127.610 ;
        RECT 22.715 127.565 23.005 127.610 ;
        RECT 20.875 127.410 21.165 127.455 ;
        RECT 23.160 127.410 23.480 127.470 ;
        RECT 20.875 127.270 23.480 127.410 ;
        RECT 20.875 127.225 21.165 127.270 ;
        RECT 23.160 127.210 23.480 127.270 ;
        RECT 23.635 127.225 23.925 127.455 ;
        RECT 17.610 127.070 17.900 127.115 ;
        RECT 20.390 127.070 20.680 127.115 ;
        RECT 22.250 127.070 22.540 127.115 ;
        RECT 23.710 127.070 23.850 127.225 ;
        RECT 17.610 126.930 22.540 127.070 ;
        RECT 17.610 126.885 17.900 126.930 ;
        RECT 20.390 126.885 20.680 126.930 ;
        RECT 22.250 126.885 22.540 126.930 ;
        RECT 23.250 126.930 23.850 127.070 ;
        RECT 18.100 126.730 18.420 126.790 ;
        RECT 23.250 126.730 23.390 126.930 ;
        RECT 29.690 126.775 29.830 127.610 ;
        RECT 36.040 127.550 36.360 127.810 ;
        RECT 46.620 127.550 46.940 127.810 ;
        RECT 49.380 127.750 49.700 127.810 ;
        RECT 49.930 127.795 50.070 127.950 ;
        RECT 52.140 127.950 56.125 128.090 ;
        RECT 52.140 127.890 52.460 127.950 ;
        RECT 55.835 127.905 56.125 127.950 ;
        RECT 63.655 128.090 63.945 128.135 ;
        RECT 67.730 128.090 68.020 128.135 ;
        RECT 70.990 128.090 71.280 128.135 ;
        RECT 63.655 127.950 71.280 128.090 ;
        RECT 63.655 127.905 63.945 127.950 ;
        RECT 67.730 127.905 68.020 127.950 ;
        RECT 70.990 127.905 71.280 127.950 ;
        RECT 71.910 128.090 72.200 128.135 ;
        RECT 73.770 128.090 74.060 128.135 ;
        RECT 71.910 127.950 74.060 128.090 ;
        RECT 71.910 127.905 72.200 127.950 ;
        RECT 73.770 127.905 74.060 127.950 ;
        RECT 82.910 128.090 83.200 128.135 ;
        RECT 86.170 128.090 86.460 128.135 ;
        RECT 86.730 128.090 86.870 128.290 ;
        RECT 91.255 128.245 91.545 128.290 ;
        RECT 98.600 128.430 98.920 128.490 ;
        RECT 99.075 128.430 99.365 128.475 ;
        RECT 98.600 128.290 99.365 128.430 ;
        RECT 98.600 128.230 98.920 128.290 ;
        RECT 99.075 128.245 99.365 128.290 ;
        RECT 100.455 128.430 100.745 128.475 ;
        RECT 100.900 128.430 101.220 128.490 ;
        RECT 100.455 128.290 101.220 128.430 ;
        RECT 100.455 128.245 100.745 128.290 ;
        RECT 100.900 128.230 101.220 128.290 ;
        RECT 105.960 128.230 106.280 128.490 ;
        RECT 107.340 128.430 107.660 128.490 ;
        RECT 107.815 128.430 108.105 128.475 ;
        RECT 107.340 128.290 108.105 128.430 ;
        RECT 107.340 128.230 107.660 128.290 ;
        RECT 107.815 128.245 108.105 128.290 ;
        RECT 113.780 128.230 114.100 128.490 ;
        RECT 82.910 127.950 86.870 128.090 ;
        RECT 87.090 128.090 87.380 128.135 ;
        RECT 88.950 128.090 89.240 128.135 ;
        RECT 87.090 127.950 89.240 128.090 ;
        RECT 82.910 127.905 83.200 127.950 ;
        RECT 86.170 127.905 86.460 127.950 ;
        RECT 87.090 127.905 87.380 127.950 ;
        RECT 88.950 127.905 89.240 127.950 ;
        RECT 98.230 127.950 109.870 128.090 ;
        RECT 47.170 127.610 49.700 127.750 ;
        RECT 45.240 127.410 45.560 127.470 ;
        RECT 47.170 127.410 47.310 127.610 ;
        RECT 49.380 127.550 49.700 127.610 ;
        RECT 49.855 127.565 50.145 127.795 ;
        RECT 50.315 127.750 50.605 127.795 ;
        RECT 50.315 127.610 50.990 127.750 ;
        RECT 50.315 127.565 50.605 127.610 ;
        RECT 45.240 127.270 47.310 127.410 ;
        RECT 45.240 127.210 45.560 127.270 ;
        RECT 47.540 127.210 47.860 127.470 ;
        RECT 50.850 127.070 50.990 127.610 ;
        RECT 51.220 127.550 51.540 127.810 ;
        RECT 59.960 127.750 60.280 127.810 ;
        RECT 54.530 127.610 60.280 127.750 ;
        RECT 52.140 127.410 52.460 127.470 ;
        RECT 54.530 127.455 54.670 127.610 ;
        RECT 59.960 127.550 60.280 127.610 ;
        RECT 60.880 127.750 61.200 127.810 ;
        RECT 63.195 127.750 63.485 127.795 ;
        RECT 60.880 127.610 63.485 127.750 ;
        RECT 60.880 127.550 61.200 127.610 ;
        RECT 63.195 127.565 63.485 127.610 ;
        RECT 69.590 127.750 69.880 127.795 ;
        RECT 71.910 127.750 72.125 127.905 ;
        RECT 69.590 127.610 72.125 127.750 ;
        RECT 69.590 127.565 69.880 127.610 ;
        RECT 72.840 127.550 73.160 127.810 ;
        RECT 77.900 127.750 78.220 127.810 ;
        RECT 78.835 127.750 79.125 127.795 ;
        RECT 77.900 127.610 79.125 127.750 ;
        RECT 77.900 127.550 78.220 127.610 ;
        RECT 78.835 127.565 79.125 127.610 ;
        RECT 80.200 127.550 80.520 127.810 ;
        RECT 84.770 127.750 85.060 127.795 ;
        RECT 87.090 127.750 87.305 127.905 ;
        RECT 98.230 127.810 98.370 127.950 ;
        RECT 84.770 127.610 87.305 127.750 ;
        RECT 88.035 127.750 88.325 127.795 ;
        RECT 89.400 127.750 89.720 127.810 ;
        RECT 88.035 127.610 89.720 127.750 ;
        RECT 84.770 127.565 85.060 127.610 ;
        RECT 88.035 127.565 88.325 127.610 ;
        RECT 89.400 127.550 89.720 127.610 ;
        RECT 90.320 127.750 90.640 127.810 ;
        RECT 91.715 127.750 92.005 127.795 ;
        RECT 90.320 127.610 97.450 127.750 ;
        RECT 90.320 127.550 90.640 127.610 ;
        RECT 91.715 127.565 92.005 127.610 ;
        RECT 54.455 127.410 54.745 127.455 ;
        RECT 52.140 127.270 54.745 127.410 ;
        RECT 52.140 127.210 52.460 127.270 ;
        RECT 54.455 127.225 54.745 127.270 ;
        RECT 55.375 127.410 55.665 127.455 ;
        RECT 58.580 127.410 58.900 127.470 ;
        RECT 55.375 127.270 58.900 127.410 ;
        RECT 55.375 127.225 55.665 127.270 ;
        RECT 55.450 127.070 55.590 127.225 ;
        RECT 58.580 127.210 58.900 127.270 ;
        RECT 74.695 127.225 74.985 127.455 ;
        RECT 75.140 127.410 75.460 127.470 ;
        RECT 79.295 127.410 79.585 127.455 ;
        RECT 80.660 127.410 80.980 127.470 ;
        RECT 89.860 127.410 90.180 127.470 ;
        RECT 92.620 127.410 92.940 127.470 ;
        RECT 75.140 127.270 79.585 127.410 ;
        RECT 50.850 126.930 55.590 127.070 ;
        RECT 69.590 127.070 69.880 127.115 ;
        RECT 72.370 127.070 72.660 127.115 ;
        RECT 74.230 127.070 74.520 127.115 ;
        RECT 69.590 126.930 74.520 127.070 ;
        RECT 74.770 127.070 74.910 127.225 ;
        RECT 75.140 127.210 75.460 127.270 ;
        RECT 79.295 127.225 79.585 127.270 ;
        RECT 80.290 127.270 92.940 127.410 ;
        RECT 80.290 127.070 80.430 127.270 ;
        RECT 80.660 127.210 80.980 127.270 ;
        RECT 89.860 127.210 90.180 127.270 ;
        RECT 92.620 127.210 92.940 127.270 ;
        RECT 74.770 126.930 80.430 127.070 ;
        RECT 84.770 127.070 85.060 127.115 ;
        RECT 87.550 127.070 87.840 127.115 ;
        RECT 89.410 127.070 89.700 127.115 ;
        RECT 84.770 126.930 89.700 127.070 ;
        RECT 97.310 127.070 97.450 127.610 ;
        RECT 97.680 127.550 98.000 127.810 ;
        RECT 98.140 127.550 98.460 127.810 ;
        RECT 101.360 127.550 101.680 127.810 ;
        RECT 105.130 127.795 105.270 127.950 ;
        RECT 105.055 127.565 105.345 127.795 ;
        RECT 107.355 127.750 107.645 127.795 ;
        RECT 106.510 127.610 107.645 127.750 ;
        RECT 104.135 127.410 104.425 127.455 ;
        RECT 105.960 127.410 106.280 127.470 ;
        RECT 104.135 127.270 106.280 127.410 ;
        RECT 104.135 127.225 104.425 127.270 ;
        RECT 105.960 127.210 106.280 127.270 ;
        RECT 104.580 127.070 104.900 127.130 ;
        RECT 106.510 127.070 106.650 127.610 ;
        RECT 107.355 127.565 107.645 127.610 ;
        RECT 107.800 127.750 108.120 127.810 ;
        RECT 109.730 127.795 109.870 127.950 ;
        RECT 108.735 127.750 109.025 127.795 ;
        RECT 107.800 127.610 109.025 127.750 ;
        RECT 107.800 127.550 108.120 127.610 ;
        RECT 108.735 127.565 109.025 127.610 ;
        RECT 109.655 127.750 109.945 127.795 ;
        RECT 112.400 127.750 112.720 127.810 ;
        RECT 112.875 127.750 113.165 127.795 ;
        RECT 109.655 127.610 113.165 127.750 ;
        RECT 109.655 127.565 109.945 127.610 ;
        RECT 112.400 127.550 112.720 127.610 ;
        RECT 112.875 127.565 113.165 127.610 ;
        RECT 110.560 127.210 110.880 127.470 ;
        RECT 111.955 127.410 112.245 127.455 ;
        RECT 114.240 127.410 114.560 127.470 ;
        RECT 111.955 127.270 114.560 127.410 ;
        RECT 111.955 127.225 112.245 127.270 ;
        RECT 114.240 127.210 114.560 127.270 ;
        RECT 97.310 126.930 106.650 127.070 ;
        RECT 69.590 126.885 69.880 126.930 ;
        RECT 72.370 126.885 72.660 126.930 ;
        RECT 74.230 126.885 74.520 126.930 ;
        RECT 84.770 126.885 85.060 126.930 ;
        RECT 87.550 126.885 87.840 126.930 ;
        RECT 89.410 126.885 89.700 126.930 ;
        RECT 104.580 126.870 104.900 126.930 ;
        RECT 18.100 126.590 23.390 126.730 ;
        RECT 29.615 126.730 29.905 126.775 ;
        RECT 36.500 126.730 36.820 126.790 ;
        RECT 29.615 126.590 36.820 126.730 ;
        RECT 18.100 126.530 18.420 126.590 ;
        RECT 29.615 126.545 29.905 126.590 ;
        RECT 36.500 126.530 36.820 126.590 ;
        RECT 48.000 126.730 48.320 126.790 ;
        RECT 51.220 126.730 51.540 126.790 ;
        RECT 48.000 126.590 51.540 126.730 ;
        RECT 48.000 126.530 48.320 126.590 ;
        RECT 51.220 126.530 51.540 126.590 ;
        RECT 57.660 126.530 57.980 126.790 ;
        RECT 75.600 126.730 75.920 126.790 ;
        RECT 77.915 126.730 78.205 126.775 ;
        RECT 75.600 126.590 78.205 126.730 ;
        RECT 75.600 126.530 75.920 126.590 ;
        RECT 77.915 126.545 78.205 126.590 ;
        RECT 80.215 126.730 80.505 126.775 ;
        RECT 81.120 126.730 81.440 126.790 ;
        RECT 80.215 126.590 81.440 126.730 ;
        RECT 80.215 126.545 80.505 126.590 ;
        RECT 81.120 126.530 81.440 126.590 ;
        RECT 9.290 125.910 129.350 126.390 ;
        RECT 15.800 125.510 16.120 125.770 ;
        RECT 20.415 125.710 20.705 125.755 ;
        RECT 24.080 125.710 24.400 125.770 ;
        RECT 20.415 125.570 24.400 125.710 ;
        RECT 20.415 125.525 20.705 125.570 ;
        RECT 24.080 125.510 24.400 125.570 ;
        RECT 25.000 125.710 25.320 125.770 ;
        RECT 26.625 125.710 26.915 125.755 ;
        RECT 35.580 125.710 35.900 125.770 ;
        RECT 25.000 125.570 35.900 125.710 ;
        RECT 25.000 125.510 25.320 125.570 ;
        RECT 26.625 125.525 26.915 125.570 ;
        RECT 35.580 125.510 35.900 125.570 ;
        RECT 46.620 125.710 46.940 125.770 ;
        RECT 65.020 125.710 65.340 125.770 ;
        RECT 46.620 125.570 65.340 125.710 ;
        RECT 46.620 125.510 46.940 125.570 ;
        RECT 65.020 125.510 65.340 125.570 ;
        RECT 106.420 125.710 106.740 125.770 ;
        RECT 106.895 125.710 107.185 125.755 ;
        RECT 106.420 125.570 107.185 125.710 ;
        RECT 106.420 125.510 106.740 125.570 ;
        RECT 106.895 125.525 107.185 125.570 ;
        RECT 30.490 125.370 30.780 125.415 ;
        RECT 33.270 125.370 33.560 125.415 ;
        RECT 35.130 125.370 35.420 125.415 ;
        RECT 30.490 125.230 35.420 125.370 ;
        RECT 30.490 125.185 30.780 125.230 ;
        RECT 33.270 125.185 33.560 125.230 ;
        RECT 35.130 125.185 35.420 125.230 ;
        RECT 36.960 125.370 37.280 125.430 ;
        RECT 67.795 125.370 68.085 125.415 ;
        RECT 98.140 125.370 98.460 125.430 ;
        RECT 36.960 125.230 98.460 125.370 ;
        RECT 36.960 125.170 37.280 125.230 ;
        RECT 67.795 125.185 68.085 125.230 ;
        RECT 98.140 125.170 98.460 125.230 ;
        RECT 103.660 125.370 103.980 125.430 ;
        RECT 111.035 125.370 111.325 125.415 ;
        RECT 103.660 125.230 111.325 125.370 ;
        RECT 103.660 125.170 103.980 125.230 ;
        RECT 111.035 125.185 111.325 125.230 ;
        RECT 121.570 125.370 121.860 125.415 ;
        RECT 124.350 125.370 124.640 125.415 ;
        RECT 126.210 125.370 126.500 125.415 ;
        RECT 121.570 125.230 126.500 125.370 ;
        RECT 121.570 125.185 121.860 125.230 ;
        RECT 124.350 125.185 124.640 125.230 ;
        RECT 126.210 125.185 126.500 125.230 ;
        RECT 17.640 124.830 17.960 125.090 ;
        RECT 18.115 125.030 18.405 125.075 ;
        RECT 20.400 125.030 20.720 125.090 ;
        RECT 18.115 124.890 20.720 125.030 ;
        RECT 18.115 124.845 18.405 124.890 ;
        RECT 20.400 124.830 20.720 124.890 ;
        RECT 31.900 125.030 32.220 125.090 ;
        RECT 33.755 125.030 34.045 125.075 ;
        RECT 31.900 124.890 34.045 125.030 ;
        RECT 31.900 124.830 32.220 124.890 ;
        RECT 33.755 124.845 34.045 124.890 ;
        RECT 49.855 125.030 50.145 125.075 ;
        RECT 50.760 125.030 51.080 125.090 ;
        RECT 49.855 124.890 51.080 125.030 ;
        RECT 49.855 124.845 50.145 124.890 ;
        RECT 50.760 124.830 51.080 124.890 ;
        RECT 59.960 124.830 60.280 125.090 ;
        RECT 60.895 125.030 61.185 125.075 ;
        RECT 61.800 125.030 62.120 125.090 ;
        RECT 60.895 124.890 62.120 125.030 ;
        RECT 60.895 124.845 61.185 124.890 ;
        RECT 61.800 124.830 62.120 124.890 ;
        RECT 66.400 125.030 66.720 125.090 ;
        RECT 70.080 125.030 70.400 125.090 ;
        RECT 66.400 124.890 70.400 125.030 ;
        RECT 66.400 124.830 66.720 124.890 ;
        RECT 70.080 124.830 70.400 124.890 ;
        RECT 89.415 125.030 89.705 125.075 ;
        RECT 89.860 125.030 90.180 125.090 ;
        RECT 89.415 124.890 90.180 125.030 ;
        RECT 89.415 124.845 89.705 124.890 ;
        RECT 89.860 124.830 90.180 124.890 ;
        RECT 102.740 124.830 103.060 125.090 ;
        RECT 112.875 125.030 113.165 125.075 ;
        RECT 117.000 125.030 117.320 125.090 ;
        RECT 107.890 124.890 112.170 125.030 ;
        RECT 12.580 124.690 12.900 124.750 ;
        RECT 15.355 124.690 15.645 124.735 ;
        RECT 24.555 124.690 24.845 124.735 ;
        RECT 12.580 124.550 24.845 124.690 ;
        RECT 12.580 124.490 12.900 124.550 ;
        RECT 15.355 124.505 15.645 124.550 ;
        RECT 24.555 124.505 24.845 124.550 ;
        RECT 30.490 124.690 30.780 124.735 ;
        RECT 35.595 124.690 35.885 124.735 ;
        RECT 36.500 124.690 36.820 124.750 ;
        RECT 30.490 124.550 33.025 124.690 ;
        RECT 30.490 124.505 30.780 124.550 ;
        RECT 32.810 124.395 33.025 124.550 ;
        RECT 35.595 124.550 36.820 124.690 ;
        RECT 35.595 124.505 35.885 124.550 ;
        RECT 36.500 124.490 36.820 124.550 ;
        RECT 38.340 124.690 38.660 124.750 ;
        RECT 38.815 124.690 39.105 124.735 ;
        RECT 38.340 124.550 39.105 124.690 ;
        RECT 38.340 124.490 38.660 124.550 ;
        RECT 38.815 124.505 39.105 124.550 ;
        RECT 57.660 124.690 57.980 124.750 ;
        RECT 58.135 124.690 58.425 124.735 ;
        RECT 57.660 124.550 58.425 124.690 ;
        RECT 57.660 124.490 57.980 124.550 ;
        RECT 58.135 124.505 58.425 124.550 ;
        RECT 58.580 124.690 58.900 124.750 ;
        RECT 61.355 124.690 61.645 124.735 ;
        RECT 58.580 124.550 61.645 124.690 ;
        RECT 58.580 124.490 58.900 124.550 ;
        RECT 61.355 124.505 61.645 124.550 ;
        RECT 65.495 124.690 65.785 124.735 ;
        RECT 66.875 124.690 67.165 124.735 ;
        RECT 69.175 124.690 69.465 124.735 ;
        RECT 71.000 124.690 71.320 124.750 ;
        RECT 65.495 124.550 71.320 124.690 ;
        RECT 65.495 124.505 65.785 124.550 ;
        RECT 66.875 124.505 67.165 124.550 ;
        RECT 69.175 124.505 69.465 124.550 ;
        RECT 71.000 124.490 71.320 124.550 ;
        RECT 80.675 124.690 80.965 124.735 ;
        RECT 94.015 124.690 94.305 124.735 ;
        RECT 96.300 124.690 96.620 124.750 ;
        RECT 107.890 124.735 108.030 124.890 ;
        RECT 112.030 124.735 112.170 124.890 ;
        RECT 112.875 124.890 117.320 125.030 ;
        RECT 112.875 124.845 113.165 124.890 ;
        RECT 117.000 124.830 117.320 124.890 ;
        RECT 126.675 125.030 126.965 125.075 ;
        RECT 127.120 125.030 127.440 125.090 ;
        RECT 126.675 124.890 127.440 125.030 ;
        RECT 126.675 124.845 126.965 124.890 ;
        RECT 127.120 124.830 127.440 124.890 ;
        RECT 80.675 124.550 96.620 124.690 ;
        RECT 80.675 124.505 80.965 124.550 ;
        RECT 94.015 124.505 94.305 124.550 ;
        RECT 25.015 124.350 25.305 124.395 ;
        RECT 28.630 124.350 28.920 124.395 ;
        RECT 31.890 124.350 32.180 124.395 ;
        RECT 25.015 124.210 32.180 124.350 ;
        RECT 25.015 124.165 25.305 124.210 ;
        RECT 28.630 124.165 28.920 124.210 ;
        RECT 31.890 124.165 32.180 124.210 ;
        RECT 32.810 124.350 33.100 124.395 ;
        RECT 34.670 124.350 34.960 124.395 ;
        RECT 32.810 124.210 34.960 124.350 ;
        RECT 32.810 124.165 33.100 124.210 ;
        RECT 34.670 124.165 34.960 124.210 ;
        RECT 36.040 124.350 36.360 124.410 ;
        RECT 41.115 124.350 41.405 124.395 ;
        RECT 80.750 124.350 80.890 124.505 ;
        RECT 96.300 124.490 96.620 124.550 ;
        RECT 107.815 124.505 108.105 124.735 ;
        RECT 108.275 124.505 108.565 124.735 ;
        RECT 111.955 124.690 112.245 124.735 ;
        RECT 112.400 124.690 112.720 124.750 ;
        RECT 116.095 124.690 116.385 124.735 ;
        RECT 111.955 124.550 112.720 124.690 ;
        RECT 111.955 124.505 112.245 124.550 ;
        RECT 36.040 124.210 80.890 124.350 ;
        RECT 107.340 124.350 107.660 124.410 ;
        RECT 108.350 124.350 108.490 124.505 ;
        RECT 112.400 124.490 112.720 124.550 ;
        RECT 112.950 124.550 116.385 124.690 ;
        RECT 107.340 124.210 108.490 124.350 ;
        RECT 36.040 124.150 36.360 124.210 ;
        RECT 41.115 124.165 41.405 124.210 ;
        RECT 107.340 124.150 107.660 124.210 ;
        RECT 18.575 124.010 18.865 124.055 ;
        RECT 24.540 124.010 24.860 124.070 ;
        RECT 18.575 123.870 24.860 124.010 ;
        RECT 18.575 123.825 18.865 123.870 ;
        RECT 24.540 123.810 24.860 123.870 ;
        RECT 39.260 123.810 39.580 124.070 ;
        RECT 59.055 124.010 59.345 124.055 ;
        RECT 61.340 124.010 61.660 124.070 ;
        RECT 59.055 123.870 61.660 124.010 ;
        RECT 59.055 123.825 59.345 123.870 ;
        RECT 61.340 123.810 61.660 123.870 ;
        RECT 62.260 124.010 62.580 124.070 ;
        RECT 63.195 124.010 63.485 124.055 ;
        RECT 62.260 123.870 63.485 124.010 ;
        RECT 62.260 123.810 62.580 123.870 ;
        RECT 63.195 123.825 63.485 123.870 ;
        RECT 68.240 123.810 68.560 124.070 ;
        RECT 104.580 124.010 104.900 124.070 ;
        RECT 112.950 124.010 113.090 124.550 ;
        RECT 116.095 124.505 116.385 124.550 ;
        RECT 121.570 124.690 121.860 124.735 ;
        RECT 124.835 124.690 125.125 124.735 ;
        RECT 126.200 124.690 126.520 124.750 ;
        RECT 121.570 124.550 124.105 124.690 ;
        RECT 121.570 124.505 121.860 124.550 ;
        RECT 117.460 124.395 117.780 124.410 ;
        RECT 117.460 124.165 117.995 124.395 ;
        RECT 119.710 124.350 120.000 124.395 ;
        RECT 120.680 124.350 121.000 124.410 ;
        RECT 123.890 124.395 124.105 124.550 ;
        RECT 124.835 124.550 126.520 124.690 ;
        RECT 124.835 124.505 125.125 124.550 ;
        RECT 126.200 124.490 126.520 124.550 ;
        RECT 122.970 124.350 123.260 124.395 ;
        RECT 119.710 124.210 123.260 124.350 ;
        RECT 119.710 124.165 120.000 124.210 ;
        RECT 117.460 124.150 117.780 124.165 ;
        RECT 120.680 124.150 121.000 124.210 ;
        RECT 122.970 124.165 123.260 124.210 ;
        RECT 123.890 124.350 124.180 124.395 ;
        RECT 125.750 124.350 126.040 124.395 ;
        RECT 123.890 124.210 126.040 124.350 ;
        RECT 123.890 124.165 124.180 124.210 ;
        RECT 125.750 124.165 126.040 124.210 ;
        RECT 113.320 124.010 113.640 124.070 ;
        RECT 104.580 123.870 113.640 124.010 ;
        RECT 104.580 123.810 104.900 123.870 ;
        RECT 113.320 123.810 113.640 123.870 ;
        RECT 116.555 124.010 116.845 124.055 ;
        RECT 118.840 124.010 119.160 124.070 ;
        RECT 116.555 123.870 119.160 124.010 ;
        RECT 116.555 123.825 116.845 123.870 ;
        RECT 118.840 123.810 119.160 123.870 ;
        RECT 9.290 123.190 129.350 123.670 ;
        RECT 35.580 122.990 35.900 123.050 ;
        RECT 36.055 122.990 36.345 123.035 ;
        RECT 35.580 122.850 36.345 122.990 ;
        RECT 35.580 122.790 35.900 122.850 ;
        RECT 36.055 122.805 36.345 122.850 ;
        RECT 36.515 122.990 36.805 123.035 ;
        RECT 36.960 122.990 37.280 123.050 ;
        RECT 36.515 122.850 37.280 122.990 ;
        RECT 36.515 122.805 36.805 122.850 ;
        RECT 36.960 122.790 37.280 122.850 ;
        RECT 38.355 122.990 38.645 123.035 ;
        RECT 41.575 122.990 41.865 123.035 ;
        RECT 42.020 122.990 42.340 123.050 ;
        RECT 38.355 122.850 41.330 122.990 ;
        RECT 38.355 122.805 38.645 122.850 ;
        RECT 31.915 122.650 32.205 122.695 ;
        RECT 38.800 122.650 39.120 122.710 ;
        RECT 31.915 122.510 39.120 122.650 ;
        RECT 41.190 122.650 41.330 122.850 ;
        RECT 41.575 122.850 42.340 122.990 ;
        RECT 41.575 122.805 41.865 122.850 ;
        RECT 42.020 122.790 42.340 122.850 ;
        RECT 54.225 122.990 54.515 123.035 ;
        RECT 58.580 122.990 58.900 123.050 ;
        RECT 54.225 122.850 58.900 122.990 ;
        RECT 54.225 122.805 54.515 122.850 ;
        RECT 58.580 122.790 58.900 122.850 ;
        RECT 76.980 122.790 77.300 123.050 ;
        RECT 79.755 122.990 80.045 123.035 ;
        RECT 81.120 122.990 81.440 123.050 ;
        RECT 79.755 122.850 81.440 122.990 ;
        RECT 79.755 122.805 80.045 122.850 ;
        RECT 81.120 122.790 81.440 122.850 ;
        RECT 81.580 122.990 81.900 123.050 ;
        RECT 82.055 122.990 82.345 123.035 ;
        RECT 81.580 122.850 82.345 122.990 ;
        RECT 81.580 122.790 81.900 122.850 ;
        RECT 82.055 122.805 82.345 122.850 ;
        RECT 107.815 122.990 108.105 123.035 ;
        RECT 110.560 122.990 110.880 123.050 ;
        RECT 113.795 122.990 114.085 123.035 ;
        RECT 116.785 122.990 117.075 123.035 ;
        RECT 107.815 122.850 117.075 122.990 ;
        RECT 107.815 122.805 108.105 122.850 ;
        RECT 110.560 122.790 110.880 122.850 ;
        RECT 113.795 122.805 114.085 122.850 ;
        RECT 116.785 122.805 117.075 122.850 ;
        RECT 126.200 122.790 126.520 123.050 ;
        RECT 59.500 122.695 59.820 122.710 ;
        RECT 56.230 122.650 56.520 122.695 ;
        RECT 59.490 122.650 59.820 122.695 ;
        RECT 41.190 122.510 42.250 122.650 ;
        RECT 31.915 122.465 32.205 122.510 ;
        RECT 38.800 122.450 39.120 122.510 ;
        RECT 30.995 122.310 31.285 122.355 ;
        RECT 33.295 122.310 33.585 122.355 ;
        RECT 36.040 122.310 36.360 122.370 ;
        RECT 39.735 122.310 40.025 122.355 ;
        RECT 30.995 122.170 35.350 122.310 ;
        RECT 30.995 122.125 31.285 122.170 ;
        RECT 33.295 122.125 33.585 122.170 ;
        RECT 23.620 121.970 23.940 122.030 ;
        RECT 30.075 121.970 30.365 122.015 ;
        RECT 23.620 121.830 30.365 121.970 ;
        RECT 23.620 121.770 23.940 121.830 ;
        RECT 30.075 121.785 30.365 121.830 ;
        RECT 32.375 121.970 32.665 122.015 ;
        RECT 32.820 121.970 33.140 122.030 ;
        RECT 32.375 121.830 33.140 121.970 ;
        RECT 32.375 121.785 32.665 121.830 ;
        RECT 32.820 121.770 33.140 121.830 ;
        RECT 35.210 121.630 35.350 122.170 ;
        RECT 36.040 122.170 40.025 122.310 ;
        RECT 36.040 122.110 36.360 122.170 ;
        RECT 39.735 122.125 40.025 122.170 ;
        RECT 40.180 122.310 40.500 122.370 ;
        RECT 42.110 122.355 42.250 122.510 ;
        RECT 56.230 122.510 59.820 122.650 ;
        RECT 56.230 122.465 56.520 122.510 ;
        RECT 59.490 122.465 59.820 122.510 ;
        RECT 59.500 122.450 59.820 122.465 ;
        RECT 60.410 122.650 60.700 122.695 ;
        RECT 62.270 122.650 62.560 122.695 ;
        RECT 60.410 122.510 62.560 122.650 ;
        RECT 60.410 122.465 60.700 122.510 ;
        RECT 62.270 122.465 62.560 122.510 ;
        RECT 66.875 122.650 67.165 122.695 ;
        RECT 68.240 122.650 68.560 122.710 ;
        RECT 69.635 122.650 69.925 122.695 ;
        RECT 66.875 122.510 69.925 122.650 ;
        RECT 66.875 122.465 67.165 122.510 ;
        RECT 40.655 122.310 40.945 122.355 ;
        RECT 40.180 122.170 40.945 122.310 ;
        RECT 40.180 122.110 40.500 122.170 ;
        RECT 40.655 122.125 40.945 122.170 ;
        RECT 42.035 122.125 42.325 122.355 ;
        RECT 49.395 122.310 49.685 122.355 ;
        RECT 50.760 122.310 51.080 122.370 ;
        RECT 49.395 122.170 51.080 122.310 ;
        RECT 49.395 122.125 49.685 122.170 ;
        RECT 50.760 122.110 51.080 122.170 ;
        RECT 58.090 122.310 58.380 122.355 ;
        RECT 60.410 122.310 60.625 122.465 ;
        RECT 68.240 122.450 68.560 122.510 ;
        RECT 69.635 122.465 69.925 122.510 ;
        RECT 113.335 122.650 113.625 122.695 ;
        RECT 114.240 122.650 114.560 122.710 ;
        RECT 117.460 122.650 117.780 122.710 ;
        RECT 118.840 122.695 119.160 122.710 ;
        RECT 113.335 122.510 117.780 122.650 ;
        RECT 113.335 122.465 113.625 122.510 ;
        RECT 114.240 122.450 114.560 122.510 ;
        RECT 117.460 122.450 117.780 122.510 ;
        RECT 118.790 122.650 119.160 122.695 ;
        RECT 122.050 122.650 122.340 122.695 ;
        RECT 118.790 122.510 122.340 122.650 ;
        RECT 118.790 122.465 119.160 122.510 ;
        RECT 122.050 122.465 122.340 122.510 ;
        RECT 122.970 122.650 123.260 122.695 ;
        RECT 124.830 122.650 125.120 122.695 ;
        RECT 122.970 122.510 125.120 122.650 ;
        RECT 122.970 122.465 123.260 122.510 ;
        RECT 124.830 122.465 125.120 122.510 ;
        RECT 118.840 122.450 119.160 122.465 ;
        RECT 58.090 122.170 60.625 122.310 ;
        RECT 58.090 122.125 58.380 122.170 ;
        RECT 61.340 122.110 61.660 122.370 ;
        RECT 62.720 122.310 63.040 122.370 ;
        RECT 63.195 122.310 63.485 122.355 ;
        RECT 62.720 122.170 63.485 122.310 ;
        RECT 62.720 122.110 63.040 122.170 ;
        RECT 63.195 122.125 63.485 122.170 ;
        RECT 65.020 122.310 65.340 122.370 ;
        RECT 75.615 122.310 75.905 122.355 ;
        RECT 77.915 122.310 78.205 122.355 ;
        RECT 80.675 122.310 80.965 122.355 ;
        RECT 82.975 122.310 83.265 122.355 ;
        RECT 65.020 122.170 83.265 122.310 ;
        RECT 65.020 122.110 65.340 122.170 ;
        RECT 75.615 122.125 75.905 122.170 ;
        RECT 77.915 122.125 78.205 122.170 ;
        RECT 80.675 122.125 80.965 122.170 ;
        RECT 82.975 122.125 83.265 122.170 ;
        RECT 88.955 122.310 89.245 122.355 ;
        RECT 89.860 122.310 90.180 122.370 ;
        RECT 88.955 122.170 90.180 122.310 ;
        RECT 88.955 122.125 89.245 122.170 ;
        RECT 89.860 122.110 90.180 122.170 ;
        RECT 104.580 122.110 104.900 122.370 ;
        RECT 106.420 122.310 106.740 122.370 ;
        RECT 108.275 122.310 108.565 122.355 ;
        RECT 106.420 122.170 108.565 122.310 ;
        RECT 106.420 122.110 106.740 122.170 ;
        RECT 108.275 122.125 108.565 122.170 ;
        RECT 120.650 122.310 120.940 122.355 ;
        RECT 122.970 122.310 123.185 122.465 ;
        RECT 120.650 122.170 123.185 122.310 ;
        RECT 125.755 122.310 126.045 122.355 ;
        RECT 126.660 122.310 126.980 122.370 ;
        RECT 125.755 122.170 126.980 122.310 ;
        RECT 120.650 122.125 120.940 122.170 ;
        RECT 125.755 122.125 126.045 122.170 ;
        RECT 126.660 122.110 126.980 122.170 ;
        RECT 127.135 122.125 127.425 122.355 ;
        RECT 35.580 121.770 35.900 122.030 ;
        RECT 74.680 121.770 75.000 122.030 ;
        RECT 78.820 121.770 79.140 122.030 ;
        RECT 81.595 121.970 81.885 122.015 ;
        RECT 83.420 121.970 83.740 122.030 ;
        RECT 81.595 121.830 83.740 121.970 ;
        RECT 81.595 121.785 81.885 121.830 ;
        RECT 83.420 121.770 83.740 121.830 ;
        RECT 83.895 121.970 84.185 122.015 ;
        RECT 84.340 121.970 84.660 122.030 ;
        RECT 83.895 121.830 84.660 121.970 ;
        RECT 83.895 121.785 84.185 121.830 ;
        RECT 84.340 121.770 84.660 121.830 ;
        RECT 107.355 121.970 107.645 122.015 ;
        RECT 107.800 121.970 108.120 122.030 ;
        RECT 112.415 121.970 112.705 122.015 ;
        RECT 113.780 121.970 114.100 122.030 ;
        RECT 107.355 121.830 114.100 121.970 ;
        RECT 107.355 121.785 107.645 121.830 ;
        RECT 107.800 121.770 108.120 121.830 ;
        RECT 112.415 121.785 112.705 121.830 ;
        RECT 113.780 121.770 114.100 121.830 ;
        RECT 122.520 121.970 122.840 122.030 ;
        RECT 123.915 121.970 124.205 122.015 ;
        RECT 122.520 121.830 124.205 121.970 ;
        RECT 122.520 121.770 122.840 121.830 ;
        RECT 123.915 121.785 124.205 121.830 ;
        RECT 37.420 121.630 37.740 121.690 ;
        RECT 35.210 121.490 37.740 121.630 ;
        RECT 37.420 121.430 37.740 121.490 ;
        RECT 58.090 121.630 58.380 121.675 ;
        RECT 60.870 121.630 61.160 121.675 ;
        RECT 62.730 121.630 63.020 121.675 ;
        RECT 58.090 121.490 63.020 121.630 ;
        RECT 58.090 121.445 58.380 121.490 ;
        RECT 60.870 121.445 61.160 121.490 ;
        RECT 62.730 121.445 63.020 121.490 ;
        RECT 76.535 121.630 76.825 121.675 ;
        RECT 82.960 121.630 83.280 121.690 ;
        RECT 76.535 121.490 83.280 121.630 ;
        RECT 76.535 121.445 76.825 121.490 ;
        RECT 82.960 121.430 83.280 121.490 ;
        RECT 120.650 121.630 120.940 121.675 ;
        RECT 123.430 121.630 123.720 121.675 ;
        RECT 125.290 121.630 125.580 121.675 ;
        RECT 120.650 121.490 125.580 121.630 ;
        RECT 120.650 121.445 120.940 121.490 ;
        RECT 123.430 121.445 123.720 121.490 ;
        RECT 125.290 121.445 125.580 121.490 ;
        RECT 34.215 121.290 34.505 121.335 ;
        RECT 40.640 121.290 40.960 121.350 ;
        RECT 34.215 121.150 40.960 121.290 ;
        RECT 34.215 121.105 34.505 121.150 ;
        RECT 40.640 121.090 40.960 121.150 ;
        RECT 42.940 121.090 43.260 121.350 ;
        RECT 50.760 121.290 51.080 121.350 ;
        RECT 65.495 121.290 65.785 121.335 ;
        RECT 50.760 121.150 65.785 121.290 ;
        RECT 50.760 121.090 51.080 121.150 ;
        RECT 65.495 121.105 65.785 121.150 ;
        RECT 71.015 121.290 71.305 121.335 ;
        RECT 73.300 121.290 73.620 121.350 ;
        RECT 71.015 121.150 73.620 121.290 ;
        RECT 71.015 121.105 71.305 121.150 ;
        RECT 73.300 121.090 73.620 121.150 ;
        RECT 105.040 121.090 105.360 121.350 ;
        RECT 110.115 121.290 110.405 121.335 ;
        RECT 110.560 121.290 110.880 121.350 ;
        RECT 110.115 121.150 110.880 121.290 ;
        RECT 110.115 121.105 110.405 121.150 ;
        RECT 110.560 121.090 110.880 121.150 ;
        RECT 115.635 121.290 115.925 121.335 ;
        RECT 117.920 121.290 118.240 121.350 ;
        RECT 115.635 121.150 118.240 121.290 ;
        RECT 115.635 121.105 115.925 121.150 ;
        RECT 117.920 121.090 118.240 121.150 ;
        RECT 119.300 121.290 119.620 121.350 ;
        RECT 127.210 121.290 127.350 122.125 ;
        RECT 119.300 121.150 127.350 121.290 ;
        RECT 119.300 121.090 119.620 121.150 ;
        RECT 9.290 120.470 129.350 120.950 ;
        RECT 37.420 120.270 37.740 120.330 ;
        RECT 40.180 120.270 40.500 120.330 ;
        RECT 43.860 120.270 44.180 120.330 ;
        RECT 37.420 120.130 44.180 120.270 ;
        RECT 37.420 120.070 37.740 120.130 ;
        RECT 40.180 120.070 40.500 120.130 ;
        RECT 43.860 120.070 44.180 120.130 ;
        RECT 44.780 120.270 45.100 120.330 ;
        RECT 45.255 120.270 45.545 120.315 ;
        RECT 44.780 120.130 45.545 120.270 ;
        RECT 44.780 120.070 45.100 120.130 ;
        RECT 45.255 120.085 45.545 120.130 ;
        RECT 47.080 120.270 47.400 120.330 ;
        RECT 48.475 120.270 48.765 120.315 ;
        RECT 47.080 120.130 48.765 120.270 ;
        RECT 47.080 120.070 47.400 120.130 ;
        RECT 48.475 120.085 48.765 120.130 ;
        RECT 59.055 120.270 59.345 120.315 ;
        RECT 59.500 120.270 59.820 120.330 ;
        RECT 59.055 120.130 59.820 120.270 ;
        RECT 59.055 120.085 59.345 120.130 ;
        RECT 59.500 120.070 59.820 120.130 ;
        RECT 119.300 120.070 119.620 120.330 ;
        RECT 120.680 120.070 121.000 120.330 ;
        RECT 122.520 120.070 122.840 120.330 ;
        RECT 39.690 119.930 39.980 119.975 ;
        RECT 42.470 119.930 42.760 119.975 ;
        RECT 44.330 119.930 44.620 119.975 ;
        RECT 51.680 119.930 52.000 119.990 ;
        RECT 39.690 119.790 44.620 119.930 ;
        RECT 39.690 119.745 39.980 119.790 ;
        RECT 42.470 119.745 42.760 119.790 ;
        RECT 44.330 119.745 44.620 119.790 ;
        RECT 44.870 119.790 52.000 119.930 ;
        RECT 17.640 119.590 17.960 119.650 ;
        RECT 25.015 119.590 25.305 119.635 ;
        RECT 34.215 119.590 34.505 119.635 ;
        RECT 35.580 119.590 35.900 119.650 ;
        RECT 42.020 119.590 42.340 119.650 ;
        RECT 17.640 119.450 42.340 119.590 ;
        RECT 17.640 119.390 17.960 119.450 ;
        RECT 25.015 119.405 25.305 119.450 ;
        RECT 34.215 119.405 34.505 119.450 ;
        RECT 35.580 119.390 35.900 119.450 ;
        RECT 42.020 119.390 42.340 119.450 ;
        RECT 42.940 119.390 43.260 119.650 ;
        RECT 43.860 119.390 44.180 119.650 ;
        RECT 44.870 119.635 45.010 119.790 ;
        RECT 51.680 119.730 52.000 119.790 ;
        RECT 73.300 119.930 73.620 119.990 ;
        RECT 91.210 119.930 91.500 119.975 ;
        RECT 93.990 119.930 94.280 119.975 ;
        RECT 95.850 119.930 96.140 119.975 ;
        RECT 102.740 119.930 103.060 119.990 ;
        RECT 73.300 119.790 82.730 119.930 ;
        RECT 73.300 119.730 73.620 119.790 ;
        RECT 82.590 119.650 82.730 119.790 ;
        RECT 91.210 119.790 96.140 119.930 ;
        RECT 91.210 119.745 91.500 119.790 ;
        RECT 93.990 119.745 94.280 119.790 ;
        RECT 95.850 119.745 96.140 119.790 ;
        RECT 96.390 119.790 103.060 119.930 ;
        RECT 44.795 119.405 45.085 119.635 ;
        RECT 46.620 119.590 46.940 119.650 ;
        RECT 74.220 119.590 74.540 119.650 ;
        RECT 78.820 119.590 79.140 119.650 ;
        RECT 81.580 119.590 81.900 119.650 ;
        RECT 46.250 119.450 49.610 119.590 ;
        RECT 18.100 119.250 18.420 119.310 ;
        RECT 18.575 119.250 18.865 119.295 ;
        RECT 22.700 119.250 23.020 119.310 ;
        RECT 18.100 119.110 23.020 119.250 ;
        RECT 18.100 119.050 18.420 119.110 ;
        RECT 18.575 119.065 18.865 119.110 ;
        RECT 22.700 119.050 23.020 119.110 ;
        RECT 24.095 119.250 24.385 119.295 ;
        RECT 24.540 119.250 24.860 119.310 ;
        RECT 32.820 119.250 33.140 119.310 ;
        RECT 24.095 119.110 33.140 119.250 ;
        RECT 24.095 119.065 24.385 119.110 ;
        RECT 24.540 119.050 24.860 119.110 ;
        RECT 32.820 119.050 33.140 119.110 ;
        RECT 33.280 119.250 33.600 119.310 ;
        RECT 36.040 119.250 36.360 119.310 ;
        RECT 33.280 119.110 36.360 119.250 ;
        RECT 33.280 119.050 33.600 119.110 ;
        RECT 36.040 119.050 36.360 119.110 ;
        RECT 39.690 119.250 39.980 119.295 ;
        RECT 43.950 119.250 44.090 119.390 ;
        RECT 46.250 119.295 46.390 119.450 ;
        RECT 46.620 119.390 46.940 119.450 ;
        RECT 46.175 119.250 46.465 119.295 ;
        RECT 39.690 119.110 42.225 119.250 ;
        RECT 43.950 119.110 46.465 119.250 ;
        RECT 39.690 119.065 39.980 119.110 ;
        RECT 23.620 118.910 23.940 118.970 ;
        RECT 18.190 118.770 23.940 118.910 ;
        RECT 17.640 118.570 17.960 118.630 ;
        RECT 18.190 118.615 18.330 118.770 ;
        RECT 23.620 118.710 23.940 118.770 ;
        RECT 37.830 118.910 38.120 118.955 ;
        RECT 39.260 118.910 39.580 118.970 ;
        RECT 42.010 118.955 42.225 119.110 ;
        RECT 46.175 119.065 46.465 119.110 ;
        RECT 47.080 119.050 47.400 119.310 ;
        RECT 49.470 119.295 49.610 119.450 ;
        RECT 74.220 119.450 81.900 119.590 ;
        RECT 74.220 119.390 74.540 119.450 ;
        RECT 78.820 119.390 79.140 119.450 ;
        RECT 81.580 119.390 81.900 119.450 ;
        RECT 82.500 119.390 82.820 119.650 ;
        RECT 94.475 119.590 94.765 119.635 ;
        RECT 95.380 119.590 95.700 119.650 ;
        RECT 96.390 119.635 96.530 119.790 ;
        RECT 102.740 119.730 103.060 119.790 ;
        RECT 107.770 119.930 108.060 119.975 ;
        RECT 110.550 119.930 110.840 119.975 ;
        RECT 112.410 119.930 112.700 119.975 ;
        RECT 107.770 119.790 112.700 119.930 ;
        RECT 107.770 119.745 108.060 119.790 ;
        RECT 110.550 119.745 110.840 119.790 ;
        RECT 112.410 119.745 112.700 119.790 ;
        RECT 94.475 119.450 95.700 119.590 ;
        RECT 94.475 119.405 94.765 119.450 ;
        RECT 95.380 119.390 95.700 119.450 ;
        RECT 96.315 119.405 96.605 119.635 ;
        RECT 98.600 119.390 98.920 119.650 ;
        RECT 99.535 119.590 99.825 119.635 ;
        RECT 103.905 119.590 104.195 119.635 ;
        RECT 106.420 119.590 106.740 119.650 ;
        RECT 99.535 119.450 106.740 119.590 ;
        RECT 99.535 119.405 99.825 119.450 ;
        RECT 103.905 119.405 104.195 119.450 ;
        RECT 106.420 119.390 106.740 119.450 ;
        RECT 113.780 119.590 114.100 119.650 ;
        RECT 116.095 119.590 116.385 119.635 ;
        RECT 113.780 119.450 116.385 119.590 ;
        RECT 113.780 119.390 114.100 119.450 ;
        RECT 116.095 119.405 116.385 119.450 ;
        RECT 117.000 119.390 117.320 119.650 ;
        RECT 117.920 119.590 118.240 119.650 ;
        RECT 117.920 119.450 121.830 119.590 ;
        RECT 117.920 119.390 118.240 119.450 ;
        RECT 49.395 119.065 49.685 119.295 ;
        RECT 50.315 119.250 50.605 119.295 ;
        RECT 51.220 119.250 51.540 119.310 ;
        RECT 50.315 119.110 51.540 119.250 ;
        RECT 50.315 119.065 50.605 119.110 ;
        RECT 51.220 119.050 51.540 119.110 ;
        RECT 59.515 119.250 59.805 119.295 ;
        RECT 60.880 119.250 61.200 119.310 ;
        RECT 59.515 119.110 61.200 119.250 ;
        RECT 59.515 119.065 59.805 119.110 ;
        RECT 60.880 119.050 61.200 119.110 ;
        RECT 62.260 119.250 62.580 119.310 ;
        RECT 64.575 119.250 64.865 119.295 ;
        RECT 62.260 119.110 64.865 119.250 ;
        RECT 62.260 119.050 62.580 119.110 ;
        RECT 64.575 119.065 64.865 119.110 ;
        RECT 80.215 119.250 80.505 119.295 ;
        RECT 81.120 119.250 81.440 119.310 ;
        RECT 80.215 119.110 81.440 119.250 ;
        RECT 80.215 119.065 80.505 119.110 ;
        RECT 81.120 119.050 81.440 119.110 ;
        RECT 83.420 119.250 83.740 119.310 ;
        RECT 87.345 119.250 87.635 119.295 ;
        RECT 83.420 119.110 87.635 119.250 ;
        RECT 83.420 119.050 83.740 119.110 ;
        RECT 87.345 119.065 87.635 119.110 ;
        RECT 91.210 119.250 91.500 119.295 ;
        RECT 97.680 119.250 98.000 119.310 ;
        RECT 99.995 119.250 100.285 119.295 ;
        RECT 91.210 119.110 93.745 119.250 ;
        RECT 91.210 119.065 91.500 119.110 ;
        RECT 41.090 118.910 41.380 118.955 ;
        RECT 37.830 118.770 41.380 118.910 ;
        RECT 37.830 118.725 38.120 118.770 ;
        RECT 39.260 118.710 39.580 118.770 ;
        RECT 41.090 118.725 41.380 118.770 ;
        RECT 42.010 118.910 42.300 118.955 ;
        RECT 43.870 118.910 44.160 118.955 ;
        RECT 42.010 118.770 44.160 118.910 ;
        RECT 42.010 118.725 42.300 118.770 ;
        RECT 43.870 118.725 44.160 118.770 ;
        RECT 74.680 118.910 75.000 118.970 ;
        RECT 92.620 118.955 92.940 118.970 ;
        RECT 82.975 118.910 83.265 118.955 ;
        RECT 74.680 118.770 83.265 118.910 ;
        RECT 74.680 118.710 75.000 118.770 ;
        RECT 82.975 118.725 83.265 118.770 ;
        RECT 89.350 118.910 89.640 118.955 ;
        RECT 92.610 118.910 92.940 118.955 ;
        RECT 89.350 118.770 92.940 118.910 ;
        RECT 89.350 118.725 89.640 118.770 ;
        RECT 92.610 118.725 92.940 118.770 ;
        RECT 93.530 118.955 93.745 119.110 ;
        RECT 97.680 119.110 100.285 119.250 ;
        RECT 97.680 119.050 98.000 119.110 ;
        RECT 99.995 119.065 100.285 119.110 ;
        RECT 107.770 119.250 108.060 119.295 ;
        RECT 107.770 119.110 110.305 119.250 ;
        RECT 107.770 119.065 108.060 119.110 ;
        RECT 93.530 118.910 93.820 118.955 ;
        RECT 95.390 118.910 95.680 118.955 ;
        RECT 93.530 118.770 95.680 118.910 ;
        RECT 93.530 118.725 93.820 118.770 ;
        RECT 95.390 118.725 95.680 118.770 ;
        RECT 105.040 118.910 105.360 118.970 ;
        RECT 110.090 118.955 110.305 119.110 ;
        RECT 111.020 119.050 111.340 119.310 ;
        RECT 112.875 119.065 113.165 119.295 ;
        RECT 105.910 118.910 106.200 118.955 ;
        RECT 109.170 118.910 109.460 118.955 ;
        RECT 105.040 118.770 109.460 118.910 ;
        RECT 92.620 118.710 92.940 118.725 ;
        RECT 105.040 118.710 105.360 118.770 ;
        RECT 105.910 118.725 106.200 118.770 ;
        RECT 109.170 118.725 109.460 118.770 ;
        RECT 110.090 118.910 110.380 118.955 ;
        RECT 111.950 118.910 112.240 118.955 ;
        RECT 110.090 118.770 112.240 118.910 ;
        RECT 112.950 118.910 113.090 119.065 ;
        RECT 117.460 119.050 117.780 119.310 ;
        RECT 120.220 119.050 120.540 119.310 ;
        RECT 121.690 119.295 121.830 119.450 ;
        RECT 121.615 119.065 121.905 119.295 ;
        RECT 126.660 118.910 126.980 118.970 ;
        RECT 112.950 118.770 126.980 118.910 ;
        RECT 110.090 118.725 110.380 118.770 ;
        RECT 111.950 118.725 112.240 118.770 ;
        RECT 126.660 118.710 126.980 118.770 ;
        RECT 18.115 118.570 18.405 118.615 ;
        RECT 17.640 118.430 18.405 118.570 ;
        RECT 17.640 118.370 17.960 118.430 ;
        RECT 18.115 118.385 18.405 118.430 ;
        RECT 20.415 118.570 20.705 118.615 ;
        RECT 21.320 118.570 21.640 118.630 ;
        RECT 20.415 118.430 21.640 118.570 ;
        RECT 20.415 118.385 20.705 118.430 ;
        RECT 21.320 118.370 21.640 118.430 ;
        RECT 21.795 118.570 22.085 118.615 ;
        RECT 24.080 118.570 24.400 118.630 ;
        RECT 21.795 118.430 24.400 118.570 ;
        RECT 21.795 118.385 22.085 118.430 ;
        RECT 24.080 118.370 24.400 118.430 ;
        RECT 30.520 118.570 30.840 118.630 ;
        RECT 30.995 118.570 31.285 118.615 ;
        RECT 30.520 118.430 31.285 118.570 ;
        RECT 30.520 118.370 30.840 118.430 ;
        RECT 30.995 118.385 31.285 118.430 ;
        RECT 35.825 118.570 36.115 118.615 ;
        RECT 36.960 118.570 37.280 118.630 ;
        RECT 47.540 118.570 47.860 118.630 ;
        RECT 35.825 118.430 47.860 118.570 ;
        RECT 35.825 118.385 36.115 118.430 ;
        RECT 36.960 118.370 37.280 118.430 ;
        RECT 47.540 118.370 47.860 118.430 ;
        RECT 65.480 118.370 65.800 118.630 ;
        RECT 77.900 118.570 78.220 118.630 ;
        RECT 79.295 118.570 79.585 118.615 ;
        RECT 77.900 118.430 79.585 118.570 ;
        RECT 77.900 118.370 78.220 118.430 ;
        RECT 79.295 118.385 79.585 118.430 ;
        RECT 83.435 118.570 83.725 118.615 ;
        RECT 84.340 118.570 84.660 118.630 ;
        RECT 83.435 118.430 84.660 118.570 ;
        RECT 83.435 118.385 83.725 118.430 ;
        RECT 84.340 118.370 84.660 118.430 ;
        RECT 85.260 118.370 85.580 118.630 ;
        RECT 101.820 118.370 102.140 118.630 ;
        RECT 9.290 117.750 129.350 118.230 ;
        RECT 15.125 117.550 15.415 117.595 ;
        RECT 17.640 117.550 17.960 117.610 ;
        RECT 15.125 117.410 17.960 117.550 ;
        RECT 15.125 117.365 15.415 117.410 ;
        RECT 17.640 117.350 17.960 117.410 ;
        RECT 24.540 117.595 24.860 117.610 ;
        RECT 24.540 117.365 25.075 117.595 ;
        RECT 47.540 117.550 47.860 117.610 ;
        RECT 51.235 117.550 51.525 117.595 ;
        RECT 47.540 117.410 51.525 117.550 ;
        RECT 24.540 117.350 24.860 117.365 ;
        RECT 47.540 117.350 47.860 117.410 ;
        RECT 51.235 117.365 51.525 117.410 ;
        RECT 53.535 117.550 53.825 117.595 ;
        RECT 53.535 117.410 54.210 117.550 ;
        RECT 53.535 117.365 53.825 117.410 ;
        RECT 13.975 117.210 14.265 117.255 ;
        RECT 17.130 117.210 17.420 117.255 ;
        RECT 20.390 117.210 20.680 117.255 ;
        RECT 13.975 117.070 20.680 117.210 ;
        RECT 13.975 117.025 14.265 117.070 ;
        RECT 17.130 117.025 17.420 117.070 ;
        RECT 20.390 117.025 20.680 117.070 ;
        RECT 21.310 117.210 21.600 117.255 ;
        RECT 23.170 117.210 23.460 117.255 ;
        RECT 21.310 117.070 23.460 117.210 ;
        RECT 21.310 117.025 21.600 117.070 ;
        RECT 23.170 117.025 23.460 117.070 ;
        RECT 26.790 117.210 27.080 117.255 ;
        RECT 29.140 117.210 29.460 117.270 ;
        RECT 30.050 117.210 30.340 117.255 ;
        RECT 26.790 117.070 30.340 117.210 ;
        RECT 26.790 117.025 27.080 117.070 ;
        RECT 12.580 116.870 12.900 116.930 ;
        RECT 13.515 116.870 13.805 116.915 ;
        RECT 12.580 116.730 13.805 116.870 ;
        RECT 12.580 116.670 12.900 116.730 ;
        RECT 13.515 116.685 13.805 116.730 ;
        RECT 18.990 116.870 19.280 116.915 ;
        RECT 21.310 116.870 21.525 117.025 ;
        RECT 29.140 117.010 29.460 117.070 ;
        RECT 30.050 117.025 30.340 117.070 ;
        RECT 30.970 117.210 31.260 117.255 ;
        RECT 32.830 117.210 33.120 117.255 ;
        RECT 30.970 117.070 33.120 117.210 ;
        RECT 30.970 117.025 31.260 117.070 ;
        RECT 32.830 117.025 33.120 117.070 ;
        RECT 42.020 117.210 42.340 117.270 ;
        RECT 50.760 117.210 51.080 117.270 ;
        RECT 42.020 117.070 51.080 117.210 ;
        RECT 18.990 116.730 21.525 116.870 ;
        RECT 18.990 116.685 19.280 116.730 ;
        RECT 22.240 116.670 22.560 116.930 ;
        RECT 28.650 116.870 28.940 116.915 ;
        RECT 30.970 116.870 31.185 117.025 ;
        RECT 42.020 117.010 42.340 117.070 ;
        RECT 50.760 117.010 51.080 117.070 ;
        RECT 28.650 116.730 31.185 116.870 ;
        RECT 31.440 116.870 31.760 116.930 ;
        RECT 31.915 116.870 32.205 116.915 ;
        RECT 31.440 116.730 32.205 116.870 ;
        RECT 28.650 116.685 28.940 116.730 ;
        RECT 31.440 116.670 31.760 116.730 ;
        RECT 31.915 116.685 32.205 116.730 ;
        RECT 32.360 116.870 32.680 116.930 ;
        RECT 35.135 116.870 35.425 116.915 ;
        RECT 38.340 116.870 38.660 116.930 ;
        RECT 32.360 116.730 41.330 116.870 ;
        RECT 32.360 116.670 32.680 116.730 ;
        RECT 35.135 116.685 35.425 116.730 ;
        RECT 38.340 116.670 38.660 116.730 ;
        RECT 20.860 116.530 21.180 116.590 ;
        RECT 24.095 116.530 24.385 116.575 ;
        RECT 33.755 116.530 34.045 116.575 ;
        RECT 36.500 116.530 36.820 116.590 ;
        RECT 41.190 116.530 41.330 116.730 ;
        RECT 41.560 116.670 41.880 116.930 ;
        RECT 48.475 116.870 48.765 116.915 ;
        RECT 51.220 116.870 51.540 116.930 ;
        RECT 54.070 116.915 54.210 117.410 ;
        RECT 81.120 117.350 81.440 117.610 ;
        RECT 81.580 117.550 81.900 117.610 ;
        RECT 82.975 117.550 83.265 117.595 ;
        RECT 81.580 117.410 83.265 117.550 ;
        RECT 81.580 117.350 81.900 117.410 ;
        RECT 82.975 117.365 83.265 117.410 ;
        RECT 83.420 117.350 83.740 117.610 ;
        RECT 87.575 117.550 87.865 117.595 ;
        RECT 91.945 117.550 92.235 117.595 ;
        RECT 97.680 117.550 98.000 117.610 ;
        RECT 101.375 117.550 101.665 117.595 ;
        RECT 87.575 117.410 98.000 117.550 ;
        RECT 87.575 117.365 87.865 117.410 ;
        RECT 91.945 117.365 92.235 117.410 ;
        RECT 97.680 117.350 98.000 117.410 ;
        RECT 100.530 117.410 101.665 117.550 ;
        RECT 76.980 117.255 77.300 117.270 ;
        RECT 73.710 117.210 74.000 117.255 ;
        RECT 76.970 117.210 77.300 117.255 ;
        RECT 73.710 117.070 77.300 117.210 ;
        RECT 73.710 117.025 74.000 117.070 ;
        RECT 76.970 117.025 77.300 117.070 ;
        RECT 76.980 117.010 77.300 117.025 ;
        RECT 77.890 117.210 78.180 117.255 ;
        RECT 79.750 117.210 80.040 117.255 ;
        RECT 77.890 117.070 80.040 117.210 ;
        RECT 83.510 117.210 83.650 117.350 ;
        RECT 88.035 117.210 88.325 117.255 ;
        RECT 83.510 117.070 88.325 117.210 ;
        RECT 77.890 117.025 78.180 117.070 ;
        RECT 79.750 117.025 80.040 117.070 ;
        RECT 88.035 117.025 88.325 117.070 ;
        RECT 93.950 117.210 94.240 117.255 ;
        RECT 96.300 117.210 96.620 117.270 ;
        RECT 97.210 117.210 97.500 117.255 ;
        RECT 93.950 117.070 97.500 117.210 ;
        RECT 93.950 117.025 94.240 117.070 ;
        RECT 51.695 116.870 51.985 116.915 ;
        RECT 46.250 116.730 49.610 116.870 ;
        RECT 46.250 116.590 46.390 116.730 ;
        RECT 48.475 116.685 48.765 116.730 ;
        RECT 46.160 116.530 46.480 116.590 ;
        RECT 20.860 116.390 38.340 116.530 ;
        RECT 41.190 116.390 46.480 116.530 ;
        RECT 20.860 116.330 21.180 116.390 ;
        RECT 24.095 116.345 24.385 116.390 ;
        RECT 33.755 116.345 34.045 116.390 ;
        RECT 36.500 116.330 36.820 116.390 ;
        RECT 18.990 116.190 19.280 116.235 ;
        RECT 21.770 116.190 22.060 116.235 ;
        RECT 23.630 116.190 23.920 116.235 ;
        RECT 18.990 116.050 23.920 116.190 ;
        RECT 18.990 116.005 19.280 116.050 ;
        RECT 21.770 116.005 22.060 116.050 ;
        RECT 23.630 116.005 23.920 116.050 ;
        RECT 28.650 116.190 28.940 116.235 ;
        RECT 31.430 116.190 31.720 116.235 ;
        RECT 33.290 116.190 33.580 116.235 ;
        RECT 28.650 116.050 33.580 116.190 ;
        RECT 38.200 116.190 38.340 116.390 ;
        RECT 46.160 116.330 46.480 116.390 ;
        RECT 48.000 116.530 48.320 116.590 ;
        RECT 48.935 116.530 49.225 116.575 ;
        RECT 48.000 116.390 49.225 116.530 ;
        RECT 48.000 116.330 48.320 116.390 ;
        RECT 48.935 116.345 49.225 116.390 ;
        RECT 41.100 116.190 41.420 116.250 ;
        RECT 38.200 116.050 41.420 116.190 ;
        RECT 49.470 116.190 49.610 116.730 ;
        RECT 51.220 116.730 51.985 116.870 ;
        RECT 51.220 116.670 51.540 116.730 ;
        RECT 51.695 116.685 51.985 116.730 ;
        RECT 53.995 116.685 54.285 116.915 ;
        RECT 57.675 116.870 57.965 116.915 ;
        RECT 60.880 116.870 61.200 116.930 ;
        RECT 62.735 116.870 63.025 116.915 ;
        RECT 57.675 116.730 63.025 116.870 ;
        RECT 57.675 116.685 57.965 116.730 ;
        RECT 60.880 116.670 61.200 116.730 ;
        RECT 62.735 116.685 63.025 116.730 ;
        RECT 75.570 116.870 75.860 116.915 ;
        RECT 77.890 116.870 78.105 117.025 ;
        RECT 96.300 117.010 96.620 117.070 ;
        RECT 97.210 117.025 97.500 117.070 ;
        RECT 98.130 117.210 98.420 117.255 ;
        RECT 99.990 117.210 100.280 117.255 ;
        RECT 98.130 117.070 100.280 117.210 ;
        RECT 98.130 117.025 98.420 117.070 ;
        RECT 99.990 117.025 100.280 117.070 ;
        RECT 75.570 116.730 78.105 116.870 ;
        RECT 75.570 116.685 75.860 116.730 ;
        RECT 80.660 116.670 80.980 116.930 ;
        RECT 95.810 116.870 96.100 116.915 ;
        RECT 98.130 116.870 98.345 117.025 ;
        RECT 95.810 116.730 98.345 116.870 ;
        RECT 95.810 116.685 96.100 116.730 ;
        RECT 98.600 116.670 98.920 116.930 ;
        RECT 99.075 116.870 99.365 116.915 ;
        RECT 100.530 116.870 100.670 117.410 ;
        RECT 101.375 117.365 101.665 117.410 ;
        RECT 109.655 117.550 109.945 117.595 ;
        RECT 111.020 117.550 111.340 117.610 ;
        RECT 109.655 117.410 111.340 117.550 ;
        RECT 109.655 117.365 109.945 117.410 ;
        RECT 111.020 117.350 111.340 117.410 ;
        RECT 99.075 116.730 100.670 116.870 ;
        RECT 101.820 116.870 102.140 116.930 ;
        RECT 102.295 116.870 102.585 116.915 ;
        RECT 101.820 116.730 102.585 116.870 ;
        RECT 99.075 116.685 99.365 116.730 ;
        RECT 101.820 116.670 102.140 116.730 ;
        RECT 102.295 116.685 102.585 116.730 ;
        RECT 108.260 116.670 108.580 116.930 ;
        RECT 108.735 116.870 109.025 116.915 ;
        RECT 110.560 116.870 110.880 116.930 ;
        RECT 108.735 116.730 110.880 116.870 ;
        RECT 108.735 116.685 109.025 116.730 ;
        RECT 110.560 116.670 110.880 116.730 ;
        RECT 113.320 116.870 113.640 116.930 ;
        RECT 119.315 116.870 119.605 116.915 ;
        RECT 120.220 116.870 120.540 116.930 ;
        RECT 113.320 116.730 120.540 116.870 ;
        RECT 113.320 116.670 113.640 116.730 ;
        RECT 119.315 116.685 119.605 116.730 ;
        RECT 120.220 116.670 120.540 116.730 ;
        RECT 50.760 116.330 51.080 116.590 ;
        RECT 56.295 116.530 56.585 116.575 ;
        RECT 52.000 116.390 56.585 116.530 ;
        RECT 52.000 116.190 52.140 116.390 ;
        RECT 56.295 116.345 56.585 116.390 ;
        RECT 63.195 116.530 63.485 116.575 ;
        RECT 65.480 116.530 65.800 116.590 ;
        RECT 63.195 116.390 65.800 116.530 ;
        RECT 63.195 116.345 63.485 116.390 ;
        RECT 65.480 116.330 65.800 116.390 ;
        RECT 71.705 116.530 71.995 116.575 ;
        RECT 74.220 116.530 74.540 116.590 ;
        RECT 71.705 116.390 74.540 116.530 ;
        RECT 71.705 116.345 71.995 116.390 ;
        RECT 74.220 116.330 74.540 116.390 ;
        RECT 77.900 116.530 78.220 116.590 ;
        RECT 78.835 116.530 79.125 116.575 ;
        RECT 77.900 116.390 79.125 116.530 ;
        RECT 77.900 116.330 78.220 116.390 ;
        RECT 78.835 116.345 79.125 116.390 ;
        RECT 82.500 116.530 82.820 116.590 ;
        RECT 84.355 116.530 84.645 116.575 ;
        RECT 87.115 116.530 87.405 116.575 ;
        RECT 98.690 116.530 98.830 116.670 ;
        RECT 82.500 116.390 98.830 116.530 ;
        RECT 100.915 116.530 101.205 116.575 ;
        RECT 102.740 116.530 103.060 116.590 ;
        RECT 100.915 116.390 103.060 116.530 ;
        RECT 82.500 116.330 82.820 116.390 ;
        RECT 84.355 116.345 84.645 116.390 ;
        RECT 87.115 116.345 87.405 116.390 ;
        RECT 100.915 116.345 101.205 116.390 ;
        RECT 102.740 116.330 103.060 116.390 ;
        RECT 118.380 116.530 118.700 116.590 ;
        RECT 118.855 116.530 119.145 116.575 ;
        RECT 118.380 116.390 119.145 116.530 ;
        RECT 118.380 116.330 118.700 116.390 ;
        RECT 118.855 116.345 119.145 116.390 ;
        RECT 49.470 116.050 52.140 116.190 ;
        RECT 75.570 116.190 75.860 116.235 ;
        RECT 78.350 116.190 78.640 116.235 ;
        RECT 80.210 116.190 80.500 116.235 ;
        RECT 75.570 116.050 80.500 116.190 ;
        RECT 28.650 116.005 28.940 116.050 ;
        RECT 31.430 116.005 31.720 116.050 ;
        RECT 33.290 116.005 33.580 116.050 ;
        RECT 41.100 115.990 41.420 116.050 ;
        RECT 75.570 116.005 75.860 116.050 ;
        RECT 78.350 116.005 78.640 116.050 ;
        RECT 80.210 116.005 80.500 116.050 ;
        RECT 95.810 116.190 96.100 116.235 ;
        RECT 98.590 116.190 98.880 116.235 ;
        RECT 100.450 116.190 100.740 116.235 ;
        RECT 107.800 116.190 108.120 116.250 ;
        RECT 95.810 116.050 100.740 116.190 ;
        RECT 95.810 116.005 96.100 116.050 ;
        RECT 98.590 116.005 98.880 116.050 ;
        RECT 100.450 116.005 100.740 116.050 ;
        RECT 105.130 116.050 108.120 116.190 ;
        RECT 35.580 115.650 35.900 115.910 ;
        RECT 39.260 115.850 39.580 115.910 ;
        RECT 40.655 115.850 40.945 115.895 ;
        RECT 39.260 115.710 40.945 115.850 ;
        RECT 39.260 115.650 39.580 115.710 ;
        RECT 40.655 115.665 40.945 115.710 ;
        RECT 54.900 115.650 55.220 115.910 ;
        RECT 89.860 115.650 90.180 115.910 ;
        RECT 99.060 115.850 99.380 115.910 ;
        RECT 105.130 115.850 105.270 116.050 ;
        RECT 107.800 115.990 108.120 116.050 ;
        RECT 99.060 115.710 105.270 115.850 ;
        RECT 105.500 115.850 105.820 115.910 ;
        RECT 107.355 115.850 107.645 115.895 ;
        RECT 105.500 115.710 107.645 115.850 ;
        RECT 99.060 115.650 99.380 115.710 ;
        RECT 105.500 115.650 105.820 115.710 ;
        RECT 107.355 115.665 107.645 115.710 ;
        RECT 9.290 115.030 129.350 115.510 ;
        RECT 11.905 114.830 12.195 114.875 ;
        RECT 17.640 114.830 17.960 114.890 ;
        RECT 11.905 114.690 17.960 114.830 ;
        RECT 11.905 114.645 12.195 114.690 ;
        RECT 17.640 114.630 17.960 114.690 ;
        RECT 22.240 114.830 22.560 114.890 ;
        RECT 23.175 114.830 23.465 114.875 ;
        RECT 22.240 114.690 23.465 114.830 ;
        RECT 22.240 114.630 22.560 114.690 ;
        RECT 23.175 114.645 23.465 114.690 ;
        RECT 28.695 114.830 28.985 114.875 ;
        RECT 29.140 114.830 29.460 114.890 ;
        RECT 28.695 114.690 29.460 114.830 ;
        RECT 28.695 114.645 28.985 114.690 ;
        RECT 29.140 114.630 29.460 114.690 ;
        RECT 31.440 114.630 31.760 114.890 ;
        RECT 41.560 114.630 41.880 114.890 ;
        RECT 61.800 114.875 62.120 114.890 ;
        RECT 61.800 114.645 62.335 114.875 ;
        RECT 76.980 114.830 77.300 114.890 ;
        RECT 78.375 114.830 78.665 114.875 ;
        RECT 76.980 114.690 78.665 114.830 ;
        RECT 61.800 114.630 62.120 114.645 ;
        RECT 76.980 114.630 77.300 114.690 ;
        RECT 78.375 114.645 78.665 114.690 ;
        RECT 92.175 114.830 92.465 114.875 ;
        RECT 92.620 114.830 92.940 114.890 ;
        RECT 92.175 114.690 92.940 114.830 ;
        RECT 92.175 114.645 92.465 114.690 ;
        RECT 92.620 114.630 92.940 114.690 ;
        RECT 95.380 114.630 95.700 114.890 ;
        RECT 107.815 114.830 108.105 114.875 ;
        RECT 108.260 114.830 108.580 114.890 ;
        RECT 107.815 114.690 108.580 114.830 ;
        RECT 107.815 114.645 108.105 114.690 ;
        RECT 108.260 114.630 108.580 114.690 ;
        RECT 114.945 114.830 115.235 114.875 ;
        RECT 117.000 114.830 117.320 114.890 ;
        RECT 114.945 114.690 117.320 114.830 ;
        RECT 114.945 114.645 115.235 114.690 ;
        RECT 15.770 114.490 16.060 114.535 ;
        RECT 18.550 114.490 18.840 114.535 ;
        RECT 20.410 114.490 20.700 114.535 ;
        RECT 15.770 114.350 20.700 114.490 ;
        RECT 15.770 114.305 16.060 114.350 ;
        RECT 18.550 114.305 18.840 114.350 ;
        RECT 20.410 114.305 20.700 114.350 ;
        RECT 36.010 114.490 36.300 114.535 ;
        RECT 38.790 114.490 39.080 114.535 ;
        RECT 40.650 114.490 40.940 114.535 ;
        RECT 36.010 114.350 40.940 114.490 ;
        RECT 36.010 114.305 36.300 114.350 ;
        RECT 38.790 114.305 39.080 114.350 ;
        RECT 40.650 114.305 40.940 114.350 ;
        RECT 56.250 114.490 56.540 114.535 ;
        RECT 59.030 114.490 59.320 114.535 ;
        RECT 60.890 114.490 61.180 114.535 ;
        RECT 56.250 114.350 61.180 114.490 ;
        RECT 56.250 114.305 56.540 114.350 ;
        RECT 59.030 114.305 59.320 114.350 ;
        RECT 60.890 114.305 61.180 114.350 ;
        RECT 65.910 114.490 66.200 114.535 ;
        RECT 68.690 114.490 68.980 114.535 ;
        RECT 70.550 114.490 70.840 114.535 ;
        RECT 80.660 114.490 80.980 114.550 ;
        RECT 65.910 114.350 70.840 114.490 ;
        RECT 65.910 114.305 66.200 114.350 ;
        RECT 68.690 114.305 68.980 114.350 ;
        RECT 70.550 114.305 70.840 114.350 ;
        RECT 71.090 114.350 80.980 114.490 ;
        RECT 20.860 113.950 21.180 114.210 ;
        RECT 21.320 114.150 21.640 114.210 ;
        RECT 32.360 114.150 32.680 114.210 ;
        RECT 21.320 114.010 22.470 114.150 ;
        RECT 21.320 113.950 21.640 114.010 ;
        RECT 22.330 113.855 22.470 114.010 ;
        RECT 29.230 114.010 32.680 114.150 ;
        RECT 29.230 113.870 29.370 114.010 ;
        RECT 32.360 113.950 32.680 114.010 ;
        RECT 39.260 113.950 39.580 114.210 ;
        RECT 41.100 113.950 41.420 114.210 ;
        RECT 42.020 114.150 42.340 114.210 ;
        RECT 44.335 114.150 44.625 114.195 ;
        RECT 48.015 114.150 48.305 114.195 ;
        RECT 42.020 114.010 48.305 114.150 ;
        RECT 42.020 113.950 42.340 114.010 ;
        RECT 44.335 113.965 44.625 114.010 ;
        RECT 48.015 113.965 48.305 114.010 ;
        RECT 48.935 114.150 49.225 114.195 ;
        RECT 51.220 114.150 51.540 114.210 ;
        RECT 52.385 114.150 52.675 114.195 ;
        RECT 48.935 114.010 52.675 114.150 ;
        RECT 48.935 113.965 49.225 114.010 ;
        RECT 51.220 113.950 51.540 114.010 ;
        RECT 52.385 113.965 52.675 114.010 ;
        RECT 54.900 114.150 55.220 114.210 ;
        RECT 59.515 114.150 59.805 114.195 ;
        RECT 54.900 114.010 59.805 114.150 ;
        RECT 54.900 113.950 55.220 114.010 ;
        RECT 59.515 113.965 59.805 114.010 ;
        RECT 61.355 114.150 61.645 114.195 ;
        RECT 62.720 114.150 63.040 114.210 ;
        RECT 61.355 114.010 63.040 114.150 ;
        RECT 61.355 113.965 61.645 114.010 ;
        RECT 62.720 113.950 63.040 114.010 ;
        RECT 66.400 114.150 66.720 114.210 ;
        RECT 71.090 114.195 71.230 114.350 ;
        RECT 80.660 114.290 80.980 114.350 ;
        RECT 82.520 114.490 82.810 114.535 ;
        RECT 84.380 114.490 84.670 114.535 ;
        RECT 87.160 114.490 87.450 114.535 ;
        RECT 82.520 114.350 87.450 114.490 ;
        RECT 82.520 114.305 82.810 114.350 ;
        RECT 84.380 114.305 84.670 114.350 ;
        RECT 87.160 114.305 87.450 114.350 ;
        RECT 93.555 114.490 93.845 114.535 ;
        RECT 96.300 114.490 96.620 114.550 ;
        RECT 115.020 114.490 115.160 114.645 ;
        RECT 117.000 114.630 117.320 114.690 ;
        RECT 93.555 114.350 96.620 114.490 ;
        RECT 93.555 114.305 93.845 114.350 ;
        RECT 96.300 114.290 96.620 114.350 ;
        RECT 105.130 114.350 108.030 114.490 ;
        RECT 69.175 114.150 69.465 114.195 ;
        RECT 66.400 114.010 69.465 114.150 ;
        RECT 66.400 113.950 66.720 114.010 ;
        RECT 69.175 113.965 69.465 114.010 ;
        RECT 71.015 113.965 71.305 114.195 ;
        RECT 73.300 113.950 73.620 114.210 ;
        RECT 74.220 113.950 74.540 114.210 ;
        RECT 86.180 114.150 86.500 114.210 ;
        RECT 89.860 114.150 90.180 114.210 ;
        RECT 105.130 114.195 105.270 114.350 ;
        RECT 107.890 114.210 108.030 114.350 ;
        RECT 114.330 114.350 115.160 114.490 ;
        RECT 118.810 114.490 119.100 114.535 ;
        RECT 121.590 114.490 121.880 114.535 ;
        RECT 123.450 114.490 123.740 114.535 ;
        RECT 118.810 114.350 123.740 114.490 ;
        RECT 78.910 114.010 87.790 114.150 ;
        RECT 15.770 113.810 16.060 113.855 ;
        RECT 19.035 113.810 19.325 113.855 ;
        RECT 15.770 113.670 18.305 113.810 ;
        RECT 15.770 113.625 16.060 113.670 ;
        RECT 13.910 113.470 14.200 113.515 ;
        RECT 16.260 113.470 16.580 113.530 ;
        RECT 18.090 113.515 18.305 113.670 ;
        RECT 19.035 113.670 21.550 113.810 ;
        RECT 19.035 113.625 19.325 113.670 ;
        RECT 17.170 113.470 17.460 113.515 ;
        RECT 13.910 113.330 17.460 113.470 ;
        RECT 13.910 113.285 14.200 113.330 ;
        RECT 16.260 113.270 16.580 113.330 ;
        RECT 17.170 113.285 17.460 113.330 ;
        RECT 18.090 113.470 18.380 113.515 ;
        RECT 19.950 113.470 20.240 113.515 ;
        RECT 18.090 113.330 20.240 113.470 ;
        RECT 18.090 113.285 18.380 113.330 ;
        RECT 19.950 113.285 20.240 113.330 ;
        RECT 21.410 113.175 21.550 113.670 ;
        RECT 22.255 113.625 22.545 113.855 ;
        RECT 24.080 113.610 24.400 113.870 ;
        RECT 29.140 113.610 29.460 113.870 ;
        RECT 30.520 113.610 30.840 113.870 ;
        RECT 36.010 113.810 36.300 113.855 ;
        RECT 36.010 113.670 38.545 113.810 ;
        RECT 36.010 113.625 36.300 113.670 ;
        RECT 34.150 113.470 34.440 113.515 ;
        RECT 35.580 113.470 35.900 113.530 ;
        RECT 38.330 113.515 38.545 113.670 ;
        RECT 46.160 113.610 46.480 113.870 ;
        RECT 47.080 113.810 47.400 113.870 ;
        RECT 49.395 113.810 49.685 113.855 ;
        RECT 47.080 113.670 49.685 113.810 ;
        RECT 47.080 113.610 47.400 113.670 ;
        RECT 49.395 113.625 49.685 113.670 ;
        RECT 56.250 113.810 56.540 113.855 ;
        RECT 65.910 113.810 66.200 113.855 ;
        RECT 71.475 113.810 71.765 113.855 ;
        RECT 56.250 113.670 58.785 113.810 ;
        RECT 56.250 113.625 56.540 113.670 ;
        RECT 58.570 113.515 58.785 113.670 ;
        RECT 65.910 113.670 68.445 113.810 ;
        RECT 65.910 113.625 66.200 113.670 ;
        RECT 37.410 113.470 37.700 113.515 ;
        RECT 34.150 113.330 37.700 113.470 ;
        RECT 34.150 113.285 34.440 113.330 ;
        RECT 35.580 113.270 35.900 113.330 ;
        RECT 37.410 113.285 37.700 113.330 ;
        RECT 38.330 113.470 38.620 113.515 ;
        RECT 40.190 113.470 40.480 113.515 ;
        RECT 38.330 113.330 40.480 113.470 ;
        RECT 38.330 113.285 38.620 113.330 ;
        RECT 40.190 113.285 40.480 113.330 ;
        RECT 46.635 113.470 46.925 113.515 ;
        RECT 54.390 113.470 54.680 113.515 ;
        RECT 57.650 113.470 57.940 113.515 ;
        RECT 46.635 113.330 57.940 113.470 ;
        RECT 46.635 113.285 46.925 113.330 ;
        RECT 54.390 113.285 54.680 113.330 ;
        RECT 57.650 113.285 57.940 113.330 ;
        RECT 58.570 113.470 58.860 113.515 ;
        RECT 60.430 113.470 60.720 113.515 ;
        RECT 58.570 113.330 60.720 113.470 ;
        RECT 58.570 113.285 58.860 113.330 ;
        RECT 60.430 113.285 60.720 113.330 ;
        RECT 64.050 113.470 64.340 113.515 ;
        RECT 65.480 113.470 65.800 113.530 ;
        RECT 68.230 113.515 68.445 113.670 ;
        RECT 71.090 113.670 72.840 113.810 ;
        RECT 67.310 113.470 67.600 113.515 ;
        RECT 64.050 113.330 67.600 113.470 ;
        RECT 64.050 113.285 64.340 113.330 ;
        RECT 65.480 113.270 65.800 113.330 ;
        RECT 67.310 113.285 67.600 113.330 ;
        RECT 68.230 113.470 68.520 113.515 ;
        RECT 70.090 113.470 70.380 113.515 ;
        RECT 68.230 113.330 70.380 113.470 ;
        RECT 68.230 113.285 68.520 113.330 ;
        RECT 70.090 113.285 70.380 113.330 ;
        RECT 21.335 112.945 21.625 113.175 ;
        RECT 32.145 113.130 32.435 113.175 ;
        RECT 32.820 113.130 33.140 113.190 ;
        RECT 43.415 113.130 43.705 113.175 ;
        RECT 32.145 112.990 43.705 113.130 ;
        RECT 32.145 112.945 32.435 112.990 ;
        RECT 32.820 112.930 33.140 112.990 ;
        RECT 43.415 112.945 43.705 112.990 ;
        RECT 43.875 113.130 44.165 113.175 ;
        RECT 47.080 113.130 47.400 113.190 ;
        RECT 43.875 112.990 47.400 113.130 ;
        RECT 43.875 112.945 44.165 112.990 ;
        RECT 47.080 112.930 47.400 112.990 ;
        RECT 50.760 113.130 51.080 113.190 ;
        RECT 51.235 113.130 51.525 113.175 ;
        RECT 50.760 112.990 51.525 113.130 ;
        RECT 50.760 112.930 51.080 112.990 ;
        RECT 51.235 112.945 51.525 112.990 ;
        RECT 58.120 113.130 58.440 113.190 ;
        RECT 71.090 113.130 71.230 113.670 ;
        RECT 71.475 113.625 71.765 113.670 ;
        RECT 72.700 113.470 72.840 113.670 ;
        RECT 74.680 113.610 75.000 113.870 ;
        RECT 78.910 113.855 79.050 114.010 ;
        RECT 86.180 113.950 86.500 114.010 ;
        RECT 78.835 113.810 79.125 113.855 ;
        RECT 76.150 113.670 79.125 113.810 ;
        RECT 76.150 113.470 76.290 113.670 ;
        RECT 78.835 113.625 79.125 113.670 ;
        RECT 80.215 113.625 80.505 113.855 ;
        RECT 80.660 113.810 80.980 113.870 ;
        RECT 82.055 113.810 82.345 113.855 ;
        RECT 83.420 113.810 83.740 113.870 ;
        RECT 80.660 113.670 83.740 113.810 ;
        RECT 80.290 113.470 80.430 113.625 ;
        RECT 80.660 113.610 80.980 113.670 ;
        RECT 82.055 113.625 82.345 113.670 ;
        RECT 83.420 113.610 83.740 113.670 ;
        RECT 83.880 113.610 84.200 113.870 ;
        RECT 87.160 113.810 87.450 113.855 ;
        RECT 84.915 113.670 87.450 113.810 ;
        RECT 87.650 113.810 87.790 114.010 ;
        RECT 89.860 114.010 94.690 114.150 ;
        RECT 89.860 113.950 90.180 114.010 ;
        RECT 94.550 113.855 94.690 114.010 ;
        RECT 105.055 113.965 105.345 114.195 ;
        RECT 107.800 114.150 108.120 114.210 ;
        RECT 111.035 114.150 111.325 114.195 ;
        RECT 113.320 114.150 113.640 114.210 ;
        RECT 107.800 114.010 111.325 114.150 ;
        RECT 107.800 113.950 108.120 114.010 ;
        RECT 111.035 113.965 111.325 114.010 ;
        RECT 112.030 114.010 113.640 114.150 ;
        RECT 92.635 113.810 92.925 113.855 ;
        RECT 93.095 113.810 93.385 113.855 ;
        RECT 87.650 113.670 93.385 113.810 ;
        RECT 84.915 113.515 85.130 113.670 ;
        RECT 87.160 113.625 87.450 113.670 ;
        RECT 92.635 113.625 92.925 113.670 ;
        RECT 93.095 113.625 93.385 113.670 ;
        RECT 94.475 113.625 94.765 113.855 ;
        RECT 107.340 113.610 107.660 113.870 ;
        RECT 109.195 113.810 109.485 113.855 ;
        RECT 112.030 113.810 112.170 114.010 ;
        RECT 113.320 113.950 113.640 114.010 ;
        RECT 109.195 113.670 112.170 113.810 ;
        RECT 112.415 113.810 112.705 113.855 ;
        RECT 114.330 113.810 114.470 114.350 ;
        RECT 118.810 114.305 119.100 114.350 ;
        RECT 121.590 114.305 121.880 114.350 ;
        RECT 123.450 114.305 123.740 114.350 ;
        RECT 122.060 113.950 122.380 114.210 ;
        RECT 123.915 114.150 124.205 114.195 ;
        RECT 126.660 114.150 126.980 114.210 ;
        RECT 123.915 114.010 126.980 114.150 ;
        RECT 123.915 113.965 124.205 114.010 ;
        RECT 112.415 113.670 114.470 113.810 ;
        RECT 118.810 113.810 119.100 113.855 ;
        RECT 121.600 113.810 121.920 113.870 ;
        RECT 123.990 113.810 124.130 113.965 ;
        RECT 126.660 113.950 126.980 114.010 ;
        RECT 118.810 113.670 121.345 113.810 ;
        RECT 109.195 113.625 109.485 113.670 ;
        RECT 112.415 113.625 112.705 113.670 ;
        RECT 118.810 113.625 119.100 113.670 ;
        RECT 72.700 113.330 76.290 113.470 ;
        RECT 76.610 113.330 80.430 113.470 ;
        RECT 82.980 113.470 83.270 113.515 ;
        RECT 84.840 113.470 85.130 113.515 ;
        RECT 82.980 113.330 85.130 113.470 ;
        RECT 58.120 112.990 71.230 113.130 ;
        RECT 58.120 112.930 58.440 112.990 ;
        RECT 71.920 112.930 72.240 113.190 ;
        RECT 76.610 113.175 76.750 113.330 ;
        RECT 82.980 113.285 83.270 113.330 ;
        RECT 84.840 113.285 85.130 113.330 ;
        RECT 85.760 113.470 86.050 113.515 ;
        RECT 86.640 113.470 86.960 113.530 ;
        RECT 89.020 113.470 89.310 113.515 ;
        RECT 91.025 113.470 91.315 113.515 ;
        RECT 105.515 113.470 105.805 113.515 ;
        RECT 85.760 113.330 89.310 113.470 ;
        RECT 85.760 113.285 86.050 113.330 ;
        RECT 86.640 113.270 86.960 113.330 ;
        RECT 89.020 113.285 89.310 113.330 ;
        RECT 89.490 113.330 105.805 113.470 ;
        RECT 76.535 112.945 76.825 113.175 ;
        RECT 77.900 113.130 78.220 113.190 ;
        RECT 79.295 113.130 79.585 113.175 ;
        RECT 77.900 112.990 79.585 113.130 ;
        RECT 77.900 112.930 78.220 112.990 ;
        RECT 79.295 112.945 79.585 112.990 ;
        RECT 84.340 113.130 84.660 113.190 ;
        RECT 89.490 113.130 89.630 113.330 ;
        RECT 91.025 113.285 91.315 113.330 ;
        RECT 105.515 113.285 105.805 113.330 ;
        RECT 105.975 113.470 106.265 113.515 ;
        RECT 107.430 113.470 107.570 113.610 ;
        RECT 116.950 113.470 117.240 113.515 ;
        RECT 118.380 113.470 118.700 113.530 ;
        RECT 121.130 113.515 121.345 113.670 ;
        RECT 121.600 113.670 124.130 113.810 ;
        RECT 121.600 113.610 121.920 113.670 ;
        RECT 120.210 113.470 120.500 113.515 ;
        RECT 105.975 113.330 112.170 113.470 ;
        RECT 105.975 113.285 106.265 113.330 ;
        RECT 112.030 113.190 112.170 113.330 ;
        RECT 116.950 113.330 120.500 113.470 ;
        RECT 116.950 113.285 117.240 113.330 ;
        RECT 118.380 113.270 118.700 113.330 ;
        RECT 120.210 113.285 120.500 113.330 ;
        RECT 121.130 113.470 121.420 113.515 ;
        RECT 122.990 113.470 123.280 113.515 ;
        RECT 121.130 113.330 123.280 113.470 ;
        RECT 121.130 113.285 121.420 113.330 ;
        RECT 122.990 113.285 123.280 113.330 ;
        RECT 84.340 112.990 89.630 113.130 ;
        RECT 107.340 113.130 107.660 113.190 ;
        RECT 108.735 113.130 109.025 113.175 ;
        RECT 107.340 112.990 109.025 113.130 ;
        RECT 84.340 112.930 84.660 112.990 ;
        RECT 107.340 112.930 107.660 112.990 ;
        RECT 108.735 112.945 109.025 112.990 ;
        RECT 111.940 112.930 112.260 113.190 ;
        RECT 114.240 112.930 114.560 113.190 ;
        RECT 9.290 112.310 129.350 112.790 ;
        RECT 16.260 111.910 16.580 112.170 ;
        RECT 45.945 112.110 46.235 112.155 ;
        RECT 47.080 112.110 47.400 112.170 ;
        RECT 45.945 111.970 47.400 112.110 ;
        RECT 45.945 111.925 46.235 111.970 ;
        RECT 47.080 111.910 47.400 111.970 ;
        RECT 68.485 112.110 68.775 112.155 ;
        RECT 74.220 112.110 74.540 112.170 ;
        RECT 68.485 111.970 74.540 112.110 ;
        RECT 68.485 111.925 68.775 111.970 ;
        RECT 74.220 111.910 74.540 111.970 ;
        RECT 83.880 112.110 84.200 112.170 ;
        RECT 84.355 112.110 84.645 112.155 ;
        RECT 83.880 111.970 84.645 112.110 ;
        RECT 83.880 111.910 84.200 111.970 ;
        RECT 84.355 111.925 84.645 111.970 ;
        RECT 86.195 112.110 86.485 112.155 ;
        RECT 86.640 112.110 86.960 112.170 ;
        RECT 86.195 111.970 86.960 112.110 ;
        RECT 86.195 111.925 86.485 111.970 ;
        RECT 86.640 111.910 86.960 111.970 ;
        RECT 111.940 112.110 112.260 112.170 ;
        RECT 112.645 112.110 112.935 112.155 ;
        RECT 111.940 111.970 112.935 112.110 ;
        RECT 111.940 111.910 112.260 111.970 ;
        RECT 112.645 111.925 112.935 111.970 ;
        RECT 120.235 112.110 120.525 112.155 ;
        RECT 122.060 112.110 122.380 112.170 ;
        RECT 120.235 111.970 122.380 112.110 ;
        RECT 120.235 111.925 120.525 111.970 ;
        RECT 122.060 111.910 122.380 111.970 ;
        RECT 48.000 111.815 48.320 111.830 ;
        RECT 47.950 111.770 48.320 111.815 ;
        RECT 51.210 111.770 51.500 111.815 ;
        RECT 47.950 111.630 51.500 111.770 ;
        RECT 47.950 111.585 48.320 111.630 ;
        RECT 51.210 111.585 51.500 111.630 ;
        RECT 52.130 111.770 52.420 111.815 ;
        RECT 53.990 111.770 54.280 111.815 ;
        RECT 52.130 111.630 54.280 111.770 ;
        RECT 52.130 111.585 52.420 111.630 ;
        RECT 53.990 111.585 54.280 111.630 ;
        RECT 70.490 111.770 70.780 111.815 ;
        RECT 71.920 111.770 72.240 111.830 ;
        RECT 107.340 111.815 107.660 111.830 ;
        RECT 73.750 111.770 74.040 111.815 ;
        RECT 70.490 111.630 74.040 111.770 ;
        RECT 70.490 111.585 70.780 111.630 ;
        RECT 48.000 111.570 48.320 111.585 ;
        RECT 12.580 111.430 12.900 111.490 ;
        RECT 16.735 111.430 17.025 111.475 ;
        RECT 29.140 111.430 29.460 111.490 ;
        RECT 12.580 111.290 29.460 111.430 ;
        RECT 12.580 111.230 12.900 111.290 ;
        RECT 16.735 111.245 17.025 111.290 ;
        RECT 29.140 111.230 29.460 111.290 ;
        RECT 49.810 111.430 50.100 111.475 ;
        RECT 52.130 111.430 52.345 111.585 ;
        RECT 71.920 111.570 72.240 111.630 ;
        RECT 73.750 111.585 74.040 111.630 ;
        RECT 74.670 111.770 74.960 111.815 ;
        RECT 76.530 111.770 76.820 111.815 ;
        RECT 74.670 111.630 76.820 111.770 ;
        RECT 74.670 111.585 74.960 111.630 ;
        RECT 76.530 111.585 76.820 111.630 ;
        RECT 104.600 111.770 104.890 111.815 ;
        RECT 106.460 111.770 106.750 111.815 ;
        RECT 104.600 111.630 106.750 111.770 ;
        RECT 104.600 111.585 104.890 111.630 ;
        RECT 106.460 111.585 106.750 111.630 ;
        RECT 49.810 111.290 52.345 111.430 ;
        RECT 49.810 111.245 50.100 111.290 ;
        RECT 53.060 111.230 53.380 111.490 ;
        RECT 54.915 111.430 55.205 111.475 ;
        RECT 60.420 111.430 60.740 111.490 ;
        RECT 62.720 111.430 63.040 111.490 ;
        RECT 54.915 111.290 63.040 111.430 ;
        RECT 54.915 111.245 55.205 111.290 ;
        RECT 51.680 111.090 52.000 111.150 ;
        RECT 54.990 111.090 55.130 111.245 ;
        RECT 60.420 111.230 60.740 111.290 ;
        RECT 62.720 111.230 63.040 111.290 ;
        RECT 72.350 111.430 72.640 111.475 ;
        RECT 74.670 111.430 74.885 111.585 ;
        RECT 72.350 111.290 74.885 111.430 ;
        RECT 75.615 111.430 75.905 111.475 ;
        RECT 77.900 111.430 78.220 111.490 ;
        RECT 75.615 111.290 78.220 111.430 ;
        RECT 72.350 111.245 72.640 111.290 ;
        RECT 75.615 111.245 75.905 111.290 ;
        RECT 77.900 111.230 78.220 111.290 ;
        RECT 85.260 111.230 85.580 111.490 ;
        RECT 86.180 111.430 86.500 111.490 ;
        RECT 86.655 111.430 86.945 111.475 ;
        RECT 86.180 111.290 86.945 111.430 ;
        RECT 86.180 111.230 86.500 111.290 ;
        RECT 86.655 111.245 86.945 111.290 ;
        RECT 102.740 111.430 103.060 111.490 ;
        RECT 103.675 111.430 103.965 111.475 ;
        RECT 102.740 111.290 103.965 111.430 ;
        RECT 102.740 111.230 103.060 111.290 ;
        RECT 103.675 111.245 103.965 111.290 ;
        RECT 105.500 111.230 105.820 111.490 ;
        RECT 106.535 111.430 106.750 111.585 ;
        RECT 107.340 111.770 107.670 111.815 ;
        RECT 110.640 111.770 110.930 111.815 ;
        RECT 107.340 111.630 110.930 111.770 ;
        RECT 107.340 111.585 107.670 111.630 ;
        RECT 110.640 111.585 110.930 111.630 ;
        RECT 107.340 111.570 107.660 111.585 ;
        RECT 108.780 111.430 109.070 111.475 ;
        RECT 106.535 111.290 109.070 111.430 ;
        RECT 108.780 111.245 109.070 111.290 ;
        RECT 114.240 111.430 114.560 111.490 ;
        RECT 119.315 111.430 119.605 111.475 ;
        RECT 114.240 111.290 119.605 111.430 ;
        RECT 114.240 111.230 114.560 111.290 ;
        RECT 119.315 111.245 119.605 111.290 ;
        RECT 51.680 110.950 55.130 111.090 ;
        RECT 77.455 111.090 77.745 111.135 ;
        RECT 83.420 111.090 83.740 111.150 ;
        RECT 77.455 110.950 83.740 111.090 ;
        RECT 51.680 110.890 52.000 110.950 ;
        RECT 77.455 110.905 77.745 110.950 ;
        RECT 83.420 110.890 83.740 110.950 ;
        RECT 49.810 110.750 50.100 110.795 ;
        RECT 52.590 110.750 52.880 110.795 ;
        RECT 54.450 110.750 54.740 110.795 ;
        RECT 49.810 110.610 54.740 110.750 ;
        RECT 49.810 110.565 50.100 110.610 ;
        RECT 52.590 110.565 52.880 110.610 ;
        RECT 54.450 110.565 54.740 110.610 ;
        RECT 72.350 110.750 72.640 110.795 ;
        RECT 75.130 110.750 75.420 110.795 ;
        RECT 76.990 110.750 77.280 110.795 ;
        RECT 72.350 110.610 77.280 110.750 ;
        RECT 72.350 110.565 72.640 110.610 ;
        RECT 75.130 110.565 75.420 110.610 ;
        RECT 76.990 110.565 77.280 110.610 ;
        RECT 104.140 110.750 104.430 110.795 ;
        RECT 106.000 110.750 106.290 110.795 ;
        RECT 108.780 110.750 109.070 110.795 ;
        RECT 104.140 110.610 109.070 110.750 ;
        RECT 104.140 110.565 104.430 110.610 ;
        RECT 106.000 110.565 106.290 110.610 ;
        RECT 108.780 110.565 109.070 110.610 ;
        RECT 9.290 109.590 129.350 110.070 ;
        RECT 53.060 109.190 53.380 109.450 ;
        RECT 13.615 109.050 13.905 109.095 ;
        RECT 16.735 109.050 17.025 109.095 ;
        RECT 18.625 109.050 18.915 109.095 ;
        RECT 13.615 108.910 18.915 109.050 ;
        RECT 13.615 108.865 13.905 108.910 ;
        RECT 16.735 108.865 17.025 108.910 ;
        RECT 18.625 108.865 18.915 108.910 ;
        RECT 19.495 108.710 19.785 108.755 ;
        RECT 20.860 108.710 21.180 108.770 ;
        RECT 19.495 108.570 21.180 108.710 ;
        RECT 19.495 108.525 19.785 108.570 ;
        RECT 20.860 108.510 21.180 108.570 ;
        RECT 12.535 108.075 12.825 108.390 ;
        RECT 13.615 108.370 13.905 108.415 ;
        RECT 17.195 108.370 17.485 108.415 ;
        RECT 19.030 108.370 19.320 108.415 ;
        RECT 13.615 108.230 19.320 108.370 ;
        RECT 13.615 108.185 13.905 108.230 ;
        RECT 17.195 108.185 17.485 108.230 ;
        RECT 19.030 108.185 19.320 108.230 ;
        RECT 21.780 108.370 22.100 108.430 ;
        RECT 22.255 108.370 22.545 108.415 ;
        RECT 21.780 108.230 22.545 108.370 ;
        RECT 21.780 108.170 22.100 108.230 ;
        RECT 22.255 108.185 22.545 108.230 ;
        RECT 27.760 108.370 28.080 108.430 ;
        RECT 28.235 108.370 28.525 108.415 ;
        RECT 27.760 108.230 28.525 108.370 ;
        RECT 27.760 108.170 28.080 108.230 ;
        RECT 28.235 108.185 28.525 108.230 ;
        RECT 50.760 108.370 51.080 108.430 ;
        RECT 52.155 108.370 52.445 108.415 ;
        RECT 50.760 108.230 52.445 108.370 ;
        RECT 50.760 108.170 51.080 108.230 ;
        RECT 52.155 108.185 52.445 108.230 ;
        RECT 61.340 108.370 61.660 108.430 ;
        RECT 80.215 108.370 80.505 108.415 ;
        RECT 61.340 108.230 80.505 108.370 ;
        RECT 61.340 108.170 61.660 108.230 ;
        RECT 80.215 108.185 80.505 108.230 ;
        RECT 97.220 108.370 97.540 108.430 ;
        RECT 98.615 108.370 98.905 108.415 ;
        RECT 97.220 108.230 98.905 108.370 ;
        RECT 97.220 108.170 97.540 108.230 ;
        RECT 98.615 108.185 98.905 108.230 ;
        RECT 102.280 108.370 102.600 108.430 ;
        RECT 122.535 108.370 122.825 108.415 ;
        RECT 102.280 108.230 122.825 108.370 ;
        RECT 102.280 108.170 102.600 108.230 ;
        RECT 122.535 108.185 122.825 108.230 ;
        RECT 122.980 108.370 123.300 108.430 ;
        RECT 123.915 108.370 124.205 108.415 ;
        RECT 122.980 108.230 124.205 108.370 ;
        RECT 122.980 108.170 123.300 108.230 ;
        RECT 123.915 108.185 124.205 108.230 ;
        RECT 15.800 108.075 16.120 108.090 ;
        RECT 12.235 108.030 12.825 108.075 ;
        RECT 15.475 108.030 16.125 108.075 ;
        RECT 12.235 107.890 16.125 108.030 ;
        RECT 12.235 107.845 12.525 107.890 ;
        RECT 15.475 107.845 16.125 107.890 ;
        RECT 18.115 108.030 18.405 108.075 ;
        RECT 18.115 107.890 21.550 108.030 ;
        RECT 18.115 107.845 18.405 107.890 ;
        RECT 15.800 107.830 16.120 107.845 ;
        RECT 7.980 107.690 8.300 107.750 ;
        RECT 21.410 107.735 21.550 107.890 ;
        RECT 81.580 107.830 81.900 108.090 ;
        RECT 10.755 107.690 11.045 107.735 ;
        RECT 7.980 107.550 11.045 107.690 ;
        RECT 7.980 107.490 8.300 107.550 ;
        RECT 10.755 107.505 11.045 107.550 ;
        RECT 21.335 107.505 21.625 107.735 ;
        RECT 23.160 107.690 23.480 107.750 ;
        RECT 27.315 107.690 27.605 107.735 ;
        RECT 23.160 107.550 27.605 107.690 ;
        RECT 23.160 107.490 23.480 107.550 ;
        RECT 27.315 107.505 27.605 107.550 ;
        RECT 99.520 107.490 99.840 107.750 ;
        RECT 120.220 107.690 120.540 107.750 ;
        RECT 121.615 107.690 121.905 107.735 ;
        RECT 120.220 107.550 121.905 107.690 ;
        RECT 120.220 107.490 120.540 107.550 ;
        RECT 121.615 107.505 121.905 107.550 ;
        RECT 122.060 107.690 122.380 107.750 ;
        RECT 122.995 107.690 123.285 107.735 ;
        RECT 122.060 107.550 123.285 107.690 ;
        RECT 122.060 107.490 122.380 107.550 ;
        RECT 122.995 107.505 123.285 107.550 ;
        RECT 9.290 106.870 129.350 107.350 ;
        RECT 42.480 106.670 42.800 106.730 ;
        RECT 44.320 106.670 44.640 106.730 ;
        RECT 70.080 106.670 70.400 106.730 ;
        RECT 73.775 106.670 74.065 106.715 ;
        RECT 42.480 106.530 44.090 106.670 ;
        RECT 42.480 106.470 42.800 106.530 ;
        RECT 14.895 106.330 15.185 106.375 ;
        RECT 17.295 106.330 17.585 106.375 ;
        RECT 20.535 106.330 21.185 106.375 ;
        RECT 14.895 106.190 21.185 106.330 ;
        RECT 14.895 106.145 15.185 106.190 ;
        RECT 17.295 106.145 17.885 106.190 ;
        RECT 20.535 106.145 21.185 106.190 ;
        RECT 15.355 105.805 15.645 106.035 ;
        RECT 17.595 105.830 17.885 106.145 ;
        RECT 23.160 106.130 23.480 106.390 ;
        RECT 39.720 106.330 40.040 106.390 ;
        RECT 43.950 106.330 44.090 106.530 ;
        RECT 44.320 106.530 64.330 106.670 ;
        RECT 44.320 106.470 44.640 106.530 ;
        RECT 39.720 106.190 42.710 106.330 ;
        RECT 43.950 106.190 52.140 106.330 ;
        RECT 39.720 106.130 40.040 106.190 ;
        RECT 18.675 105.990 18.965 106.035 ;
        RECT 22.255 105.990 22.545 106.035 ;
        RECT 24.090 105.990 24.380 106.035 ;
        RECT 18.675 105.850 24.380 105.990 ;
        RECT 18.675 105.805 18.965 105.850 ;
        RECT 22.255 105.805 22.545 105.850 ;
        RECT 24.090 105.805 24.380 105.850 ;
        RECT 27.300 105.990 27.620 106.050 ;
        RECT 28.235 105.990 28.525 106.035 ;
        RECT 27.300 105.850 28.525 105.990 ;
        RECT 15.430 105.650 15.570 105.805 ;
        RECT 27.300 105.790 27.620 105.850 ;
        RECT 28.235 105.805 28.525 105.850 ;
        RECT 28.680 105.990 29.000 106.050 ;
        RECT 32.375 105.990 32.665 106.035 ;
        RECT 28.680 105.850 32.665 105.990 ;
        RECT 28.680 105.790 29.000 105.850 ;
        RECT 32.375 105.805 32.665 105.850 ;
        RECT 37.880 105.790 38.200 106.050 ;
        RECT 42.570 106.035 42.710 106.190 ;
        RECT 41.115 105.805 41.405 106.035 ;
        RECT 42.495 105.805 42.785 106.035 ;
        RECT 43.400 105.990 43.720 106.050 ;
        RECT 45.255 105.990 45.545 106.035 ;
        RECT 43.400 105.850 45.545 105.990 ;
        RECT 52.000 105.990 52.140 106.190 ;
        RECT 55.375 105.990 55.665 106.035 ;
        RECT 52.000 105.850 55.665 105.990 ;
        RECT 21.320 105.650 21.640 105.710 ;
        RECT 24.555 105.650 24.845 105.695 ;
        RECT 15.430 105.510 17.870 105.650 ;
        RECT 17.730 105.370 17.870 105.510 ;
        RECT 21.320 105.510 24.845 105.650 ;
        RECT 21.320 105.450 21.640 105.510 ;
        RECT 24.555 105.465 24.845 105.510 ;
        RECT 31.900 105.650 32.220 105.710 ;
        RECT 41.190 105.650 41.330 105.805 ;
        RECT 43.400 105.790 43.720 105.850 ;
        RECT 45.255 105.805 45.545 105.850 ;
        RECT 55.375 105.805 55.665 105.850 ;
        RECT 57.200 105.990 57.520 106.050 ;
        RECT 57.675 105.990 57.965 106.035 ;
        RECT 57.200 105.850 57.965 105.990 ;
        RECT 57.200 105.790 57.520 105.850 ;
        RECT 57.675 105.805 57.965 105.850 ;
        RECT 61.340 105.790 61.660 106.050 ;
        RECT 64.190 106.035 64.330 106.530 ;
        RECT 70.080 106.530 74.065 106.670 ;
        RECT 70.080 106.470 70.400 106.530 ;
        RECT 73.775 106.485 74.065 106.530 ;
        RECT 75.600 106.670 75.920 106.730 ;
        RECT 117.935 106.670 118.225 106.715 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 75.600 106.530 91.930 106.670 ;
        RECT 75.600 106.470 75.920 106.530 ;
        RECT 75.140 106.330 75.460 106.390 ;
        RECT 76.175 106.330 76.465 106.375 ;
        RECT 79.415 106.330 80.065 106.375 ;
        RECT 75.140 106.190 80.065 106.330 ;
        RECT 75.140 106.130 75.460 106.190 ;
        RECT 76.175 106.145 76.765 106.190 ;
        RECT 79.415 106.145 80.065 106.190 ;
        RECT 64.115 105.805 64.405 106.035 ;
        RECT 74.220 105.790 74.540 106.050 ;
        RECT 76.475 105.830 76.765 106.145 ;
        RECT 91.790 106.035 91.930 106.530 ;
        RECT 117.935 106.530 122.290 106.670 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 117.935 106.485 118.225 106.530 ;
        RECT 98.140 106.375 98.460 106.390 ;
        RECT 95.035 106.330 95.325 106.375 ;
        RECT 98.140 106.330 98.925 106.375 ;
        RECT 95.035 106.190 98.925 106.330 ;
        RECT 95.035 106.145 95.625 106.190 ;
        RECT 77.555 105.990 77.845 106.035 ;
        RECT 81.135 105.990 81.425 106.035 ;
        RECT 82.970 105.990 83.260 106.035 ;
        RECT 77.555 105.850 83.260 105.990 ;
        RECT 77.555 105.805 77.845 105.850 ;
        RECT 81.135 105.805 81.425 105.850 ;
        RECT 82.970 105.805 83.260 105.850 ;
        RECT 91.715 105.805 92.005 106.035 ;
        RECT 95.335 105.830 95.625 106.145 ;
        RECT 98.140 106.145 98.925 106.190 ;
        RECT 99.520 106.330 99.840 106.390 ;
        RECT 100.915 106.330 101.205 106.375 ;
        RECT 99.520 106.190 101.205 106.330 ;
        RECT 98.140 106.130 98.460 106.145 ;
        RECT 99.520 106.130 99.840 106.190 ;
        RECT 100.915 106.145 101.205 106.190 ;
        RECT 106.880 106.330 107.200 106.390 ;
        RECT 120.235 106.330 120.525 106.375 ;
        RECT 121.600 106.330 121.920 106.390 ;
        RECT 106.880 106.190 108.950 106.330 ;
        RECT 106.880 106.130 107.200 106.190 ;
        RECT 96.415 105.990 96.705 106.035 ;
        RECT 99.995 105.990 100.285 106.035 ;
        RECT 101.830 105.990 102.120 106.035 ;
        RECT 96.415 105.850 102.120 105.990 ;
        RECT 96.415 105.805 96.705 105.850 ;
        RECT 99.995 105.805 100.285 105.850 ;
        RECT 101.830 105.805 102.120 105.850 ;
        RECT 102.295 105.990 102.585 106.035 ;
        RECT 102.740 105.990 103.060 106.050 ;
        RECT 102.295 105.850 103.060 105.990 ;
        RECT 102.295 105.805 102.585 105.850 ;
        RECT 102.740 105.790 103.060 105.850 ;
        RECT 104.120 105.990 104.440 106.050 ;
        RECT 108.810 106.035 108.950 106.190 ;
        RECT 120.235 106.190 121.920 106.330 ;
        RECT 122.150 106.330 122.290 106.530 ;
        RECT 122.515 106.330 123.165 106.375 ;
        RECT 126.115 106.330 126.405 106.375 ;
        RECT 122.150 106.190 126.405 106.330 ;
        RECT 120.235 106.145 120.525 106.190 ;
        RECT 121.600 106.130 121.920 106.190 ;
        RECT 122.515 106.145 123.165 106.190 ;
        RECT 125.815 106.145 126.405 106.190 ;
        RECT 105.055 105.990 105.345 106.035 ;
        RECT 104.120 105.850 105.345 105.990 ;
        RECT 104.120 105.790 104.440 105.850 ;
        RECT 105.055 105.805 105.345 105.850 ;
        RECT 107.355 105.805 107.645 106.035 ;
        RECT 108.735 105.805 109.025 106.035 ;
        RECT 112.860 105.990 113.180 106.050 ;
        RECT 113.795 105.990 114.085 106.035 ;
        RECT 112.860 105.850 114.085 105.990 ;
        RECT 44.320 105.650 44.640 105.710 ;
        RECT 54.900 105.650 55.220 105.710 ;
        RECT 59.975 105.650 60.265 105.695 ;
        RECT 31.900 105.510 60.265 105.650 ;
        RECT 31.900 105.450 32.220 105.510 ;
        RECT 44.320 105.450 44.640 105.510 ;
        RECT 54.900 105.450 55.220 105.510 ;
        RECT 59.975 105.465 60.265 105.510 ;
        RECT 82.040 105.450 82.360 105.710 ;
        RECT 83.420 105.450 83.740 105.710 ;
        RECT 17.640 105.110 17.960 105.370 ;
        RECT 18.675 105.310 18.965 105.355 ;
        RECT 21.795 105.310 22.085 105.355 ;
        RECT 23.685 105.310 23.975 105.355 ;
        RECT 18.675 105.170 23.975 105.310 ;
        RECT 18.675 105.125 18.965 105.170 ;
        RECT 21.795 105.125 22.085 105.170 ;
        RECT 23.685 105.125 23.975 105.170 ;
        RECT 77.555 105.310 77.845 105.355 ;
        RECT 80.675 105.310 80.965 105.355 ;
        RECT 82.565 105.310 82.855 105.355 ;
        RECT 77.555 105.170 82.855 105.310 ;
        RECT 77.555 105.125 77.845 105.170 ;
        RECT 80.675 105.125 80.965 105.170 ;
        RECT 82.565 105.125 82.855 105.170 ;
        RECT 96.415 105.310 96.705 105.355 ;
        RECT 99.535 105.310 99.825 105.355 ;
        RECT 101.425 105.310 101.715 105.355 ;
        RECT 107.430 105.310 107.570 105.805 ;
        RECT 112.860 105.790 113.180 105.850 ;
        RECT 113.795 105.805 114.085 105.850 ;
        RECT 117.460 105.790 117.780 106.050 ;
        RECT 119.320 105.990 119.610 106.035 ;
        RECT 121.155 105.990 121.445 106.035 ;
        RECT 124.735 105.990 125.025 106.035 ;
        RECT 119.320 105.850 125.025 105.990 ;
        RECT 119.320 105.805 119.610 105.850 ;
        RECT 121.155 105.805 121.445 105.850 ;
        RECT 124.735 105.805 125.025 105.850 ;
        RECT 125.815 105.830 126.105 106.145 ;
        RECT 107.800 105.650 108.120 105.710 ;
        RECT 118.840 105.650 119.160 105.710 ;
        RECT 120.680 105.650 121.000 105.710 ;
        RECT 107.800 105.510 121.000 105.650 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 107.800 105.450 108.120 105.510 ;
        RECT 118.840 105.450 119.160 105.510 ;
        RECT 120.680 105.450 121.000 105.510 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 117.460 105.310 117.780 105.370 ;
        RECT 96.415 105.170 101.715 105.310 ;
        RECT 96.415 105.125 96.705 105.170 ;
        RECT 99.535 105.125 99.825 105.170 ;
        RECT 101.425 105.125 101.715 105.170 ;
        RECT 102.370 105.170 117.780 105.310 ;
        RECT 14.420 104.970 14.740 105.030 ;
        RECT 15.815 104.970 16.105 105.015 ;
        RECT 14.420 104.830 16.105 104.970 ;
        RECT 14.420 104.770 14.740 104.830 ;
        RECT 15.815 104.785 16.105 104.830 ;
        RECT 24.080 104.970 24.400 105.030 ;
        RECT 27.315 104.970 27.605 105.015 ;
        RECT 24.080 104.830 27.605 104.970 ;
        RECT 24.080 104.770 24.400 104.830 ;
        RECT 27.315 104.785 27.605 104.830 ;
        RECT 27.760 104.970 28.080 105.030 ;
        RECT 31.455 104.970 31.745 105.015 ;
        RECT 27.760 104.830 31.745 104.970 ;
        RECT 27.760 104.770 28.080 104.830 ;
        RECT 31.455 104.785 31.745 104.830 ;
        RECT 36.960 104.770 37.280 105.030 ;
        RECT 40.180 104.970 40.500 105.030 ;
        RECT 40.655 104.970 40.945 105.015 ;
        RECT 40.180 104.830 40.945 104.970 ;
        RECT 40.180 104.770 40.500 104.830 ;
        RECT 40.655 104.785 40.945 104.830 ;
        RECT 41.560 104.770 41.880 105.030 ;
        RECT 46.160 104.770 46.480 105.030 ;
        RECT 47.540 104.970 47.860 105.030 ;
        RECT 54.455 104.970 54.745 105.015 ;
        RECT 47.540 104.830 54.745 104.970 ;
        RECT 47.540 104.770 47.860 104.830 ;
        RECT 54.455 104.785 54.745 104.830 ;
        RECT 58.580 104.770 58.900 105.030 ;
        RECT 61.800 104.970 62.120 105.030 ;
        RECT 63.195 104.970 63.485 105.015 ;
        RECT 61.800 104.830 63.485 104.970 ;
        RECT 61.800 104.770 62.120 104.830 ;
        RECT 63.195 104.785 63.485 104.830 ;
        RECT 74.695 104.970 74.985 105.015 ;
        RECT 76.980 104.970 77.300 105.030 ;
        RECT 74.695 104.830 77.300 104.970 ;
        RECT 74.695 104.785 74.985 104.830 ;
        RECT 76.980 104.770 77.300 104.830 ;
        RECT 92.620 104.770 92.940 105.030 ;
        RECT 93.555 104.970 93.845 105.015 ;
        RECT 97.220 104.970 97.540 105.030 ;
        RECT 93.555 104.830 97.540 104.970 ;
        RECT 93.555 104.785 93.845 104.830 ;
        RECT 97.220 104.770 97.540 104.830 ;
        RECT 101.820 104.970 102.140 105.030 ;
        RECT 102.370 104.970 102.510 105.170 ;
        RECT 117.460 105.110 117.780 105.170 ;
        RECT 119.725 105.310 120.015 105.355 ;
        RECT 121.615 105.310 121.905 105.355 ;
        RECT 124.735 105.310 125.025 105.355 ;
        RECT 119.725 105.170 125.025 105.310 ;
        RECT 119.725 105.125 120.015 105.170 ;
        RECT 121.615 105.125 121.905 105.170 ;
        RECT 124.735 105.125 125.025 105.170 ;
        RECT 101.820 104.830 102.510 104.970 ;
        RECT 101.820 104.770 102.140 104.830 ;
        RECT 105.960 104.770 106.280 105.030 ;
        RECT 107.815 104.970 108.105 105.015 ;
        RECT 108.260 104.970 108.580 105.030 ;
        RECT 107.815 104.830 108.580 104.970 ;
        RECT 107.815 104.785 108.105 104.830 ;
        RECT 108.260 104.770 108.580 104.830 ;
        RECT 109.640 104.770 109.960 105.030 ;
        RECT 114.700 104.770 115.020 105.030 ;
        RECT 127.595 104.970 127.885 105.015 ;
        RECT 130.340 104.970 130.660 105.030 ;
        RECT 127.595 104.830 130.660 104.970 ;
        RECT 127.595 104.785 127.885 104.830 ;
        RECT 130.340 104.770 130.660 104.830 ;
        RECT 9.290 104.150 129.350 104.630 ;
        RECT 15.800 103.750 16.120 104.010 ;
        RECT 21.320 103.950 21.640 104.010 ;
        RECT 38.340 103.950 38.660 104.010 ;
        RECT 21.320 103.810 25.690 103.950 ;
        RECT 21.320 103.750 21.640 103.810 ;
        RECT 19.595 103.610 19.885 103.655 ;
        RECT 22.715 103.610 23.005 103.655 ;
        RECT 24.605 103.610 24.895 103.655 ;
        RECT 19.595 103.470 24.895 103.610 ;
        RECT 19.595 103.425 19.885 103.470 ;
        RECT 22.715 103.425 23.005 103.470 ;
        RECT 24.605 103.425 24.895 103.470 ;
        RECT 16.735 103.270 17.025 103.315 ;
        RECT 20.860 103.270 21.180 103.330 ;
        RECT 16.735 103.130 21.180 103.270 ;
        RECT 16.735 103.085 17.025 103.130 ;
        RECT 20.860 103.070 21.180 103.130 ;
        RECT 24.080 103.070 24.400 103.330 ;
        RECT 25.550 103.315 25.690 103.810 ;
        RECT 33.370 103.810 38.660 103.950 ;
        RECT 33.370 103.315 33.510 103.810 ;
        RECT 38.340 103.750 38.660 103.810 ;
        RECT 42.495 103.950 42.785 103.995 ;
        RECT 46.620 103.950 46.940 104.010 ;
        RECT 42.495 103.810 46.940 103.950 ;
        RECT 42.495 103.765 42.785 103.810 ;
        RECT 46.620 103.750 46.940 103.810 ;
        RECT 75.140 103.750 75.460 104.010 ;
        RECT 76.060 103.950 76.380 104.010 ;
        RECT 80.215 103.950 80.505 103.995 ;
        RECT 82.040 103.950 82.360 104.010 ;
        RECT 76.060 103.810 79.970 103.950 ;
        RECT 76.060 103.750 76.380 103.810 ;
        RECT 34.165 103.610 34.455 103.655 ;
        RECT 36.055 103.610 36.345 103.655 ;
        RECT 39.175 103.610 39.465 103.655 ;
        RECT 41.560 103.610 41.880 103.670 ;
        RECT 34.165 103.470 39.465 103.610 ;
        RECT 34.165 103.425 34.455 103.470 ;
        RECT 36.055 103.425 36.345 103.470 ;
        RECT 39.175 103.425 39.465 103.470 ;
        RECT 40.270 103.470 41.880 103.610 ;
        RECT 25.475 103.270 25.765 103.315 ;
        RECT 33.295 103.270 33.585 103.315 ;
        RECT 25.475 103.130 33.585 103.270 ;
        RECT 25.475 103.085 25.765 103.130 ;
        RECT 33.295 103.085 33.585 103.130 ;
        RECT 34.675 103.270 34.965 103.315 ;
        RECT 40.270 103.270 40.410 103.470 ;
        RECT 41.560 103.410 41.880 103.470 ;
        RECT 45.355 103.610 45.645 103.655 ;
        RECT 48.475 103.610 48.765 103.655 ;
        RECT 50.365 103.610 50.655 103.655 ;
        RECT 45.355 103.470 50.655 103.610 ;
        RECT 45.355 103.425 45.645 103.470 ;
        RECT 48.475 103.425 48.765 103.470 ;
        RECT 50.365 103.425 50.655 103.470 ;
        RECT 61.305 103.610 61.595 103.655 ;
        RECT 63.195 103.610 63.485 103.655 ;
        RECT 66.315 103.610 66.605 103.655 ;
        RECT 61.305 103.470 66.605 103.610 ;
        RECT 61.305 103.425 61.595 103.470 ;
        RECT 63.195 103.425 63.485 103.470 ;
        RECT 66.315 103.425 66.605 103.470 ;
        RECT 76.520 103.610 76.840 103.670 ;
        RECT 79.280 103.610 79.600 103.670 ;
        RECT 76.520 103.470 79.600 103.610 ;
        RECT 79.830 103.610 79.970 103.810 ;
        RECT 80.215 103.810 82.360 103.950 ;
        RECT 80.215 103.765 80.505 103.810 ;
        RECT 82.040 103.750 82.360 103.810 ;
        RECT 87.190 103.810 96.990 103.950 ;
        RECT 85.720 103.610 86.040 103.670 ;
        RECT 79.830 103.470 86.040 103.610 ;
        RECT 76.520 103.410 76.840 103.470 ;
        RECT 79.280 103.410 79.600 103.470 ;
        RECT 85.720 103.410 86.040 103.470 ;
        RECT 34.675 103.130 40.410 103.270 ;
        RECT 40.640 103.270 40.960 103.330 ;
        RECT 42.035 103.270 42.325 103.315 ;
        RECT 40.640 103.130 42.325 103.270 ;
        RECT 34.675 103.085 34.965 103.130 ;
        RECT 40.640 103.070 40.960 103.130 ;
        RECT 42.035 103.085 42.325 103.130 ;
        RECT 46.160 103.270 46.480 103.330 ;
        RECT 49.855 103.270 50.145 103.315 ;
        RECT 60.420 103.270 60.740 103.330 ;
        RECT 46.160 103.130 50.145 103.270 ;
        RECT 46.160 103.070 46.480 103.130 ;
        RECT 49.855 103.085 50.145 103.130 ;
        RECT 52.000 103.130 60.740 103.270 ;
        RECT 16.275 102.930 16.565 102.975 ;
        RECT 16.275 102.790 17.870 102.930 ;
        RECT 16.275 102.745 16.565 102.790 ;
        RECT 17.730 102.310 17.870 102.790 ;
        RECT 18.515 102.635 18.805 102.950 ;
        RECT 19.595 102.930 19.885 102.975 ;
        RECT 23.175 102.930 23.465 102.975 ;
        RECT 25.010 102.930 25.300 102.975 ;
        RECT 19.595 102.790 25.300 102.930 ;
        RECT 19.595 102.745 19.885 102.790 ;
        RECT 23.175 102.745 23.465 102.790 ;
        RECT 25.010 102.745 25.300 102.790 ;
        RECT 27.300 102.730 27.620 102.990 ;
        RECT 27.775 102.930 28.065 102.975 ;
        RECT 31.900 102.930 32.220 102.990 ;
        RECT 27.775 102.790 32.220 102.930 ;
        RECT 27.775 102.745 28.065 102.790 ;
        RECT 18.215 102.590 18.805 102.635 ;
        RECT 20.400 102.590 20.720 102.650 ;
        RECT 21.455 102.590 22.105 102.635 ;
        RECT 27.850 102.590 27.990 102.745 ;
        RECT 31.900 102.730 32.220 102.790 ;
        RECT 33.760 102.930 34.050 102.975 ;
        RECT 35.595 102.930 35.885 102.975 ;
        RECT 39.175 102.930 39.465 102.975 ;
        RECT 33.760 102.790 39.465 102.930 ;
        RECT 33.760 102.745 34.050 102.790 ;
        RECT 35.595 102.745 35.885 102.790 ;
        RECT 39.175 102.745 39.465 102.790 ;
        RECT 40.180 102.950 40.500 102.990 ;
        RECT 40.180 102.730 40.545 102.950 ;
        RECT 40.255 102.635 40.545 102.730 ;
        RECT 44.275 102.635 44.565 102.950 ;
        RECT 45.355 102.930 45.645 102.975 ;
        RECT 48.935 102.930 49.225 102.975 ;
        RECT 50.770 102.930 51.060 102.975 ;
        RECT 45.355 102.790 51.060 102.930 ;
        RECT 45.355 102.745 45.645 102.790 ;
        RECT 48.935 102.745 49.225 102.790 ;
        RECT 50.770 102.745 51.060 102.790 ;
        RECT 51.220 102.930 51.540 102.990 ;
        RECT 52.000 102.930 52.140 103.130 ;
        RECT 60.420 103.070 60.740 103.130 ;
        RECT 61.800 103.070 62.120 103.330 ;
        RECT 66.860 103.270 67.180 103.330 ;
        RECT 69.175 103.270 69.465 103.315 ;
        RECT 81.580 103.270 81.900 103.330 ;
        RECT 87.190 103.270 87.330 103.810 ;
        RECT 91.355 103.610 91.645 103.655 ;
        RECT 94.475 103.610 94.765 103.655 ;
        RECT 96.365 103.610 96.655 103.655 ;
        RECT 91.355 103.470 96.655 103.610 ;
        RECT 96.850 103.610 96.990 103.810 ;
        RECT 98.140 103.750 98.460 104.010 ;
        RECT 107.800 103.950 108.120 104.010 ;
        RECT 104.670 103.810 108.120 103.950 ;
        RECT 101.820 103.610 102.140 103.670 ;
        RECT 96.850 103.470 102.140 103.610 ;
        RECT 91.355 103.425 91.645 103.470 ;
        RECT 94.475 103.425 94.765 103.470 ;
        RECT 96.365 103.425 96.655 103.470 ;
        RECT 101.820 103.410 102.140 103.470 ;
        RECT 66.860 103.130 69.465 103.270 ;
        RECT 66.860 103.070 67.180 103.130 ;
        RECT 69.175 103.085 69.465 103.130 ;
        RECT 75.690 103.130 87.330 103.270 ;
        RECT 51.220 102.790 52.140 102.930 ;
        RECT 51.220 102.730 51.540 102.790 ;
        RECT 54.440 102.730 54.760 102.990 ;
        RECT 54.900 102.930 55.220 102.990 ;
        RECT 75.690 102.975 75.830 103.130 ;
        RECT 57.675 102.930 57.965 102.975 ;
        RECT 59.055 102.930 59.345 102.975 ;
        RECT 54.900 102.790 59.345 102.930 ;
        RECT 54.900 102.730 55.220 102.790 ;
        RECT 57.675 102.745 57.965 102.790 ;
        RECT 59.055 102.745 59.345 102.790 ;
        RECT 59.515 102.930 59.805 102.975 ;
        RECT 60.900 102.930 61.190 102.975 ;
        RECT 62.735 102.930 63.025 102.975 ;
        RECT 66.315 102.930 66.605 102.975 ;
        RECT 59.515 102.790 60.650 102.930 ;
        RECT 59.515 102.745 59.805 102.790 ;
        RECT 18.215 102.450 22.105 102.590 ;
        RECT 18.215 102.405 18.505 102.450 ;
        RECT 20.400 102.390 20.720 102.450 ;
        RECT 21.455 102.405 22.105 102.450 ;
        RECT 22.330 102.450 27.990 102.590 ;
        RECT 36.955 102.590 37.605 102.635 ;
        RECT 40.255 102.590 40.845 102.635 ;
        RECT 36.955 102.450 40.845 102.590 ;
        RECT 17.640 102.250 17.960 102.310 ;
        RECT 22.330 102.250 22.470 102.450 ;
        RECT 36.955 102.405 37.605 102.450 ;
        RECT 40.555 102.405 40.845 102.450 ;
        RECT 43.975 102.590 44.565 102.635 ;
        RECT 44.780 102.590 45.100 102.650 ;
        RECT 47.215 102.590 47.865 102.635 ;
        RECT 43.975 102.450 47.865 102.590 ;
        RECT 60.510 102.590 60.650 102.790 ;
        RECT 60.900 102.790 66.605 102.930 ;
        RECT 60.900 102.745 61.190 102.790 ;
        RECT 62.735 102.745 63.025 102.790 ;
        RECT 66.315 102.745 66.605 102.790 ;
        RECT 67.395 102.635 67.685 102.950 ;
        RECT 75.615 102.745 75.905 102.975 ;
        RECT 76.520 102.730 76.840 102.990 ;
        RECT 77.070 102.975 77.210 103.130 ;
        RECT 81.580 103.070 81.900 103.130 ;
        RECT 76.995 102.745 77.285 102.975 ;
        RECT 77.440 102.930 77.760 102.990 ;
        RECT 77.915 102.930 78.205 102.975 ;
        RECT 77.440 102.790 78.205 102.930 ;
        RECT 77.440 102.730 77.760 102.790 ;
        RECT 77.915 102.745 78.205 102.790 ;
        RECT 79.280 102.730 79.600 102.990 ;
        RECT 84.800 102.730 85.120 102.990 ;
        RECT 85.350 102.975 85.490 103.130 ;
        RECT 85.275 102.745 85.565 102.975 ;
        RECT 85.720 102.730 86.040 102.990 ;
        RECT 87.190 102.975 87.330 103.130 ;
        RECT 88.495 103.270 88.785 103.315 ;
        RECT 90.780 103.270 91.100 103.330 ;
        RECT 88.495 103.130 91.100 103.270 ;
        RECT 88.495 103.085 88.785 103.130 ;
        RECT 90.780 103.070 91.100 103.130 ;
        RECT 92.620 103.270 92.940 103.330 ;
        RECT 95.855 103.270 96.145 103.315 ;
        RECT 102.740 103.270 103.060 103.330 ;
        RECT 104.670 103.315 104.810 103.810 ;
        RECT 107.800 103.750 108.120 103.810 ;
        RECT 105.465 103.610 105.755 103.655 ;
        RECT 107.355 103.610 107.645 103.655 ;
        RECT 110.475 103.610 110.765 103.655 ;
        RECT 105.465 103.470 110.765 103.610 ;
        RECT 105.465 103.425 105.755 103.470 ;
        RECT 107.355 103.425 107.645 103.470 ;
        RECT 110.475 103.425 110.765 103.470 ;
        RECT 119.725 103.610 120.015 103.655 ;
        RECT 121.615 103.610 121.905 103.655 ;
        RECT 124.735 103.610 125.025 103.655 ;
        RECT 119.725 103.470 125.025 103.610 ;
        RECT 119.725 103.425 120.015 103.470 ;
        RECT 121.615 103.425 121.905 103.470 ;
        RECT 124.735 103.425 125.025 103.470 ;
        RECT 125.740 103.610 126.060 103.670 ;
        RECT 127.595 103.610 127.885 103.655 ;
        RECT 125.740 103.470 127.885 103.610 ;
        RECT 125.740 103.410 126.060 103.470 ;
        RECT 127.595 103.425 127.885 103.470 ;
        RECT 104.595 103.270 104.885 103.315 ;
        RECT 92.620 103.130 96.145 103.270 ;
        RECT 92.620 103.070 92.940 103.130 ;
        RECT 95.855 103.085 96.145 103.130 ;
        RECT 97.770 103.130 104.885 103.270 ;
        RECT 87.115 102.745 87.405 102.975 ;
        RECT 87.575 102.930 87.865 102.975 ;
        RECT 90.275 102.930 90.565 102.950 ;
        RECT 87.575 102.790 90.565 102.930 ;
        RECT 87.575 102.745 87.865 102.790 ;
        RECT 64.095 102.590 64.745 102.635 ;
        RECT 67.395 102.590 67.985 102.635 ;
        RECT 60.510 102.450 67.985 102.590 ;
        RECT 43.975 102.405 44.265 102.450 ;
        RECT 44.780 102.390 45.100 102.450 ;
        RECT 47.215 102.405 47.865 102.450 ;
        RECT 64.095 102.405 64.745 102.450 ;
        RECT 67.695 102.405 67.985 102.450 ;
        RECT 74.220 102.590 74.540 102.650 ;
        RECT 90.275 102.635 90.565 102.790 ;
        RECT 91.355 102.930 91.645 102.975 ;
        RECT 94.935 102.930 95.225 102.975 ;
        RECT 96.770 102.930 97.060 102.975 ;
        RECT 91.355 102.790 97.060 102.930 ;
        RECT 91.355 102.745 91.645 102.790 ;
        RECT 94.935 102.745 95.225 102.790 ;
        RECT 96.770 102.745 97.060 102.790 ;
        RECT 97.235 102.930 97.525 102.975 ;
        RECT 97.770 102.930 97.910 103.130 ;
        RECT 102.740 103.070 103.060 103.130 ;
        RECT 104.595 103.085 104.885 103.130 ;
        RECT 105.975 103.270 106.265 103.315 ;
        RECT 109.640 103.270 109.960 103.330 ;
        RECT 105.975 103.130 109.960 103.270 ;
        RECT 105.975 103.085 106.265 103.130 ;
        RECT 109.640 103.070 109.960 103.130 ;
        RECT 111.020 103.270 111.340 103.330 ;
        RECT 113.335 103.270 113.625 103.315 ;
        RECT 111.020 103.130 113.625 103.270 ;
        RECT 111.020 103.070 111.340 103.130 ;
        RECT 113.335 103.085 113.625 103.130 ;
        RECT 115.710 103.130 117.690 103.270 ;
        RECT 97.235 102.790 97.910 102.930 ;
        RECT 98.615 102.930 98.905 102.975 ;
        RECT 101.820 102.930 102.140 102.990 ;
        RECT 98.615 102.790 102.140 102.930 ;
        RECT 97.235 102.745 97.525 102.790 ;
        RECT 98.615 102.745 98.905 102.790 ;
        RECT 101.820 102.730 102.140 102.790 ;
        RECT 102.280 102.730 102.600 102.990 ;
        RECT 115.710 102.975 115.850 103.130 ;
        RECT 117.550 102.990 117.690 103.130 ;
        RECT 118.840 103.070 119.160 103.330 ;
        RECT 120.220 103.070 120.540 103.330 ;
        RECT 105.060 102.930 105.350 102.975 ;
        RECT 106.895 102.930 107.185 102.975 ;
        RECT 110.475 102.930 110.765 102.975 ;
        RECT 105.060 102.790 110.765 102.930 ;
        RECT 105.060 102.745 105.350 102.790 ;
        RECT 106.895 102.745 107.185 102.790 ;
        RECT 110.475 102.745 110.765 102.790 ;
        RECT 108.260 102.635 108.580 102.650 ;
        RECT 111.555 102.635 111.845 102.950 ;
        RECT 115.635 102.745 115.925 102.975 ;
        RECT 116.080 102.730 116.400 102.990 ;
        RECT 117.460 102.730 117.780 102.990 ;
        RECT 117.935 102.930 118.225 102.975 ;
        RECT 119.320 102.930 119.610 102.975 ;
        RECT 121.155 102.930 121.445 102.975 ;
        RECT 124.735 102.930 125.025 102.975 ;
        RECT 117.935 102.790 119.070 102.930 ;
        RECT 117.935 102.745 118.225 102.790 ;
        RECT 89.975 102.590 90.565 102.635 ;
        RECT 93.215 102.590 93.865 102.635 ;
        RECT 74.220 102.450 89.630 102.590 ;
        RECT 74.220 102.390 74.540 102.450 ;
        RECT 17.640 102.110 22.470 102.250 ;
        RECT 31.900 102.250 32.220 102.310 ;
        RECT 32.375 102.250 32.665 102.295 ;
        RECT 31.900 102.110 32.665 102.250 ;
        RECT 17.640 102.050 17.960 102.110 ;
        RECT 31.900 102.050 32.220 102.110 ;
        RECT 32.375 102.065 32.665 102.110 ;
        RECT 57.660 102.250 57.980 102.310 ;
        RECT 58.135 102.250 58.425 102.295 ;
        RECT 57.660 102.110 58.425 102.250 ;
        RECT 57.660 102.050 57.980 102.110 ;
        RECT 58.135 102.065 58.425 102.110 ;
        RECT 77.900 102.250 78.220 102.310 ;
        RECT 78.835 102.250 79.125 102.295 ;
        RECT 77.900 102.110 79.125 102.250 ;
        RECT 77.900 102.050 78.220 102.110 ;
        RECT 78.835 102.065 79.125 102.110 ;
        RECT 86.655 102.250 86.945 102.295 ;
        RECT 88.480 102.250 88.800 102.310 ;
        RECT 86.655 102.110 88.800 102.250 ;
        RECT 89.490 102.250 89.630 102.450 ;
        RECT 89.975 102.450 93.865 102.590 ;
        RECT 89.975 102.405 90.265 102.450 ;
        RECT 93.215 102.405 93.865 102.450 ;
        RECT 108.255 102.590 108.905 102.635 ;
        RECT 111.555 102.590 112.145 102.635 ;
        RECT 108.255 102.450 112.145 102.590 ;
        RECT 118.930 102.590 119.070 102.790 ;
        RECT 119.320 102.790 125.025 102.930 ;
        RECT 119.320 102.745 119.610 102.790 ;
        RECT 121.155 102.745 121.445 102.790 ;
        RECT 124.735 102.745 125.025 102.790 ;
        RECT 125.815 102.635 126.105 102.950 ;
        RECT 122.515 102.590 123.165 102.635 ;
        RECT 125.815 102.590 126.405 102.635 ;
        RECT 118.930 102.450 126.405 102.590 ;
        RECT 108.255 102.405 108.905 102.450 ;
        RECT 111.855 102.405 112.145 102.450 ;
        RECT 122.515 102.405 123.165 102.450 ;
        RECT 126.115 102.405 126.405 102.450 ;
        RECT 108.260 102.390 108.580 102.405 ;
        RECT 126.660 102.250 126.980 102.310 ;
        RECT 89.490 102.110 126.980 102.250 ;
        RECT 86.655 102.065 86.945 102.110 ;
        RECT 88.480 102.050 88.800 102.110 ;
        RECT 126.660 102.050 126.980 102.110 ;
        RECT 9.290 101.430 129.350 101.910 ;
        RECT 19.495 101.230 19.785 101.275 ;
        RECT 20.400 101.230 20.720 101.290 ;
        RECT 19.495 101.090 20.720 101.230 ;
        RECT 19.495 101.045 19.785 101.090 ;
        RECT 20.400 101.030 20.720 101.090 ;
        RECT 44.780 101.230 45.100 101.290 ;
        RECT 45.255 101.230 45.545 101.275 ;
        RECT 44.780 101.090 45.545 101.230 ;
        RECT 44.780 101.030 45.100 101.090 ;
        RECT 45.255 101.045 45.545 101.090 ;
        RECT 58.580 101.230 58.900 101.290 ;
        RECT 77.900 101.230 78.220 101.290 ;
        RECT 114.700 101.230 115.020 101.290 ;
        RECT 58.580 101.090 62.950 101.230 ;
        RECT 58.580 101.030 58.900 101.090 ;
        RECT 21.320 100.890 21.640 100.950 ;
        RECT 20.490 100.750 21.640 100.890 ;
        RECT 17.640 100.550 17.960 100.610 ;
        RECT 20.490 100.595 20.630 100.750 ;
        RECT 21.320 100.690 21.640 100.750 ;
        RECT 24.075 100.890 24.725 100.935 ;
        RECT 27.675 100.890 27.965 100.935 ;
        RECT 24.075 100.750 27.965 100.890 ;
        RECT 24.075 100.705 24.725 100.750 ;
        RECT 27.375 100.705 27.965 100.750 ;
        RECT 31.095 100.890 31.385 100.935 ;
        RECT 31.900 100.890 32.220 100.950 ;
        RECT 34.335 100.890 34.985 100.935 ;
        RECT 31.095 100.750 34.985 100.890 ;
        RECT 31.095 100.705 31.685 100.750 ;
        RECT 27.375 100.610 27.665 100.705 ;
        RECT 19.035 100.550 19.325 100.595 ;
        RECT 17.640 100.410 19.325 100.550 ;
        RECT 17.640 100.350 17.960 100.410 ;
        RECT 19.035 100.365 19.325 100.410 ;
        RECT 20.415 100.365 20.705 100.595 ;
        RECT 20.880 100.550 21.170 100.595 ;
        RECT 22.715 100.550 23.005 100.595 ;
        RECT 26.295 100.550 26.585 100.595 ;
        RECT 20.880 100.410 26.585 100.550 ;
        RECT 20.880 100.365 21.170 100.410 ;
        RECT 22.715 100.365 23.005 100.410 ;
        RECT 26.295 100.365 26.585 100.410 ;
        RECT 27.300 100.390 27.665 100.610 ;
        RECT 31.395 100.390 31.685 100.705 ;
        RECT 31.900 100.690 32.220 100.750 ;
        RECT 34.335 100.705 34.985 100.750 ;
        RECT 36.960 100.690 37.280 100.950 ;
        RECT 47.540 100.690 47.860 100.950 ;
        RECT 49.835 100.890 50.485 100.935 ;
        RECT 53.435 100.890 53.725 100.935 ;
        RECT 54.440 100.890 54.760 100.950 ;
        RECT 49.835 100.750 54.760 100.890 ;
        RECT 49.835 100.705 50.485 100.750 ;
        RECT 53.135 100.705 53.725 100.750 ;
        RECT 32.475 100.550 32.765 100.595 ;
        RECT 36.055 100.550 36.345 100.595 ;
        RECT 37.890 100.550 38.180 100.595 ;
        RECT 32.475 100.410 38.180 100.550 ;
        RECT 27.300 100.350 27.620 100.390 ;
        RECT 32.475 100.365 32.765 100.410 ;
        RECT 36.055 100.365 36.345 100.410 ;
        RECT 37.890 100.365 38.180 100.410 ;
        RECT 38.340 100.350 38.660 100.610 ;
        RECT 44.320 100.550 44.640 100.610 ;
        RECT 44.795 100.550 45.085 100.595 ;
        RECT 44.320 100.410 45.085 100.550 ;
        RECT 44.320 100.350 44.640 100.410 ;
        RECT 44.795 100.365 45.085 100.410 ;
        RECT 46.640 100.550 46.930 100.595 ;
        RECT 48.475 100.550 48.765 100.595 ;
        RECT 52.055 100.550 52.345 100.595 ;
        RECT 46.640 100.410 52.345 100.550 ;
        RECT 46.640 100.365 46.930 100.410 ;
        RECT 48.475 100.365 48.765 100.410 ;
        RECT 52.055 100.365 52.345 100.410 ;
        RECT 53.135 100.390 53.425 100.705 ;
        RECT 54.440 100.690 54.760 100.750 ;
        RECT 56.855 100.890 57.145 100.935 ;
        RECT 57.660 100.890 57.980 100.950 ;
        RECT 62.810 100.935 62.950 101.090 ;
        RECT 77.900 101.090 79.050 101.230 ;
        RECT 77.900 101.030 78.220 101.090 ;
        RECT 76.520 100.935 76.840 100.950 ;
        RECT 78.910 100.935 79.050 101.090 ;
        RECT 114.700 101.090 124.130 101.230 ;
        RECT 114.700 101.030 115.020 101.090 ;
        RECT 60.095 100.890 60.745 100.935 ;
        RECT 56.855 100.750 60.745 100.890 ;
        RECT 56.855 100.705 57.445 100.750 ;
        RECT 57.155 100.390 57.445 100.705 ;
        RECT 57.660 100.690 57.980 100.750 ;
        RECT 60.095 100.705 60.745 100.750 ;
        RECT 62.735 100.705 63.025 100.935 ;
        RECT 72.955 100.890 73.245 100.935 ;
        RECT 76.195 100.890 76.845 100.935 ;
        RECT 72.955 100.750 76.845 100.890 ;
        RECT 72.955 100.705 73.545 100.750 ;
        RECT 76.195 100.705 76.845 100.750 ;
        RECT 78.835 100.705 79.125 100.935 ;
        RECT 82.615 100.890 82.905 100.935 ;
        RECT 84.800 100.890 85.120 100.950 ;
        RECT 85.855 100.890 86.505 100.935 ;
        RECT 82.615 100.750 86.505 100.890 ;
        RECT 82.615 100.705 83.205 100.750 ;
        RECT 58.235 100.550 58.525 100.595 ;
        RECT 61.815 100.550 62.105 100.595 ;
        RECT 63.650 100.550 63.940 100.595 ;
        RECT 58.235 100.410 63.940 100.550 ;
        RECT 58.235 100.365 58.525 100.410 ;
        RECT 61.815 100.365 62.105 100.410 ;
        RECT 63.650 100.365 63.940 100.410 ;
        RECT 73.255 100.390 73.545 100.705 ;
        RECT 76.520 100.690 76.840 100.705 ;
        RECT 74.335 100.550 74.625 100.595 ;
        RECT 77.915 100.550 78.205 100.595 ;
        RECT 79.750 100.550 80.040 100.595 ;
        RECT 74.335 100.410 80.040 100.550 ;
        RECT 74.335 100.365 74.625 100.410 ;
        RECT 77.915 100.365 78.205 100.410 ;
        RECT 79.750 100.365 80.040 100.410 ;
        RECT 82.915 100.390 83.205 100.705 ;
        RECT 84.800 100.690 85.120 100.750 ;
        RECT 85.855 100.705 86.505 100.750 ;
        RECT 88.480 100.690 88.800 100.950 ;
        RECT 101.475 100.890 101.765 100.935 ;
        RECT 102.280 100.890 102.600 100.950 ;
        RECT 104.715 100.890 105.365 100.935 ;
        RECT 101.475 100.750 105.365 100.890 ;
        RECT 101.475 100.705 102.065 100.750 ;
        RECT 83.995 100.550 84.285 100.595 ;
        RECT 87.575 100.550 87.865 100.595 ;
        RECT 89.410 100.550 89.700 100.595 ;
        RECT 83.995 100.410 89.700 100.550 ;
        RECT 83.995 100.365 84.285 100.410 ;
        RECT 87.575 100.365 87.865 100.410 ;
        RECT 89.410 100.365 89.700 100.410 ;
        RECT 101.775 100.390 102.065 100.705 ;
        RECT 102.280 100.690 102.600 100.750 ;
        RECT 104.715 100.705 105.365 100.750 ;
        RECT 105.960 100.890 106.280 100.950 ;
        RECT 107.355 100.890 107.645 100.935 ;
        RECT 105.960 100.750 107.645 100.890 ;
        RECT 105.960 100.690 106.280 100.750 ;
        RECT 107.355 100.705 107.645 100.750 ;
        RECT 107.800 100.890 108.120 100.950 ;
        RECT 116.080 100.890 116.400 100.950 ;
        RECT 123.990 100.935 124.130 101.090 ;
        RECT 126.660 101.030 126.980 101.290 ;
        RECT 118.035 100.890 118.325 100.935 ;
        RECT 121.275 100.890 121.925 100.935 ;
        RECT 107.800 100.750 108.950 100.890 ;
        RECT 107.800 100.690 108.120 100.750 ;
        RECT 108.810 100.595 108.950 100.750 ;
        RECT 116.080 100.750 121.925 100.890 ;
        RECT 116.080 100.690 116.400 100.750 ;
        RECT 118.035 100.705 118.625 100.750 ;
        RECT 121.275 100.705 121.925 100.750 ;
        RECT 123.915 100.705 124.205 100.935 ;
        RECT 102.855 100.550 103.145 100.595 ;
        RECT 106.435 100.550 106.725 100.595 ;
        RECT 108.270 100.550 108.560 100.595 ;
        RECT 102.855 100.410 108.560 100.550 ;
        RECT 102.855 100.365 103.145 100.410 ;
        RECT 106.435 100.365 106.725 100.410 ;
        RECT 108.270 100.365 108.560 100.410 ;
        RECT 108.735 100.365 109.025 100.595 ;
        RECT 118.335 100.390 118.625 100.705 ;
        RECT 119.415 100.550 119.705 100.595 ;
        RECT 122.995 100.550 123.285 100.595 ;
        RECT 124.830 100.550 125.120 100.595 ;
        RECT 119.415 100.410 125.120 100.550 ;
        RECT 119.415 100.365 119.705 100.410 ;
        RECT 122.995 100.365 123.285 100.410 ;
        RECT 124.830 100.365 125.120 100.410 ;
        RECT 127.580 100.350 127.900 100.610 ;
        RECT 21.795 100.210 22.085 100.255 ;
        RECT 27.760 100.210 28.080 100.270 ;
        RECT 21.795 100.070 28.080 100.210 ;
        RECT 21.795 100.025 22.085 100.070 ;
        RECT 27.760 100.010 28.080 100.070 ;
        RECT 46.175 100.210 46.465 100.255 ;
        RECT 51.220 100.210 51.540 100.270 ;
        RECT 46.175 100.070 51.540 100.210 ;
        RECT 46.175 100.025 46.465 100.070 ;
        RECT 51.220 100.010 51.540 100.070 ;
        RECT 60.420 100.210 60.740 100.270 ;
        RECT 64.115 100.210 64.405 100.255 ;
        RECT 60.420 100.070 64.405 100.210 ;
        RECT 60.420 100.010 60.740 100.070 ;
        RECT 64.115 100.025 64.405 100.070 ;
        RECT 80.215 100.210 80.505 100.255 ;
        RECT 83.420 100.210 83.740 100.270 ;
        RECT 89.875 100.210 90.165 100.255 ;
        RECT 80.215 100.070 90.165 100.210 ;
        RECT 80.215 100.025 80.505 100.070 ;
        RECT 83.420 100.010 83.740 100.070 ;
        RECT 89.875 100.025 90.165 100.070 ;
        RECT 118.840 100.210 119.160 100.270 ;
        RECT 125.295 100.210 125.585 100.255 ;
        RECT 118.840 100.070 125.585 100.210 ;
        RECT 118.840 100.010 119.160 100.070 ;
        RECT 125.295 100.025 125.585 100.070 ;
        RECT 21.285 99.870 21.575 99.915 ;
        RECT 23.175 99.870 23.465 99.915 ;
        RECT 26.295 99.870 26.585 99.915 ;
        RECT 21.285 99.730 26.585 99.870 ;
        RECT 21.285 99.685 21.575 99.730 ;
        RECT 23.175 99.685 23.465 99.730 ;
        RECT 26.295 99.685 26.585 99.730 ;
        RECT 32.475 99.870 32.765 99.915 ;
        RECT 35.595 99.870 35.885 99.915 ;
        RECT 37.485 99.870 37.775 99.915 ;
        RECT 32.475 99.730 37.775 99.870 ;
        RECT 32.475 99.685 32.765 99.730 ;
        RECT 35.595 99.685 35.885 99.730 ;
        RECT 37.485 99.685 37.775 99.730 ;
        RECT 47.045 99.870 47.335 99.915 ;
        RECT 48.935 99.870 49.225 99.915 ;
        RECT 52.055 99.870 52.345 99.915 ;
        RECT 47.045 99.730 52.345 99.870 ;
        RECT 47.045 99.685 47.335 99.730 ;
        RECT 48.935 99.685 49.225 99.730 ;
        RECT 52.055 99.685 52.345 99.730 ;
        RECT 58.235 99.870 58.525 99.915 ;
        RECT 61.355 99.870 61.645 99.915 ;
        RECT 63.245 99.870 63.535 99.915 ;
        RECT 58.235 99.730 63.535 99.870 ;
        RECT 58.235 99.685 58.525 99.730 ;
        RECT 61.355 99.685 61.645 99.730 ;
        RECT 63.245 99.685 63.535 99.730 ;
        RECT 74.335 99.870 74.625 99.915 ;
        RECT 77.455 99.870 77.745 99.915 ;
        RECT 79.345 99.870 79.635 99.915 ;
        RECT 74.335 99.730 79.635 99.870 ;
        RECT 74.335 99.685 74.625 99.730 ;
        RECT 77.455 99.685 77.745 99.730 ;
        RECT 79.345 99.685 79.635 99.730 ;
        RECT 83.995 99.870 84.285 99.915 ;
        RECT 87.115 99.870 87.405 99.915 ;
        RECT 89.005 99.870 89.295 99.915 ;
        RECT 83.995 99.730 89.295 99.870 ;
        RECT 83.995 99.685 84.285 99.730 ;
        RECT 87.115 99.685 87.405 99.730 ;
        RECT 89.005 99.685 89.295 99.730 ;
        RECT 102.855 99.870 103.145 99.915 ;
        RECT 105.975 99.870 106.265 99.915 ;
        RECT 107.865 99.870 108.155 99.915 ;
        RECT 102.855 99.730 108.155 99.870 ;
        RECT 102.855 99.685 103.145 99.730 ;
        RECT 105.975 99.685 106.265 99.730 ;
        RECT 107.865 99.685 108.155 99.730 ;
        RECT 119.415 99.870 119.705 99.915 ;
        RECT 122.535 99.870 122.825 99.915 ;
        RECT 124.425 99.870 124.715 99.915 ;
        RECT 119.415 99.730 124.715 99.870 ;
        RECT 119.415 99.685 119.705 99.730 ;
        RECT 122.535 99.685 122.825 99.730 ;
        RECT 124.425 99.685 124.715 99.730 ;
        RECT 27.300 99.530 27.620 99.590 ;
        RECT 29.155 99.530 29.445 99.575 ;
        RECT 27.300 99.390 29.445 99.530 ;
        RECT 27.300 99.330 27.620 99.390 ;
        RECT 29.155 99.345 29.445 99.390 ;
        RECT 29.615 99.530 29.905 99.575 ;
        RECT 31.900 99.530 32.220 99.590 ;
        RECT 29.615 99.390 32.220 99.530 ;
        RECT 29.615 99.345 29.905 99.390 ;
        RECT 31.900 99.330 32.220 99.390 ;
        RECT 53.060 99.530 53.380 99.590 ;
        RECT 54.915 99.530 55.205 99.575 ;
        RECT 53.060 99.390 55.205 99.530 ;
        RECT 53.060 99.330 53.380 99.390 ;
        RECT 54.915 99.345 55.205 99.390 ;
        RECT 55.375 99.530 55.665 99.575 ;
        RECT 59.500 99.530 59.820 99.590 ;
        RECT 55.375 99.390 59.820 99.530 ;
        RECT 55.375 99.345 55.665 99.390 ;
        RECT 59.500 99.330 59.820 99.390 ;
        RECT 71.460 99.330 71.780 99.590 ;
        RECT 81.135 99.530 81.425 99.575 ;
        RECT 85.260 99.530 85.580 99.590 ;
        RECT 81.135 99.390 85.580 99.530 ;
        RECT 81.135 99.345 81.425 99.390 ;
        RECT 85.260 99.330 85.580 99.390 ;
        RECT 99.995 99.530 100.285 99.575 ;
        RECT 104.580 99.530 104.900 99.590 ;
        RECT 99.995 99.390 104.900 99.530 ;
        RECT 99.995 99.345 100.285 99.390 ;
        RECT 104.580 99.330 104.900 99.390 ;
        RECT 116.555 99.530 116.845 99.575 ;
        RECT 117.460 99.530 117.780 99.590 ;
        RECT 116.555 99.390 117.780 99.530 ;
        RECT 116.555 99.345 116.845 99.390 ;
        RECT 117.460 99.330 117.780 99.390 ;
        RECT 9.290 98.710 129.350 99.190 ;
        RECT 9.290 95.990 129.350 96.470 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 18.410 215.725 20.290 216.095 ;
        RECT 48.410 215.725 50.290 216.095 ;
        RECT 78.410 215.725 80.290 216.095 ;
        RECT 108.410 215.725 110.290 216.095 ;
        RECT 33.410 213.005 35.290 213.375 ;
        RECT 63.410 213.005 65.290 213.375 ;
        RECT 93.410 213.005 95.290 213.375 ;
        RECT 123.410 213.005 125.290 213.375 ;
        RECT 18.410 210.285 20.290 210.655 ;
        RECT 48.410 210.285 50.290 210.655 ;
        RECT 78.410 210.285 80.290 210.655 ;
        RECT 108.410 210.285 110.290 210.655 ;
        RECT 33.410 207.565 35.290 207.935 ;
        RECT 63.410 207.565 65.290 207.935 ;
        RECT 93.410 207.565 95.290 207.935 ;
        RECT 123.410 207.565 125.290 207.935 ;
        RECT 18.410 204.845 20.290 205.215 ;
        RECT 48.410 204.845 50.290 205.215 ;
        RECT 78.410 204.845 80.290 205.215 ;
        RECT 108.410 204.845 110.290 205.215 ;
        RECT 33.410 202.125 35.290 202.495 ;
        RECT 63.410 202.125 65.290 202.495 ;
        RECT 93.410 202.125 95.290 202.495 ;
        RECT 123.410 202.125 125.290 202.495 ;
        RECT 18.410 199.405 20.290 199.775 ;
        RECT 48.410 199.405 50.290 199.775 ;
        RECT 78.410 199.405 80.290 199.775 ;
        RECT 108.410 199.405 110.290 199.775 ;
        RECT 62.750 198.240 63.010 198.560 ;
        RECT 66.430 198.240 66.690 198.560 ;
        RECT 100.470 198.240 100.730 198.560 ;
        RECT 116.110 198.240 116.370 198.560 ;
        RECT 54.930 197.900 55.190 198.220 ;
        RECT 33.410 196.685 35.290 197.055 ;
        RECT 54.990 195.840 55.130 197.900 ;
        RECT 54.930 195.520 55.190 195.840 ;
        RECT 56.770 195.520 57.030 195.840 ;
        RECT 38.370 195.180 38.630 195.500 ;
        RECT 51.710 195.180 51.970 195.500 ;
        RECT 54.010 195.180 54.270 195.500 ;
        RECT 18.410 193.965 20.290 194.335 ;
        RECT 36.070 192.800 36.330 193.120 ;
        RECT 35.610 192.460 35.870 192.780 ;
        RECT 33.410 191.245 35.290 191.615 ;
        RECT 31.470 190.080 31.730 190.400 ;
        RECT 22.730 189.740 22.990 190.060 ;
        RECT 18.410 188.525 20.290 188.895 ;
        RECT 22.790 187.680 22.930 189.740 ;
        RECT 31.530 188.020 31.670 190.080 ;
        RECT 31.470 187.700 31.730 188.020 ;
        RECT 35.670 187.760 35.810 192.460 ;
        RECT 36.130 189.380 36.270 192.800 ;
        RECT 38.430 192.440 38.570 195.180 ;
        RECT 40.670 194.500 40.930 194.820 ;
        RECT 46.190 194.500 46.450 194.820 ;
        RECT 50.790 194.500 51.050 194.820 ;
        RECT 40.730 193.460 40.870 194.500 ;
        RECT 40.670 193.140 40.930 193.460 ;
        RECT 46.250 193.120 46.390 194.500 ;
        RECT 48.410 193.965 50.290 194.335 ;
        RECT 50.850 193.120 50.990 194.500 ;
        RECT 46.190 192.800 46.450 193.120 ;
        RECT 50.790 192.800 51.050 193.120 ;
        RECT 38.830 192.460 39.090 192.780 ;
        RECT 38.370 192.120 38.630 192.440 ;
        RECT 38.890 190.400 39.030 192.460 ;
        RECT 46.650 191.780 46.910 192.100 ;
        RECT 50.790 191.780 51.050 192.100 ;
        RECT 38.830 190.080 39.090 190.400 ;
        RECT 41.590 189.740 41.850 190.060 ;
        RECT 36.070 189.060 36.330 189.380 ;
        RECT 41.130 189.060 41.390 189.380 ;
        RECT 22.730 187.360 22.990 187.680 ;
        RECT 31.010 187.360 31.270 187.680 ;
        RECT 18.410 183.085 20.290 183.455 ;
        RECT 22.790 181.900 22.930 187.360 ;
        RECT 27.330 187.020 27.590 187.340 ;
        RECT 27.390 183.850 27.530 187.020 ;
        RECT 31.070 185.640 31.210 187.360 ;
        RECT 31.010 185.320 31.270 185.640 ;
        RECT 27.790 183.850 28.050 183.940 ;
        RECT 27.390 183.710 28.050 183.850 ;
        RECT 27.790 183.620 28.050 183.710 ;
        RECT 28.250 183.620 28.510 183.940 ;
        RECT 27.330 181.920 27.590 182.240 ;
        RECT 22.730 181.580 22.990 181.900 ;
        RECT 21.810 180.900 22.070 181.220 ;
        RECT 16.750 178.860 17.010 179.180 ;
        RECT 16.290 165.940 16.550 166.260 ;
        RECT 16.350 163.880 16.490 165.940 ;
        RECT 16.810 165.580 16.950 178.860 ;
        RECT 21.870 178.840 22.010 180.900 ;
        RECT 21.810 178.520 22.070 178.840 ;
        RECT 18.410 177.645 20.290 178.015 ;
        RECT 22.790 176.800 22.930 181.580 ;
        RECT 26.410 180.900 26.670 181.220 ;
        RECT 26.470 179.520 26.610 180.900 ;
        RECT 27.390 180.200 27.530 181.920 ;
        RECT 27.330 179.880 27.590 180.200 ;
        RECT 26.410 179.200 26.670 179.520 ;
        RECT 22.730 176.480 22.990 176.800 ;
        RECT 18.410 172.205 20.290 172.575 ;
        RECT 18.410 166.765 20.290 167.135 ;
        RECT 17.670 165.940 17.930 166.260 ;
        RECT 16.750 165.260 17.010 165.580 ;
        RECT 16.290 163.560 16.550 163.880 ;
        RECT 16.810 162.860 16.950 165.260 ;
        RECT 15.370 162.540 15.630 162.860 ;
        RECT 16.750 162.540 17.010 162.860 ;
        RECT 15.430 160.820 15.570 162.540 ;
        RECT 15.370 160.500 15.630 160.820 ;
        RECT 16.810 159.460 16.950 162.540 ;
        RECT 17.730 161.160 17.870 165.940 ;
        RECT 22.790 165.920 22.930 176.480 ;
        RECT 27.850 171.020 27.990 183.620 ;
        RECT 28.310 179.860 28.450 183.620 ;
        RECT 28.250 179.540 28.510 179.860 ;
        RECT 28.250 178.520 28.510 178.840 ;
        RECT 30.550 178.520 30.810 178.840 ;
        RECT 28.310 177.480 28.450 178.520 ;
        RECT 28.250 177.160 28.510 177.480 ;
        RECT 28.310 174.080 28.450 177.160 ;
        RECT 30.090 176.140 30.350 176.460 ;
        RECT 30.150 174.760 30.290 176.140 ;
        RECT 30.090 174.440 30.350 174.760 ;
        RECT 28.250 173.760 28.510 174.080 ;
        RECT 27.790 170.700 28.050 171.020 ;
        RECT 22.730 165.600 22.990 165.920 ;
        RECT 21.350 165.260 21.610 165.580 ;
        RECT 18.410 161.325 20.290 161.695 ;
        RECT 17.670 160.840 17.930 161.160 ;
        RECT 21.410 160.140 21.550 165.260 ;
        RECT 22.790 160.480 22.930 165.600 ;
        RECT 23.650 164.580 23.910 164.900 ;
        RECT 28.710 164.580 28.970 164.900 ;
        RECT 23.710 162.860 23.850 164.580 ;
        RECT 23.650 162.540 23.910 162.860 ;
        RECT 28.770 162.180 28.910 164.580 ;
        RECT 29.170 162.880 29.430 163.200 ;
        RECT 29.230 162.180 29.370 162.880 ;
        RECT 26.410 161.860 26.670 162.180 ;
        RECT 26.870 161.860 27.130 162.180 ;
        RECT 28.710 161.860 28.970 162.180 ;
        RECT 29.170 161.860 29.430 162.180 ;
        RECT 26.470 161.160 26.610 161.860 ;
        RECT 26.410 160.840 26.670 161.160 ;
        RECT 26.930 160.480 27.070 161.860 ;
        RECT 22.730 160.160 22.990 160.480 ;
        RECT 26.870 160.160 27.130 160.480 ;
        RECT 21.350 159.820 21.610 160.140 ;
        RECT 22.270 159.820 22.530 160.140 ;
        RECT 26.410 159.820 26.670 160.140 ;
        RECT 16.750 159.140 17.010 159.460 ;
        RECT 20.430 159.140 20.690 159.460 ;
        RECT 17.670 157.440 17.930 157.760 ;
        RECT 15.830 156.760 16.090 157.080 ;
        RECT 15.890 155.720 16.030 156.760 ;
        RECT 16.290 156.420 16.550 156.740 ;
        RECT 15.830 155.400 16.090 155.720 ;
        RECT 16.350 152.660 16.490 156.420 ;
        RECT 17.730 155.720 17.870 157.440 ;
        RECT 20.490 157.420 20.630 159.140 ;
        RECT 20.430 157.100 20.690 157.420 ;
        RECT 18.410 155.885 20.290 156.255 ;
        RECT 17.670 155.400 17.930 155.720 ;
        RECT 19.510 154.720 19.770 155.040 ;
        RECT 19.570 153.000 19.710 154.720 ;
        RECT 19.510 152.680 19.770 153.000 ;
        RECT 16.290 152.340 16.550 152.660 ;
        RECT 17.670 150.980 17.930 151.300 ;
        RECT 13.990 148.260 14.250 148.580 ;
        RECT 15.830 148.260 16.090 148.580 ;
        RECT 14.050 146.200 14.190 148.260 ;
        RECT 15.890 146.880 16.030 148.260 ;
        RECT 15.830 146.560 16.090 146.880 ;
        RECT 13.990 145.880 14.250 146.200 ;
        RECT 17.730 143.820 17.870 150.980 ;
        RECT 18.410 150.445 20.290 150.815 ;
        RECT 19.970 149.280 20.230 149.600 ;
        RECT 18.590 148.940 18.850 149.260 ;
        RECT 18.650 147.560 18.790 148.940 ;
        RECT 18.590 147.240 18.850 147.560 ;
        RECT 20.030 146.280 20.170 149.280 ;
        RECT 20.490 147.220 20.630 157.100 ;
        RECT 20.890 154.380 21.150 154.700 ;
        RECT 20.950 149.600 21.090 154.380 ;
        RECT 21.410 149.940 21.550 159.820 ;
        RECT 22.330 151.980 22.470 159.820 ;
        RECT 26.470 158.100 26.610 159.820 ;
        RECT 26.410 157.780 26.670 158.100 ;
        RECT 28.770 157.760 28.910 161.860 ;
        RECT 29.230 160.820 29.370 161.860 ;
        RECT 29.170 160.500 29.430 160.820 ;
        RECT 28.710 157.440 28.970 157.760 ;
        RECT 24.110 157.100 24.370 157.420 ;
        RECT 27.790 157.100 28.050 157.420 ;
        RECT 24.170 154.700 24.310 157.100 ;
        RECT 25.030 156.420 25.290 156.740 ;
        RECT 25.090 155.380 25.230 156.420 ;
        RECT 27.850 155.720 27.990 157.100 ;
        RECT 27.790 155.400 28.050 155.720 ;
        RECT 25.030 155.060 25.290 155.380 ;
        RECT 24.110 154.380 24.370 154.700 ;
        RECT 29.230 152.320 29.370 160.500 ;
        RECT 29.630 156.420 29.890 156.740 ;
        RECT 29.170 152.000 29.430 152.320 ;
        RECT 29.690 151.980 29.830 156.420 ;
        RECT 30.090 154.380 30.350 154.700 ;
        RECT 30.150 153.000 30.290 154.380 ;
        RECT 30.090 152.680 30.350 153.000 ;
        RECT 22.270 151.660 22.530 151.980 ;
        RECT 29.630 151.660 29.890 151.980 ;
        RECT 21.350 149.620 21.610 149.940 ;
        RECT 20.890 149.280 21.150 149.600 ;
        RECT 22.330 149.260 22.470 151.660 ;
        RECT 22.270 148.940 22.530 149.260 ;
        RECT 20.430 146.900 20.690 147.220 ;
        RECT 22.330 146.880 22.470 148.940 ;
        RECT 22.270 146.560 22.530 146.880 ;
        RECT 20.430 146.280 20.690 146.540 ;
        RECT 20.030 146.220 20.690 146.280 ;
        RECT 20.030 146.140 20.630 146.220 ;
        RECT 18.410 145.005 20.290 145.375 ;
        RECT 17.670 143.500 17.930 143.820 ;
        RECT 16.290 142.820 16.550 143.140 ;
        RECT 16.350 141.440 16.490 142.820 ;
        RECT 17.730 142.120 17.870 143.500 ;
        RECT 17.670 141.800 17.930 142.120 ;
        RECT 16.290 141.120 16.550 141.440 ;
        RECT 17.670 140.100 17.930 140.420 ;
        RECT 17.730 139.400 17.870 140.100 ;
        RECT 18.410 139.565 20.290 139.935 ;
        RECT 17.670 139.080 17.930 139.400 ;
        RECT 20.490 138.720 20.630 146.140 ;
        RECT 21.810 145.880 22.070 146.200 ;
        RECT 21.350 143.500 21.610 143.820 ;
        RECT 21.410 141.520 21.550 143.500 ;
        RECT 20.950 141.440 21.550 141.520 ;
        RECT 20.950 141.380 21.610 141.440 ;
        RECT 20.430 138.400 20.690 138.720 ;
        RECT 18.410 134.125 20.290 134.495 ;
        RECT 20.430 132.960 20.690 133.280 ;
        RECT 17.670 132.620 17.930 132.940 ;
        RECT 12.150 129.560 12.410 129.880 ;
        RECT 12.210 128.520 12.350 129.560 ;
        RECT 12.150 128.200 12.410 128.520 ;
        RECT 15.830 127.860 16.090 128.180 ;
        RECT 12.610 127.520 12.870 127.840 ;
        RECT 12.670 124.780 12.810 127.520 ;
        RECT 15.890 125.800 16.030 127.860 ;
        RECT 17.730 126.560 17.870 132.620 ;
        RECT 20.490 129.540 20.630 132.960 ;
        RECT 20.950 130.220 21.090 141.380 ;
        RECT 21.350 141.120 21.610 141.380 ;
        RECT 20.890 129.900 21.150 130.220 ;
        RECT 20.430 129.220 20.690 129.540 ;
        RECT 18.410 128.685 20.290 129.055 ;
        RECT 18.130 126.560 18.390 126.820 ;
        RECT 17.730 126.500 18.390 126.560 ;
        RECT 17.730 126.420 18.330 126.500 ;
        RECT 15.830 125.480 16.090 125.800 ;
        RECT 17.730 125.120 17.870 126.420 ;
        RECT 20.490 125.120 20.630 129.220 ;
        RECT 20.950 127.920 21.090 129.900 ;
        RECT 20.950 127.840 21.550 127.920 ;
        RECT 20.950 127.780 21.610 127.840 ;
        RECT 21.350 127.520 21.610 127.780 ;
        RECT 17.670 124.800 17.930 125.120 ;
        RECT 20.430 124.800 20.690 125.120 ;
        RECT 12.610 124.460 12.870 124.780 ;
        RECT 12.670 116.960 12.810 124.460 ;
        RECT 17.730 119.680 17.870 124.800 ;
        RECT 18.410 123.245 20.290 123.615 ;
        RECT 17.670 119.360 17.930 119.680 ;
        RECT 18.130 119.080 18.390 119.340 ;
        RECT 17.270 119.020 18.390 119.080 ;
        RECT 17.270 118.940 18.330 119.020 ;
        RECT 17.270 117.040 17.410 118.940 ;
        RECT 17.670 118.340 17.930 118.660 ;
        RECT 21.350 118.340 21.610 118.660 ;
        RECT 17.730 117.640 17.870 118.340 ;
        RECT 18.410 117.805 20.290 118.175 ;
        RECT 17.670 117.320 17.930 117.640 ;
        RECT 12.610 116.640 12.870 116.960 ;
        RECT 17.270 116.900 17.870 117.040 ;
        RECT 12.670 111.520 12.810 116.640 ;
        RECT 17.730 114.920 17.870 116.900 ;
        RECT 20.890 116.300 21.150 116.620 ;
        RECT 17.670 114.600 17.930 114.920 ;
        RECT 20.950 114.240 21.090 116.300 ;
        RECT 21.410 114.240 21.550 118.340 ;
        RECT 20.890 113.920 21.150 114.240 ;
        RECT 21.350 113.920 21.610 114.240 ;
        RECT 16.290 113.240 16.550 113.560 ;
        RECT 16.350 112.200 16.490 113.240 ;
        RECT 18.410 112.365 20.290 112.735 ;
        RECT 16.290 111.880 16.550 112.200 ;
        RECT 12.610 111.200 12.870 111.520 ;
        RECT 20.950 108.800 21.090 113.920 ;
        RECT 20.890 108.480 21.150 108.800 ;
        RECT 15.830 107.800 16.090 108.120 ;
        RECT 8.010 107.460 8.270 107.780 ;
        RECT 8.070 86.920 8.210 107.460 ;
        RECT 14.450 104.740 14.710 105.060 ;
        RECT 14.510 89.420 14.650 104.740 ;
        RECT 15.890 104.040 16.030 107.800 ;
        RECT 18.410 106.925 20.290 107.295 ;
        RECT 20.950 106.840 21.090 108.480 ;
        RECT 21.870 108.460 22.010 145.880 ;
        RECT 22.330 143.480 22.470 146.560 ;
        RECT 22.730 145.540 22.990 145.860 ;
        RECT 23.190 145.540 23.450 145.860 ;
        RECT 27.790 145.540 28.050 145.860 ;
        RECT 22.790 144.500 22.930 145.540 ;
        RECT 23.250 144.840 23.390 145.540 ;
        RECT 23.190 144.520 23.450 144.840 ;
        RECT 22.730 144.180 22.990 144.500 ;
        RECT 27.850 144.160 27.990 145.540 ;
        RECT 27.790 143.840 28.050 144.160 ;
        RECT 22.270 143.160 22.530 143.480 ;
        RECT 28.250 140.100 28.510 140.420 ;
        RECT 27.790 138.740 28.050 139.060 ;
        RECT 27.330 137.380 27.590 137.700 ;
        RECT 22.730 133.300 22.990 133.620 ;
        RECT 22.270 131.940 22.530 132.260 ;
        RECT 22.330 130.220 22.470 131.940 ;
        RECT 22.270 129.900 22.530 130.220 ;
        RECT 22.790 119.340 22.930 133.300 ;
        RECT 26.870 132.960 27.130 133.280 ;
        RECT 26.930 132.600 27.070 132.960 ;
        RECT 26.870 132.280 27.130 132.600 ;
        RECT 24.570 130.920 24.830 131.240 ;
        RECT 24.110 129.900 24.370 130.220 ;
        RECT 23.190 129.220 23.450 129.540 ;
        RECT 23.250 127.500 23.390 129.220 ;
        RECT 23.190 127.180 23.450 127.500 ;
        RECT 24.170 125.800 24.310 129.900 ;
        RECT 24.630 128.520 24.770 130.920 ;
        RECT 24.570 128.200 24.830 128.520 ;
        RECT 24.110 125.480 24.370 125.800 ;
        RECT 24.630 124.100 24.770 128.200 ;
        RECT 25.030 127.860 25.290 128.180 ;
        RECT 25.090 125.800 25.230 127.860 ;
        RECT 25.030 125.480 25.290 125.800 ;
        RECT 24.570 123.780 24.830 124.100 ;
        RECT 23.650 121.740 23.910 122.060 ;
        RECT 22.730 119.020 22.990 119.340 ;
        RECT 23.710 119.000 23.850 121.740 ;
        RECT 24.570 119.020 24.830 119.340 ;
        RECT 23.650 118.680 23.910 119.000 ;
        RECT 24.110 118.340 24.370 118.660 ;
        RECT 22.270 116.640 22.530 116.960 ;
        RECT 22.330 114.920 22.470 116.640 ;
        RECT 22.270 114.600 22.530 114.920 ;
        RECT 24.170 113.900 24.310 118.340 ;
        RECT 24.630 117.640 24.770 119.020 ;
        RECT 24.570 117.320 24.830 117.640 ;
        RECT 24.110 113.580 24.370 113.900 ;
        RECT 21.810 108.140 22.070 108.460 ;
        RECT 23.190 107.460 23.450 107.780 ;
        RECT 20.950 106.700 21.550 106.840 ;
        RECT 21.410 105.740 21.550 106.700 ;
        RECT 23.250 106.420 23.390 107.460 ;
        RECT 23.190 106.100 23.450 106.420 ;
        RECT 27.390 106.080 27.530 137.380 ;
        RECT 27.850 108.460 27.990 138.740 ;
        RECT 28.310 138.720 28.450 140.100 ;
        RECT 28.710 139.080 28.970 139.400 ;
        RECT 28.250 138.400 28.510 138.720 ;
        RECT 28.250 137.380 28.510 137.700 ;
        RECT 28.310 133.960 28.450 137.380 ;
        RECT 28.250 133.640 28.510 133.960 ;
        RECT 27.790 108.140 28.050 108.460 ;
        RECT 28.770 106.080 28.910 139.080 ;
        RECT 29.630 138.400 29.890 138.720 ;
        RECT 29.690 136.340 29.830 138.400 ;
        RECT 30.610 138.380 30.750 178.520 ;
        RECT 31.530 176.800 31.670 187.700 ;
        RECT 35.210 187.620 35.810 187.760 ;
        RECT 35.210 187.340 35.350 187.620 ;
        RECT 35.150 187.020 35.410 187.340 ;
        RECT 33.410 185.805 35.290 186.175 ;
        RECT 35.670 184.960 35.810 187.620 ;
        RECT 36.130 187.340 36.270 189.060 ;
        RECT 36.070 187.020 36.330 187.340 ;
        RECT 32.390 184.640 32.650 184.960 ;
        RECT 35.610 184.640 35.870 184.960 ;
        RECT 32.450 181.220 32.590 184.640 ;
        RECT 32.850 183.620 33.110 183.940 ;
        RECT 32.910 182.580 33.050 183.620 ;
        RECT 32.850 182.260 33.110 182.580 ;
        RECT 36.130 182.320 36.270 187.020 ;
        RECT 41.190 184.960 41.330 189.060 ;
        RECT 41.650 188.360 41.790 189.740 ;
        RECT 41.590 188.040 41.850 188.360 ;
        RECT 46.710 188.020 46.850 191.780 ;
        RECT 48.030 189.060 48.290 189.380 ;
        RECT 48.090 188.360 48.230 189.060 ;
        RECT 48.410 188.525 50.290 188.895 ;
        RECT 48.030 188.040 48.290 188.360 ;
        RECT 46.650 187.700 46.910 188.020 ;
        RECT 41.130 184.640 41.390 184.960 ;
        RECT 36.530 183.960 36.790 184.280 ;
        RECT 40.210 183.960 40.470 184.280 ;
        RECT 36.590 182.920 36.730 183.960 ;
        RECT 40.270 182.920 40.410 183.960 ;
        RECT 41.190 182.920 41.330 184.640 ;
        RECT 45.730 184.300 45.990 184.620 ;
        RECT 42.970 183.620 43.230 183.940 ;
        RECT 36.530 182.600 36.790 182.920 ;
        RECT 40.210 182.600 40.470 182.920 ;
        RECT 41.130 182.600 41.390 182.920 ;
        RECT 32.390 180.900 32.650 181.220 ;
        RECT 32.450 180.200 32.590 180.900 ;
        RECT 32.390 179.880 32.650 180.200 ;
        RECT 31.930 179.540 32.190 179.860 ;
        RECT 31.990 179.180 32.130 179.540 ;
        RECT 31.930 178.860 32.190 179.180 ;
        RECT 31.470 176.480 31.730 176.800 ;
        RECT 31.530 165.580 31.670 176.480 ;
        RECT 32.450 176.460 32.590 179.880 ;
        RECT 32.910 177.480 33.050 182.260 ;
        RECT 36.130 182.180 36.730 182.320 ;
        RECT 33.410 180.365 35.290 180.735 ;
        RECT 35.610 179.540 35.870 179.860 ;
        RECT 35.670 179.180 35.810 179.540 ;
        RECT 36.590 179.180 36.730 182.180 ;
        RECT 35.610 178.860 35.870 179.180 ;
        RECT 36.070 178.860 36.330 179.180 ;
        RECT 36.530 178.860 36.790 179.180 ;
        RECT 36.990 178.860 37.250 179.180 ;
        RECT 33.310 178.520 33.570 178.840 ;
        RECT 32.850 177.160 33.110 177.480 ;
        RECT 32.390 176.140 32.650 176.460 ;
        RECT 33.370 176.200 33.510 178.520 ;
        RECT 36.130 178.500 36.270 178.860 ;
        RECT 36.070 178.180 36.330 178.500 ;
        RECT 32.910 176.060 33.510 176.200 ;
        RECT 31.930 175.460 32.190 175.780 ;
        RECT 31.990 173.740 32.130 175.460 ;
        RECT 31.930 173.420 32.190 173.740 ;
        RECT 32.390 172.740 32.650 173.060 ;
        RECT 31.470 165.260 31.730 165.580 ;
        RECT 31.530 164.760 31.670 165.260 ;
        RECT 31.530 164.620 32.130 164.760 ;
        RECT 31.470 163.220 31.730 163.540 ;
        RECT 31.010 159.820 31.270 160.140 ;
        RECT 31.070 157.420 31.210 159.820 ;
        RECT 31.010 157.100 31.270 157.420 ;
        RECT 31.530 154.440 31.670 163.220 ;
        RECT 31.990 159.460 32.130 164.620 ;
        RECT 32.450 163.540 32.590 172.740 ;
        RECT 32.390 163.220 32.650 163.540 ;
        RECT 32.910 162.600 33.050 176.060 ;
        RECT 33.410 174.925 35.290 175.295 ;
        RECT 34.230 174.100 34.490 174.420 ;
        RECT 34.290 173.740 34.430 174.100 ;
        RECT 34.230 173.420 34.490 173.740 ;
        RECT 35.610 173.420 35.870 173.740 ;
        RECT 35.670 172.120 35.810 173.420 ;
        RECT 36.130 173.060 36.270 178.180 ;
        RECT 37.050 173.740 37.190 178.860 ;
        RECT 37.450 178.180 37.710 178.500 ;
        RECT 37.510 177.140 37.650 178.180 ;
        RECT 37.910 177.160 38.170 177.480 ;
        RECT 37.450 176.820 37.710 177.140 ;
        RECT 37.510 174.420 37.650 176.820 ;
        RECT 37.450 174.100 37.710 174.420 ;
        RECT 37.510 173.740 37.650 174.100 ;
        RECT 37.970 174.080 38.110 177.160 ;
        RECT 41.190 177.140 41.330 182.600 ;
        RECT 43.030 181.220 43.170 183.620 ;
        RECT 45.790 181.900 45.930 184.300 ;
        RECT 45.730 181.580 45.990 181.900 ;
        RECT 42.970 180.900 43.230 181.220 ;
        RECT 43.030 178.840 43.170 180.900 ;
        RECT 45.790 179.520 45.930 181.580 ;
        RECT 45.730 179.200 45.990 179.520 ;
        RECT 42.970 178.520 43.230 178.840 ;
        RECT 41.130 176.820 41.390 177.140 ;
        RECT 40.670 176.480 40.930 176.800 ;
        RECT 37.910 173.760 38.170 174.080 ;
        RECT 40.730 173.740 40.870 176.480 ;
        RECT 42.510 176.140 42.770 176.460 ;
        RECT 41.130 175.460 41.390 175.780 ;
        RECT 36.990 173.420 37.250 173.740 ;
        RECT 37.450 173.420 37.710 173.740 ;
        RECT 40.670 173.420 40.930 173.740 ;
        RECT 36.070 172.740 36.330 173.060 ;
        RECT 37.450 172.740 37.710 173.060 ;
        RECT 35.670 171.980 36.270 172.120 ;
        RECT 35.610 170.020 35.870 170.340 ;
        RECT 33.410 169.485 35.290 169.855 ;
        RECT 33.410 164.045 35.290 164.415 ;
        RECT 32.450 162.460 33.050 162.600 ;
        RECT 33.310 162.540 33.570 162.860 ;
        RECT 31.930 159.140 32.190 159.460 ;
        RECT 31.990 157.420 32.130 159.140 ;
        RECT 31.930 157.100 32.190 157.420 ;
        RECT 31.990 155.040 32.130 157.100 ;
        RECT 31.930 154.720 32.190 155.040 ;
        RECT 31.530 154.300 32.130 154.440 ;
        RECT 31.470 149.280 31.730 149.600 ;
        RECT 31.530 149.000 31.670 149.280 ;
        RECT 31.070 148.860 31.670 149.000 ;
        RECT 31.070 145.770 31.210 148.860 ;
        RECT 31.470 148.260 31.730 148.580 ;
        RECT 31.530 146.540 31.670 148.260 ;
        RECT 31.470 146.220 31.730 146.540 ;
        RECT 31.070 145.630 31.670 145.770 ;
        RECT 31.010 144.180 31.270 144.500 ;
        RECT 31.070 138.720 31.210 144.180 ;
        RECT 31.530 143.480 31.670 145.630 ;
        RECT 31.470 143.160 31.730 143.480 ;
        RECT 31.010 138.400 31.270 138.720 ;
        RECT 31.990 138.380 32.130 154.300 ;
        RECT 32.450 146.880 32.590 162.460 ;
        RECT 32.850 161.860 33.110 162.180 ;
        RECT 32.910 158.440 33.050 161.860 ;
        RECT 33.370 159.460 33.510 162.540 ;
        RECT 34.690 162.200 34.950 162.520 ;
        RECT 34.750 161.160 34.890 162.200 ;
        RECT 34.690 160.840 34.950 161.160 ;
        RECT 33.310 159.140 33.570 159.460 ;
        RECT 33.410 158.605 35.290 158.975 ;
        RECT 32.850 158.120 33.110 158.440 ;
        RECT 32.850 155.400 33.110 155.720 ;
        RECT 32.910 152.570 33.050 155.400 ;
        RECT 35.670 154.440 35.810 170.020 ;
        RECT 36.130 163.280 36.270 171.980 ;
        RECT 36.530 165.940 36.790 166.260 ;
        RECT 36.590 163.880 36.730 165.940 ;
        RECT 36.530 163.560 36.790 163.880 ;
        RECT 36.990 163.560 37.250 163.880 ;
        RECT 37.050 163.280 37.190 163.560 ;
        RECT 36.130 163.140 37.190 163.280 ;
        RECT 36.130 155.720 36.270 163.140 ;
        RECT 36.530 160.160 36.790 160.480 ;
        RECT 36.590 159.995 36.730 160.160 ;
        RECT 36.520 159.625 36.800 159.995 ;
        RECT 36.990 156.760 37.250 157.080 ;
        RECT 36.070 155.400 36.330 155.720 ;
        RECT 36.130 155.040 36.730 155.120 ;
        RECT 37.050 155.040 37.190 156.760 ;
        RECT 36.070 154.980 36.730 155.040 ;
        RECT 36.070 154.720 36.330 154.980 ;
        RECT 35.670 154.300 36.270 154.440 ;
        RECT 35.610 153.700 35.870 154.020 ;
        RECT 33.410 153.165 35.290 153.535 ;
        RECT 34.230 152.680 34.490 153.000 ;
        RECT 32.910 152.430 33.970 152.570 ;
        RECT 33.830 149.600 33.970 152.430 ;
        RECT 34.290 151.980 34.430 152.680 ;
        RECT 34.230 151.890 34.490 151.980 ;
        RECT 34.230 151.750 35.350 151.890 ;
        RECT 34.230 151.660 34.490 151.750 ;
        RECT 35.210 149.600 35.350 151.750 ;
        RECT 33.770 149.280 34.030 149.600 ;
        RECT 35.150 149.280 35.410 149.600 ;
        RECT 35.210 149.115 35.350 149.280 ;
        RECT 35.140 148.745 35.420 149.115 ;
        RECT 33.410 147.725 35.290 148.095 ;
        RECT 32.850 147.240 33.110 147.560 ;
        RECT 32.390 146.560 32.650 146.880 ;
        RECT 32.390 143.160 32.650 143.480 ;
        RECT 32.450 141.100 32.590 143.160 ;
        RECT 32.390 140.780 32.650 141.100 ;
        RECT 30.550 138.060 30.810 138.380 ;
        RECT 31.930 138.060 32.190 138.380 ;
        RECT 30.090 137.380 30.350 137.700 ;
        RECT 32.390 137.380 32.650 137.700 ;
        RECT 29.630 136.020 29.890 136.340 ;
        RECT 30.150 133.960 30.290 137.380 ;
        RECT 32.450 133.960 32.590 137.380 ;
        RECT 30.090 133.640 30.350 133.960 ;
        RECT 32.390 133.640 32.650 133.960 ;
        RECT 31.470 132.960 31.730 133.280 ;
        RECT 30.550 132.620 30.810 132.940 ;
        RECT 30.610 131.240 30.750 132.620 ;
        RECT 30.550 130.920 30.810 131.240 ;
        RECT 31.530 130.220 31.670 132.960 ;
        RECT 31.010 129.900 31.270 130.220 ;
        RECT 31.470 129.900 31.730 130.220 ;
        RECT 31.070 128.520 31.210 129.900 ;
        RECT 32.910 129.880 33.050 147.240 ;
        RECT 35.140 146.705 35.420 147.075 ;
        RECT 35.210 146.540 35.350 146.705 ;
        RECT 35.150 146.220 35.410 146.540 ;
        RECT 33.410 142.285 35.290 142.655 ;
        RECT 35.670 138.380 35.810 153.700 ;
        RECT 36.130 139.060 36.270 154.300 ;
        RECT 36.590 151.550 36.730 154.980 ;
        RECT 36.990 154.720 37.250 155.040 ;
        RECT 36.990 154.040 37.250 154.360 ;
        RECT 37.050 152.320 37.190 154.040 ;
        RECT 36.990 152.000 37.250 152.320 ;
        RECT 36.990 151.550 37.250 151.640 ;
        RECT 36.590 151.410 37.250 151.550 ;
        RECT 36.990 151.320 37.250 151.410 ;
        RECT 37.050 149.600 37.190 151.320 ;
        RECT 36.990 149.280 37.250 149.600 ;
        RECT 36.530 148.600 36.790 148.920 ;
        RECT 36.590 144.160 36.730 148.600 ;
        RECT 36.990 148.260 37.250 148.580 ;
        RECT 37.050 147.220 37.190 148.260 ;
        RECT 36.990 146.900 37.250 147.220 ;
        RECT 36.530 143.840 36.790 144.160 ;
        RECT 36.590 141.100 36.730 143.840 ;
        RECT 37.050 143.820 37.190 146.900 ;
        RECT 36.990 143.500 37.250 143.820 ;
        RECT 36.530 140.780 36.790 141.100 ;
        RECT 36.590 139.060 36.730 140.780 ;
        RECT 37.050 140.760 37.190 143.500 ;
        RECT 36.990 140.440 37.250 140.760 ;
        RECT 36.070 138.740 36.330 139.060 ;
        RECT 36.530 138.740 36.790 139.060 ;
        RECT 35.610 138.060 35.870 138.380 ;
        RECT 33.410 136.845 35.290 137.215 ;
        RECT 33.410 131.405 35.290 131.775 ;
        RECT 35.610 130.240 35.870 130.560 ;
        RECT 32.850 129.560 33.110 129.880 ;
        RECT 31.930 129.220 32.190 129.540 ;
        RECT 31.010 128.200 31.270 128.520 ;
        RECT 31.990 125.120 32.130 129.220 ;
        RECT 33.410 125.965 35.290 126.335 ;
        RECT 35.670 125.800 35.810 130.240 ;
        RECT 36.990 129.900 37.250 130.220 ;
        RECT 37.510 130.130 37.650 172.740 ;
        RECT 40.730 171.360 40.870 173.420 ;
        RECT 40.670 171.040 40.930 171.360 ;
        RECT 40.670 167.980 40.930 168.300 ;
        RECT 40.210 167.300 40.470 167.620 ;
        RECT 38.370 165.600 38.630 165.920 ;
        RECT 38.430 164.760 38.570 165.600 ;
        RECT 37.970 164.620 38.570 164.760 ;
        RECT 37.970 160.480 38.110 164.620 ;
        RECT 38.370 162.880 38.630 163.200 ;
        RECT 37.910 160.160 38.170 160.480 ;
        RECT 38.430 159.880 38.570 162.880 ;
        RECT 40.270 162.860 40.410 167.300 ;
        RECT 40.730 166.600 40.870 167.980 ;
        RECT 40.670 166.280 40.930 166.600 ;
        RECT 40.730 165.920 40.870 166.280 ;
        RECT 40.670 165.600 40.930 165.920 ;
        RECT 40.210 162.540 40.470 162.860 ;
        RECT 37.970 159.800 38.570 159.880 ;
        RECT 37.910 159.740 38.570 159.800 ;
        RECT 37.910 159.480 38.170 159.740 ;
        RECT 37.970 158.440 38.110 159.480 ;
        RECT 37.910 158.120 38.170 158.440 ;
        RECT 37.970 157.760 38.110 158.120 ;
        RECT 37.910 157.440 38.170 157.760 ;
        RECT 38.830 157.440 39.090 157.760 ;
        RECT 37.910 154.040 38.170 154.360 ;
        RECT 37.970 153.080 38.110 154.040 ;
        RECT 37.970 153.000 38.570 153.080 ;
        RECT 37.970 152.940 38.630 153.000 ;
        RECT 38.370 152.680 38.630 152.940 ;
        RECT 38.430 151.980 38.570 152.680 ;
        RECT 38.890 151.980 39.030 157.440 ;
        RECT 39.750 154.720 40.010 155.040 ;
        RECT 39.810 151.980 39.950 154.720 ;
        RECT 38.370 151.660 38.630 151.980 ;
        RECT 38.830 151.660 39.090 151.980 ;
        RECT 39.290 151.660 39.550 151.980 ;
        RECT 39.750 151.660 40.010 151.980 ;
        RECT 38.830 150.980 39.090 151.300 ;
        RECT 37.910 146.220 38.170 146.540 ;
        RECT 37.970 143.480 38.110 146.220 ;
        RECT 38.370 145.540 38.630 145.860 ;
        RECT 37.910 143.160 38.170 143.480 ;
        RECT 37.910 130.130 38.170 130.220 ;
        RECT 37.510 129.990 38.170 130.130 ;
        RECT 37.910 129.900 38.170 129.990 ;
        RECT 36.070 127.520 36.330 127.840 ;
        RECT 35.610 125.480 35.870 125.800 ;
        RECT 31.930 124.800 32.190 125.120 ;
        RECT 35.670 123.080 35.810 125.480 ;
        RECT 36.130 124.440 36.270 127.520 ;
        RECT 36.530 126.500 36.790 126.820 ;
        RECT 36.590 124.780 36.730 126.500 ;
        RECT 37.050 125.460 37.190 129.900 ;
        RECT 38.430 129.880 38.570 145.540 ;
        RECT 38.890 133.280 39.030 150.980 ;
        RECT 39.350 149.940 39.490 151.660 ;
        RECT 39.290 149.620 39.550 149.940 ;
        RECT 40.210 148.260 40.470 148.580 ;
        RECT 38.830 132.960 39.090 133.280 ;
        RECT 38.830 130.920 39.090 131.240 ;
        RECT 38.370 129.560 38.630 129.880 ;
        RECT 37.910 129.220 38.170 129.540 ;
        RECT 36.990 125.140 37.250 125.460 ;
        RECT 36.530 124.460 36.790 124.780 ;
        RECT 36.070 124.120 36.330 124.440 ;
        RECT 35.610 122.760 35.870 123.080 ;
        RECT 36.070 122.080 36.330 122.400 ;
        RECT 32.850 121.740 33.110 122.060 ;
        RECT 35.610 121.740 35.870 122.060 ;
        RECT 32.910 119.340 33.050 121.740 ;
        RECT 33.410 120.525 35.290 120.895 ;
        RECT 35.670 119.680 35.810 121.740 ;
        RECT 35.610 119.360 35.870 119.680 ;
        RECT 36.130 119.340 36.270 122.080 ;
        RECT 32.850 119.020 33.110 119.340 ;
        RECT 33.310 119.020 33.570 119.340 ;
        RECT 36.070 119.020 36.330 119.340 ;
        RECT 30.550 118.340 30.810 118.660 ;
        RECT 29.170 116.980 29.430 117.300 ;
        RECT 29.230 114.920 29.370 116.980 ;
        RECT 29.170 114.600 29.430 114.920 ;
        RECT 30.610 113.900 30.750 118.340 ;
        RECT 31.470 116.640 31.730 116.960 ;
        RECT 32.390 116.640 32.650 116.960 ;
        RECT 31.530 114.920 31.670 116.640 ;
        RECT 31.470 114.600 31.730 114.920 ;
        RECT 32.450 114.240 32.590 116.640 ;
        RECT 33.370 116.460 33.510 119.020 ;
        RECT 36.590 116.620 36.730 124.460 ;
        RECT 36.990 122.760 37.250 123.080 ;
        RECT 37.050 118.660 37.190 122.760 ;
        RECT 37.450 121.400 37.710 121.720 ;
        RECT 37.510 120.360 37.650 121.400 ;
        RECT 37.450 120.040 37.710 120.360 ;
        RECT 36.990 118.340 37.250 118.660 ;
        RECT 32.910 116.320 33.510 116.460 ;
        RECT 32.390 113.920 32.650 114.240 ;
        RECT 29.170 113.580 29.430 113.900 ;
        RECT 30.550 113.580 30.810 113.900 ;
        RECT 29.230 111.520 29.370 113.580 ;
        RECT 32.910 113.220 33.050 116.320 ;
        RECT 36.530 116.300 36.790 116.620 ;
        RECT 35.610 115.620 35.870 115.940 ;
        RECT 33.410 115.085 35.290 115.455 ;
        RECT 35.670 113.560 35.810 115.620 ;
        RECT 35.610 113.240 35.870 113.560 ;
        RECT 32.850 112.900 33.110 113.220 ;
        RECT 29.170 111.200 29.430 111.520 ;
        RECT 33.410 109.645 35.290 110.015 ;
        RECT 37.970 106.080 38.110 129.220 ;
        RECT 38.370 124.460 38.630 124.780 ;
        RECT 38.430 116.960 38.570 124.460 ;
        RECT 38.890 122.740 39.030 130.920 ;
        RECT 40.270 130.220 40.410 148.260 ;
        RECT 40.670 130.920 40.930 131.240 ;
        RECT 40.210 129.900 40.470 130.220 ;
        RECT 39.750 129.220 40.010 129.540 ;
        RECT 39.290 123.780 39.550 124.100 ;
        RECT 38.830 122.420 39.090 122.740 ;
        RECT 39.350 119.000 39.490 123.780 ;
        RECT 39.290 118.680 39.550 119.000 ;
        RECT 38.370 116.640 38.630 116.960 ;
        RECT 39.290 115.620 39.550 115.940 ;
        RECT 39.350 114.240 39.490 115.620 ;
        RECT 39.290 113.920 39.550 114.240 ;
        RECT 39.810 106.420 39.950 129.220 ;
        RECT 40.210 122.080 40.470 122.400 ;
        RECT 40.270 120.360 40.410 122.080 ;
        RECT 40.730 121.380 40.870 130.920 ;
        RECT 41.190 130.220 41.330 175.460 ;
        RECT 42.570 173.740 42.710 176.140 ;
        RECT 43.030 173.740 43.170 178.520 ;
        RECT 45.270 176.480 45.530 176.800 ;
        RECT 45.330 174.420 45.470 176.480 ;
        RECT 45.790 176.460 45.930 179.200 ;
        RECT 45.730 176.140 45.990 176.460 ;
        RECT 45.270 174.100 45.530 174.420 ;
        RECT 46.710 173.740 46.850 187.700 ;
        RECT 48.030 187.360 48.290 187.680 ;
        RECT 48.090 185.640 48.230 187.360 ;
        RECT 50.850 187.340 50.990 191.780 ;
        RECT 51.770 190.060 51.910 195.180 ;
        RECT 51.250 189.740 51.510 190.060 ;
        RECT 51.710 189.740 51.970 190.060 ;
        RECT 53.550 189.740 53.810 190.060 ;
        RECT 49.870 187.020 50.130 187.340 ;
        RECT 50.790 187.020 51.050 187.340 ;
        RECT 48.030 185.320 48.290 185.640 ;
        RECT 49.930 184.960 50.070 187.020 ;
        RECT 49.870 184.640 50.130 184.960 ;
        RECT 48.410 183.085 50.290 183.455 ;
        RECT 48.030 178.180 48.290 178.500 ;
        RECT 48.090 176.120 48.230 178.180 ;
        RECT 48.410 177.645 50.290 178.015 ;
        RECT 50.850 176.880 50.990 187.020 ;
        RECT 51.310 184.280 51.450 189.740 ;
        RECT 53.610 184.620 53.750 189.740 ;
        RECT 54.070 188.360 54.210 195.180 ;
        RECT 56.310 194.500 56.570 194.820 ;
        RECT 56.370 193.460 56.510 194.500 ;
        RECT 56.830 193.460 56.970 195.520 ;
        RECT 56.310 193.140 56.570 193.460 ;
        RECT 56.770 193.140 57.030 193.460 ;
        RECT 62.810 193.120 62.950 198.240 ;
        RECT 66.490 197.540 66.630 198.240 ;
        RECT 68.270 197.900 68.530 198.220 ;
        RECT 72.870 197.900 73.130 198.220 ;
        RECT 66.430 197.220 66.690 197.540 ;
        RECT 63.410 196.685 65.290 197.055 ;
        RECT 65.510 195.180 65.770 195.500 ;
        RECT 63.210 194.840 63.470 195.160 ;
        RECT 63.270 193.800 63.410 194.840 ;
        RECT 65.570 193.800 65.710 195.180 ;
        RECT 63.210 193.480 63.470 193.800 ;
        RECT 65.510 193.480 65.770 193.800 ;
        RECT 58.150 192.800 58.410 193.120 ;
        RECT 62.750 192.800 63.010 193.120 ;
        RECT 65.510 192.800 65.770 193.120 ;
        RECT 54.010 188.040 54.270 188.360 ;
        RECT 53.550 184.300 53.810 184.620 ;
        RECT 51.250 183.960 51.510 184.280 ;
        RECT 51.310 178.840 51.450 183.960 ;
        RECT 53.090 183.620 53.350 183.940 ;
        RECT 53.150 182.580 53.290 183.620 ;
        RECT 53.090 182.260 53.350 182.580 ;
        RECT 51.250 178.520 51.510 178.840 ;
        RECT 50.390 176.800 50.990 176.880 ;
        RECT 50.330 176.740 50.990 176.800 ;
        RECT 50.330 176.480 50.590 176.740 ;
        RECT 48.030 175.800 48.290 176.120 ;
        RECT 47.570 174.100 47.830 174.420 ;
        RECT 47.630 173.740 47.770 174.100 ;
        RECT 42.510 173.650 42.770 173.740 ;
        RECT 42.110 173.510 42.770 173.650 ;
        RECT 42.110 171.700 42.250 173.510 ;
        RECT 42.510 173.420 42.770 173.510 ;
        RECT 42.970 173.420 43.230 173.740 ;
        RECT 43.430 173.650 43.690 173.740 ;
        RECT 44.810 173.650 45.070 173.740 ;
        RECT 43.430 173.510 45.070 173.650 ;
        RECT 43.430 173.420 43.690 173.510 ;
        RECT 44.810 173.420 45.070 173.510 ;
        RECT 46.650 173.420 46.910 173.740 ;
        RECT 47.570 173.420 47.830 173.740 ;
        RECT 42.510 172.740 42.770 173.060 ;
        RECT 44.350 172.740 44.610 173.060 ;
        RECT 42.050 171.380 42.310 171.700 ;
        RECT 42.570 164.760 42.710 172.740 ;
        RECT 43.890 171.040 44.150 171.360 ;
        RECT 43.430 170.020 43.690 170.340 ;
        RECT 42.570 164.620 43.170 164.760 ;
        RECT 42.050 154.040 42.310 154.360 ;
        RECT 42.110 151.980 42.250 154.040 ;
        RECT 42.050 151.660 42.310 151.980 ;
        RECT 42.510 144.520 42.770 144.840 ;
        RECT 42.050 131.940 42.310 132.260 ;
        RECT 41.130 129.900 41.390 130.220 ;
        RECT 42.110 123.080 42.250 131.940 ;
        RECT 42.050 122.760 42.310 123.080 ;
        RECT 40.670 121.060 40.930 121.380 ;
        RECT 40.210 120.040 40.470 120.360 ;
        RECT 42.050 119.360 42.310 119.680 ;
        RECT 42.110 117.300 42.250 119.360 ;
        RECT 42.050 116.980 42.310 117.300 ;
        RECT 41.590 116.640 41.850 116.960 ;
        RECT 41.130 115.960 41.390 116.280 ;
        RECT 41.190 114.240 41.330 115.960 ;
        RECT 41.650 114.920 41.790 116.640 ;
        RECT 41.590 114.600 41.850 114.920 ;
        RECT 42.110 114.240 42.250 116.980 ;
        RECT 41.130 113.920 41.390 114.240 ;
        RECT 42.050 113.920 42.310 114.240 ;
        RECT 42.570 106.760 42.710 144.520 ;
        RECT 43.030 132.940 43.170 164.620 ;
        RECT 43.490 143.820 43.630 170.020 ;
        RECT 43.950 166.600 44.090 171.040 ;
        RECT 43.890 166.280 44.150 166.600 ;
        RECT 43.890 162.880 44.150 163.200 ;
        RECT 43.950 160.140 44.090 162.880 ;
        RECT 43.890 159.820 44.150 160.140 ;
        RECT 43.950 157.420 44.090 159.820 ;
        RECT 43.890 157.100 44.150 157.420 ;
        RECT 43.950 152.660 44.090 157.100 ;
        RECT 43.890 152.340 44.150 152.660 ;
        RECT 43.890 150.980 44.150 151.300 ;
        RECT 43.950 144.160 44.090 150.980 ;
        RECT 44.410 149.260 44.550 172.740 ;
        RECT 44.870 171.360 45.010 173.420 ;
        RECT 47.570 172.740 47.830 173.060 ;
        RECT 44.810 171.040 45.070 171.360 ;
        RECT 44.810 164.580 45.070 164.900 ;
        RECT 47.630 164.760 47.770 172.740 ;
        RECT 48.090 171.440 48.230 175.800 ;
        RECT 50.390 173.740 50.530 176.480 ;
        RECT 49.410 173.420 49.670 173.740 ;
        RECT 50.330 173.420 50.590 173.740 ;
        RECT 50.790 173.420 51.050 173.740 ;
        RECT 49.470 173.060 49.610 173.420 ;
        RECT 49.410 172.740 49.670 173.060 ;
        RECT 48.410 172.205 50.290 172.575 ;
        RECT 48.090 171.360 48.690 171.440 ;
        RECT 50.850 171.360 50.990 173.420 ;
        RECT 48.090 171.300 48.750 171.360 ;
        RECT 48.490 171.040 48.750 171.300 ;
        RECT 49.410 171.040 49.670 171.360 ;
        RECT 50.790 171.040 51.050 171.360 ;
        RECT 49.470 169.320 49.610 171.040 ;
        RECT 49.410 169.000 49.670 169.320 ;
        RECT 48.030 167.980 48.290 168.300 ;
        RECT 48.090 165.580 48.230 167.980 ;
        RECT 48.410 166.765 50.290 167.135 ;
        RECT 51.310 165.580 51.450 178.520 ;
        RECT 53.090 176.820 53.350 177.140 ;
        RECT 53.150 174.760 53.290 176.820 ;
        RECT 53.090 174.440 53.350 174.760 ;
        RECT 53.610 173.740 53.750 184.300 ;
        RECT 58.210 182.240 58.350 192.800 ;
        RECT 63.410 191.245 65.290 191.615 ;
        RECT 65.570 191.080 65.710 192.800 ;
        RECT 66.490 192.360 66.630 197.220 ;
        RECT 66.890 194.840 67.150 195.160 ;
        RECT 66.950 193.120 67.090 194.840 ;
        RECT 68.330 193.800 68.470 197.900 ;
        RECT 72.930 195.500 73.070 197.900 ;
        RECT 98.630 197.220 98.890 197.540 ;
        RECT 93.410 196.685 95.290 197.055 ;
        RECT 83.450 196.200 83.710 196.520 ;
        RECT 91.270 196.200 91.530 196.520 ;
        RECT 74.710 195.520 74.970 195.840 ;
        RECT 72.870 195.180 73.130 195.500 ;
        RECT 69.190 194.840 69.450 195.160 ;
        RECT 71.490 194.840 71.750 195.160 ;
        RECT 69.250 193.800 69.390 194.840 ;
        RECT 68.270 193.480 68.530 193.800 ;
        RECT 69.190 193.480 69.450 193.800 ;
        RECT 67.350 193.140 67.610 193.460 ;
        RECT 66.890 192.800 67.150 193.120 ;
        RECT 66.490 192.220 67.090 192.360 ;
        RECT 66.950 191.080 67.090 192.220 ;
        RECT 65.510 190.760 65.770 191.080 ;
        RECT 66.890 190.760 67.150 191.080 ;
        RECT 66.430 190.080 66.690 190.400 ;
        RECT 65.970 189.740 66.230 190.060 ;
        RECT 63.410 185.805 65.290 186.175 ;
        RECT 66.030 182.580 66.170 189.740 ;
        RECT 66.490 189.380 66.630 190.080 ;
        RECT 66.430 189.060 66.690 189.380 ;
        RECT 66.490 183.940 66.630 189.060 ;
        RECT 66.430 183.620 66.690 183.940 ;
        RECT 65.970 182.260 66.230 182.580 ;
        RECT 58.150 181.920 58.410 182.240 ;
        RECT 56.770 181.580 57.030 181.900 ;
        RECT 56.830 180.200 56.970 181.580 ;
        RECT 56.770 179.880 57.030 180.200 ;
        RECT 58.210 178.840 58.350 181.920 ;
        RECT 63.410 180.365 65.290 180.735 ;
        RECT 58.150 178.520 58.410 178.840 ;
        RECT 58.210 176.800 58.350 178.520 ;
        RECT 60.910 178.180 61.170 178.500 ;
        RECT 58.150 176.480 58.410 176.800 ;
        RECT 56.770 176.140 57.030 176.460 ;
        RECT 54.930 175.460 55.190 175.780 ;
        RECT 54.990 173.740 55.130 175.460 ;
        RECT 56.830 174.760 56.970 176.140 ;
        RECT 56.770 174.440 57.030 174.760 ;
        RECT 59.990 174.100 60.250 174.420 ;
        RECT 53.550 173.420 53.810 173.740 ;
        RECT 54.930 173.420 55.190 173.740 ;
        RECT 58.150 173.080 58.410 173.400 ;
        RECT 58.210 165.580 58.350 173.080 ;
        RECT 60.050 172.040 60.190 174.100 ;
        RECT 59.990 171.720 60.250 172.040 ;
        RECT 59.070 165.600 59.330 165.920 ;
        RECT 48.030 165.260 48.290 165.580 ;
        RECT 51.250 165.260 51.510 165.580 ;
        RECT 58.150 165.260 58.410 165.580 ;
        RECT 47.630 164.620 48.230 164.760 ;
        RECT 44.870 162.520 45.010 164.580 ;
        RECT 44.810 162.200 45.070 162.520 ;
        RECT 45.270 161.860 45.530 162.180 ;
        RECT 45.330 160.480 45.470 161.860 ;
        RECT 45.270 160.160 45.530 160.480 ;
        RECT 47.570 159.820 47.830 160.140 ;
        RECT 46.190 157.100 46.450 157.420 ;
        RECT 46.250 154.700 46.390 157.100 ;
        RECT 46.640 154.865 46.920 155.235 ;
        RECT 47.630 155.040 47.770 159.820 ;
        RECT 46.650 154.720 46.910 154.865 ;
        RECT 47.110 154.720 47.370 155.040 ;
        RECT 47.570 154.720 47.830 155.040 ;
        RECT 46.190 154.380 46.450 154.700 ;
        RECT 44.810 153.700 45.070 154.020 ;
        RECT 44.870 149.600 45.010 153.700 ;
        RECT 45.270 151.320 45.530 151.640 ;
        RECT 44.810 149.280 45.070 149.600 ;
        RECT 44.350 148.940 44.610 149.260 ;
        RECT 44.350 148.260 44.610 148.580 ;
        RECT 43.890 143.840 44.150 144.160 ;
        RECT 43.430 143.500 43.690 143.820 ;
        RECT 43.890 139.080 44.150 139.400 ;
        RECT 43.950 135.660 44.090 139.080 ;
        RECT 43.890 135.340 44.150 135.660 ;
        RECT 42.970 132.620 43.230 132.940 ;
        RECT 43.430 132.280 43.690 132.600 ;
        RECT 42.970 121.060 43.230 121.380 ;
        RECT 43.030 119.680 43.170 121.060 ;
        RECT 42.970 119.360 43.230 119.680 ;
        RECT 42.510 106.440 42.770 106.760 ;
        RECT 39.750 106.100 40.010 106.420 ;
        RECT 43.490 106.080 43.630 132.280 ;
        RECT 43.890 120.040 44.150 120.360 ;
        RECT 43.950 119.680 44.090 120.040 ;
        RECT 43.890 119.360 44.150 119.680 ;
        RECT 44.410 106.760 44.550 148.260 ;
        RECT 45.330 146.880 45.470 151.320 ;
        RECT 45.730 148.260 45.990 148.580 ;
        RECT 45.270 146.560 45.530 146.880 ;
        RECT 44.810 145.880 45.070 146.200 ;
        RECT 45.270 145.880 45.530 146.200 ;
        RECT 44.870 144.840 45.010 145.880 ;
        RECT 44.810 144.520 45.070 144.840 ;
        RECT 44.810 142.820 45.070 143.140 ;
        RECT 44.870 120.360 45.010 142.820 ;
        RECT 45.330 141.100 45.470 145.880 ;
        RECT 45.270 140.780 45.530 141.100 ;
        RECT 45.330 133.280 45.470 140.780 ;
        RECT 45.270 132.960 45.530 133.280 ;
        RECT 45.330 130.220 45.470 132.960 ;
        RECT 45.270 129.900 45.530 130.220 ;
        RECT 45.330 127.500 45.470 129.900 ;
        RECT 45.790 128.520 45.930 148.260 ;
        RECT 46.250 146.540 46.390 154.380 ;
        RECT 46.710 152.320 46.850 154.720 ;
        RECT 47.170 153.000 47.310 154.720 ;
        RECT 47.110 152.680 47.370 153.000 ;
        RECT 46.650 152.000 46.910 152.320 ;
        RECT 47.570 150.980 47.830 151.300 ;
        RECT 47.630 149.600 47.770 150.980 ;
        RECT 48.090 149.600 48.230 164.620 ;
        RECT 51.310 163.200 51.450 165.260 ;
        RECT 51.250 162.880 51.510 163.200 ;
        RECT 50.790 161.860 51.050 162.180 ;
        RECT 48.410 161.325 50.290 161.695 ;
        RECT 50.850 161.160 50.990 161.860 ;
        RECT 50.790 160.840 51.050 161.160 ;
        RECT 48.410 155.885 50.290 156.255 ;
        RECT 51.310 154.700 51.450 162.880 ;
        RECT 54.470 156.420 54.730 156.740 ;
        RECT 55.850 156.420 56.110 156.740 ;
        RECT 54.530 155.380 54.670 156.420 ;
        RECT 54.470 155.060 54.730 155.380 ;
        RECT 55.390 154.720 55.650 155.040 ;
        RECT 51.250 154.380 51.510 154.700 ;
        RECT 55.450 154.555 55.590 154.720 ;
        RECT 50.790 154.040 51.050 154.360 ;
        RECT 55.380 154.185 55.660 154.555 ;
        RECT 48.410 150.445 50.290 150.815 ;
        RECT 47.570 149.280 47.830 149.600 ;
        RECT 48.030 149.280 48.290 149.600 ;
        RECT 47.110 148.260 47.370 148.580 ;
        RECT 46.190 146.220 46.450 146.540 ;
        RECT 46.250 139.400 46.390 146.220 ;
        RECT 46.650 143.840 46.910 144.160 ;
        RECT 46.710 142.120 46.850 143.840 ;
        RECT 46.650 141.800 46.910 142.120 ;
        RECT 46.650 141.120 46.910 141.440 ;
        RECT 46.190 139.080 46.450 139.400 ;
        RECT 46.190 138.060 46.450 138.380 ;
        RECT 46.250 134.980 46.390 138.060 ;
        RECT 46.190 134.660 46.450 134.980 ;
        RECT 46.250 132.940 46.390 134.660 ;
        RECT 46.190 132.620 46.450 132.940 ;
        RECT 46.710 132.600 46.850 141.120 ;
        RECT 46.650 132.280 46.910 132.600 ;
        RECT 46.710 130.560 46.850 132.280 ;
        RECT 46.650 130.240 46.910 130.560 ;
        RECT 46.710 128.520 46.850 130.240 ;
        RECT 45.730 128.200 45.990 128.520 ;
        RECT 46.650 128.200 46.910 128.520 ;
        RECT 46.650 127.520 46.910 127.840 ;
        RECT 45.270 127.180 45.530 127.500 ;
        RECT 46.710 125.800 46.850 127.520 ;
        RECT 46.650 125.480 46.910 125.800 ;
        RECT 44.810 120.040 45.070 120.360 ;
        RECT 46.710 119.680 46.850 125.480 ;
        RECT 47.170 120.360 47.310 148.260 ;
        RECT 50.850 147.220 50.990 154.040 ;
        RECT 54.470 153.700 54.730 154.020 ;
        RECT 54.530 151.300 54.670 153.700 ;
        RECT 55.910 151.300 56.050 156.420 ;
        RECT 56.310 152.000 56.570 152.320 ;
        RECT 54.470 150.980 54.730 151.300 ;
        RECT 55.850 150.980 56.110 151.300 ;
        RECT 52.170 149.280 52.430 149.600 ;
        RECT 51.710 148.940 51.970 149.260 ;
        RECT 50.790 146.900 51.050 147.220 ;
        RECT 51.250 146.900 51.510 147.220 ;
        RECT 47.570 145.880 47.830 146.200 ;
        RECT 47.630 143.560 47.770 145.880 ;
        RECT 48.030 145.540 48.290 145.860 ;
        RECT 48.090 144.500 48.230 145.540 ;
        RECT 48.410 145.005 50.290 145.375 ;
        RECT 48.030 144.180 48.290 144.500 ;
        RECT 47.630 143.420 48.230 143.560 ;
        RECT 50.330 143.500 50.590 143.820 ;
        RECT 48.090 143.140 48.230 143.420 ;
        RECT 48.030 142.820 48.290 143.140 ;
        RECT 48.090 140.420 48.230 142.820 ;
        RECT 50.390 141.100 50.530 143.500 ;
        RECT 50.790 142.820 51.050 143.140 ;
        RECT 50.330 140.780 50.590 141.100 ;
        RECT 48.030 140.100 48.290 140.420 ;
        RECT 48.090 139.400 48.230 140.100 ;
        RECT 48.410 139.565 50.290 139.935 ;
        RECT 48.030 139.080 48.290 139.400 ;
        RECT 47.570 137.380 47.830 137.700 ;
        RECT 47.630 133.960 47.770 137.380 ;
        RECT 50.850 136.000 50.990 142.820 ;
        RECT 51.310 141.780 51.450 146.900 ;
        RECT 51.770 146.540 51.910 148.940 ;
        RECT 52.230 147.560 52.370 149.280 ;
        RECT 54.010 148.940 54.270 149.260 ;
        RECT 54.070 147.560 54.210 148.940 ;
        RECT 52.170 147.240 52.430 147.560 ;
        RECT 54.010 147.240 54.270 147.560 ;
        RECT 54.070 146.540 54.210 147.240 ;
        RECT 54.530 146.540 54.670 150.980 ;
        RECT 55.910 150.280 56.050 150.980 ;
        RECT 55.850 149.960 56.110 150.280 ;
        RECT 56.370 149.940 56.510 152.000 ;
        RECT 56.310 149.620 56.570 149.940 ;
        RECT 55.390 149.280 55.650 149.600 ;
        RECT 55.450 146.540 55.590 149.280 ;
        RECT 56.370 146.880 56.510 149.620 ;
        RECT 57.230 148.600 57.490 148.920 ;
        RECT 56.310 146.560 56.570 146.880 ;
        RECT 51.710 146.220 51.970 146.540 ;
        RECT 54.010 146.220 54.270 146.540 ;
        RECT 54.470 146.220 54.730 146.540 ;
        RECT 55.390 146.220 55.650 146.540 ;
        RECT 51.710 145.540 51.970 145.860 ;
        RECT 51.250 141.460 51.510 141.780 ;
        RECT 51.770 141.100 51.910 145.540 ;
        RECT 55.450 144.160 55.590 146.220 ;
        RECT 55.390 143.840 55.650 144.160 ;
        RECT 53.090 143.500 53.350 143.820 ;
        RECT 53.150 142.120 53.290 143.500 ;
        RECT 53.090 141.800 53.350 142.120 ;
        RECT 56.370 141.100 56.510 146.560 ;
        RECT 51.250 140.780 51.510 141.100 ;
        RECT 51.710 140.780 51.970 141.100 ;
        RECT 56.310 140.780 56.570 141.100 ;
        RECT 50.790 135.680 51.050 136.000 ;
        RECT 48.030 135.340 48.290 135.660 ;
        RECT 48.090 133.960 48.230 135.340 ;
        RECT 48.410 134.125 50.290 134.495 ;
        RECT 47.570 133.640 47.830 133.960 ;
        RECT 48.030 133.640 48.290 133.960 ;
        RECT 47.570 132.960 47.830 133.280 ;
        RECT 48.950 132.960 49.210 133.280 ;
        RECT 47.630 132.600 47.770 132.960 ;
        RECT 47.570 132.280 47.830 132.600 ;
        RECT 49.010 130.220 49.150 132.960 ;
        RECT 49.410 132.620 49.670 132.940 ;
        RECT 49.470 130.220 49.610 132.620 ;
        RECT 47.570 129.900 47.830 130.220 ;
        RECT 48.950 129.900 49.210 130.220 ;
        RECT 49.410 129.900 49.670 130.220 ;
        RECT 47.630 127.920 47.770 129.900 ;
        RECT 48.030 129.220 48.290 129.540 ;
        RECT 48.090 128.520 48.230 129.220 ;
        RECT 48.410 128.685 50.290 129.055 ;
        RECT 48.030 128.200 48.290 128.520 ;
        RECT 49.410 128.200 49.670 128.520 ;
        RECT 47.630 127.780 48.230 127.920 ;
        RECT 49.470 127.840 49.610 128.200 ;
        RECT 47.570 127.180 47.830 127.500 ;
        RECT 47.110 120.040 47.370 120.360 ;
        RECT 46.650 119.360 46.910 119.680 ;
        RECT 47.110 119.020 47.370 119.340 ;
        RECT 46.190 116.300 46.450 116.620 ;
        RECT 46.250 113.900 46.390 116.300 ;
        RECT 47.170 113.900 47.310 119.020 ;
        RECT 47.630 118.660 47.770 127.180 ;
        RECT 48.090 126.820 48.230 127.780 ;
        RECT 49.410 127.520 49.670 127.840 ;
        RECT 48.030 126.500 48.290 126.820 ;
        RECT 50.850 125.120 50.990 135.680 ;
        RECT 51.310 133.620 51.450 140.780 ;
        RECT 56.370 138.380 56.510 140.780 ;
        RECT 56.770 140.100 57.030 140.420 ;
        RECT 51.710 138.060 51.970 138.380 ;
        RECT 56.310 138.060 56.570 138.380 ;
        RECT 51.250 133.300 51.510 133.620 ;
        RECT 51.250 132.620 51.510 132.940 ;
        RECT 51.310 131.240 51.450 132.620 ;
        RECT 51.250 130.920 51.510 131.240 ;
        RECT 51.770 130.560 51.910 138.060 ;
        RECT 56.370 136.000 56.510 138.060 ;
        RECT 56.830 137.700 56.970 140.100 ;
        RECT 56.770 137.380 57.030 137.700 ;
        RECT 56.310 135.680 56.570 136.000 ;
        RECT 55.390 135.340 55.650 135.660 ;
        RECT 55.450 133.280 55.590 135.340 ;
        RECT 55.390 132.960 55.650 133.280 ;
        RECT 55.850 131.940 56.110 132.260 ;
        RECT 51.710 130.240 51.970 130.560 ;
        RECT 51.240 129.705 51.520 130.075 ;
        RECT 51.310 128.520 51.450 129.705 ;
        RECT 51.250 128.200 51.510 128.520 ;
        RECT 51.250 127.520 51.510 127.840 ;
        RECT 51.310 126.820 51.450 127.520 ;
        RECT 51.770 127.410 51.910 130.240 ;
        RECT 55.910 129.880 56.050 131.940 ;
        RECT 55.850 129.560 56.110 129.880 ;
        RECT 52.170 129.220 52.430 129.540 ;
        RECT 52.230 128.180 52.370 129.220 ;
        RECT 52.170 127.860 52.430 128.180 ;
        RECT 52.170 127.410 52.430 127.500 ;
        RECT 51.770 127.270 52.430 127.410 ;
        RECT 52.170 127.180 52.430 127.270 ;
        RECT 51.250 126.500 51.510 126.820 ;
        RECT 50.790 124.800 51.050 125.120 ;
        RECT 48.410 123.245 50.290 123.615 ;
        RECT 50.850 122.400 50.990 124.800 ;
        RECT 50.790 122.310 51.050 122.400 ;
        RECT 50.790 122.170 51.910 122.310 ;
        RECT 50.790 122.080 51.050 122.170 ;
        RECT 50.790 121.060 51.050 121.380 ;
        RECT 47.570 118.340 47.830 118.660 ;
        RECT 47.630 117.640 47.770 118.340 ;
        RECT 48.410 117.805 50.290 118.175 ;
        RECT 47.570 117.320 47.830 117.640 ;
        RECT 50.850 117.300 50.990 121.060 ;
        RECT 51.770 120.020 51.910 122.170 ;
        RECT 51.710 119.700 51.970 120.020 ;
        RECT 51.250 119.020 51.510 119.340 ;
        RECT 50.790 116.980 51.050 117.300 ;
        RECT 50.850 116.620 50.990 116.980 ;
        RECT 51.310 116.960 51.450 119.020 ;
        RECT 51.250 116.640 51.510 116.960 ;
        RECT 48.030 116.300 48.290 116.620 ;
        RECT 50.790 116.300 51.050 116.620 ;
        RECT 46.190 113.580 46.450 113.900 ;
        RECT 47.110 113.580 47.370 113.900 ;
        RECT 47.170 113.220 47.310 113.580 ;
        RECT 47.110 112.900 47.370 113.220 ;
        RECT 47.170 112.200 47.310 112.900 ;
        RECT 47.110 111.880 47.370 112.200 ;
        RECT 48.090 111.860 48.230 116.300 ;
        RECT 51.310 114.240 51.450 116.640 ;
        RECT 51.250 113.920 51.510 114.240 ;
        RECT 50.790 112.900 51.050 113.220 ;
        RECT 48.410 112.365 50.290 112.735 ;
        RECT 48.030 111.540 48.290 111.860 ;
        RECT 50.850 108.460 50.990 112.900 ;
        RECT 51.770 111.180 51.910 119.700 ;
        RECT 54.930 115.620 55.190 115.940 ;
        RECT 54.990 114.240 55.130 115.620 ;
        RECT 54.930 113.920 55.190 114.240 ;
        RECT 53.090 111.200 53.350 111.520 ;
        RECT 51.710 110.860 51.970 111.180 ;
        RECT 53.150 109.480 53.290 111.200 ;
        RECT 53.090 109.160 53.350 109.480 ;
        RECT 50.790 108.140 51.050 108.460 ;
        RECT 48.410 106.925 50.290 107.295 ;
        RECT 44.350 106.440 44.610 106.760 ;
        RECT 57.290 106.080 57.430 148.600 ;
        RECT 57.690 140.780 57.950 141.100 ;
        RECT 57.750 138.720 57.890 140.780 ;
        RECT 57.690 138.400 57.950 138.720 ;
        RECT 57.690 131.940 57.950 132.260 ;
        RECT 57.750 130.560 57.890 131.940 ;
        RECT 57.690 130.240 57.950 130.560 ;
        RECT 57.690 126.500 57.950 126.820 ;
        RECT 57.750 124.780 57.890 126.500 ;
        RECT 57.690 124.460 57.950 124.780 ;
        RECT 58.210 113.220 58.350 165.260 ;
        RECT 59.130 162.860 59.270 165.600 ;
        RECT 60.970 163.200 61.110 178.180 ;
        RECT 66.030 177.560 66.170 182.260 ;
        RECT 66.430 180.900 66.690 181.220 ;
        RECT 65.570 177.420 66.170 177.560 ;
        RECT 62.280 175.945 62.560 176.315 ;
        RECT 62.750 176.140 63.010 176.460 ;
        RECT 61.370 173.420 61.630 173.740 ;
        RECT 61.430 171.360 61.570 173.420 ;
        RECT 61.370 171.040 61.630 171.360 ;
        RECT 62.350 163.880 62.490 175.945 ;
        RECT 62.810 173.650 62.950 176.140 ;
        RECT 63.410 174.925 65.290 175.295 ;
        RECT 65.570 174.760 65.710 177.420 ;
        RECT 65.970 176.480 66.230 176.800 ;
        RECT 65.510 174.440 65.770 174.760 ;
        RECT 63.670 174.100 63.930 174.420 ;
        RECT 66.030 174.160 66.170 176.480 ;
        RECT 63.210 173.650 63.470 173.740 ;
        RECT 62.810 173.510 63.470 173.650 ;
        RECT 63.210 173.420 63.470 173.510 ;
        RECT 63.270 171.700 63.410 173.420 ;
        RECT 63.210 171.380 63.470 171.700 ;
        RECT 63.730 171.020 63.870 174.100 ;
        RECT 64.190 174.080 66.170 174.160 ;
        RECT 64.130 174.020 66.170 174.080 ;
        RECT 64.130 173.760 64.390 174.020 ;
        RECT 64.120 171.865 64.400 172.235 ;
        RECT 64.130 171.720 64.390 171.865 ;
        RECT 63.670 170.700 63.930 171.020 ;
        RECT 63.410 169.485 65.290 169.855 ;
        RECT 66.490 164.760 66.630 180.900 ;
        RECT 66.950 173.650 67.090 190.760 ;
        RECT 67.410 189.380 67.550 193.140 ;
        RECT 67.810 192.460 68.070 192.780 ;
        RECT 67.870 190.480 68.010 192.460 ;
        RECT 68.330 192.100 68.470 193.480 ;
        RECT 69.650 192.800 69.910 193.120 ;
        RECT 69.710 192.520 69.850 192.800 ;
        RECT 69.710 192.380 71.230 192.520 ;
        RECT 68.270 191.780 68.530 192.100 ;
        RECT 67.870 190.400 68.470 190.480 ;
        RECT 67.870 190.340 68.530 190.400 ;
        RECT 68.270 190.080 68.530 190.340 ;
        RECT 69.710 189.720 69.850 192.380 ;
        RECT 70.110 191.780 70.370 192.100 ;
        RECT 69.650 189.400 69.910 189.720 ;
        RECT 67.350 189.060 67.610 189.380 ;
        RECT 70.170 187.680 70.310 191.780 ;
        RECT 71.090 190.060 71.230 192.380 ;
        RECT 71.550 191.080 71.690 194.840 ;
        RECT 71.950 193.140 72.210 193.460 ;
        RECT 71.490 190.760 71.750 191.080 ;
        RECT 71.030 189.740 71.290 190.060 ;
        RECT 70.110 187.360 70.370 187.680 ;
        RECT 69.190 186.340 69.450 186.660 ;
        RECT 69.250 184.960 69.390 186.340 ;
        RECT 70.170 184.960 70.310 187.360 ;
        RECT 71.090 184.960 71.230 189.740 ;
        RECT 71.550 188.360 71.690 190.760 ;
        RECT 72.010 190.060 72.150 193.140 ;
        RECT 71.950 189.740 72.210 190.060 ;
        RECT 72.410 189.740 72.670 190.060 ;
        RECT 71.490 188.040 71.750 188.360 ;
        RECT 69.190 184.640 69.450 184.960 ;
        RECT 70.110 184.640 70.370 184.960 ;
        RECT 71.030 184.640 71.290 184.960 ;
        RECT 67.810 183.620 68.070 183.940 ;
        RECT 68.270 183.620 68.530 183.940 ;
        RECT 68.730 183.620 68.990 183.940 ;
        RECT 67.350 181.240 67.610 181.560 ;
        RECT 67.410 176.710 67.550 181.240 ;
        RECT 67.870 179.180 68.010 183.620 ;
        RECT 67.810 178.860 68.070 179.180 ;
        RECT 67.810 176.710 68.070 176.800 ;
        RECT 67.410 176.570 68.070 176.710 ;
        RECT 67.810 176.480 68.070 176.570 ;
        RECT 67.870 174.760 68.010 176.480 ;
        RECT 67.810 174.440 68.070 174.760 ;
        RECT 67.810 173.650 68.070 173.740 ;
        RECT 66.950 173.510 68.070 173.650 ;
        RECT 67.810 173.420 68.070 173.510 ;
        RECT 67.870 168.640 68.010 173.420 ;
        RECT 67.810 168.320 68.070 168.640 ;
        RECT 67.350 166.280 67.610 166.600 ;
        RECT 66.490 164.620 67.090 164.760 ;
        RECT 63.410 164.045 65.290 164.415 ;
        RECT 62.290 163.560 62.550 163.880 ;
        RECT 60.910 162.880 61.170 163.200 ;
        RECT 59.070 162.540 59.330 162.860 ;
        RECT 59.130 157.840 59.270 162.540 ;
        RECT 59.990 158.120 60.250 158.440 ;
        RECT 58.670 157.760 59.270 157.840 ;
        RECT 58.610 157.700 59.270 157.760 ;
        RECT 58.610 157.440 58.870 157.700 ;
        RECT 60.050 155.040 60.190 158.120 ;
        RECT 59.530 154.720 59.790 155.040 ;
        RECT 59.990 154.720 60.250 155.040 ;
        RECT 59.590 153.000 59.730 154.720 ;
        RECT 59.530 152.680 59.790 153.000 ;
        RECT 60.970 143.820 61.110 162.880 ;
        RECT 62.350 161.160 62.490 163.560 ;
        RECT 65.510 162.540 65.770 162.860 ;
        RECT 62.290 160.840 62.550 161.160 ;
        RECT 63.410 158.605 65.290 158.975 ;
        RECT 65.050 157.100 65.310 157.420 ;
        RECT 61.370 156.760 61.630 157.080 ;
        RECT 61.430 155.720 61.570 156.760 ;
        RECT 62.750 156.420 63.010 156.740 ;
        RECT 61.370 155.400 61.630 155.720 ;
        RECT 62.810 153.000 62.950 156.420 ;
        RECT 65.110 154.700 65.250 157.100 ;
        RECT 65.050 154.380 65.310 154.700 ;
        RECT 63.410 153.165 65.290 153.535 ;
        RECT 62.750 152.680 63.010 153.000 ;
        RECT 65.570 152.660 65.710 162.540 ;
        RECT 65.970 157.440 66.230 157.760 ;
        RECT 65.510 152.340 65.770 152.660 ;
        RECT 66.030 152.320 66.170 157.440 ;
        RECT 65.970 152.000 66.230 152.320 ;
        RECT 62.750 151.660 63.010 151.980 ;
        RECT 62.810 150.280 62.950 151.660 ;
        RECT 62.750 149.960 63.010 150.280 ;
        RECT 66.950 149.600 67.090 164.620 ;
        RECT 61.370 149.280 61.630 149.600 ;
        RECT 66.890 149.280 67.150 149.600 ;
        RECT 61.430 143.820 61.570 149.280 ;
        RECT 61.830 148.600 62.090 148.920 ;
        RECT 61.890 144.160 62.030 148.600 ;
        RECT 62.750 148.260 63.010 148.580 ;
        RECT 62.290 147.075 62.550 147.220 ;
        RECT 62.280 146.705 62.560 147.075 ;
        RECT 62.810 144.160 62.950 148.260 ;
        RECT 63.410 147.725 65.290 148.095 ;
        RECT 63.670 144.180 63.930 144.500 ;
        RECT 61.830 143.840 62.090 144.160 ;
        RECT 62.750 143.840 63.010 144.160 ;
        RECT 59.070 143.500 59.330 143.820 ;
        RECT 60.910 143.500 61.170 143.820 ;
        RECT 61.370 143.500 61.630 143.820 ;
        RECT 59.130 141.440 59.270 143.500 ;
        RECT 59.070 141.120 59.330 141.440 ;
        RECT 60.970 127.840 61.110 143.500 ;
        RECT 61.890 141.440 62.030 143.840 ;
        RECT 62.810 143.560 62.950 143.840 ;
        RECT 62.350 143.420 62.950 143.560 ;
        RECT 61.830 141.120 62.090 141.440 ;
        RECT 61.890 139.060 62.030 141.120 ;
        RECT 62.350 139.400 62.490 143.420 ;
        RECT 63.730 143.140 63.870 144.180 ;
        RECT 67.410 144.160 67.550 166.280 ;
        RECT 68.330 163.880 68.470 183.620 ;
        RECT 68.790 181.900 68.930 183.620 ;
        RECT 69.250 182.920 69.390 184.640 ;
        RECT 69.190 182.600 69.450 182.920 ;
        RECT 71.090 182.580 71.230 184.640 ;
        RECT 71.030 182.260 71.290 182.580 ;
        RECT 69.190 181.920 69.450 182.240 ;
        RECT 68.730 181.580 68.990 181.900 ;
        RECT 68.790 180.200 68.930 181.580 ;
        RECT 68.730 179.880 68.990 180.200 ;
        RECT 68.730 178.860 68.990 179.180 ;
        RECT 68.790 176.120 68.930 178.860 ;
        RECT 69.250 176.800 69.390 181.920 ;
        RECT 69.650 179.880 69.910 180.200 ;
        RECT 69.710 179.520 69.850 179.880 ;
        RECT 69.650 179.200 69.910 179.520 ;
        RECT 69.190 176.480 69.450 176.800 ;
        RECT 68.730 175.800 68.990 176.120 ;
        RECT 68.790 174.080 68.930 175.800 ;
        RECT 69.190 174.440 69.450 174.760 ;
        RECT 69.250 174.080 69.390 174.440 ;
        RECT 68.730 173.760 68.990 174.080 ;
        RECT 69.190 173.760 69.450 174.080 ;
        RECT 68.790 171.020 68.930 173.760 ;
        RECT 69.250 172.040 69.390 173.760 ;
        RECT 69.190 171.720 69.450 172.040 ;
        RECT 68.730 170.700 68.990 171.020 ;
        RECT 69.250 168.640 69.390 171.720 ;
        RECT 69.710 171.700 69.850 179.200 ;
        RECT 71.090 177.140 71.230 182.260 ;
        RECT 71.550 181.560 71.690 188.040 ;
        RECT 72.470 184.280 72.610 189.740 ;
        RECT 72.930 184.960 73.070 195.180 ;
        RECT 73.330 194.500 73.590 194.820 ;
        RECT 73.390 193.120 73.530 194.500 ;
        RECT 74.770 193.800 74.910 195.520 ;
        RECT 77.470 194.500 77.730 194.820 ;
        RECT 74.710 193.480 74.970 193.800 ;
        RECT 73.330 192.800 73.590 193.120 ;
        RECT 74.770 192.360 74.910 193.480 ;
        RECT 77.530 193.460 77.670 194.500 ;
        RECT 78.410 193.965 80.290 194.335 ;
        RECT 77.470 193.140 77.730 193.460 ;
        RECT 80.690 192.460 80.950 192.780 ;
        RECT 74.770 192.220 75.370 192.360 ;
        RECT 75.230 189.720 75.370 192.220 ;
        RECT 75.170 189.400 75.430 189.720 ;
        RECT 73.790 189.060 74.050 189.380 ;
        RECT 72.870 184.640 73.130 184.960 ;
        RECT 73.850 184.620 73.990 189.060 ;
        RECT 78.410 188.525 80.290 188.895 ;
        RECT 75.630 187.700 75.890 188.020 ;
        RECT 75.690 185.300 75.830 187.700 ;
        RECT 80.750 187.340 80.890 192.460 ;
        RECT 83.510 192.360 83.650 196.200 ;
        RECT 90.810 195.180 91.070 195.500 ;
        RECT 90.350 193.140 90.610 193.460 ;
        RECT 86.670 192.460 86.930 192.780 ;
        RECT 83.050 192.220 83.650 192.360 ;
        RECT 78.850 187.020 79.110 187.340 ;
        RECT 80.690 187.020 80.950 187.340 ;
        RECT 78.910 185.640 79.050 187.020 ;
        RECT 78.850 185.320 79.110 185.640 ;
        RECT 75.630 184.980 75.890 185.300 ;
        RECT 73.790 184.300 74.050 184.620 ;
        RECT 75.630 184.300 75.890 184.620 ;
        RECT 72.410 183.960 72.670 184.280 ;
        RECT 75.690 182.240 75.830 184.300 ;
        RECT 78.410 183.085 80.290 183.455 ;
        RECT 75.630 181.920 75.890 182.240 ;
        RECT 71.490 181.240 71.750 181.560 ;
        RECT 73.790 180.900 74.050 181.220 ;
        RECT 75.170 180.900 75.430 181.220 ;
        RECT 73.850 179.520 73.990 180.900 ;
        RECT 73.790 179.200 74.050 179.520 ;
        RECT 75.230 178.840 75.370 180.900 ;
        RECT 75.170 178.520 75.430 178.840 ;
        RECT 75.690 177.140 75.830 181.920 ;
        RECT 80.750 179.520 80.890 187.020 ;
        RECT 82.530 183.620 82.790 183.940 ;
        RECT 82.590 181.220 82.730 183.620 ;
        RECT 82.530 180.900 82.790 181.220 ;
        RECT 80.690 179.200 80.950 179.520 ;
        RECT 77.470 178.180 77.730 178.500 ;
        RECT 71.030 176.820 71.290 177.140 ;
        RECT 75.630 176.820 75.890 177.140 ;
        RECT 70.110 176.480 70.370 176.800 ;
        RECT 69.650 171.380 69.910 171.700 ;
        RECT 70.170 170.680 70.310 176.480 ;
        RECT 70.570 176.140 70.830 176.460 ;
        RECT 70.630 172.235 70.770 176.140 ;
        RECT 71.090 173.740 71.230 176.820 ;
        RECT 77.530 176.800 77.670 178.180 ;
        RECT 78.410 177.645 80.290 178.015 ;
        RECT 77.470 176.480 77.730 176.800 ;
        RECT 81.610 176.480 81.870 176.800 ;
        RECT 82.070 176.480 82.330 176.800 ;
        RECT 77.470 175.460 77.730 175.780 ;
        RECT 75.630 174.440 75.890 174.760 ;
        RECT 71.030 173.420 71.290 173.740 ;
        RECT 70.560 171.865 70.840 172.235 ;
        RECT 71.090 171.700 71.230 173.420 ;
        RECT 71.490 173.080 71.750 173.400 ;
        RECT 71.030 171.380 71.290 171.700 ;
        RECT 70.570 171.040 70.830 171.360 ;
        RECT 69.650 170.360 69.910 170.680 ;
        RECT 70.110 170.360 70.370 170.680 ;
        RECT 69.710 170.080 69.850 170.360 ;
        RECT 69.710 169.940 70.310 170.080 ;
        RECT 69.190 168.320 69.450 168.640 ;
        RECT 69.190 167.640 69.450 167.960 ;
        RECT 68.270 163.560 68.530 163.880 ;
        RECT 68.330 157.330 68.470 163.560 ;
        RECT 69.250 162.860 69.390 167.640 ;
        RECT 70.170 167.620 70.310 169.940 ;
        RECT 70.110 167.300 70.370 167.620 ;
        RECT 70.170 165.920 70.310 167.300 ;
        RECT 70.110 165.600 70.370 165.920 ;
        RECT 70.170 162.860 70.310 165.600 ;
        RECT 70.630 163.200 70.770 171.040 ;
        RECT 71.090 168.980 71.230 171.380 ;
        RECT 71.030 168.660 71.290 168.980 ;
        RECT 70.570 162.880 70.830 163.200 ;
        RECT 69.190 162.540 69.450 162.860 ;
        RECT 70.110 162.540 70.370 162.860 ;
        RECT 69.250 157.760 69.390 162.540 ;
        RECT 70.170 160.480 70.310 162.540 ;
        RECT 70.110 160.160 70.370 160.480 ;
        RECT 69.190 157.440 69.450 157.760 ;
        RECT 68.730 157.330 68.990 157.420 ;
        RECT 68.330 157.190 68.990 157.330 ;
        RECT 68.330 155.040 68.470 157.190 ;
        RECT 68.730 157.100 68.990 157.190 ;
        RECT 69.650 156.420 69.910 156.740 ;
        RECT 69.710 155.380 69.850 156.420 ;
        RECT 69.650 155.060 69.910 155.380 ;
        RECT 70.170 155.040 70.310 160.160 ;
        RECT 68.270 154.720 68.530 155.040 ;
        RECT 70.110 154.720 70.370 155.040 ;
        RECT 69.180 154.185 69.460 154.555 ;
        RECT 69.190 154.040 69.450 154.185 ;
        RECT 67.810 152.000 68.070 152.320 ;
        RECT 67.350 143.840 67.610 144.160 ;
        RECT 65.510 143.160 65.770 143.480 ;
        RECT 62.750 142.820 63.010 143.140 ;
        RECT 63.670 142.820 63.930 143.140 ;
        RECT 62.810 140.760 62.950 142.820 ;
        RECT 63.410 142.285 65.290 142.655 ;
        RECT 65.570 142.120 65.710 143.160 ;
        RECT 65.510 141.800 65.770 142.120 ;
        RECT 67.410 141.780 67.550 143.840 ;
        RECT 67.350 141.460 67.610 141.780 ;
        RECT 65.510 141.120 65.770 141.440 ;
        RECT 62.750 140.440 63.010 140.760 ;
        RECT 62.290 139.080 62.550 139.400 ;
        RECT 61.830 138.740 62.090 139.060 ;
        RECT 61.830 138.060 62.090 138.380 ;
        RECT 61.890 129.880 62.030 138.060 ;
        RECT 63.410 136.845 65.290 137.215 ;
        RECT 65.050 135.680 65.310 136.000 ;
        RECT 65.110 132.170 65.250 135.680 ;
        RECT 65.570 135.660 65.710 141.120 ;
        RECT 65.970 138.740 66.230 139.060 ;
        RECT 66.030 135.660 66.170 138.740 ;
        RECT 67.410 138.720 67.550 141.460 ;
        RECT 67.350 138.400 67.610 138.720 ;
        RECT 66.430 137.380 66.690 137.700 ;
        RECT 65.510 135.340 65.770 135.660 ;
        RECT 65.970 135.340 66.230 135.660 ;
        RECT 65.110 132.030 65.710 132.170 ;
        RECT 63.410 131.405 65.290 131.775 ;
        RECT 65.570 130.560 65.710 132.030 ;
        RECT 65.510 130.240 65.770 130.560 ;
        RECT 62.750 129.900 63.010 130.220 ;
        RECT 61.830 129.560 62.090 129.880 ;
        RECT 59.990 127.520 60.250 127.840 ;
        RECT 60.910 127.520 61.170 127.840 ;
        RECT 58.610 127.180 58.870 127.500 ;
        RECT 58.670 124.780 58.810 127.180 ;
        RECT 60.050 125.120 60.190 127.520 ;
        RECT 59.990 124.800 60.250 125.120 ;
        RECT 58.610 124.460 58.870 124.780 ;
        RECT 58.670 123.080 58.810 124.460 ;
        RECT 58.610 122.760 58.870 123.080 ;
        RECT 59.530 122.420 59.790 122.740 ;
        RECT 59.590 120.360 59.730 122.420 ;
        RECT 59.530 120.040 59.790 120.360 ;
        RECT 60.970 119.340 61.110 127.520 ;
        RECT 61.890 125.120 62.030 129.560 ;
        RECT 61.830 124.800 62.090 125.120 ;
        RECT 61.370 123.780 61.630 124.100 ;
        RECT 61.430 122.400 61.570 123.780 ;
        RECT 61.370 122.080 61.630 122.400 ;
        RECT 60.910 119.020 61.170 119.340 ;
        RECT 60.970 116.960 61.110 119.020 ;
        RECT 60.910 116.640 61.170 116.960 ;
        RECT 60.970 116.460 61.110 116.640 ;
        RECT 60.970 116.320 61.570 116.460 ;
        RECT 58.150 112.900 58.410 113.220 ;
        RECT 60.450 111.200 60.710 111.520 ;
        RECT 27.330 105.760 27.590 106.080 ;
        RECT 28.710 105.760 28.970 106.080 ;
        RECT 37.910 105.760 38.170 106.080 ;
        RECT 43.430 105.760 43.690 106.080 ;
        RECT 57.230 105.760 57.490 106.080 ;
        RECT 21.350 105.420 21.610 105.740 ;
        RECT 31.930 105.420 32.190 105.740 ;
        RECT 44.350 105.420 44.610 105.740 ;
        RECT 54.930 105.420 55.190 105.740 ;
        RECT 17.670 105.080 17.930 105.400 ;
        RECT 15.830 103.720 16.090 104.040 ;
        RECT 17.730 102.340 17.870 105.080 ;
        RECT 21.410 104.040 21.550 105.420 ;
        RECT 24.110 104.740 24.370 105.060 ;
        RECT 27.790 104.740 28.050 105.060 ;
        RECT 21.350 103.720 21.610 104.040 ;
        RECT 20.890 103.040 21.150 103.360 ;
        RECT 20.430 102.360 20.690 102.680 ;
        RECT 17.670 102.020 17.930 102.340 ;
        RECT 17.730 100.640 17.870 102.020 ;
        RECT 18.410 101.485 20.290 101.855 ;
        RECT 20.490 101.320 20.630 102.360 ;
        RECT 20.430 101.000 20.690 101.320 ;
        RECT 17.670 100.320 17.930 100.640 ;
        RECT 18.410 96.045 20.290 96.415 ;
        RECT 20.950 89.850 21.090 103.040 ;
        RECT 21.410 100.980 21.550 103.720 ;
        RECT 24.170 103.360 24.310 104.740 ;
        RECT 24.110 103.040 24.370 103.360 ;
        RECT 27.330 102.700 27.590 103.020 ;
        RECT 21.350 100.660 21.610 100.980 ;
        RECT 27.390 100.640 27.530 102.700 ;
        RECT 27.330 100.320 27.590 100.640 ;
        RECT 27.850 100.300 27.990 104.740 ;
        RECT 31.990 103.020 32.130 105.420 ;
        RECT 36.990 104.740 37.250 105.060 ;
        RECT 40.210 104.740 40.470 105.060 ;
        RECT 41.590 104.740 41.850 105.060 ;
        RECT 33.410 104.205 35.290 104.575 ;
        RECT 31.930 102.700 32.190 103.020 ;
        RECT 31.930 102.020 32.190 102.340 ;
        RECT 31.990 100.980 32.130 102.020 ;
        RECT 37.050 100.980 37.190 104.740 ;
        RECT 38.370 103.720 38.630 104.040 ;
        RECT 31.930 100.660 32.190 100.980 ;
        RECT 36.990 100.660 37.250 100.980 ;
        RECT 38.430 100.640 38.570 103.720 ;
        RECT 40.270 103.020 40.410 104.740 ;
        RECT 41.650 103.700 41.790 104.740 ;
        RECT 41.590 103.380 41.850 103.700 ;
        RECT 40.670 103.040 40.930 103.360 ;
        RECT 40.210 102.700 40.470 103.020 ;
        RECT 38.370 100.320 38.630 100.640 ;
        RECT 27.790 99.980 28.050 100.300 ;
        RECT 27.330 99.300 27.590 99.620 ;
        RECT 31.930 99.300 32.190 99.620 ;
        RECT 8.000 84.920 8.280 86.920 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 86.920 21.130 89.850 ;
        RECT 19.910 85.980 21.160 86.920 ;
        RECT 14.440 84.920 14.720 85.550 ;
        RECT 20.880 84.920 21.160 85.980 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 27.390 86.920 27.530 99.300 ;
        RECT 31.990 89.380 32.130 99.300 ;
        RECT 33.410 98.765 35.290 99.135 ;
        RECT 27.320 84.920 27.600 86.920 ;
        RECT 31.780 86.440 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 33.760 86.440 34.040 86.920 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 31.780 86.300 34.040 86.440 ;
        RECT 31.780 85.510 33.000 86.300 ;
        RECT 33.760 84.920 34.040 86.300 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 40.200 86.440 40.480 86.920 ;
        RECT 40.730 86.440 40.870 103.040 ;
        RECT 44.410 100.640 44.550 105.420 ;
        RECT 46.190 104.740 46.450 105.060 ;
        RECT 47.570 104.740 47.830 105.060 ;
        RECT 46.250 103.360 46.390 104.740 ;
        RECT 46.650 103.720 46.910 104.040 ;
        RECT 46.190 103.040 46.450 103.360 ;
        RECT 44.810 102.360 45.070 102.680 ;
        RECT 44.870 101.320 45.010 102.360 ;
        RECT 44.810 101.000 45.070 101.320 ;
        RECT 44.350 100.320 44.610 100.640 ;
        RECT 40.200 86.300 40.870 86.440 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 46.710 86.920 46.850 103.720 ;
        RECT 47.630 100.980 47.770 104.740 ;
        RECT 54.990 103.020 55.130 105.420 ;
        RECT 58.610 104.740 58.870 105.060 ;
        RECT 51.250 102.700 51.510 103.020 ;
        RECT 54.470 102.700 54.730 103.020 ;
        RECT 54.930 102.700 55.190 103.020 ;
        RECT 48.410 101.485 50.290 101.855 ;
        RECT 47.570 100.660 47.830 100.980 ;
        RECT 51.310 100.300 51.450 102.700 ;
        RECT 54.530 100.980 54.670 102.700 ;
        RECT 57.690 102.020 57.950 102.340 ;
        RECT 57.750 100.980 57.890 102.020 ;
        RECT 58.670 101.320 58.810 104.740 ;
        RECT 60.510 103.360 60.650 111.200 ;
        RECT 61.430 108.460 61.570 116.320 ;
        RECT 61.890 114.920 62.030 124.800 ;
        RECT 62.290 123.780 62.550 124.100 ;
        RECT 62.350 119.340 62.490 123.780 ;
        RECT 62.810 122.400 62.950 129.900 ;
        RECT 63.410 125.965 65.290 126.335 ;
        RECT 65.050 125.480 65.310 125.800 ;
        RECT 65.110 122.400 65.250 125.480 ;
        RECT 66.490 125.120 66.630 137.380 ;
        RECT 67.410 135.660 67.550 138.400 ;
        RECT 67.870 137.700 68.010 152.000 ;
        RECT 70.170 151.980 70.310 154.720 ;
        RECT 70.630 152.320 70.770 162.880 ;
        RECT 71.030 161.860 71.290 162.180 ;
        RECT 71.090 160.820 71.230 161.860 ;
        RECT 71.030 160.500 71.290 160.820 ;
        RECT 71.030 156.420 71.290 156.740 ;
        RECT 71.090 155.235 71.230 156.420 ;
        RECT 71.020 154.865 71.300 155.235 ;
        RECT 70.570 152.000 70.830 152.320 ;
        RECT 70.110 151.660 70.370 151.980 ;
        RECT 71.030 151.660 71.290 151.980 ;
        RECT 68.270 150.980 68.530 151.300 ;
        RECT 70.110 150.980 70.370 151.300 ;
        RECT 68.330 150.280 68.470 150.980 ;
        RECT 68.270 149.960 68.530 150.280 ;
        RECT 68.330 138.380 68.470 149.960 ;
        RECT 70.170 146.880 70.310 150.980 ;
        RECT 71.090 149.600 71.230 151.660 ;
        RECT 71.030 149.280 71.290 149.600 ;
        RECT 71.550 149.000 71.690 173.080 ;
        RECT 72.870 170.700 73.130 171.020 ;
        RECT 71.950 170.360 72.210 170.680 ;
        RECT 72.010 168.640 72.150 170.360 ;
        RECT 72.410 170.020 72.670 170.340 ;
        RECT 71.950 168.320 72.210 168.640 ;
        RECT 72.470 153.000 72.610 170.020 ;
        RECT 72.930 168.300 73.070 170.700 ;
        RECT 72.870 167.980 73.130 168.300 ;
        RECT 75.690 164.760 75.830 174.440 ;
        RECT 76.550 172.740 76.810 173.060 ;
        RECT 76.090 170.020 76.350 170.340 ;
        RECT 75.230 164.620 75.830 164.760 ;
        RECT 74.710 161.860 74.970 162.180 ;
        RECT 72.860 154.865 73.140 155.235 ;
        RECT 74.250 155.060 74.510 155.380 ;
        RECT 72.410 152.680 72.670 153.000 ;
        RECT 71.090 148.860 71.690 149.000 ;
        RECT 71.950 149.170 72.210 149.260 ;
        RECT 72.470 149.170 72.610 152.680 ;
        RECT 72.930 151.300 73.070 154.865 ;
        RECT 73.780 154.185 74.060 154.555 ;
        RECT 73.850 152.660 73.990 154.185 ;
        RECT 73.790 152.340 74.050 152.660 ;
        RECT 73.850 151.980 73.990 152.340 ;
        RECT 73.790 151.660 74.050 151.980 ;
        RECT 74.310 151.640 74.450 155.060 ;
        RECT 74.770 151.980 74.910 161.860 ;
        RECT 74.710 151.660 74.970 151.980 ;
        RECT 73.330 151.320 73.590 151.640 ;
        RECT 74.250 151.320 74.510 151.640 ;
        RECT 72.870 150.980 73.130 151.300 ;
        RECT 72.930 149.600 73.070 150.980 ;
        RECT 73.390 149.940 73.530 151.320 ;
        RECT 73.330 149.620 73.590 149.940 ;
        RECT 72.870 149.280 73.130 149.600 ;
        RECT 71.950 149.030 72.610 149.170 ;
        RECT 71.950 148.940 72.210 149.030 ;
        RECT 70.110 146.560 70.370 146.880 ;
        RECT 68.730 145.880 68.990 146.200 ;
        RECT 68.790 138.915 68.930 145.880 ;
        RECT 70.170 143.820 70.310 146.560 ;
        RECT 70.110 143.500 70.370 143.820 ;
        RECT 70.570 140.780 70.830 141.100 ;
        RECT 69.190 140.440 69.450 140.760 ;
        RECT 68.720 138.545 69.000 138.915 ;
        RECT 68.270 138.060 68.530 138.380 ;
        RECT 69.250 137.700 69.390 140.440 ;
        RECT 70.630 137.700 70.770 140.780 ;
        RECT 67.810 137.380 68.070 137.700 ;
        RECT 69.190 137.380 69.450 137.700 ;
        RECT 70.570 137.380 70.830 137.700 ;
        RECT 69.250 136.000 69.390 137.380 ;
        RECT 69.190 135.680 69.450 136.000 ;
        RECT 66.890 135.340 67.150 135.660 ;
        RECT 67.350 135.340 67.610 135.660 ;
        RECT 66.950 129.540 67.090 135.340 ;
        RECT 70.630 134.980 70.770 137.380 ;
        RECT 70.570 134.660 70.830 134.980 ;
        RECT 66.890 129.220 67.150 129.540 ;
        RECT 66.950 128.520 67.090 129.220 ;
        RECT 66.890 128.200 67.150 128.520 ;
        RECT 66.430 124.800 66.690 125.120 ;
        RECT 70.110 124.800 70.370 125.120 ;
        RECT 68.270 123.780 68.530 124.100 ;
        RECT 68.330 122.740 68.470 123.780 ;
        RECT 68.270 122.420 68.530 122.740 ;
        RECT 62.750 122.080 63.010 122.400 ;
        RECT 65.050 122.080 65.310 122.400 ;
        RECT 62.290 119.020 62.550 119.340 ;
        RECT 61.830 114.600 62.090 114.920 ;
        RECT 62.810 114.240 62.950 122.080 ;
        RECT 63.410 120.525 65.290 120.895 ;
        RECT 65.510 118.340 65.770 118.660 ;
        RECT 65.570 117.040 65.710 118.340 ;
        RECT 65.570 116.900 66.630 117.040 ;
        RECT 65.510 116.300 65.770 116.620 ;
        RECT 63.410 115.085 65.290 115.455 ;
        RECT 62.750 113.920 63.010 114.240 ;
        RECT 62.810 111.520 62.950 113.920 ;
        RECT 65.570 113.560 65.710 116.300 ;
        RECT 66.490 114.240 66.630 116.900 ;
        RECT 66.430 113.920 66.690 114.240 ;
        RECT 65.510 113.240 65.770 113.560 ;
        RECT 62.750 111.200 63.010 111.520 ;
        RECT 63.410 109.645 65.290 110.015 ;
        RECT 61.370 108.140 61.630 108.460 ;
        RECT 61.430 106.080 61.570 108.140 ;
        RECT 70.170 106.760 70.310 124.800 ;
        RECT 71.090 124.780 71.230 148.860 ;
        RECT 72.470 146.540 72.610 149.030 ;
        RECT 74.710 146.900 74.970 147.220 ;
        RECT 72.410 146.220 72.670 146.540 ;
        RECT 74.770 144.500 74.910 146.900 ;
        RECT 74.710 144.180 74.970 144.500 ;
        RECT 72.410 142.820 72.670 143.140 ;
        RECT 72.470 141.780 72.610 142.820 ;
        RECT 72.410 141.460 72.670 141.780 ;
        RECT 71.490 141.120 71.750 141.440 ;
        RECT 71.550 139.400 71.690 141.120 ;
        RECT 71.950 140.780 72.210 141.100 ;
        RECT 71.490 139.080 71.750 139.400 ;
        RECT 72.010 138.380 72.150 140.780 ;
        RECT 72.870 140.100 73.130 140.420 ;
        RECT 72.930 139.060 73.070 140.100 ;
        RECT 72.870 138.740 73.130 139.060 ;
        RECT 71.950 138.060 72.210 138.380 ;
        RECT 74.250 138.060 74.510 138.380 ;
        RECT 74.310 136.680 74.450 138.060 ;
        RECT 74.250 136.360 74.510 136.680 ;
        RECT 72.870 129.220 73.130 129.540 ;
        RECT 72.930 127.840 73.070 129.220 ;
        RECT 72.870 127.520 73.130 127.840 ;
        RECT 75.230 127.500 75.370 164.620 ;
        RECT 75.630 153.700 75.890 154.020 ;
        RECT 75.690 130.220 75.830 153.700 ;
        RECT 76.150 130.220 76.290 170.020 ;
        RECT 76.610 141.440 76.750 172.740 ;
        RECT 77.010 162.540 77.270 162.860 ;
        RECT 77.070 160.820 77.210 162.540 ;
        RECT 77.010 160.500 77.270 160.820 ;
        RECT 77.010 150.980 77.270 151.300 ;
        RECT 76.550 141.120 76.810 141.440 ;
        RECT 77.070 141.100 77.210 150.980 ;
        RECT 77.530 146.880 77.670 175.460 ;
        RECT 81.670 173.740 81.810 176.480 ;
        RECT 82.130 173.740 82.270 176.480 ;
        RECT 81.610 173.420 81.870 173.740 ;
        RECT 82.070 173.420 82.330 173.740 ;
        RECT 78.410 172.205 80.290 172.575 ;
        RECT 81.670 171.360 81.810 173.420 ;
        RECT 82.130 171.360 82.270 173.420 ;
        RECT 82.590 171.360 82.730 180.900 ;
        RECT 83.050 176.800 83.190 192.220 ;
        RECT 84.370 192.010 84.630 192.100 ;
        RECT 84.370 191.870 85.030 192.010 ;
        RECT 84.370 191.780 84.630 191.870 ;
        RECT 84.890 189.380 85.030 191.870 ;
        RECT 84.830 189.060 85.090 189.380 ;
        RECT 84.890 187.680 85.030 189.060 ;
        RECT 84.830 187.360 85.090 187.680 ;
        RECT 82.990 176.480 83.250 176.800 ;
        RECT 83.450 176.480 83.710 176.800 ;
        RECT 83.510 173.740 83.650 176.480 ;
        RECT 84.890 174.080 85.030 187.360 ;
        RECT 86.730 181.900 86.870 192.460 ;
        RECT 90.410 191.080 90.550 193.140 ;
        RECT 90.870 193.120 91.010 195.180 ;
        RECT 90.810 192.800 91.070 193.120 ;
        RECT 91.330 192.440 91.470 196.200 ;
        RECT 93.570 195.520 93.830 195.840 ;
        RECT 92.650 195.180 92.910 195.500 ;
        RECT 91.730 194.500 91.990 194.820 ;
        RECT 91.790 193.800 91.930 194.500 ;
        RECT 91.730 193.480 91.990 193.800 ;
        RECT 92.190 192.460 92.450 192.780 ;
        RECT 91.270 192.360 91.530 192.440 ;
        RECT 90.870 192.220 91.530 192.360 ;
        RECT 90.350 190.760 90.610 191.080 ;
        RECT 90.870 190.400 91.010 192.220 ;
        RECT 91.270 192.120 91.530 192.220 ;
        RECT 92.250 190.740 92.390 192.460 ;
        RECT 92.190 190.420 92.450 190.740 ;
        RECT 92.710 190.400 92.850 195.180 ;
        RECT 93.630 193.800 93.770 195.520 ;
        RECT 98.690 195.160 98.830 197.220 ;
        RECT 98.630 194.840 98.890 195.160 ;
        RECT 96.790 194.500 97.050 194.820 ;
        RECT 93.570 193.480 93.830 193.800 ;
        RECT 95.870 193.140 96.130 193.460 ;
        RECT 93.410 191.245 95.290 191.615 ;
        RECT 87.130 190.080 87.390 190.400 ;
        RECT 90.810 190.080 91.070 190.400 ;
        RECT 92.650 190.080 92.910 190.400 ;
        RECT 87.190 187.000 87.330 190.080 ;
        RECT 91.270 189.740 91.530 190.060 ;
        RECT 91.330 188.360 91.470 189.740 ;
        RECT 95.410 189.400 95.670 189.720 ;
        RECT 95.470 188.360 95.610 189.400 ;
        RECT 91.270 188.040 91.530 188.360 ;
        RECT 95.410 188.040 95.670 188.360 ;
        RECT 87.590 187.360 87.850 187.680 ;
        RECT 87.130 186.680 87.390 187.000 ;
        RECT 87.190 184.960 87.330 186.680 ;
        RECT 87.130 184.640 87.390 184.960 ;
        RECT 86.670 181.580 86.930 181.900 ;
        RECT 87.190 180.200 87.330 184.640 ;
        RECT 87.650 183.940 87.790 187.360 ;
        RECT 93.410 185.805 95.290 186.175 ;
        RECT 87.590 183.620 87.850 183.940 ;
        RECT 88.510 183.620 88.770 183.940 ;
        RECT 90.350 183.620 90.610 183.940 ;
        RECT 88.050 182.260 88.310 182.580 ;
        RECT 88.110 180.200 88.250 182.260 ;
        RECT 88.570 181.220 88.710 183.620 ;
        RECT 90.410 182.240 90.550 183.620 ;
        RECT 90.350 181.920 90.610 182.240 ;
        RECT 91.270 181.580 91.530 181.900 ;
        RECT 88.510 180.900 88.770 181.220 ;
        RECT 87.130 179.880 87.390 180.200 ;
        RECT 88.050 179.880 88.310 180.200 ;
        RECT 88.570 174.080 88.710 180.900 ;
        RECT 84.830 173.760 85.090 174.080 ;
        RECT 88.510 173.760 88.770 174.080 ;
        RECT 83.450 173.420 83.710 173.740 ;
        RECT 83.510 173.060 83.650 173.420 ;
        RECT 83.450 172.740 83.710 173.060 ;
        RECT 83.510 171.360 83.650 172.740 ;
        RECT 91.330 171.360 91.470 181.580 ;
        RECT 93.410 180.365 95.290 180.735 ;
        RECT 95.930 179.180 96.070 193.140 ;
        RECT 96.850 192.780 96.990 194.500 ;
        RECT 100.530 193.800 100.670 198.240 ;
        RECT 111.050 197.900 111.310 198.220 ;
        RECT 101.390 197.220 101.650 197.540 ;
        RECT 101.450 195.840 101.590 197.220 ;
        RECT 101.390 195.520 101.650 195.840 ;
        RECT 111.110 195.500 111.250 197.900 ;
        RECT 115.190 197.220 115.450 197.540 ;
        RECT 102.770 195.180 103.030 195.500 ;
        RECT 111.050 195.180 111.310 195.500 ;
        RECT 100.470 193.480 100.730 193.800 ;
        RECT 102.830 192.780 102.970 195.180 ;
        RECT 115.250 195.160 115.390 197.220 ;
        RECT 115.190 194.840 115.450 195.160 ;
        RECT 110.590 194.500 110.850 194.820 ;
        RECT 111.510 194.500 111.770 194.820 ;
        RECT 108.410 193.965 110.290 194.335 ;
        RECT 110.650 193.460 110.790 194.500 ;
        RECT 110.590 193.140 110.850 193.460 ;
        RECT 107.830 192.800 108.090 193.120 ;
        RECT 96.330 192.460 96.590 192.780 ;
        RECT 96.790 192.460 97.050 192.780 ;
        RECT 100.930 192.460 101.190 192.780 ;
        RECT 102.770 192.460 103.030 192.780 ;
        RECT 96.390 184.960 96.530 192.460 ;
        RECT 100.990 190.060 101.130 192.460 ;
        RECT 100.930 189.740 101.190 190.060 ;
        RECT 102.310 189.060 102.570 189.380 ;
        RECT 102.370 188.360 102.510 189.060 ;
        RECT 102.310 188.040 102.570 188.360 ;
        RECT 96.330 184.640 96.590 184.960 ;
        RECT 102.370 184.280 102.510 188.040 ;
        RECT 100.930 183.960 101.190 184.280 ;
        RECT 102.310 183.960 102.570 184.280 ;
        RECT 99.550 183.620 99.810 183.940 ;
        RECT 96.330 182.260 96.590 182.580 ;
        RECT 96.390 180.200 96.530 182.260 ;
        RECT 96.330 179.880 96.590 180.200 ;
        RECT 99.610 179.180 99.750 183.620 ;
        RECT 100.010 181.580 100.270 181.900 ;
        RECT 100.070 180.200 100.210 181.580 ;
        RECT 100.010 179.880 100.270 180.200 ;
        RECT 95.870 178.860 96.130 179.180 ;
        RECT 99.550 178.860 99.810 179.180 ;
        RECT 95.930 177.140 96.070 178.860 ;
        RECT 95.870 176.820 96.130 177.140 ;
        RECT 93.410 174.925 95.290 175.295 ;
        RECT 95.930 173.740 96.070 176.820 ;
        RECT 100.990 176.800 101.130 183.960 ;
        RECT 102.830 182.240 102.970 192.460 ;
        RECT 106.910 191.780 107.170 192.100 ;
        RECT 106.970 187.680 107.110 191.780 ;
        RECT 107.890 189.380 108.030 192.800 ;
        RECT 110.590 190.080 110.850 190.400 ;
        RECT 107.830 189.060 108.090 189.380 ;
        RECT 106.910 187.360 107.170 187.680 ;
        RECT 102.770 181.920 103.030 182.240 ;
        RECT 100.930 176.480 101.190 176.800 ;
        RECT 101.850 176.480 102.110 176.800 ;
        RECT 101.910 176.315 102.050 176.480 ;
        RECT 101.840 175.945 102.120 176.315 ;
        RECT 98.630 175.460 98.890 175.780 ;
        RECT 95.870 173.420 96.130 173.740 ;
        RECT 94.950 172.740 95.210 173.060 ;
        RECT 95.010 171.700 95.150 172.740 ;
        RECT 95.930 172.040 96.070 173.420 ;
        RECT 95.870 171.720 96.130 172.040 ;
        RECT 94.950 171.380 95.210 171.700 ;
        RECT 81.610 171.040 81.870 171.360 ;
        RECT 82.070 171.040 82.330 171.360 ;
        RECT 82.530 171.040 82.790 171.360 ;
        RECT 83.450 171.040 83.710 171.360 ;
        RECT 91.270 171.040 91.530 171.360 ;
        RECT 83.510 169.320 83.650 171.040 ;
        RECT 83.450 169.000 83.710 169.320 ;
        RECT 82.070 168.320 82.330 168.640 ;
        RECT 81.610 167.300 81.870 167.620 ;
        RECT 78.410 166.765 80.290 167.135 ;
        RECT 77.930 165.600 78.190 165.920 ;
        RECT 77.990 161.160 78.130 165.600 ;
        RECT 81.670 165.240 81.810 167.300 ;
        RECT 81.610 164.920 81.870 165.240 ;
        RECT 81.150 161.860 81.410 162.180 ;
        RECT 78.410 161.325 80.290 161.695 ;
        RECT 81.210 161.160 81.350 161.860 ;
        RECT 77.930 160.840 78.190 161.160 ;
        RECT 81.150 160.840 81.410 161.160 ;
        RECT 80.690 160.160 80.950 160.480 ;
        RECT 80.750 157.420 80.890 160.160 ;
        RECT 80.690 157.100 80.950 157.420 ;
        RECT 78.410 155.885 80.290 156.255 ;
        RECT 80.750 155.380 80.890 157.100 ;
        RECT 80.690 155.060 80.950 155.380 ;
        RECT 78.390 154.720 78.650 155.040 ;
        RECT 80.230 154.720 80.490 155.040 ;
        RECT 81.150 154.720 81.410 155.040 ;
        RECT 78.450 151.980 78.590 154.720 ;
        RECT 79.770 154.380 80.030 154.700 ;
        RECT 78.850 153.700 79.110 154.020 ;
        RECT 78.910 152.320 79.050 153.700 ;
        RECT 78.850 152.000 79.110 152.320 ;
        RECT 79.830 151.980 79.970 154.380 ;
        RECT 80.290 152.660 80.430 154.720 ;
        RECT 80.230 152.340 80.490 152.660 ;
        RECT 78.390 151.660 78.650 151.980 ;
        RECT 79.770 151.890 80.030 151.980 ;
        RECT 79.770 151.750 80.890 151.890 ;
        RECT 79.770 151.660 80.030 151.750 ;
        RECT 77.930 150.980 78.190 151.300 ;
        RECT 77.470 146.560 77.730 146.880 ;
        RECT 77.990 146.540 78.130 150.980 ;
        RECT 78.410 150.445 80.290 150.815 ;
        RECT 80.230 149.510 80.490 149.600 ;
        RECT 80.750 149.510 80.890 151.750 ;
        RECT 81.210 149.600 81.350 154.720 ;
        RECT 81.670 152.320 81.810 164.920 ;
        RECT 82.130 164.760 82.270 168.320 ;
        RECT 87.130 167.980 87.390 168.300 ;
        RECT 82.990 167.300 83.250 167.620 ;
        RECT 84.830 167.300 85.090 167.620 ;
        RECT 86.210 167.300 86.470 167.620 ;
        RECT 82.130 164.620 82.730 164.760 ;
        RECT 82.590 163.200 82.730 164.620 ;
        RECT 82.530 162.880 82.790 163.200 ;
        RECT 82.590 160.140 82.730 162.880 ;
        RECT 83.050 162.180 83.190 167.300 ;
        RECT 84.890 166.600 85.030 167.300 ;
        RECT 84.830 166.280 85.090 166.600 ;
        RECT 86.270 166.260 86.410 167.300 ;
        RECT 86.210 165.940 86.470 166.260 ;
        RECT 85.290 164.580 85.550 164.900 ;
        RECT 85.350 163.200 85.490 164.580 ;
        RECT 85.290 162.880 85.550 163.200 ;
        RECT 82.990 161.860 83.250 162.180 ;
        RECT 87.190 160.820 87.330 167.980 ;
        RECT 91.330 165.920 91.470 171.040 ;
        RECT 92.650 170.700 92.910 171.020 ;
        RECT 92.710 169.320 92.850 170.700 ;
        RECT 95.410 170.020 95.670 170.340 ;
        RECT 93.410 169.485 95.290 169.855 ;
        RECT 92.650 169.000 92.910 169.320 ;
        RECT 95.470 168.640 95.610 170.020 ;
        RECT 95.410 168.320 95.670 168.640 ;
        RECT 91.270 165.600 91.530 165.920 ;
        RECT 96.330 165.600 96.590 165.920 ;
        RECT 91.330 163.880 91.470 165.600 ;
        RECT 93.410 164.045 95.290 164.415 ;
        RECT 91.270 163.560 91.530 163.880 ;
        RECT 89.430 162.880 89.690 163.200 ;
        RECT 87.130 160.500 87.390 160.820 ;
        RECT 89.490 160.480 89.630 162.880 ;
        RECT 96.390 162.860 96.530 165.600 ;
        RECT 96.330 162.540 96.590 162.860 ;
        RECT 85.750 160.160 86.010 160.480 ;
        RECT 89.430 160.160 89.690 160.480 ;
        RECT 95.410 160.160 95.670 160.480 ;
        RECT 82.530 159.820 82.790 160.140 ;
        RECT 82.590 154.700 82.730 159.820 ;
        RECT 84.830 159.140 85.090 159.460 ;
        RECT 84.890 157.080 85.030 159.140 ;
        RECT 85.810 157.840 85.950 160.160 ;
        RECT 87.590 159.140 87.850 159.460 ;
        RECT 85.350 157.700 85.950 157.840 ;
        RECT 87.650 157.760 87.790 159.140 ;
        RECT 89.490 157.760 89.630 160.160 ;
        RECT 93.410 158.605 95.290 158.975 ;
        RECT 84.830 156.760 85.090 157.080 ;
        RECT 83.450 156.420 83.710 156.740 ;
        RECT 83.510 155.040 83.650 156.420 ;
        RECT 85.350 155.720 85.490 157.700 ;
        RECT 86.670 157.440 86.930 157.760 ;
        RECT 87.590 157.440 87.850 157.760 ;
        RECT 89.430 157.440 89.690 157.760 ;
        RECT 85.290 155.400 85.550 155.720 ;
        RECT 83.450 154.720 83.710 155.040 ;
        RECT 82.530 154.380 82.790 154.700 ;
        RECT 82.990 152.680 83.250 153.000 ;
        RECT 81.610 152.000 81.870 152.320 ;
        RECT 82.070 151.660 82.330 151.980 ;
        RECT 82.130 149.600 82.270 151.660 ;
        RECT 83.050 150.280 83.190 152.680 ;
        RECT 86.730 151.980 86.870 157.440 ;
        RECT 95.470 156.740 95.610 160.160 ;
        RECT 95.870 159.140 96.130 159.460 ;
        RECT 95.930 157.080 96.070 159.140 ;
        RECT 95.870 156.760 96.130 157.080 ;
        RECT 95.410 156.420 95.670 156.740 ;
        RECT 89.890 155.060 90.150 155.380 ;
        RECT 86.670 151.660 86.930 151.980 ;
        RECT 82.990 149.960 83.250 150.280 ;
        RECT 80.230 149.370 80.890 149.510 ;
        RECT 80.230 149.280 80.490 149.370 ;
        RECT 81.150 149.280 81.410 149.600 ;
        RECT 82.070 149.280 82.330 149.600 ;
        RECT 86.210 149.280 86.470 149.600 ;
        RECT 82.070 148.600 82.330 148.920 ;
        RECT 78.390 148.260 78.650 148.580 ;
        RECT 77.930 146.220 78.190 146.540 ;
        RECT 77.470 145.540 77.730 145.860 ;
        RECT 78.450 145.770 78.590 148.260 ;
        RECT 81.610 147.240 81.870 147.560 ;
        RECT 80.690 145.880 80.950 146.200 ;
        RECT 77.990 145.630 78.590 145.770 ;
        RECT 77.010 140.780 77.270 141.100 ;
        RECT 76.550 140.100 76.810 140.420 ;
        RECT 75.630 129.900 75.890 130.220 ;
        RECT 76.090 129.900 76.350 130.220 ;
        RECT 76.090 129.220 76.350 129.540 ;
        RECT 75.170 127.180 75.430 127.500 ;
        RECT 75.630 126.500 75.890 126.820 ;
        RECT 71.030 124.460 71.290 124.780 ;
        RECT 74.710 121.740 74.970 122.060 ;
        RECT 73.330 121.060 73.590 121.380 ;
        RECT 73.390 120.020 73.530 121.060 ;
        RECT 73.330 119.700 73.590 120.020 ;
        RECT 73.390 114.240 73.530 119.700 ;
        RECT 74.250 119.360 74.510 119.680 ;
        RECT 74.310 116.620 74.450 119.360 ;
        RECT 74.770 119.000 74.910 121.740 ;
        RECT 74.710 118.680 74.970 119.000 ;
        RECT 74.250 116.300 74.510 116.620 ;
        RECT 74.310 114.240 74.450 116.300 ;
        RECT 73.330 113.920 73.590 114.240 ;
        RECT 74.250 113.920 74.510 114.240 ;
        RECT 74.770 113.900 74.910 118.680 ;
        RECT 74.710 113.580 74.970 113.900 ;
        RECT 71.950 112.900 72.210 113.220 ;
        RECT 72.010 111.860 72.150 112.900 ;
        RECT 74.250 112.110 74.510 112.200 ;
        RECT 74.770 112.110 74.910 113.580 ;
        RECT 74.250 111.970 74.910 112.110 ;
        RECT 74.250 111.880 74.510 111.970 ;
        RECT 71.950 111.540 72.210 111.860 ;
        RECT 75.690 106.760 75.830 126.500 ;
        RECT 70.110 106.440 70.370 106.760 ;
        RECT 75.630 106.440 75.890 106.760 ;
        RECT 75.170 106.100 75.430 106.420 ;
        RECT 61.370 105.760 61.630 106.080 ;
        RECT 74.250 105.760 74.510 106.080 ;
        RECT 61.830 104.740 62.090 105.060 ;
        RECT 61.890 103.360 62.030 104.740 ;
        RECT 63.410 104.205 65.290 104.575 ;
        RECT 60.450 103.040 60.710 103.360 ;
        RECT 61.830 103.040 62.090 103.360 ;
        RECT 66.890 103.040 67.150 103.360 ;
        RECT 58.610 101.000 58.870 101.320 ;
        RECT 54.470 100.660 54.730 100.980 ;
        RECT 57.690 100.660 57.950 100.980 ;
        RECT 60.510 100.300 60.650 103.040 ;
        RECT 51.250 99.980 51.510 100.300 ;
        RECT 60.450 99.980 60.710 100.300 ;
        RECT 53.090 99.300 53.350 99.620 ;
        RECT 59.530 99.300 59.790 99.620 ;
        RECT 48.410 96.045 50.290 96.415 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 53.150 86.920 53.290 99.300 ;
        RECT 40.200 84.920 40.480 86.300 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 46.640 84.920 46.920 86.920 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 53.080 84.920 53.360 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 59.590 86.920 59.730 99.300 ;
        RECT 63.410 98.765 65.290 99.135 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 59.520 84.920 59.800 86.920 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 65.960 86.440 66.240 86.920 ;
        RECT 66.950 86.440 67.090 103.040 ;
        RECT 74.310 102.680 74.450 105.760 ;
        RECT 75.230 104.040 75.370 106.100 ;
        RECT 76.150 104.040 76.290 129.220 ;
        RECT 75.170 103.720 75.430 104.040 ;
        RECT 76.090 103.720 76.350 104.040 ;
        RECT 76.610 103.700 76.750 140.100 ;
        RECT 77.010 130.920 77.270 131.240 ;
        RECT 77.070 123.080 77.210 130.920 ;
        RECT 77.010 122.760 77.270 123.080 ;
        RECT 77.010 116.980 77.270 117.300 ;
        RECT 77.070 114.920 77.210 116.980 ;
        RECT 77.010 114.600 77.270 114.920 ;
        RECT 77.010 104.740 77.270 105.060 ;
        RECT 76.550 103.380 76.810 103.700 ;
        RECT 76.550 102.700 76.810 103.020 ;
        RECT 74.250 102.360 74.510 102.680 ;
        RECT 76.610 100.980 76.750 102.700 ;
        RECT 76.550 100.660 76.810 100.980 ;
        RECT 71.490 99.300 71.750 99.620 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 65.960 86.300 67.090 86.440 ;
        RECT 65.960 84.920 66.240 86.300 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 71.550 86.440 71.690 99.300 ;
        RECT 77.070 95.280 77.210 104.740 ;
        RECT 77.530 103.020 77.670 145.540 ;
        RECT 77.990 127.840 78.130 145.630 ;
        RECT 78.410 145.005 80.290 145.375 ;
        RECT 79.830 144.160 80.430 144.240 ;
        RECT 80.750 144.160 80.890 145.880 ;
        RECT 81.150 144.520 81.410 144.840 ;
        RECT 79.770 144.100 80.430 144.160 ;
        RECT 79.770 143.840 80.030 144.100 ;
        RECT 79.770 143.160 80.030 143.480 ;
        RECT 79.830 140.420 79.970 143.160 ;
        RECT 80.290 141.440 80.430 144.100 ;
        RECT 80.690 143.840 80.950 144.160 ;
        RECT 80.230 141.120 80.490 141.440 ;
        RECT 80.690 140.440 80.950 140.760 ;
        RECT 79.770 140.100 80.030 140.420 ;
        RECT 78.410 139.565 80.290 139.935 ;
        RECT 80.750 139.400 80.890 140.440 ;
        RECT 80.690 139.080 80.950 139.400 ;
        RECT 81.210 138.720 81.350 144.520 ;
        RECT 80.690 138.400 80.950 138.720 ;
        RECT 81.150 138.400 81.410 138.720 ;
        RECT 80.750 138.040 80.890 138.400 ;
        RECT 80.690 137.720 80.950 138.040 ;
        RECT 78.410 134.125 80.290 134.495 ;
        RECT 80.750 133.360 80.890 137.720 ;
        RECT 81.210 133.620 81.350 138.400 ;
        RECT 80.290 133.280 80.890 133.360 ;
        RECT 81.150 133.300 81.410 133.620 ;
        RECT 80.230 133.220 80.890 133.280 ;
        RECT 80.230 132.960 80.490 133.220 ;
        RECT 80.290 130.220 80.430 132.960 ;
        RECT 80.690 131.940 80.950 132.260 ;
        RECT 80.230 130.075 80.490 130.220 ;
        RECT 80.220 129.705 80.500 130.075 ;
        RECT 78.410 128.685 80.290 129.055 ;
        RECT 80.750 127.920 80.890 131.940 ;
        RECT 81.210 130.900 81.350 133.300 ;
        RECT 81.150 130.580 81.410 130.900 ;
        RECT 80.290 127.840 80.890 127.920 ;
        RECT 77.930 127.520 78.190 127.840 ;
        RECT 80.230 127.780 80.890 127.840 ;
        RECT 80.230 127.520 80.490 127.780 ;
        RECT 80.690 127.180 80.950 127.500 ;
        RECT 78.410 123.245 80.290 123.615 ;
        RECT 78.850 121.740 79.110 122.060 ;
        RECT 78.910 119.680 79.050 121.740 ;
        RECT 78.850 119.360 79.110 119.680 ;
        RECT 77.930 118.340 78.190 118.660 ;
        RECT 77.990 116.620 78.130 118.340 ;
        RECT 78.410 117.805 80.290 118.175 ;
        RECT 80.750 116.960 80.890 127.180 ;
        RECT 81.150 126.500 81.410 126.820 ;
        RECT 81.210 123.080 81.350 126.500 ;
        RECT 81.670 123.080 81.810 147.240 ;
        RECT 82.130 141.440 82.270 148.600 ;
        RECT 86.270 146.200 86.410 149.280 ;
        RECT 86.670 148.940 86.930 149.260 ;
        RECT 87.590 148.940 87.850 149.260 ;
        RECT 86.730 146.880 86.870 148.940 ;
        RECT 87.650 147.560 87.790 148.940 ;
        RECT 87.590 147.240 87.850 147.560 ;
        RECT 86.670 146.560 86.930 146.880 ;
        RECT 86.210 145.880 86.470 146.200 ;
        RECT 84.370 145.540 84.630 145.860 ;
        RECT 85.750 145.540 86.010 145.860 ;
        RECT 84.430 144.500 84.570 145.540 ;
        RECT 84.370 144.180 84.630 144.500 ;
        RECT 82.990 141.800 83.250 142.120 ;
        RECT 82.070 141.120 82.330 141.440 ;
        RECT 82.130 138.040 82.270 141.120 ;
        RECT 82.530 140.100 82.790 140.420 ;
        RECT 82.590 138.720 82.730 140.100 ;
        RECT 82.530 138.400 82.790 138.720 ;
        RECT 82.070 137.720 82.330 138.040 ;
        RECT 82.590 133.960 82.730 138.400 ;
        RECT 82.530 133.640 82.790 133.960 ;
        RECT 82.530 132.960 82.790 133.280 ;
        RECT 82.590 131.240 82.730 132.960 ;
        RECT 82.530 130.920 82.790 131.240 ;
        RECT 82.070 129.900 82.330 130.220 ;
        RECT 82.130 128.520 82.270 129.900 ;
        RECT 82.070 128.200 82.330 128.520 ;
        RECT 81.150 122.760 81.410 123.080 ;
        RECT 81.610 122.760 81.870 123.080 ;
        RECT 83.050 121.720 83.190 141.800 ;
        RECT 85.810 139.060 85.950 145.540 ;
        RECT 86.270 143.140 86.410 145.880 ;
        RECT 86.210 142.820 86.470 143.140 ;
        RECT 85.750 138.740 86.010 139.060 ;
        RECT 85.810 136.680 85.950 138.740 ;
        RECT 85.750 136.360 86.010 136.680 ;
        RECT 85.810 133.960 85.950 136.360 ;
        RECT 85.750 133.640 86.010 133.960 ;
        RECT 86.730 133.620 86.870 146.560 ;
        RECT 89.950 146.540 90.090 155.060 ;
        RECT 93.410 153.165 95.290 153.535 ;
        RECT 95.470 149.940 95.610 156.420 ;
        RECT 95.870 154.720 96.130 155.040 ;
        RECT 95.930 152.320 96.070 154.720 ;
        RECT 95.870 152.000 96.130 152.320 ;
        RECT 95.410 149.620 95.670 149.940 ;
        RECT 92.190 148.260 92.450 148.580 ;
        RECT 95.410 148.260 95.670 148.580 ;
        RECT 89.890 146.220 90.150 146.540 ;
        RECT 89.950 138.720 90.090 146.220 ;
        RECT 92.250 146.200 92.390 148.260 ;
        RECT 93.410 147.725 95.290 148.095 ;
        RECT 95.470 146.880 95.610 148.260 ;
        RECT 96.390 147.075 96.530 162.540 ;
        RECT 97.710 150.980 97.970 151.300 ;
        RECT 95.410 146.560 95.670 146.880 ;
        RECT 96.320 146.705 96.600 147.075 ;
        RECT 92.190 145.880 92.450 146.200 ;
        RECT 90.810 145.770 91.070 145.860 ;
        RECT 90.810 145.630 91.470 145.770 ;
        RECT 90.810 145.540 91.070 145.630 ;
        RECT 91.330 144.160 91.470 145.630 ;
        RECT 91.270 143.840 91.530 144.160 ;
        RECT 92.650 143.500 92.910 143.820 ;
        RECT 89.890 138.400 90.150 138.720 ;
        RECT 89.950 138.120 90.090 138.400 ;
        RECT 92.710 138.380 92.850 143.500 ;
        RECT 93.410 142.285 95.290 142.655 ;
        RECT 89.950 137.980 90.550 138.120 ;
        RECT 92.650 138.060 92.910 138.380 ;
        RECT 89.890 137.380 90.150 137.700 ;
        RECT 89.950 135.320 90.090 137.380 ;
        RECT 89.890 135.000 90.150 135.320 ;
        RECT 86.670 133.300 86.930 133.620 ;
        RECT 83.450 132.960 83.710 133.280 ;
        RECT 86.210 132.960 86.470 133.280 ;
        RECT 83.510 130.220 83.650 132.960 ;
        RECT 83.450 129.900 83.710 130.220 ;
        RECT 86.270 129.880 86.410 132.960 ;
        RECT 86.730 132.940 86.870 133.300 ;
        RECT 90.410 133.280 90.550 137.980 ;
        RECT 92.710 136.000 92.850 138.060 ;
        RECT 93.410 136.845 95.290 137.215 ;
        RECT 92.650 135.680 92.910 136.000 ;
        RECT 91.730 135.340 91.990 135.660 ;
        RECT 91.790 133.960 91.930 135.340 ;
        RECT 91.730 133.640 91.990 133.960 ;
        RECT 90.350 132.960 90.610 133.280 ;
        RECT 86.670 132.620 86.930 132.940 ;
        RECT 86.730 130.560 86.870 132.620 ;
        RECT 86.670 130.240 86.930 130.560 ;
        RECT 86.210 129.560 86.470 129.880 ;
        RECT 89.430 129.220 89.690 129.540 ;
        RECT 89.490 127.840 89.630 129.220 ;
        RECT 90.410 127.840 90.550 132.960 ;
        RECT 89.430 127.520 89.690 127.840 ;
        RECT 90.350 127.520 90.610 127.840 ;
        RECT 92.710 127.500 92.850 135.680 ;
        RECT 93.410 131.405 95.290 131.775 ;
        RECT 89.890 127.180 90.150 127.500 ;
        RECT 92.650 127.180 92.910 127.500 ;
        RECT 89.950 125.120 90.090 127.180 ;
        RECT 93.410 125.965 95.290 126.335 ;
        RECT 89.890 124.800 90.150 125.120 ;
        RECT 89.950 122.400 90.090 124.800 ;
        RECT 96.390 124.780 96.530 146.705 ;
        RECT 97.770 138.720 97.910 150.980 ;
        RECT 97.710 138.400 97.970 138.720 ;
        RECT 98.690 138.380 98.830 175.460 ;
        RECT 102.310 170.020 102.570 170.340 ;
        RECT 102.370 167.960 102.510 170.020 ;
        RECT 102.310 167.640 102.570 167.960 ;
        RECT 102.830 167.620 102.970 181.920 ;
        RECT 105.990 178.860 106.250 179.180 ;
        RECT 105.070 178.520 105.330 178.840 ;
        RECT 104.150 175.460 104.410 175.780 ;
        RECT 103.690 168.320 103.950 168.640 ;
        RECT 102.770 167.300 103.030 167.620 ;
        RECT 102.830 166.600 102.970 167.300 ;
        RECT 102.770 166.280 103.030 166.600 ;
        RECT 100.470 162.880 100.730 163.200 ;
        RECT 100.010 161.860 100.270 162.180 ;
        RECT 100.070 159.460 100.210 161.860 ;
        RECT 100.010 159.140 100.270 159.460 ;
        RECT 99.550 157.100 99.810 157.420 ;
        RECT 99.090 154.040 99.350 154.360 ;
        RECT 99.150 151.980 99.290 154.040 ;
        RECT 99.090 151.660 99.350 151.980 ;
        RECT 99.150 149.940 99.290 151.660 ;
        RECT 99.090 149.620 99.350 149.940 ;
        RECT 99.610 146.880 99.750 157.100 ;
        RECT 100.070 152.320 100.210 159.140 ;
        RECT 100.530 154.700 100.670 162.880 ;
        RECT 102.830 160.140 102.970 166.280 ;
        RECT 103.750 162.180 103.890 168.320 ;
        RECT 103.690 161.860 103.950 162.180 ;
        RECT 103.230 160.500 103.490 160.820 ;
        RECT 102.770 159.820 103.030 160.140 ;
        RECT 102.830 157.420 102.970 159.820 ;
        RECT 103.290 157.420 103.430 160.500 ;
        RECT 100.930 157.100 101.190 157.420 ;
        RECT 102.770 157.100 103.030 157.420 ;
        RECT 103.230 157.100 103.490 157.420 ;
        RECT 100.990 155.720 101.130 157.100 ;
        RECT 100.930 155.400 101.190 155.720 ;
        RECT 100.470 154.380 100.730 154.700 ;
        RECT 100.010 152.000 100.270 152.320 ;
        RECT 102.770 151.660 103.030 151.980 ;
        RECT 102.830 149.600 102.970 151.660 ;
        RECT 103.750 149.600 103.890 161.860 ;
        RECT 102.770 149.280 103.030 149.600 ;
        RECT 103.690 149.280 103.950 149.600 ;
        RECT 103.690 147.240 103.950 147.560 ;
        RECT 99.550 146.560 99.810 146.880 ;
        RECT 102.310 145.540 102.570 145.860 ;
        RECT 101.850 138.400 102.110 138.720 ;
        RECT 98.630 138.060 98.890 138.380 ;
        RECT 97.250 137.380 97.510 137.700 ;
        RECT 98.630 137.380 98.890 137.700 ;
        RECT 96.790 131.940 97.050 132.260 ;
        RECT 96.850 129.880 96.990 131.940 ;
        RECT 96.790 129.560 97.050 129.880 ;
        RECT 96.330 124.460 96.590 124.780 ;
        RECT 89.890 122.080 90.150 122.400 ;
        RECT 83.450 121.740 83.710 122.060 ;
        RECT 84.370 121.740 84.630 122.060 ;
        RECT 82.990 121.400 83.250 121.720 ;
        RECT 81.610 119.360 81.870 119.680 ;
        RECT 82.530 119.360 82.790 119.680 ;
        RECT 81.150 119.020 81.410 119.340 ;
        RECT 81.210 117.640 81.350 119.020 ;
        RECT 81.670 117.640 81.810 119.360 ;
        RECT 81.150 117.320 81.410 117.640 ;
        RECT 81.610 117.320 81.870 117.640 ;
        RECT 80.690 116.640 80.950 116.960 ;
        RECT 77.930 116.300 78.190 116.620 ;
        RECT 80.750 114.580 80.890 116.640 ;
        RECT 82.590 116.620 82.730 119.360 ;
        RECT 83.510 119.340 83.650 121.740 ;
        RECT 83.450 119.020 83.710 119.340 ;
        RECT 83.510 117.640 83.650 119.020 ;
        RECT 84.430 118.660 84.570 121.740 ;
        RECT 93.410 120.525 95.290 120.895 ;
        RECT 95.410 119.360 95.670 119.680 ;
        RECT 92.650 118.680 92.910 119.000 ;
        RECT 84.370 118.340 84.630 118.660 ;
        RECT 85.290 118.340 85.550 118.660 ;
        RECT 83.450 117.320 83.710 117.640 ;
        RECT 82.530 116.300 82.790 116.620 ;
        RECT 80.690 114.260 80.950 114.580 ;
        RECT 80.750 113.900 80.890 114.260 ;
        RECT 80.690 113.580 80.950 113.900 ;
        RECT 83.450 113.580 83.710 113.900 ;
        RECT 83.910 113.580 84.170 113.900 ;
        RECT 77.930 112.900 78.190 113.220 ;
        RECT 77.990 111.520 78.130 112.900 ;
        RECT 78.410 112.365 80.290 112.735 ;
        RECT 77.930 111.200 78.190 111.520 ;
        RECT 83.510 111.180 83.650 113.580 ;
        RECT 83.970 112.200 84.110 113.580 ;
        RECT 84.430 113.220 84.570 118.340 ;
        RECT 84.370 112.900 84.630 113.220 ;
        RECT 83.910 111.880 84.170 112.200 ;
        RECT 85.350 111.520 85.490 118.340 ;
        RECT 89.890 115.620 90.150 115.940 ;
        RECT 89.950 114.240 90.090 115.620 ;
        RECT 92.710 114.920 92.850 118.680 ;
        RECT 93.410 115.085 95.290 115.455 ;
        RECT 95.470 114.920 95.610 119.360 ;
        RECT 96.330 116.980 96.590 117.300 ;
        RECT 92.650 114.600 92.910 114.920 ;
        RECT 95.410 114.600 95.670 114.920 ;
        RECT 96.390 114.580 96.530 116.980 ;
        RECT 96.330 114.260 96.590 114.580 ;
        RECT 86.210 113.920 86.470 114.240 ;
        RECT 89.890 113.920 90.150 114.240 ;
        RECT 86.270 111.520 86.410 113.920 ;
        RECT 86.670 113.240 86.930 113.560 ;
        RECT 86.730 112.200 86.870 113.240 ;
        RECT 86.670 111.880 86.930 112.200 ;
        RECT 85.290 111.200 85.550 111.520 ;
        RECT 86.210 111.200 86.470 111.520 ;
        RECT 83.450 110.860 83.710 111.180 ;
        RECT 81.610 107.800 81.870 108.120 ;
        RECT 78.410 106.925 80.290 107.295 ;
        RECT 79.310 103.380 79.570 103.700 ;
        RECT 79.370 103.020 79.510 103.380 ;
        RECT 81.670 103.360 81.810 107.800 ;
        RECT 83.510 105.740 83.650 110.860 ;
        RECT 93.410 109.645 95.290 110.015 ;
        RECT 97.310 108.460 97.450 137.380 ;
        RECT 98.690 128.520 98.830 137.380 ;
        RECT 101.910 133.280 102.050 138.400 ;
        RECT 101.850 132.960 102.110 133.280 ;
        RECT 99.090 132.620 99.350 132.940 ;
        RECT 99.150 131.240 99.290 132.620 ;
        RECT 101.390 131.940 101.650 132.260 ;
        RECT 99.090 130.920 99.350 131.240 ;
        RECT 100.930 129.900 101.190 130.220 ;
        RECT 100.990 128.520 101.130 129.900 ;
        RECT 98.630 128.200 98.890 128.520 ;
        RECT 100.930 128.200 101.190 128.520 ;
        RECT 101.450 127.840 101.590 131.940 ;
        RECT 97.710 127.520 97.970 127.840 ;
        RECT 98.170 127.520 98.430 127.840 ;
        RECT 101.390 127.520 101.650 127.840 ;
        RECT 97.770 119.340 97.910 127.520 ;
        RECT 98.230 125.460 98.370 127.520 ;
        RECT 98.170 125.140 98.430 125.460 ;
        RECT 98.630 119.360 98.890 119.680 ;
        RECT 97.710 119.020 97.970 119.340 ;
        RECT 97.770 117.640 97.910 119.020 ;
        RECT 97.710 117.320 97.970 117.640 ;
        RECT 98.690 116.960 98.830 119.360 ;
        RECT 101.850 118.340 102.110 118.660 ;
        RECT 101.910 116.960 102.050 118.340 ;
        RECT 98.630 116.640 98.890 116.960 ;
        RECT 101.850 116.640 102.110 116.960 ;
        RECT 98.690 116.460 98.830 116.640 ;
        RECT 98.690 116.320 99.290 116.460 ;
        RECT 99.150 115.940 99.290 116.320 ;
        RECT 99.090 115.620 99.350 115.940 ;
        RECT 102.370 108.460 102.510 145.540 ;
        RECT 102.770 140.780 103.030 141.100 ;
        RECT 102.830 139.400 102.970 140.780 ;
        RECT 102.770 139.080 103.030 139.400 ;
        RECT 102.830 138.720 102.970 139.080 ;
        RECT 102.770 138.400 103.030 138.720 ;
        RECT 102.770 129.900 103.030 130.220 ;
        RECT 102.830 125.120 102.970 129.900 ;
        RECT 103.750 125.460 103.890 147.240 ;
        RECT 104.210 138.380 104.350 175.460 ;
        RECT 104.610 167.980 104.870 168.300 ;
        RECT 104.670 164.900 104.810 167.980 ;
        RECT 104.610 164.580 104.870 164.900 ;
        RECT 104.670 163.540 104.810 164.580 ;
        RECT 104.610 163.220 104.870 163.540 ;
        RECT 104.670 152.320 104.810 163.220 ;
        RECT 105.130 154.440 105.270 178.520 ;
        RECT 106.050 177.480 106.190 178.860 ;
        RECT 105.990 177.160 106.250 177.480 ;
        RECT 106.050 176.800 106.190 177.160 ;
        RECT 106.970 176.800 107.110 187.360 ;
        RECT 107.370 187.020 107.630 187.340 ;
        RECT 107.430 184.960 107.570 187.020 ;
        RECT 107.370 184.640 107.630 184.960 ;
        RECT 107.890 179.180 108.030 189.060 ;
        RECT 108.410 188.525 110.290 188.895 ;
        RECT 110.650 187.340 110.790 190.080 ;
        RECT 111.570 189.720 111.710 194.500 ;
        RECT 115.190 191.780 115.450 192.100 ;
        RECT 115.250 191.080 115.390 191.780 ;
        RECT 115.190 190.760 115.450 191.080 ;
        RECT 115.650 189.740 115.910 190.060 ;
        RECT 111.510 189.400 111.770 189.720 ;
        RECT 113.810 189.400 114.070 189.720 ;
        RECT 111.050 188.040 111.310 188.360 ;
        RECT 110.590 187.020 110.850 187.340 ;
        RECT 108.410 183.085 110.290 183.455 ;
        RECT 110.650 181.900 110.790 187.020 ;
        RECT 111.110 182.240 111.250 188.040 ;
        RECT 112.890 182.260 113.150 182.580 ;
        RECT 111.050 181.920 111.310 182.240 ;
        RECT 110.590 181.580 110.850 181.900 ;
        RECT 107.370 178.860 107.630 179.180 ;
        RECT 107.830 178.860 108.090 179.180 ;
        RECT 105.990 176.480 106.250 176.800 ;
        RECT 106.910 176.480 107.170 176.800 ;
        RECT 106.050 173.740 106.190 176.480 ;
        RECT 107.430 176.460 107.570 178.860 ;
        RECT 107.830 178.180 108.090 178.500 ;
        RECT 107.890 176.800 108.030 178.180 ;
        RECT 108.410 177.645 110.290 178.015 ;
        RECT 111.110 176.800 111.250 181.920 ;
        RECT 112.430 181.580 112.690 181.900 ;
        RECT 112.490 179.520 112.630 181.580 ;
        RECT 112.430 179.200 112.690 179.520 ;
        RECT 111.510 178.520 111.770 178.840 ;
        RECT 111.570 176.800 111.710 178.520 ;
        RECT 112.950 178.500 113.090 182.260 ;
        RECT 113.870 178.500 114.010 189.400 ;
        RECT 115.710 188.360 115.850 189.740 ;
        RECT 115.650 188.040 115.910 188.360 ;
        RECT 116.170 184.620 116.310 198.240 ;
        RECT 123.410 196.685 125.290 197.055 ;
        RECT 120.250 195.180 120.510 195.500 ;
        RECT 117.490 194.840 117.750 195.160 ;
        RECT 117.550 193.800 117.690 194.840 ;
        RECT 117.490 193.480 117.750 193.800 ;
        RECT 116.570 192.800 116.830 193.120 ;
        RECT 116.630 190.740 116.770 192.800 ;
        RECT 120.310 192.780 120.450 195.180 ;
        RECT 120.250 192.520 120.510 192.780 ;
        RECT 120.250 192.460 121.370 192.520 ;
        RECT 120.310 192.380 121.370 192.460 ;
        RECT 116.570 190.420 116.830 190.740 ;
        RECT 116.110 184.300 116.370 184.620 ;
        RECT 115.650 183.960 115.910 184.280 ;
        RECT 115.710 182.920 115.850 183.960 ;
        RECT 117.030 183.620 117.290 183.940 ;
        RECT 118.410 183.620 118.670 183.940 ;
        RECT 115.650 182.600 115.910 182.920 ;
        RECT 117.090 182.580 117.230 183.620 ;
        RECT 117.030 182.260 117.290 182.580 ;
        RECT 118.470 178.840 118.610 183.620 ;
        RECT 121.230 181.900 121.370 192.380 ;
        RECT 123.410 191.245 125.290 191.615 ;
        RECT 123.410 185.805 125.290 186.175 ;
        RECT 123.930 183.620 124.190 183.940 ;
        RECT 123.990 182.580 124.130 183.620 ;
        RECT 123.930 182.260 124.190 182.580 ;
        RECT 121.170 181.580 121.430 181.900 ;
        RECT 125.770 181.580 126.030 181.900 ;
        RECT 123.410 180.365 125.290 180.735 ;
        RECT 125.830 179.520 125.970 181.580 ;
        RECT 125.770 179.200 126.030 179.520 ;
        RECT 118.410 178.520 118.670 178.840 ;
        RECT 123.470 178.520 123.730 178.840 ;
        RECT 112.890 178.180 113.150 178.500 ;
        RECT 113.810 178.180 114.070 178.500 ;
        RECT 115.650 178.180 115.910 178.500 ;
        RECT 112.950 176.800 113.090 178.180 ;
        RECT 107.830 176.480 108.090 176.800 ;
        RECT 110.130 176.480 110.390 176.800 ;
        RECT 111.050 176.480 111.310 176.800 ;
        RECT 111.510 176.480 111.770 176.800 ;
        RECT 112.890 176.480 113.150 176.800 ;
        RECT 107.370 176.140 107.630 176.460 ;
        RECT 107.830 175.460 108.090 175.780 ;
        RECT 105.990 173.420 106.250 173.740 ;
        RECT 106.450 172.740 106.710 173.060 ;
        RECT 105.990 168.660 106.250 168.980 ;
        RECT 106.050 162.860 106.190 168.660 ;
        RECT 105.990 162.540 106.250 162.860 ;
        RECT 105.530 161.860 105.790 162.180 ;
        RECT 105.590 160.480 105.730 161.860 ;
        RECT 105.530 160.160 105.790 160.480 ;
        RECT 106.510 155.800 106.650 172.740 ;
        RECT 106.970 168.640 107.570 168.720 ;
        RECT 106.970 168.580 107.630 168.640 ;
        RECT 106.970 163.880 107.110 168.580 ;
        RECT 107.370 168.320 107.630 168.580 ;
        RECT 106.910 163.560 107.170 163.880 ;
        RECT 106.050 155.660 106.650 155.800 ;
        RECT 105.130 154.300 105.730 154.440 ;
        RECT 104.610 152.000 104.870 152.320 ;
        RECT 104.610 151.320 104.870 151.640 ;
        RECT 104.670 149.600 104.810 151.320 ;
        RECT 104.610 149.280 104.870 149.600 ;
        RECT 104.610 148.260 104.870 148.580 ;
        RECT 104.670 138.720 104.810 148.260 ;
        RECT 105.070 145.540 105.330 145.860 ;
        RECT 105.130 144.500 105.270 145.540 ;
        RECT 105.070 144.180 105.330 144.500 ;
        RECT 105.590 143.820 105.730 154.300 ;
        RECT 106.050 146.880 106.190 155.660 ;
        RECT 107.370 154.380 107.630 154.700 ;
        RECT 106.910 153.700 107.170 154.020 ;
        RECT 106.450 148.260 106.710 148.580 ;
        RECT 105.990 146.560 106.250 146.880 ;
        RECT 106.510 144.160 106.650 148.260 ;
        RECT 106.970 146.540 107.110 153.700 ;
        RECT 107.430 151.980 107.570 154.380 ;
        RECT 107.370 151.660 107.630 151.980 ;
        RECT 107.430 149.940 107.570 151.660 ;
        RECT 107.370 149.620 107.630 149.940 ;
        RECT 107.370 147.240 107.630 147.560 ;
        RECT 107.430 146.540 107.570 147.240 ;
        RECT 106.910 146.220 107.170 146.540 ;
        RECT 107.370 146.220 107.630 146.540 ;
        RECT 107.370 145.540 107.630 145.860 ;
        RECT 107.430 144.840 107.570 145.540 ;
        RECT 107.370 144.520 107.630 144.840 ;
        RECT 106.450 143.840 106.710 144.160 ;
        RECT 105.530 143.500 105.790 143.820 ;
        RECT 106.450 142.820 106.710 143.140 ;
        RECT 104.610 138.400 104.870 138.720 ;
        RECT 104.150 138.060 104.410 138.380 ;
        RECT 104.150 137.380 104.410 137.700 ;
        RECT 105.990 137.380 106.250 137.700 ;
        RECT 103.690 125.140 103.950 125.460 ;
        RECT 102.770 124.800 103.030 125.120 ;
        RECT 102.830 120.020 102.970 124.800 ;
        RECT 102.770 119.700 103.030 120.020 ;
        RECT 102.830 116.620 102.970 119.700 ;
        RECT 102.770 116.300 103.030 116.620 ;
        RECT 102.830 111.520 102.970 116.300 ;
        RECT 102.770 111.200 103.030 111.520 ;
        RECT 97.250 108.140 97.510 108.460 ;
        RECT 102.310 108.140 102.570 108.460 ;
        RECT 99.550 107.460 99.810 107.780 ;
        RECT 99.610 106.420 99.750 107.460 ;
        RECT 98.170 106.100 98.430 106.420 ;
        RECT 99.550 106.100 99.810 106.420 ;
        RECT 82.070 105.420 82.330 105.740 ;
        RECT 83.450 105.420 83.710 105.740 ;
        RECT 82.130 104.040 82.270 105.420 ;
        RECT 82.070 103.720 82.330 104.040 ;
        RECT 81.610 103.040 81.870 103.360 ;
        RECT 77.470 102.700 77.730 103.020 ;
        RECT 79.310 102.700 79.570 103.020 ;
        RECT 77.930 102.020 78.190 102.340 ;
        RECT 77.990 101.320 78.130 102.020 ;
        RECT 78.410 101.485 80.290 101.855 ;
        RECT 77.930 101.000 78.190 101.320 ;
        RECT 83.510 100.300 83.650 105.420 ;
        RECT 92.650 104.740 92.910 105.060 ;
        RECT 97.250 104.740 97.510 105.060 ;
        RECT 85.750 103.380 86.010 103.700 ;
        RECT 85.810 103.020 85.950 103.380 ;
        RECT 92.710 103.360 92.850 104.740 ;
        RECT 93.410 104.205 95.290 104.575 ;
        RECT 90.810 103.040 91.070 103.360 ;
        RECT 92.650 103.040 92.910 103.360 ;
        RECT 84.830 102.700 85.090 103.020 ;
        RECT 85.750 102.700 86.010 103.020 ;
        RECT 90.870 102.760 91.010 103.040 ;
        RECT 84.890 100.980 85.030 102.700 ;
        RECT 90.870 102.620 91.930 102.760 ;
        RECT 88.510 102.020 88.770 102.340 ;
        RECT 88.570 100.980 88.710 102.020 ;
        RECT 84.830 100.660 85.090 100.980 ;
        RECT 88.510 100.660 88.770 100.980 ;
        RECT 83.450 99.980 83.710 100.300 ;
        RECT 85.290 99.300 85.550 99.620 ;
        RECT 78.410 96.045 80.290 96.415 ;
        RECT 77.070 95.140 79.050 95.280 ;
        RECT 72.400 86.440 72.680 86.920 ;
        RECT 71.550 86.300 72.680 86.440 ;
        RECT 72.400 84.920 72.680 86.300 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 78.910 86.920 79.050 95.140 ;
        RECT 78.840 84.920 79.120 86.920 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 85.350 87.970 85.490 99.300 ;
        RECT 91.790 88.320 91.930 102.620 ;
        RECT 93.410 98.765 95.290 99.135 ;
        RECT 85.350 86.920 86.690 87.970 ;
        RECT 85.280 84.920 86.690 86.920 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 84.920 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.310 86.440 97.450 104.740 ;
        RECT 98.230 104.040 98.370 106.100 ;
        RECT 102.830 106.080 102.970 111.200 ;
        RECT 104.210 106.080 104.350 137.380 ;
        RECT 105.530 132.960 105.790 133.280 ;
        RECT 105.590 130.220 105.730 132.960 ;
        RECT 105.530 129.900 105.790 130.220 ;
        RECT 106.050 128.520 106.190 137.380 ;
        RECT 105.990 128.200 106.250 128.520 ;
        RECT 105.990 127.180 106.250 127.500 ;
        RECT 104.610 126.840 104.870 127.160 ;
        RECT 104.670 124.100 104.810 126.840 ;
        RECT 106.050 125.200 106.190 127.180 ;
        RECT 106.510 125.800 106.650 142.820 ;
        RECT 107.370 140.780 107.630 141.100 ;
        RECT 107.430 138.720 107.570 140.780 ;
        RECT 107.890 139.310 108.030 175.460 ;
        RECT 110.190 173.740 110.330 176.480 ;
        RECT 111.570 173.740 111.710 176.480 ;
        RECT 112.890 175.460 113.150 175.780 ;
        RECT 110.130 173.420 110.390 173.740 ;
        RECT 111.510 173.420 111.770 173.740 ;
        RECT 108.410 172.205 110.290 172.575 ;
        RECT 111.050 170.360 111.310 170.680 ;
        RECT 110.590 170.020 110.850 170.340 ;
        RECT 108.410 166.765 110.290 167.135 ;
        RECT 110.650 166.260 110.790 170.020 ;
        RECT 110.590 165.940 110.850 166.260 ;
        RECT 110.590 161.860 110.850 162.180 ;
        RECT 108.410 161.325 110.290 161.695 ;
        RECT 108.410 155.885 110.290 156.255 ;
        RECT 108.290 154.720 108.550 155.040 ;
        RECT 108.350 151.980 108.490 154.720 ;
        RECT 110.130 154.040 110.390 154.360 ;
        RECT 110.190 151.980 110.330 154.040 ;
        RECT 110.650 151.980 110.790 161.860 ;
        RECT 108.290 151.660 108.550 151.980 ;
        RECT 110.130 151.660 110.390 151.980 ;
        RECT 110.590 151.660 110.850 151.980 ;
        RECT 108.350 151.300 108.490 151.660 ;
        RECT 108.290 150.980 108.550 151.300 ;
        RECT 110.190 151.210 110.330 151.660 ;
        RECT 110.190 151.070 110.790 151.210 ;
        RECT 108.410 150.445 110.290 150.815 ;
        RECT 110.130 149.280 110.390 149.600 ;
        RECT 109.210 146.960 109.470 147.220 ;
        RECT 108.350 146.900 109.470 146.960 ;
        RECT 108.350 146.820 109.410 146.900 ;
        RECT 110.190 146.880 110.330 149.280 ;
        RECT 110.650 149.260 110.790 151.070 ;
        RECT 111.110 149.940 111.250 170.360 ;
        RECT 111.510 150.980 111.770 151.300 ;
        RECT 111.050 149.620 111.310 149.940 ;
        RECT 110.590 148.940 110.850 149.260 ;
        RECT 111.050 147.240 111.310 147.560 ;
        RECT 108.350 146.540 108.490 146.820 ;
        RECT 110.130 146.560 110.390 146.880 ;
        RECT 111.110 146.540 111.250 147.240 ;
        RECT 108.290 146.220 108.550 146.540 ;
        RECT 110.590 146.220 110.850 146.540 ;
        RECT 111.050 146.220 111.310 146.540 ;
        RECT 108.410 145.005 110.290 145.375 ;
        RECT 109.670 143.500 109.930 143.820 ;
        RECT 109.730 140.760 109.870 143.500 ;
        RECT 110.650 143.480 110.790 146.220 ;
        RECT 111.110 144.160 111.250 146.220 ;
        RECT 111.050 143.840 111.310 144.160 ;
        RECT 110.590 143.160 110.850 143.480 ;
        RECT 111.110 141.780 111.250 143.840 ;
        RECT 111.050 141.460 111.310 141.780 ;
        RECT 111.050 140.780 111.310 141.100 ;
        RECT 109.670 140.440 109.930 140.760 ;
        RECT 110.590 140.100 110.850 140.420 ;
        RECT 108.410 139.565 110.290 139.935 ;
        RECT 107.890 139.170 108.490 139.310 ;
        RECT 107.370 138.400 107.630 138.720 ;
        RECT 107.830 136.360 108.090 136.680 ;
        RECT 106.910 134.660 107.170 134.980 ;
        RECT 106.450 125.480 106.710 125.800 ;
        RECT 106.050 125.060 106.650 125.200 ;
        RECT 104.610 123.780 104.870 124.100 ;
        RECT 104.670 122.400 104.810 123.780 ;
        RECT 106.510 122.400 106.650 125.060 ;
        RECT 104.610 122.080 104.870 122.400 ;
        RECT 106.450 122.080 106.710 122.400 ;
        RECT 105.070 121.060 105.330 121.380 ;
        RECT 105.130 119.000 105.270 121.060 ;
        RECT 106.510 119.680 106.650 122.080 ;
        RECT 106.450 119.360 106.710 119.680 ;
        RECT 105.070 118.680 105.330 119.000 ;
        RECT 105.530 115.620 105.790 115.940 ;
        RECT 105.590 111.520 105.730 115.620 ;
        RECT 105.530 111.200 105.790 111.520 ;
        RECT 106.970 106.420 107.110 134.660 ;
        RECT 107.370 129.560 107.630 129.880 ;
        RECT 107.430 128.520 107.570 129.560 ;
        RECT 107.370 128.200 107.630 128.520 ;
        RECT 107.890 127.840 108.030 136.360 ;
        RECT 108.350 136.000 108.490 139.170 ;
        RECT 108.290 135.680 108.550 136.000 ;
        RECT 110.650 135.660 110.790 140.100 ;
        RECT 111.110 139.060 111.250 140.780 ;
        RECT 111.050 138.740 111.310 139.060 ;
        RECT 111.050 138.060 111.310 138.380 ;
        RECT 110.590 135.340 110.850 135.660 ;
        RECT 108.410 134.125 110.290 134.495 ;
        RECT 111.110 132.940 111.250 138.060 ;
        RECT 111.570 136.000 111.710 150.980 ;
        RECT 111.970 146.450 112.230 146.540 ;
        RECT 111.970 146.310 112.630 146.450 ;
        RECT 111.970 146.220 112.230 146.310 ;
        RECT 111.970 143.160 112.230 143.480 ;
        RECT 112.030 141.100 112.170 143.160 ;
        RECT 111.970 140.780 112.230 141.100 ;
        RECT 112.030 139.400 112.170 140.780 ;
        RECT 112.490 140.760 112.630 146.310 ;
        RECT 112.950 143.820 113.090 175.460 ;
        RECT 113.870 174.080 114.010 178.180 ;
        RECT 115.710 176.800 115.850 178.180 ;
        RECT 123.530 177.480 123.670 178.520 ;
        RECT 123.470 177.160 123.730 177.480 ;
        RECT 115.650 176.480 115.910 176.800 ;
        RECT 123.410 174.925 125.290 175.295 ;
        RECT 113.810 173.760 114.070 174.080 ;
        RECT 113.810 170.360 114.070 170.680 ;
        RECT 120.710 170.360 120.970 170.680 ;
        RECT 113.870 167.620 114.010 170.360 ;
        RECT 117.490 170.020 117.750 170.340 ;
        RECT 118.410 170.020 118.670 170.340 ;
        RECT 117.030 168.320 117.290 168.640 ;
        RECT 114.270 167.640 114.530 167.960 ;
        RECT 113.810 167.300 114.070 167.620 ;
        RECT 113.810 165.260 114.070 165.580 ;
        RECT 113.870 163.880 114.010 165.260 ;
        RECT 113.810 163.560 114.070 163.880 ;
        RECT 114.330 163.540 114.470 167.640 ;
        RECT 116.570 164.580 116.830 164.900 ;
        RECT 114.270 163.220 114.530 163.540 ;
        RECT 116.630 162.860 116.770 164.580 ;
        RECT 116.570 162.540 116.830 162.860 ;
        RECT 117.090 162.180 117.230 168.320 ;
        RECT 117.550 167.960 117.690 170.020 ;
        RECT 117.490 167.640 117.750 167.960 ;
        RECT 118.470 165.920 118.610 170.020 ;
        RECT 118.410 165.600 118.670 165.920 ;
        RECT 114.270 161.860 114.530 162.180 ;
        RECT 117.030 161.860 117.290 162.180 ;
        RECT 114.330 155.380 114.470 161.860 ;
        RECT 120.770 160.480 120.910 170.360 ;
        RECT 123.410 169.485 125.290 169.855 ;
        RECT 125.830 168.640 125.970 179.200 ;
        RECT 127.600 174.585 127.880 174.955 ;
        RECT 127.670 171.700 127.810 174.585 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 127.610 171.380 127.870 171.700 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 125.770 168.320 126.030 168.640 ;
        RECT 124.390 167.640 124.650 167.960 ;
        RECT 124.450 166.600 124.590 167.640 ;
        RECT 124.390 166.280 124.650 166.600 ;
        RECT 122.550 165.940 122.810 166.260 ;
        RECT 122.610 163.880 122.750 165.940 ;
        RECT 125.830 165.920 125.970 168.320 ;
        RECT 126.690 167.300 126.950 167.620 ;
        RECT 126.750 165.920 126.890 167.300 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 125.770 165.600 126.030 165.920 ;
        RECT 126.690 165.600 126.950 165.920 ;
        RECT 123.410 164.045 125.290 164.415 ;
        RECT 122.550 163.560 122.810 163.880 ;
        RECT 117.950 160.160 118.210 160.480 ;
        RECT 120.710 160.160 120.970 160.480 ;
        RECT 116.570 157.100 116.830 157.420 ;
        RECT 114.270 155.060 114.530 155.380 ;
        RECT 116.110 151.660 116.370 151.980 ;
        RECT 113.350 150.980 113.610 151.300 ;
        RECT 113.410 144.500 113.550 150.980 ;
        RECT 116.170 150.280 116.310 151.660 ;
        RECT 116.110 149.960 116.370 150.280 ;
        RECT 114.270 149.680 114.530 149.940 ;
        RECT 113.870 149.620 114.530 149.680 ;
        RECT 113.870 149.540 114.470 149.620 ;
        RECT 113.870 148.920 114.010 149.540 ;
        RECT 114.270 148.940 114.530 149.260 ;
        RECT 113.810 148.600 114.070 148.920 ;
        RECT 113.870 145.600 114.010 148.600 ;
        RECT 114.330 146.880 114.470 148.940 ;
        RECT 114.270 146.560 114.530 146.880 ;
        RECT 113.870 145.460 114.470 145.600 ;
        RECT 113.810 144.520 114.070 144.840 ;
        RECT 113.350 144.180 113.610 144.500 ;
        RECT 112.890 143.500 113.150 143.820 ;
        RECT 113.870 143.560 114.010 144.520 ;
        RECT 113.410 143.420 114.010 143.560 ;
        RECT 113.410 143.050 113.550 143.420 ;
        RECT 112.950 142.910 113.550 143.050 ;
        RECT 112.430 140.440 112.690 140.760 ;
        RECT 111.970 139.080 112.230 139.400 ;
        RECT 112.490 137.700 112.630 140.440 ;
        RECT 112.430 137.380 112.690 137.700 ;
        RECT 111.510 135.680 111.770 136.000 ;
        RECT 111.050 132.620 111.310 132.940 ;
        RECT 108.410 128.685 110.290 129.055 ;
        RECT 107.830 127.520 108.090 127.840 ;
        RECT 112.430 127.520 112.690 127.840 ;
        RECT 110.590 127.180 110.850 127.500 ;
        RECT 107.370 124.120 107.630 124.440 ;
        RECT 107.430 113.900 107.570 124.120 ;
        RECT 108.410 123.245 110.290 123.615 ;
        RECT 110.650 123.080 110.790 127.180 ;
        RECT 112.490 124.780 112.630 127.520 ;
        RECT 112.430 124.460 112.690 124.780 ;
        RECT 110.590 122.760 110.850 123.080 ;
        RECT 107.830 121.740 108.090 122.060 ;
        RECT 107.890 116.280 108.030 121.740 ;
        RECT 110.590 121.060 110.850 121.380 ;
        RECT 108.410 117.805 110.290 118.175 ;
        RECT 110.650 116.960 110.790 121.060 ;
        RECT 111.050 119.020 111.310 119.340 ;
        RECT 111.110 117.640 111.250 119.020 ;
        RECT 111.050 117.320 111.310 117.640 ;
        RECT 108.290 116.640 108.550 116.960 ;
        RECT 110.590 116.640 110.850 116.960 ;
        RECT 107.830 115.960 108.090 116.280 ;
        RECT 107.890 114.240 108.030 115.960 ;
        RECT 108.350 114.920 108.490 116.640 ;
        RECT 108.290 114.600 108.550 114.920 ;
        RECT 107.830 113.920 108.090 114.240 ;
        RECT 107.370 113.580 107.630 113.900 ;
        RECT 107.370 112.900 107.630 113.220 ;
        RECT 111.970 112.900 112.230 113.220 ;
        RECT 107.430 111.860 107.570 112.900 ;
        RECT 108.410 112.365 110.290 112.735 ;
        RECT 112.030 112.200 112.170 112.900 ;
        RECT 111.970 111.880 112.230 112.200 ;
        RECT 107.370 111.540 107.630 111.860 ;
        RECT 108.410 106.925 110.290 107.295 ;
        RECT 106.910 106.100 107.170 106.420 ;
        RECT 112.950 106.080 113.090 142.910 ;
        RECT 113.810 142.820 114.070 143.140 ;
        RECT 113.350 138.060 113.610 138.380 ;
        RECT 113.410 136.680 113.550 138.060 ;
        RECT 113.350 136.360 113.610 136.680 ;
        RECT 113.410 133.960 113.550 136.360 ;
        RECT 113.350 133.640 113.610 133.960 ;
        RECT 113.350 131.940 113.610 132.260 ;
        RECT 113.410 130.560 113.550 131.940 ;
        RECT 113.350 130.240 113.610 130.560 ;
        RECT 113.870 128.520 114.010 142.820 ;
        RECT 114.330 141.440 114.470 145.460 ;
        RECT 114.270 141.120 114.530 141.440 ;
        RECT 114.330 138.720 114.470 141.120 ;
        RECT 116.630 141.100 116.770 157.100 ;
        RECT 118.010 155.040 118.150 160.160 ;
        RECT 119.330 159.820 119.590 160.140 ;
        RECT 119.390 157.420 119.530 159.820 ;
        RECT 123.410 158.605 125.290 158.975 ;
        RECT 119.330 157.100 119.590 157.420 ;
        RECT 119.790 156.420 120.050 156.740 ;
        RECT 120.710 156.420 120.970 156.740 ;
        RECT 117.950 154.720 118.210 155.040 ;
        RECT 117.030 153.700 117.290 154.020 ;
        RECT 117.090 149.260 117.230 153.700 ;
        RECT 119.850 151.640 119.990 156.420 ;
        RECT 120.770 155.380 120.910 156.420 ;
        RECT 120.710 155.060 120.970 155.380 ;
        RECT 125.830 155.040 125.970 165.600 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 125.770 154.720 126.030 155.040 ;
        RECT 122.550 154.380 122.810 154.700 ;
        RECT 119.790 151.320 120.050 151.640 ;
        RECT 118.870 150.980 119.130 151.300 ;
        RECT 117.030 148.940 117.290 149.260 ;
        RECT 118.930 149.170 119.070 150.980 ;
        RECT 122.610 150.280 122.750 154.380 ;
        RECT 123.410 153.165 125.290 153.535 ;
        RECT 125.830 152.320 125.970 154.720 ;
        RECT 125.770 152.000 126.030 152.320 ;
        RECT 122.550 149.960 122.810 150.280 ;
        RECT 119.790 149.170 120.050 149.260 ;
        RECT 118.930 149.030 120.050 149.170 ;
        RECT 119.790 148.940 120.050 149.030 ;
        RECT 119.850 143.820 119.990 148.940 ;
        RECT 123.410 147.725 125.290 148.095 ;
        RECT 123.010 145.540 123.270 145.860 ;
        RECT 119.790 143.500 120.050 143.820 ;
        RECT 119.850 141.100 119.990 143.500 ;
        RECT 116.570 140.780 116.830 141.100 ;
        RECT 119.790 140.780 120.050 141.100 ;
        RECT 116.630 138.720 116.770 140.780 ;
        RECT 117.030 140.100 117.290 140.420 ;
        RECT 119.330 140.100 119.590 140.420 ;
        RECT 117.090 139.060 117.230 140.100 ;
        RECT 119.390 139.400 119.530 140.100 ;
        RECT 119.330 139.080 119.590 139.400 ;
        RECT 117.030 138.740 117.290 139.060 ;
        RECT 114.270 138.400 114.530 138.720 ;
        RECT 116.570 138.400 116.830 138.720 ;
        RECT 115.650 137.380 115.910 137.700 ;
        RECT 117.030 137.380 117.290 137.700 ;
        RECT 115.710 133.280 115.850 137.380 ;
        RECT 117.090 135.320 117.230 137.380 ;
        RECT 117.030 135.000 117.290 135.320 ;
        RECT 115.650 132.960 115.910 133.280 ;
        RECT 113.810 128.200 114.070 128.520 ;
        RECT 114.270 127.180 114.530 127.500 ;
        RECT 113.350 123.780 113.610 124.100 ;
        RECT 113.410 116.960 113.550 123.780 ;
        RECT 114.330 122.740 114.470 127.180 ;
        RECT 117.030 124.800 117.290 125.120 ;
        RECT 114.270 122.420 114.530 122.740 ;
        RECT 113.810 121.740 114.070 122.060 ;
        RECT 113.870 119.680 114.010 121.740 ;
        RECT 117.090 119.680 117.230 124.800 ;
        RECT 117.490 124.120 117.750 124.440 ;
        RECT 120.710 124.120 120.970 124.440 ;
        RECT 117.550 122.740 117.690 124.120 ;
        RECT 118.870 123.780 119.130 124.100 ;
        RECT 118.930 122.740 119.070 123.780 ;
        RECT 117.490 122.420 117.750 122.740 ;
        RECT 118.870 122.420 119.130 122.740 ;
        RECT 113.810 119.360 114.070 119.680 ;
        RECT 117.030 119.360 117.290 119.680 ;
        RECT 113.350 116.640 113.610 116.960 ;
        RECT 113.410 114.240 113.550 116.640 ;
        RECT 117.090 114.920 117.230 119.360 ;
        RECT 117.550 119.340 117.690 122.420 ;
        RECT 117.950 121.060 118.210 121.380 ;
        RECT 119.330 121.060 119.590 121.380 ;
        RECT 118.010 119.680 118.150 121.060 ;
        RECT 119.390 120.360 119.530 121.060 ;
        RECT 120.770 120.360 120.910 124.120 ;
        RECT 122.550 121.740 122.810 122.060 ;
        RECT 122.610 120.360 122.750 121.740 ;
        RECT 119.330 120.040 119.590 120.360 ;
        RECT 120.710 120.040 120.970 120.360 ;
        RECT 122.550 120.040 122.810 120.360 ;
        RECT 117.950 119.360 118.210 119.680 ;
        RECT 117.490 119.020 117.750 119.340 ;
        RECT 120.250 119.020 120.510 119.340 ;
        RECT 120.310 116.960 120.450 119.020 ;
        RECT 120.250 116.640 120.510 116.960 ;
        RECT 118.410 116.300 118.670 116.620 ;
        RECT 117.030 114.600 117.290 114.920 ;
        RECT 113.350 113.920 113.610 114.240 ;
        RECT 118.470 113.560 118.610 116.300 ;
        RECT 122.090 113.920 122.350 114.240 ;
        RECT 121.630 113.580 121.890 113.900 ;
        RECT 118.410 113.240 118.670 113.560 ;
        RECT 114.270 112.900 114.530 113.220 ;
        RECT 114.330 111.520 114.470 112.900 ;
        RECT 114.270 111.200 114.530 111.520 ;
        RECT 121.690 109.560 121.830 113.580 ;
        RECT 122.150 112.200 122.290 113.920 ;
        RECT 122.090 111.880 122.350 112.200 ;
        RECT 120.770 109.420 121.830 109.560 ;
        RECT 120.250 107.460 120.510 107.780 ;
        RECT 102.770 105.760 103.030 106.080 ;
        RECT 104.150 105.760 104.410 106.080 ;
        RECT 112.890 105.760 113.150 106.080 ;
        RECT 117.490 105.760 117.750 106.080 ;
        RECT 101.850 104.740 102.110 105.060 ;
        RECT 98.170 103.720 98.430 104.040 ;
        RECT 101.910 103.700 102.050 104.740 ;
        RECT 101.850 103.380 102.110 103.700 ;
        RECT 101.910 103.020 102.050 103.380 ;
        RECT 102.830 103.360 102.970 105.760 ;
        RECT 107.830 105.420 108.090 105.740 ;
        RECT 105.990 104.740 106.250 105.060 ;
        RECT 102.770 103.040 103.030 103.360 ;
        RECT 101.850 102.700 102.110 103.020 ;
        RECT 102.310 102.700 102.570 103.020 ;
        RECT 102.370 100.980 102.510 102.700 ;
        RECT 106.050 100.980 106.190 104.740 ;
        RECT 107.890 104.040 108.030 105.420 ;
        RECT 117.550 105.400 117.690 105.760 ;
        RECT 118.870 105.420 119.130 105.740 ;
        RECT 117.490 105.080 117.750 105.400 ;
        RECT 108.290 104.740 108.550 105.060 ;
        RECT 109.670 104.740 109.930 105.060 ;
        RECT 114.730 104.740 114.990 105.060 ;
        RECT 107.830 103.720 108.090 104.040 ;
        RECT 107.890 100.980 108.030 103.720 ;
        RECT 108.350 102.680 108.490 104.740 ;
        RECT 109.730 103.360 109.870 104.740 ;
        RECT 109.670 103.040 109.930 103.360 ;
        RECT 111.050 103.040 111.310 103.360 ;
        RECT 108.290 102.360 108.550 102.680 ;
        RECT 108.410 101.485 110.290 101.855 ;
        RECT 102.310 100.660 102.570 100.980 ;
        RECT 105.990 100.660 106.250 100.980 ;
        RECT 107.830 100.660 108.090 100.980 ;
        RECT 104.610 99.300 104.870 99.620 ;
        RECT 104.670 88.610 104.810 99.300 ;
        RECT 108.410 96.045 110.290 96.415 ;
        RECT 97.600 86.440 98.820 88.240 ;
        RECT 97.310 86.300 98.820 86.440 ;
        RECT 97.600 84.630 98.820 86.300 ;
        RECT 103.650 86.920 104.870 88.610 ;
        RECT 103.650 84.920 104.880 86.920 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 111.110 86.920 111.250 103.040 ;
        RECT 114.790 101.320 114.930 104.740 ;
        RECT 117.550 103.020 117.690 105.080 ;
        RECT 118.930 103.360 119.070 105.420 ;
        RECT 120.310 103.360 120.450 107.460 ;
        RECT 120.770 105.740 120.910 109.420 ;
        RECT 123.070 108.460 123.210 145.540 ;
        RECT 123.410 142.285 125.290 142.655 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 125.310 140.100 125.570 140.420 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 125.370 138.720 125.510 140.100 ;
        RECT 125.310 138.400 125.570 138.720 ;
        RECT 127.150 138.060 127.410 138.380 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 123.410 136.845 125.290 137.215 ;
        RECT 127.210 136.000 127.350 138.060 ;
        RECT 127.150 135.680 127.410 136.000 ;
        RECT 124.390 135.340 124.650 135.660 ;
        RECT 124.450 133.960 124.590 135.340 ;
        RECT 124.390 133.640 124.650 133.960 ;
        RECT 123.410 131.405 125.290 131.775 ;
        RECT 127.210 130.220 127.350 135.680 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 127.150 129.900 127.410 130.220 ;
        RECT 123.410 125.965 125.290 126.335 ;
        RECT 127.210 125.120 127.350 129.900 ;
        RECT 127.150 124.800 127.410 125.120 ;
        RECT 126.230 124.460 126.490 124.780 ;
        RECT 126.290 123.080 126.430 124.460 ;
        RECT 126.230 122.760 126.490 123.080 ;
        RECT 127.210 122.480 127.350 124.800 ;
        RECT 126.750 122.400 127.350 122.480 ;
        RECT 126.690 122.340 127.350 122.400 ;
        RECT 126.690 122.080 126.950 122.340 ;
        RECT 123.410 120.525 125.290 120.895 ;
        RECT 126.750 119.000 126.890 122.080 ;
        RECT 126.690 118.680 126.950 119.000 ;
        RECT 123.410 115.085 125.290 115.455 ;
        RECT 126.750 114.240 126.890 118.680 ;
        RECT 126.690 113.920 126.950 114.240 ;
        RECT 123.410 109.645 125.290 110.015 ;
        RECT 123.010 108.140 123.270 108.460 ;
        RECT 122.090 107.690 122.350 107.780 ;
        RECT 121.690 107.550 122.350 107.690 ;
        RECT 121.690 106.420 121.830 107.550 ;
        RECT 122.090 107.460 122.350 107.550 ;
        RECT 121.630 106.100 121.890 106.420 ;
        RECT 120.710 105.420 120.970 105.740 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 130.370 104.740 130.630 105.060 ;
        RECT 123.410 104.205 125.290 104.575 ;
        RECT 127.600 103.865 127.880 104.235 ;
        RECT 125.770 103.380 126.030 103.700 ;
        RECT 118.870 103.040 119.130 103.360 ;
        RECT 120.250 103.040 120.510 103.360 ;
        RECT 116.110 102.700 116.370 103.020 ;
        RECT 117.490 102.700 117.750 103.020 ;
        RECT 114.730 101.000 114.990 101.320 ;
        RECT 116.170 100.980 116.310 102.700 ;
        RECT 116.110 100.660 116.370 100.980 ;
        RECT 118.930 100.300 119.070 103.040 ;
        RECT 118.870 99.980 119.130 100.300 ;
        RECT 117.490 99.300 117.750 99.620 ;
        RECT 103.650 84.740 104.870 84.920 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 111.040 84.920 111.320 86.920 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 117.550 86.920 117.690 99.300 ;
        RECT 123.410 98.765 125.290 99.135 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 117.480 84.920 117.760 86.920 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 123.920 86.440 124.200 86.920 ;
        RECT 125.830 86.440 125.970 103.380 ;
        RECT 126.690 102.020 126.950 102.340 ;
        RECT 126.750 101.320 126.890 102.020 ;
        RECT 126.690 101.000 126.950 101.320 ;
        RECT 127.670 100.640 127.810 103.865 ;
        RECT 127.610 100.320 127.870 100.640 ;
        RECT 123.920 86.300 125.970 86.440 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 123.920 84.920 124.200 86.300 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 130.430 86.920 130.570 104.740 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 130.360 84.920 130.640 86.920 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 18.360 215.745 20.340 216.075 ;
        RECT 48.360 215.745 50.340 216.075 ;
        RECT 78.360 215.745 80.340 216.075 ;
        RECT 108.360 215.745 110.340 216.075 ;
        RECT 33.360 213.025 35.340 213.355 ;
        RECT 63.360 213.025 65.340 213.355 ;
        RECT 93.360 213.025 95.340 213.355 ;
        RECT 123.360 213.025 125.340 213.355 ;
        RECT 18.360 210.305 20.340 210.635 ;
        RECT 48.360 210.305 50.340 210.635 ;
        RECT 78.360 210.305 80.340 210.635 ;
        RECT 108.360 210.305 110.340 210.635 ;
        RECT 33.360 207.585 35.340 207.915 ;
        RECT 63.360 207.585 65.340 207.915 ;
        RECT 93.360 207.585 95.340 207.915 ;
        RECT 123.360 207.585 125.340 207.915 ;
        RECT 18.360 204.865 20.340 205.195 ;
        RECT 48.360 204.865 50.340 205.195 ;
        RECT 78.360 204.865 80.340 205.195 ;
        RECT 108.360 204.865 110.340 205.195 ;
        RECT 33.360 202.145 35.340 202.475 ;
        RECT 63.360 202.145 65.340 202.475 ;
        RECT 93.360 202.145 95.340 202.475 ;
        RECT 123.360 202.145 125.340 202.475 ;
        RECT 18.360 199.425 20.340 199.755 ;
        RECT 48.360 199.425 50.340 199.755 ;
        RECT 78.360 199.425 80.340 199.755 ;
        RECT 108.360 199.425 110.340 199.755 ;
        RECT 33.360 196.705 35.340 197.035 ;
        RECT 63.360 196.705 65.340 197.035 ;
        RECT 93.360 196.705 95.340 197.035 ;
        RECT 123.360 196.705 125.340 197.035 ;
        RECT 18.360 193.985 20.340 194.315 ;
        RECT 48.360 193.985 50.340 194.315 ;
        RECT 78.360 193.985 80.340 194.315 ;
        RECT 108.360 193.985 110.340 194.315 ;
        RECT 33.360 191.265 35.340 191.595 ;
        RECT 63.360 191.265 65.340 191.595 ;
        RECT 93.360 191.265 95.340 191.595 ;
        RECT 123.360 191.265 125.340 191.595 ;
        RECT 18.360 188.545 20.340 188.875 ;
        RECT 48.360 188.545 50.340 188.875 ;
        RECT 78.360 188.545 80.340 188.875 ;
        RECT 108.360 188.545 110.340 188.875 ;
        RECT 33.360 185.825 35.340 186.155 ;
        RECT 63.360 185.825 65.340 186.155 ;
        RECT 93.360 185.825 95.340 186.155 ;
        RECT 123.360 185.825 125.340 186.155 ;
        RECT 18.360 183.105 20.340 183.435 ;
        RECT 48.360 183.105 50.340 183.435 ;
        RECT 78.360 183.105 80.340 183.435 ;
        RECT 108.360 183.105 110.340 183.435 ;
        RECT 33.360 180.385 35.340 180.715 ;
        RECT 63.360 180.385 65.340 180.715 ;
        RECT 93.360 180.385 95.340 180.715 ;
        RECT 123.360 180.385 125.340 180.715 ;
        RECT 18.360 177.665 20.340 177.995 ;
        RECT 48.360 177.665 50.340 177.995 ;
        RECT 78.360 177.665 80.340 177.995 ;
        RECT 108.360 177.665 110.340 177.995 ;
        RECT 62.255 176.280 62.585 176.295 ;
        RECT 101.815 176.280 102.145 176.295 ;
        RECT 62.255 175.980 102.145 176.280 ;
        RECT 62.255 175.965 62.585 175.980 ;
        RECT 101.815 175.965 102.145 175.980 ;
        RECT 33.360 174.945 35.340 175.275 ;
        RECT 63.360 174.945 65.340 175.275 ;
        RECT 93.360 174.945 95.340 175.275 ;
        RECT 123.360 174.945 125.340 175.275 ;
        RECT 127.575 174.920 127.905 174.935 ;
        RECT 132.870 174.920 134.870 175.070 ;
        RECT 127.575 174.620 134.870 174.920 ;
        RECT 127.575 174.605 127.905 174.620 ;
        RECT 132.870 174.470 134.870 174.620 ;
        RECT 18.360 172.225 20.340 172.555 ;
        RECT 48.360 172.225 50.340 172.555 ;
        RECT 78.360 172.225 80.340 172.555 ;
        RECT 108.360 172.225 110.340 172.555 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 64.095 172.200 64.425 172.215 ;
        RECT 70.535 172.200 70.865 172.215 ;
        RECT 64.095 171.900 70.865 172.200 ;
        RECT 64.095 171.885 64.425 171.900 ;
        RECT 70.535 171.885 70.865 171.900 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 33.360 169.505 35.340 169.835 ;
        RECT 63.360 169.505 65.340 169.835 ;
        RECT 93.360 169.505 95.340 169.835 ;
        RECT 123.360 169.505 125.340 169.835 ;
        RECT 18.360 166.785 20.340 167.115 ;
        RECT 48.360 166.785 50.340 167.115 ;
        RECT 78.360 166.785 80.340 167.115 ;
        RECT 108.360 166.785 110.340 167.115 ;
        RECT 33.360 164.065 35.340 164.395 ;
        RECT 63.360 164.065 65.340 164.395 ;
        RECT 93.360 164.065 95.340 164.395 ;
        RECT 123.360 164.065 125.340 164.395 ;
        RECT 18.360 161.345 20.340 161.675 ;
        RECT 48.360 161.345 50.340 161.675 ;
        RECT 78.360 161.345 80.340 161.675 ;
        RECT 108.360 161.345 110.340 161.675 ;
        RECT 36.495 159.960 36.825 159.975 ;
        RECT 38.540 159.960 38.920 159.970 ;
        RECT 36.495 159.660 38.920 159.960 ;
        RECT 36.495 159.645 36.825 159.660 ;
        RECT 38.540 159.650 38.920 159.660 ;
        RECT 33.360 158.625 35.340 158.955 ;
        RECT 63.360 158.625 65.340 158.955 ;
        RECT 93.360 158.625 95.340 158.955 ;
        RECT 123.360 158.625 125.340 158.955 ;
        RECT 18.360 155.905 20.340 156.235 ;
        RECT 48.360 155.905 50.340 156.235 ;
        RECT 78.360 155.905 80.340 156.235 ;
        RECT 108.360 155.905 110.340 156.235 ;
        RECT 46.615 155.200 46.945 155.215 ;
        RECT 70.995 155.200 71.325 155.215 ;
        RECT 72.835 155.200 73.165 155.215 ;
        RECT 46.615 154.900 73.165 155.200 ;
        RECT 46.615 154.885 46.945 154.900 ;
        RECT 70.995 154.885 71.325 154.900 ;
        RECT 72.835 154.885 73.165 154.900 ;
        RECT 55.355 154.520 55.685 154.535 ;
        RECT 69.155 154.520 69.485 154.535 ;
        RECT 73.755 154.520 74.085 154.535 ;
        RECT 55.355 154.220 74.085 154.520 ;
        RECT 55.355 154.205 55.685 154.220 ;
        RECT 69.155 154.205 69.485 154.220 ;
        RECT 73.755 154.205 74.085 154.220 ;
        RECT 33.360 153.185 35.340 153.515 ;
        RECT 63.360 153.185 65.340 153.515 ;
        RECT 93.360 153.185 95.340 153.515 ;
        RECT 123.360 153.185 125.340 153.515 ;
        RECT 18.360 150.465 20.340 150.795 ;
        RECT 48.360 150.465 50.340 150.795 ;
        RECT 78.360 150.465 80.340 150.795 ;
        RECT 108.360 150.465 110.340 150.795 ;
        RECT 35.115 149.080 35.445 149.095 ;
        RECT 35.115 148.780 36.120 149.080 ;
        RECT 35.115 148.765 35.445 148.780 ;
        RECT 33.360 147.745 35.340 148.075 ;
        RECT 35.115 147.040 35.445 147.055 ;
        RECT 35.820 147.040 36.120 148.780 ;
        RECT 63.360 147.745 65.340 148.075 ;
        RECT 93.360 147.745 95.340 148.075 ;
        RECT 123.360 147.745 125.340 148.075 ;
        RECT 35.115 146.740 36.120 147.040 ;
        RECT 38.540 147.040 38.920 147.050 ;
        RECT 62.255 147.040 62.585 147.055 ;
        RECT 96.295 147.040 96.625 147.055 ;
        RECT 38.540 146.740 96.625 147.040 ;
        RECT 35.115 146.725 35.445 146.740 ;
        RECT 38.540 146.730 38.920 146.740 ;
        RECT 62.255 146.725 62.585 146.740 ;
        RECT 96.295 146.725 96.625 146.740 ;
        RECT 18.360 145.025 20.340 145.355 ;
        RECT 48.360 145.025 50.340 145.355 ;
        RECT 78.360 145.025 80.340 145.355 ;
        RECT 108.360 145.025 110.340 145.355 ;
        RECT 33.360 142.305 35.340 142.635 ;
        RECT 63.360 142.305 65.340 142.635 ;
        RECT 93.360 142.305 95.340 142.635 ;
        RECT 123.360 142.305 125.340 142.635 ;
        RECT 18.360 139.585 20.340 139.915 ;
        RECT 48.360 139.585 50.340 139.915 ;
        RECT 78.360 139.585 80.340 139.915 ;
        RECT 108.360 139.585 110.340 139.915 ;
        RECT 132.510 139.560 135.210 140.035 ;
        RECT 120.920 139.260 135.210 139.560 ;
        RECT 68.695 138.880 69.025 138.895 ;
        RECT 120.920 138.880 121.220 139.260 ;
        RECT 68.695 138.580 121.220 138.880 ;
        RECT 68.695 138.565 69.025 138.580 ;
        RECT 132.510 138.165 135.210 139.260 ;
        RECT 33.360 136.865 35.340 137.195 ;
        RECT 63.360 136.865 65.340 137.195 ;
        RECT 93.360 136.865 95.340 137.195 ;
        RECT 123.360 136.865 125.340 137.195 ;
        RECT 18.360 134.145 20.340 134.475 ;
        RECT 48.360 134.145 50.340 134.475 ;
        RECT 78.360 134.145 80.340 134.475 ;
        RECT 108.360 134.145 110.340 134.475 ;
        RECT 33.360 131.425 35.340 131.755 ;
        RECT 63.360 131.425 65.340 131.755 ;
        RECT 93.360 131.425 95.340 131.755 ;
        RECT 123.360 131.425 125.340 131.755 ;
        RECT 51.215 130.040 51.545 130.055 ;
        RECT 80.195 130.040 80.525 130.055 ;
        RECT 51.215 129.740 80.525 130.040 ;
        RECT 51.215 129.725 51.545 129.740 ;
        RECT 80.195 129.725 80.525 129.740 ;
        RECT 18.360 128.705 20.340 129.035 ;
        RECT 48.360 128.705 50.340 129.035 ;
        RECT 78.360 128.705 80.340 129.035 ;
        RECT 108.360 128.705 110.340 129.035 ;
        RECT 33.360 125.985 35.340 126.315 ;
        RECT 63.360 125.985 65.340 126.315 ;
        RECT 93.360 125.985 95.340 126.315 ;
        RECT 123.360 125.985 125.340 126.315 ;
        RECT 18.360 123.265 20.340 123.595 ;
        RECT 48.360 123.265 50.340 123.595 ;
        RECT 78.360 123.265 80.340 123.595 ;
        RECT 108.360 123.265 110.340 123.595 ;
        RECT 33.360 120.545 35.340 120.875 ;
        RECT 63.360 120.545 65.340 120.875 ;
        RECT 93.360 120.545 95.340 120.875 ;
        RECT 123.360 120.545 125.340 120.875 ;
        RECT 18.360 117.825 20.340 118.155 ;
        RECT 48.360 117.825 50.340 118.155 ;
        RECT 78.360 117.825 80.340 118.155 ;
        RECT 108.360 117.825 110.340 118.155 ;
        RECT 33.360 115.105 35.340 115.435 ;
        RECT 63.360 115.105 65.340 115.435 ;
        RECT 93.360 115.105 95.340 115.435 ;
        RECT 123.360 115.105 125.340 115.435 ;
        RECT 18.360 112.385 20.340 112.715 ;
        RECT 48.360 112.385 50.340 112.715 ;
        RECT 78.360 112.385 80.340 112.715 ;
        RECT 108.360 112.385 110.340 112.715 ;
        RECT 33.360 109.665 35.340 109.995 ;
        RECT 63.360 109.665 65.340 109.995 ;
        RECT 93.360 109.665 95.340 109.995 ;
        RECT 123.360 109.665 125.340 109.995 ;
        RECT 18.360 106.945 20.340 107.275 ;
        RECT 48.360 106.945 50.340 107.275 ;
        RECT 78.360 106.945 80.340 107.275 ;
        RECT 108.360 106.945 110.340 107.275 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 33.360 104.225 35.340 104.555 ;
        RECT 63.360 104.225 65.340 104.555 ;
        RECT 93.360 104.225 95.340 104.555 ;
        RECT 123.360 104.225 125.340 104.555 ;
        RECT 127.575 104.200 127.905 104.215 ;
        RECT 132.870 104.200 134.870 104.350 ;
        RECT 127.575 103.900 134.870 104.200 ;
        RECT 127.575 103.885 127.905 103.900 ;
        RECT 132.870 103.750 134.870 103.900 ;
        RECT 18.360 101.505 20.340 101.835 ;
        RECT 48.360 101.505 50.340 101.835 ;
        RECT 78.360 101.505 80.340 101.835 ;
        RECT 108.360 101.505 110.340 101.835 ;
        RECT 33.360 98.785 35.340 99.115 ;
        RECT 63.360 98.785 65.340 99.115 ;
        RECT 93.360 98.785 95.340 99.115 ;
        RECT 123.360 98.785 125.340 99.115 ;
        RECT 18.360 96.065 20.340 96.395 ;
        RECT 48.360 96.065 50.340 96.395 ;
        RECT 78.360 96.065 80.340 96.395 ;
        RECT 108.360 96.065 110.340 96.395 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 18.350 95.990 20.350 216.150 ;
        RECT 33.350 95.990 35.350 216.150 ;
        RECT 38.565 159.645 38.895 159.975 ;
        RECT 38.580 147.055 38.880 159.645 ;
        RECT 38.565 146.725 38.895 147.055 ;
        RECT 48.350 95.990 50.350 216.150 ;
        RECT 63.350 95.990 65.350 216.150 ;
        RECT 78.350 95.990 80.350 216.150 ;
        RECT 93.350 95.990 95.350 216.150 ;
        RECT 108.350 95.990 110.350 216.150 ;
        RECT 123.350 99.720 125.350 216.150 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 125.350 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 125.350 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

